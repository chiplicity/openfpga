magic
tech EFS8A
magscale 1 2
timestamp 1604337270
<< locali >>
rect 949 12087 983 15861
rect 6469 13855 6503 13957
rect 10701 12155 10735 12325
rect 20453 12155 20487 12325
rect 3249 11543 3283 11849
rect 12817 10591 12851 10761
rect 15209 9367 15243 9469
rect 12817 4471 12851 4777
rect 15209 2839 15243 2941
rect 19349 2839 19383 3145
<< viali >>
rect 24593 19805 24627 19839
rect 24593 19261 24627 19295
rect 25145 19261 25179 19295
rect 24777 19125 24811 19159
rect 23489 18785 23523 18819
rect 24593 18785 24627 18819
rect 22477 18717 22511 18751
rect 23673 18581 23707 18615
rect 24777 18581 24811 18615
rect 25145 18377 25179 18411
rect 1409 18173 1443 18207
rect 24593 18173 24627 18207
rect 1593 18037 1627 18071
rect 2053 18037 2087 18071
rect 20177 18037 20211 18071
rect 22569 18037 22603 18071
rect 23857 18037 23891 18071
rect 24409 18037 24443 18071
rect 24777 18037 24811 18071
rect 22937 17833 22971 17867
rect 1409 17697 1443 17731
rect 2513 17697 2547 17731
rect 22753 17697 22787 17731
rect 24593 17697 24627 17731
rect 2053 17629 2087 17663
rect 19533 17629 19567 17663
rect 21373 17629 21407 17663
rect 23029 17629 23063 17663
rect 1593 17493 1627 17527
rect 2697 17493 2731 17527
rect 22109 17493 22143 17527
rect 22477 17493 22511 17527
rect 24777 17493 24811 17527
rect 2421 17289 2455 17323
rect 23029 17289 23063 17323
rect 2697 17221 2731 17255
rect 22109 17221 22143 17255
rect 23397 17221 23431 17255
rect 25145 17221 25179 17255
rect 21557 17153 21591 17187
rect 1409 17085 1443 17119
rect 2513 17085 2547 17119
rect 20913 17085 20947 17119
rect 23673 17085 23707 17119
rect 24961 17085 24995 17119
rect 25513 17085 25547 17119
rect 22385 17017 22419 17051
rect 22661 17017 22695 17051
rect 23949 17017 23983 17051
rect 1593 16949 1627 16983
rect 2053 16949 2087 16983
rect 3157 16949 3191 16983
rect 19901 16949 19935 16983
rect 20821 16949 20855 16983
rect 21097 16949 21131 16983
rect 21833 16949 21867 16983
rect 22569 16949 22603 16983
rect 24593 16949 24627 16983
rect 2053 16745 2087 16779
rect 2697 16745 2731 16779
rect 19809 16745 19843 16779
rect 22109 16745 22143 16779
rect 23949 16745 23983 16779
rect 25237 16745 25271 16779
rect 4629 16677 4663 16711
rect 22836 16677 22870 16711
rect 1409 16609 1443 16643
rect 2513 16609 2547 16643
rect 4445 16609 4479 16643
rect 9965 16609 9999 16643
rect 16313 16609 16347 16643
rect 17601 16609 17635 16643
rect 18797 16609 18831 16643
rect 21465 16609 21499 16643
rect 22477 16609 22511 16643
rect 25053 16609 25087 16643
rect 4721 16541 4755 16575
rect 22569 16541 22603 16575
rect 21189 16473 21223 16507
rect 1593 16405 1627 16439
rect 2421 16405 2455 16439
rect 3157 16405 3191 16439
rect 4169 16405 4203 16439
rect 10517 16405 10551 16439
rect 14289 16405 14323 16439
rect 21649 16405 21683 16439
rect 3985 16201 4019 16235
rect 22477 16201 22511 16235
rect 2697 16133 2731 16167
rect 4169 16133 4203 16167
rect 10517 16133 10551 16167
rect 14289 16133 14323 16167
rect 2053 16065 2087 16099
rect 14841 16065 14875 16099
rect 1409 15997 1443 16031
rect 2513 15997 2547 16031
rect 5825 15997 5859 16031
rect 10333 15997 10367 16031
rect 11069 15997 11103 16031
rect 14105 15997 14139 16031
rect 19993 15997 20027 16031
rect 21097 15997 21131 16031
rect 23673 15997 23707 16031
rect 23940 15997 23974 16031
rect 3157 15929 3191 15963
rect 4445 15929 4479 15963
rect 4629 15929 4663 15963
rect 4721 15929 4755 15963
rect 5089 15929 5123 15963
rect 9965 15929 9999 15963
rect 10793 15929 10827 15963
rect 10977 15929 11011 15963
rect 14565 15929 14599 15963
rect 14749 15929 14783 15963
rect 21364 15929 21398 15963
rect 949 15861 983 15895
rect 1593 15861 1627 15895
rect 2421 15861 2455 15895
rect 3617 15861 3651 15895
rect 5457 15861 5491 15895
rect 6285 15861 6319 15895
rect 6653 15861 6687 15895
rect 16313 15861 16347 15895
rect 18981 15861 19015 15895
rect 20177 15861 20211 15895
rect 20637 15861 20671 15895
rect 20913 15861 20947 15895
rect 23121 15861 23155 15895
rect 23397 15861 23431 15895
rect 25053 15861 25087 15895
rect 25605 15861 25639 15895
rect 2973 15657 3007 15691
rect 11897 15657 11931 15691
rect 14289 15657 14323 15691
rect 19809 15657 19843 15691
rect 22937 15657 22971 15691
rect 23765 15657 23799 15691
rect 4905 15589 4939 15623
rect 9965 15589 9999 15623
rect 10762 15589 10796 15623
rect 15669 15589 15703 15623
rect 15853 15589 15887 15623
rect 20729 15589 20763 15623
rect 18153 15521 18187 15555
rect 19901 15521 19935 15555
rect 21169 15521 21203 15555
rect 24216 15521 24250 15555
rect 2973 15453 3007 15487
rect 3065 15453 3099 15487
rect 4905 15453 4939 15487
rect 4997 15453 5031 15487
rect 5917 15453 5951 15487
rect 7021 15453 7055 15487
rect 8493 15453 8527 15487
rect 10517 15453 10551 15487
rect 13001 15453 13035 15487
rect 15945 15453 15979 15487
rect 17141 15453 17175 15487
rect 19717 15453 19751 15487
rect 20913 15453 20947 15487
rect 23949 15453 23983 15487
rect 2329 15385 2363 15419
rect 3525 15385 3559 15419
rect 4445 15385 4479 15419
rect 6745 15385 6779 15419
rect 19349 15385 19383 15419
rect 1869 15317 1903 15351
rect 2513 15317 2547 15351
rect 3893 15317 3927 15351
rect 5365 15317 5399 15351
rect 5825 15317 5859 15351
rect 6469 15317 6503 15351
rect 12541 15317 12575 15351
rect 15393 15317 15427 15351
rect 18337 15317 18371 15351
rect 20361 15317 20395 15351
rect 22293 15317 22327 15351
rect 23213 15317 23247 15351
rect 25329 15317 25363 15351
rect 2881 15113 2915 15147
rect 4353 15113 4387 15147
rect 5365 15113 5399 15147
rect 9689 15113 9723 15147
rect 9965 15113 9999 15147
rect 11805 15113 11839 15147
rect 14657 15113 14691 15147
rect 16497 15113 16531 15147
rect 17049 15113 17083 15147
rect 18429 15113 18463 15147
rect 19349 15113 19383 15147
rect 21005 15113 21039 15147
rect 21925 15113 21959 15147
rect 12541 15045 12575 15079
rect 24501 15045 24535 15079
rect 2973 14977 3007 15011
rect 10517 14977 10551 15011
rect 11253 14977 11287 15011
rect 13001 14977 13035 15011
rect 14105 14977 14139 15011
rect 23121 14977 23155 15011
rect 25053 14977 25087 15011
rect 1409 14909 1443 14943
rect 5457 14909 5491 14943
rect 6193 14909 6227 14943
rect 6837 14909 6871 14943
rect 10241 14909 10275 14943
rect 12265 14909 12299 14943
rect 13093 14909 13127 14943
rect 15117 14909 15151 14943
rect 18521 14909 18555 14943
rect 19625 14909 19659 14943
rect 22109 14909 22143 14943
rect 23949 14909 23983 14943
rect 2053 14841 2087 14875
rect 2513 14841 2547 14875
rect 3218 14841 3252 14875
rect 5733 14841 5767 14875
rect 7082 14841 7116 14875
rect 10425 14841 10459 14875
rect 10977 14841 11011 14875
rect 13001 14841 13035 14875
rect 15362 14841 15396 14875
rect 17877 14841 17911 14875
rect 19892 14841 19926 14875
rect 22385 14841 22419 14875
rect 24317 14841 24351 14875
rect 24777 14841 24811 14875
rect 24961 14841 24995 14875
rect 1593 14773 1627 14807
rect 4997 14773 5031 14807
rect 6653 14773 6687 14807
rect 8217 14773 8251 14807
rect 9321 14773 9355 14807
rect 15025 14773 15059 14807
rect 18705 14773 18739 14807
rect 21649 14773 21683 14807
rect 23397 14773 23431 14807
rect 3893 14569 3927 14603
rect 7757 14569 7791 14603
rect 9965 14569 9999 14603
rect 10517 14569 10551 14603
rect 15761 14569 15795 14603
rect 19349 14569 19383 14603
rect 20729 14569 20763 14603
rect 21465 14569 21499 14603
rect 22109 14569 22143 14603
rect 24593 14569 24627 14603
rect 2789 14501 2823 14535
rect 2973 14501 3007 14535
rect 3065 14501 3099 14535
rect 4966 14501 5000 14535
rect 7573 14501 7607 14535
rect 7849 14501 7883 14535
rect 10977 14501 11011 14535
rect 11161 14501 11195 14535
rect 12725 14501 12759 14535
rect 16558 14501 16592 14535
rect 21281 14501 21315 14535
rect 25329 14501 25363 14535
rect 12817 14433 12851 14467
rect 16313 14433 16347 14467
rect 19717 14433 19751 14467
rect 22569 14433 22603 14467
rect 22836 14433 22870 14467
rect 25053 14433 25087 14467
rect 1409 14365 1443 14399
rect 4721 14365 4755 14399
rect 11253 14365 11287 14399
rect 12725 14365 12759 14399
rect 13737 14365 13771 14399
rect 15301 14365 15335 14399
rect 21557 14365 21591 14399
rect 2329 14297 2363 14331
rect 7297 14297 7331 14331
rect 10701 14297 10735 14331
rect 16129 14297 16163 14331
rect 21005 14297 21039 14331
rect 1961 14229 1995 14263
rect 2513 14229 2547 14263
rect 3433 14229 3467 14263
rect 4261 14229 4295 14263
rect 6101 14229 6135 14263
rect 6837 14229 6871 14263
rect 8309 14229 8343 14263
rect 8585 14229 8619 14263
rect 8953 14229 8987 14263
rect 9413 14229 9447 14263
rect 11621 14229 11655 14263
rect 11989 14229 12023 14263
rect 12265 14229 12299 14263
rect 13185 14229 13219 14263
rect 17693 14229 17727 14263
rect 18521 14229 18555 14263
rect 19901 14229 19935 14263
rect 20269 14229 20303 14263
rect 23949 14229 23983 14263
rect 1685 14025 1719 14059
rect 3709 14025 3743 14059
rect 4353 14025 4387 14059
rect 5641 14025 5675 14059
rect 7205 14025 7239 14059
rect 10793 14025 10827 14059
rect 11805 14025 11839 14059
rect 12265 14025 12299 14059
rect 13829 14025 13863 14059
rect 14841 14025 14875 14059
rect 16313 14025 16347 14059
rect 21373 14025 21407 14059
rect 21833 14025 21867 14059
rect 25513 14025 25547 14059
rect 3157 13957 3191 13991
rect 5273 13957 5307 13991
rect 6469 13957 6503 13991
rect 6561 13957 6595 13991
rect 9873 13957 9907 13991
rect 18521 13957 18555 13991
rect 20821 13957 20855 13991
rect 22109 13957 22143 13991
rect 1777 13889 1811 13923
rect 4905 13889 4939 13923
rect 6285 13889 6319 13923
rect 11253 13889 11287 13923
rect 14933 13889 14967 13923
rect 22477 13889 22511 13923
rect 22661 13889 22695 13923
rect 2044 13821 2078 13855
rect 4629 13821 4663 13855
rect 6469 13821 6503 13855
rect 7297 13821 7331 13855
rect 7564 13821 7598 13855
rect 9505 13821 9539 13855
rect 12449 13821 12483 13855
rect 12716 13821 12750 13855
rect 15189 13821 15223 13855
rect 18337 13821 18371 13855
rect 18889 13821 18923 13855
rect 19441 13821 19475 13855
rect 24133 13821 24167 13855
rect 24400 13821 24434 13855
rect 10241 13753 10275 13787
rect 11253 13753 11287 13787
rect 11345 13753 11379 13787
rect 19686 13753 19720 13787
rect 22569 13753 22603 13787
rect 23489 13753 23523 13787
rect 4169 13685 4203 13719
rect 4813 13685 4847 13719
rect 8677 13685 8711 13719
rect 10609 13685 10643 13719
rect 14381 13685 14415 13719
rect 16957 13685 16991 13719
rect 19349 13685 19383 13719
rect 23029 13685 23063 13719
rect 23949 13685 23983 13719
rect 1777 13481 1811 13515
rect 3709 13481 3743 13515
rect 5089 13481 5123 13515
rect 6653 13481 6687 13515
rect 7021 13481 7055 13515
rect 8953 13481 8987 13515
rect 11069 13481 11103 13515
rect 11621 13481 11655 13515
rect 12081 13481 12115 13515
rect 16129 13481 16163 13515
rect 16589 13481 16623 13515
rect 20269 13481 20303 13515
rect 20729 13481 20763 13515
rect 21465 13481 21499 13515
rect 24685 13481 24719 13515
rect 2789 13413 2823 13447
rect 4629 13413 4663 13447
rect 6009 13413 6043 13447
rect 6193 13413 6227 13447
rect 7757 13413 7791 13447
rect 8585 13413 8619 13447
rect 16221 13413 16255 13447
rect 17049 13413 17083 13447
rect 17408 13413 17442 13447
rect 23020 13413 23054 13447
rect 2605 13345 2639 13379
rect 4445 13345 4479 13379
rect 7573 13345 7607 13379
rect 7849 13345 7883 13379
rect 9945 13345 9979 13379
rect 12541 13345 12575 13379
rect 12725 13345 12759 13379
rect 12981 13345 13015 13379
rect 17141 13345 17175 13379
rect 19717 13345 19751 13379
rect 21281 13345 21315 13379
rect 22109 13345 22143 13379
rect 25237 13345 25271 13379
rect 2881 13277 2915 13311
rect 4721 13277 4755 13311
rect 6285 13277 6319 13311
rect 9689 13277 9723 13311
rect 16129 13277 16163 13311
rect 21557 13277 21591 13311
rect 22753 13277 22787 13311
rect 4169 13209 4203 13243
rect 5733 13209 5767 13243
rect 7297 13209 7331 13243
rect 15669 13209 15703 13243
rect 2329 13141 2363 13175
rect 3249 13141 3283 13175
rect 5457 13141 5491 13175
rect 8309 13141 8343 13175
rect 9505 13141 9539 13175
rect 14105 13141 14139 13175
rect 14933 13141 14967 13175
rect 18521 13141 18555 13175
rect 19441 13141 19475 13175
rect 19901 13141 19935 13175
rect 21005 13141 21039 13175
rect 22661 13141 22695 13175
rect 24133 13141 24167 13175
rect 25053 13141 25087 13175
rect 25421 13141 25455 13175
rect 1685 12937 1719 12971
rect 1961 12937 1995 12971
rect 3525 12937 3559 12971
rect 4629 12937 4663 12971
rect 5273 12937 5307 12971
rect 7481 12937 7515 12971
rect 9413 12937 9447 12971
rect 10885 12937 10919 12971
rect 13553 12937 13587 12971
rect 14381 12937 14415 12971
rect 15945 12937 15979 12971
rect 21833 12937 21867 12971
rect 22201 12937 22235 12971
rect 23397 12937 23431 12971
rect 24041 12937 24075 12971
rect 25237 12937 25271 12971
rect 25697 12937 25731 12971
rect 3709 12869 3743 12903
rect 12541 12869 12575 12903
rect 15669 12869 15703 12903
rect 16221 12869 16255 12903
rect 18429 12869 18463 12903
rect 2421 12801 2455 12835
rect 4169 12801 4203 12835
rect 4261 12801 4295 12835
rect 5641 12801 5675 12835
rect 7849 12801 7883 12835
rect 8033 12801 8067 12835
rect 11437 12801 11471 12835
rect 11897 12801 11931 12835
rect 13001 12801 13035 12835
rect 14197 12801 14231 12835
rect 14749 12801 14783 12835
rect 16589 12801 16623 12835
rect 16773 12801 16807 12835
rect 18797 12801 18831 12835
rect 22937 12801 22971 12835
rect 24593 12801 24627 12835
rect 5089 12733 5123 12767
rect 5825 12733 5859 12767
rect 6837 12733 6871 12767
rect 14933 12733 14967 12767
rect 19809 12733 19843 12767
rect 19901 12733 19935 12767
rect 20168 12733 20202 12767
rect 22385 12733 22419 12767
rect 24317 12733 24351 12767
rect 25513 12733 25547 12767
rect 26065 12733 26099 12767
rect 2513 12665 2547 12699
rect 4169 12665 4203 12699
rect 5733 12665 5767 12699
rect 6285 12665 6319 12699
rect 6653 12665 6687 12699
rect 8278 12665 8312 12699
rect 10057 12665 10091 12699
rect 11161 12665 11195 12699
rect 13093 12665 13127 12699
rect 14841 12665 14875 12699
rect 16681 12665 16715 12699
rect 17785 12665 17819 12699
rect 18889 12665 18923 12699
rect 18981 12665 19015 12699
rect 19441 12665 19475 12699
rect 2421 12597 2455 12631
rect 2973 12597 3007 12631
rect 7021 12597 7055 12631
rect 10701 12597 10735 12631
rect 11345 12597 11379 12631
rect 12265 12597 12299 12631
rect 13001 12597 13035 12631
rect 17233 12597 17267 12631
rect 21281 12597 21315 12631
rect 22569 12597 22603 12631
rect 24501 12597 24535 12631
rect 2789 12393 2823 12427
rect 3893 12393 3927 12427
rect 7021 12393 7055 12427
rect 8309 12393 8343 12427
rect 9321 12393 9355 12427
rect 12909 12393 12943 12427
rect 13461 12393 13495 12427
rect 14749 12393 14783 12427
rect 16405 12393 16439 12427
rect 18797 12393 18831 12427
rect 19165 12393 19199 12427
rect 21465 12393 21499 12427
rect 22845 12393 22879 12427
rect 24501 12393 24535 12427
rect 4629 12325 4663 12359
rect 6193 12325 6227 12359
rect 7757 12325 7791 12359
rect 7849 12325 7883 12359
rect 9965 12325 9999 12359
rect 10701 12325 10735 12359
rect 14197 12325 14231 12359
rect 17040 12325 17074 12359
rect 19809 12325 19843 12359
rect 20453 12325 20487 12359
rect 21557 12325 21591 12359
rect 23949 12325 23983 12359
rect 25237 12325 25271 12359
rect 1409 12257 1443 12291
rect 1676 12257 1710 12291
rect 4445 12257 4479 12291
rect 5549 12257 5583 12291
rect 6009 12257 6043 12291
rect 9689 12257 9723 12291
rect 4721 12189 4755 12223
rect 5181 12189 5215 12223
rect 6285 12189 6319 12223
rect 7757 12189 7791 12223
rect 11244 12257 11278 12291
rect 15025 12257 15059 12291
rect 15301 12257 15335 12291
rect 16773 12257 16807 12291
rect 19901 12257 19935 12291
rect 10977 12189 11011 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 15577 12189 15611 12223
rect 19809 12189 19843 12223
rect 21281 12257 21315 12291
rect 23305 12257 23339 12291
rect 24961 12257 24995 12291
rect 23857 12189 23891 12223
rect 24041 12189 24075 12223
rect 4169 12121 4203 12155
rect 5733 12121 5767 12155
rect 7297 12121 7331 12155
rect 8585 12121 8619 12155
rect 10701 12121 10735 12155
rect 10793 12121 10827 12155
rect 13737 12121 13771 12155
rect 20453 12121 20487 12155
rect 21005 12121 21039 12155
rect 22017 12121 22051 12155
rect 23489 12121 23523 12155
rect 949 12053 983 12087
rect 3433 12053 3467 12087
rect 6653 12053 6687 12087
rect 8953 12053 8987 12087
rect 10425 12053 10459 12087
rect 12357 12053 12391 12087
rect 16037 12053 16071 12087
rect 18153 12053 18187 12087
rect 19349 12053 19383 12087
rect 20361 12053 20395 12087
rect 20729 12053 20763 12087
rect 22293 12053 22327 12087
rect 1593 11849 1627 11883
rect 3157 11849 3191 11883
rect 3249 11849 3283 11883
rect 3525 11849 3559 11883
rect 7389 11849 7423 11883
rect 10885 11849 10919 11883
rect 11805 11849 11839 11883
rect 12909 11849 12943 11883
rect 14749 11849 14783 11883
rect 15669 11849 15703 11883
rect 17785 11849 17819 11883
rect 18981 11849 19015 11883
rect 21189 11849 21223 11883
rect 21741 11849 21775 11883
rect 22109 11849 22143 11883
rect 24777 11849 24811 11883
rect 25421 11849 25455 11883
rect 1869 11781 1903 11815
rect 2237 11713 2271 11747
rect 2329 11577 2363 11611
rect 2421 11577 2455 11611
rect 8953 11781 8987 11815
rect 16497 11781 16531 11815
rect 23765 11781 23799 11815
rect 25145 11781 25179 11815
rect 7757 11713 7791 11747
rect 7941 11713 7975 11747
rect 9321 11713 9355 11747
rect 9505 11713 9539 11747
rect 9965 11713 9999 11747
rect 11345 11713 11379 11747
rect 16957 11713 16991 11747
rect 24317 11713 24351 11747
rect 3985 11645 4019 11679
rect 4241 11645 4275 11679
rect 7205 11645 7239 11679
rect 8401 11645 8435 11679
rect 8769 11645 8803 11679
rect 13369 11645 13403 11679
rect 13636 11645 13670 11679
rect 18061 11645 18095 11679
rect 19625 11645 19659 11679
rect 19809 11645 19843 11679
rect 22293 11645 22327 11679
rect 23489 11645 23523 11679
rect 25237 11645 25271 11679
rect 25789 11645 25823 11679
rect 3893 11577 3927 11611
rect 6561 11577 6595 11611
rect 7849 11577 7883 11611
rect 10701 11577 10735 11611
rect 11437 11577 11471 11611
rect 13277 11577 13311 11611
rect 16313 11577 16347 11611
rect 17049 11577 17083 11611
rect 20054 11577 20088 11611
rect 23121 11577 23155 11611
rect 24041 11577 24075 11611
rect 3249 11509 3283 11543
rect 5365 11509 5399 11543
rect 5917 11509 5951 11543
rect 9413 11509 9447 11543
rect 10333 11509 10367 11543
rect 11345 11509 11379 11543
rect 12265 11509 12299 11543
rect 16957 11509 16991 11543
rect 17509 11509 17543 11543
rect 18245 11509 18279 11543
rect 19349 11509 19383 11543
rect 22477 11509 22511 11543
rect 24225 11509 24259 11543
rect 1961 11305 1995 11339
rect 3525 11305 3559 11339
rect 7021 11305 7055 11339
rect 8861 11305 8895 11339
rect 11437 11305 11471 11339
rect 13185 11305 13219 11339
rect 14105 11305 14139 11339
rect 17141 11305 17175 11339
rect 17969 11305 18003 11339
rect 18889 11305 18923 11339
rect 19349 11305 19383 11339
rect 20269 11305 20303 11339
rect 20729 11305 20763 11339
rect 21649 11305 21683 11339
rect 24685 11305 24719 11339
rect 25053 11305 25087 11339
rect 25421 11305 25455 11339
rect 2973 11237 3007 11271
rect 3801 11237 3835 11271
rect 4261 11237 4295 11271
rect 4721 11237 4755 11271
rect 5264 11237 5298 11271
rect 7389 11237 7423 11271
rect 8033 11237 8067 11271
rect 8125 11237 8159 11271
rect 10241 11237 10275 11271
rect 15577 11237 15611 11271
rect 16221 11237 16255 11271
rect 17233 11237 17267 11271
rect 21189 11237 21223 11271
rect 22661 11237 22695 11271
rect 23020 11237 23054 11271
rect 2329 11169 2363 11203
rect 3065 11169 3099 11203
rect 10057 11169 10091 11203
rect 12061 11169 12095 11203
rect 15301 11169 15335 11203
rect 18153 11169 18187 11203
rect 19717 11169 19751 11203
rect 20913 11169 20947 11203
rect 25237 11169 25271 11203
rect 1409 11101 1443 11135
rect 2973 11101 3007 11135
rect 4997 11101 5031 11135
rect 8033 11101 8067 11135
rect 9505 11101 9539 11135
rect 10333 11101 10367 11135
rect 11069 11101 11103 11135
rect 11805 11101 11839 11135
rect 13829 11101 13863 11135
rect 17141 11101 17175 11135
rect 18337 11101 18371 11135
rect 22753 11101 22787 11135
rect 2513 11033 2547 11067
rect 6377 11033 6411 11067
rect 7573 11033 7607 11067
rect 9781 11033 9815 11067
rect 14473 11033 14507 11067
rect 15117 11033 15151 11067
rect 16681 11033 16715 11067
rect 17601 11033 17635 11067
rect 19901 11033 19935 11067
rect 8585 10965 8619 10999
rect 22109 10965 22143 10999
rect 24133 10965 24167 10999
rect 2237 10761 2271 10795
rect 3985 10761 4019 10795
rect 4997 10761 5031 10795
rect 6193 10761 6227 10795
rect 6653 10761 6687 10795
rect 7849 10761 7883 10795
rect 10885 10761 10919 10795
rect 12817 10761 12851 10795
rect 12909 10761 12943 10795
rect 14565 10761 14599 10795
rect 16497 10761 16531 10795
rect 20729 10761 20763 10795
rect 2421 10693 2455 10727
rect 8125 10693 8159 10727
rect 11897 10693 11931 10727
rect 2789 10625 2823 10659
rect 2973 10625 3007 10659
rect 4537 10625 4571 10659
rect 5733 10625 5767 10659
rect 11437 10625 11471 10659
rect 13185 10693 13219 10727
rect 15117 10693 15151 10727
rect 22109 10693 22143 10727
rect 13737 10625 13771 10659
rect 14105 10625 14139 10659
rect 15669 10625 15703 10659
rect 22661 10625 22695 10659
rect 3801 10557 3835 10591
rect 4261 10557 4295 10591
rect 5457 10557 5491 10591
rect 7021 10557 7055 10591
rect 8309 10557 8343 10591
rect 8576 10557 8610 10591
rect 12817 10557 12851 10591
rect 13461 10557 13495 10591
rect 15393 10557 15427 10591
rect 16589 10557 16623 10591
rect 18061 10557 18095 10591
rect 18317 10557 18351 10591
rect 20085 10557 20119 10591
rect 20821 10557 20855 10591
rect 21925 10557 21959 10591
rect 23673 10557 23707 10591
rect 23929 10557 23963 10591
rect 2881 10489 2915 10523
rect 7297 10489 7331 10523
rect 11161 10489 11195 10523
rect 13645 10489 13679 10523
rect 16037 10489 16071 10523
rect 16865 10489 16899 10523
rect 22385 10489 22419 10523
rect 22569 10489 22603 10523
rect 1777 10421 1811 10455
rect 3433 10421 3467 10455
rect 4445 10421 4479 10455
rect 9689 10421 9723 10455
rect 10241 10421 10275 10455
rect 10701 10421 10735 10455
rect 11345 10421 11379 10455
rect 12265 10421 12299 10455
rect 14933 10421 14967 10455
rect 15577 10421 15611 10455
rect 17325 10421 17359 10455
rect 17785 10421 17819 10455
rect 19441 10421 19475 10455
rect 21005 10421 21039 10455
rect 21465 10421 21499 10455
rect 23029 10421 23063 10455
rect 23489 10421 23523 10455
rect 25053 10421 25087 10455
rect 25605 10421 25639 10455
rect 1685 10217 1719 10251
rect 2329 10217 2363 10251
rect 2789 10217 2823 10251
rect 3249 10217 3283 10251
rect 4261 10217 4295 10251
rect 4997 10217 5031 10251
rect 5457 10217 5491 10251
rect 8033 10217 8067 10251
rect 8309 10217 8343 10251
rect 14013 10217 14047 10251
rect 15025 10217 15059 10251
rect 17325 10217 17359 10251
rect 17693 10217 17727 10251
rect 18429 10217 18463 10251
rect 20729 10217 20763 10251
rect 22845 10217 22879 10251
rect 23765 10217 23799 10251
rect 4813 10149 4847 10183
rect 5089 10149 5123 10183
rect 6254 10149 6288 10183
rect 10241 10149 10275 10183
rect 11529 10149 11563 10183
rect 13185 10149 13219 10183
rect 15660 10149 15694 10183
rect 18521 10149 18555 10183
rect 2145 10081 2179 10115
rect 6009 10081 6043 10115
rect 8493 10081 8527 10115
rect 10333 10081 10367 10115
rect 11253 10081 11287 10115
rect 13001 10081 13035 10115
rect 13645 10081 13679 10115
rect 14197 10081 14231 10115
rect 15393 10081 15427 10115
rect 18245 10081 18279 10115
rect 19533 10081 19567 10115
rect 21373 10081 21407 10115
rect 21732 10081 21766 10115
rect 23949 10081 23983 10115
rect 24216 10081 24250 10115
rect 2421 10013 2455 10047
rect 3525 10013 3559 10047
rect 10149 10013 10183 10047
rect 13277 10013 13311 10047
rect 21465 10013 21499 10047
rect 4537 9945 4571 9979
rect 8677 9945 8711 9979
rect 9137 9945 9171 9979
rect 9781 9945 9815 9979
rect 12725 9945 12759 9979
rect 14657 9945 14691 9979
rect 18889 9945 18923 9979
rect 1869 9877 1903 9911
rect 5825 9877 5859 9911
rect 7389 9877 7423 9911
rect 9413 9877 9447 9911
rect 10885 9877 10919 9911
rect 11989 9877 12023 9911
rect 12449 9877 12483 9911
rect 16773 9877 16807 9911
rect 17969 9877 18003 9911
rect 19349 9877 19383 9911
rect 19717 9877 19751 9911
rect 25329 9877 25363 9911
rect 6101 9673 6135 9707
rect 6469 9673 6503 9707
rect 8677 9673 8711 9707
rect 10333 9673 10367 9707
rect 18613 9673 18647 9707
rect 23857 9673 23891 9707
rect 4077 9605 4111 9639
rect 7113 9605 7147 9639
rect 10885 9605 10919 9639
rect 12265 9605 12299 9639
rect 13185 9605 13219 9639
rect 14105 9605 14139 9639
rect 17877 9605 17911 9639
rect 20269 9605 20303 9639
rect 23489 9605 23523 9639
rect 24133 9605 24167 9639
rect 1685 9537 1719 9571
rect 3709 9537 3743 9571
rect 4169 9537 4203 9571
rect 7297 9537 7331 9571
rect 11437 9537 11471 9571
rect 11897 9537 11931 9571
rect 13553 9537 13587 9571
rect 18245 9537 18279 9571
rect 21281 9537 21315 9571
rect 22017 9537 22051 9571
rect 22753 9537 22787 9571
rect 24593 9537 24627 9571
rect 25605 9537 25639 9571
rect 1952 9469 1986 9503
rect 13001 9469 13035 9503
rect 13737 9469 13771 9503
rect 15209 9469 15243 9503
rect 15485 9469 15519 9503
rect 15752 9469 15786 9503
rect 18889 9469 18923 9503
rect 19156 9469 19190 9503
rect 21741 9469 21775 9503
rect 22385 9469 22419 9503
rect 25421 9469 25455 9503
rect 4436 9401 4470 9435
rect 7542 9401 7576 9435
rect 9689 9401 9723 9435
rect 10701 9401 10735 9435
rect 11161 9401 11195 9435
rect 13645 9401 13679 9435
rect 14657 9401 14691 9435
rect 17417 9401 17451 9435
rect 21925 9401 21959 9435
rect 24593 9401 24627 9435
rect 24685 9401 24719 9435
rect 3065 9333 3099 9367
rect 5549 9333 5583 9367
rect 9229 9333 9263 9367
rect 9781 9333 9815 9367
rect 11345 9333 11379 9367
rect 14933 9333 14967 9367
rect 15209 9333 15243 9367
rect 15301 9333 15335 9367
rect 16865 9333 16899 9367
rect 20913 9333 20947 9367
rect 21455 9333 21489 9367
rect 25053 9333 25087 9367
rect 1593 9129 1627 9163
rect 3065 9129 3099 9163
rect 3433 9129 3467 9163
rect 3893 9129 3927 9163
rect 5089 9129 5123 9163
rect 5549 9129 5583 9163
rect 6377 9129 6411 9163
rect 6929 9129 6963 9163
rect 14105 9129 14139 9163
rect 14749 9129 14783 9163
rect 15853 9129 15887 9163
rect 19073 9129 19107 9163
rect 20085 9129 20119 9163
rect 23673 9129 23707 9163
rect 24133 9129 24167 9163
rect 24869 9129 24903 9163
rect 2283 9061 2317 9095
rect 2421 9061 2455 9095
rect 4629 9061 4663 9095
rect 6193 9061 6227 9095
rect 8401 9061 8435 9095
rect 8585 9061 8619 9095
rect 9045 9061 9079 9095
rect 12970 9061 13004 9095
rect 15117 9061 15151 9095
rect 15669 9061 15703 9095
rect 15945 9061 15979 9095
rect 17960 9061 17994 9095
rect 21180 9061 21214 9095
rect 4721 8993 4755 9027
rect 10508 8993 10542 9027
rect 12725 8993 12759 9027
rect 16313 8993 16347 9027
rect 24685 8993 24719 9027
rect 2329 8925 2363 8959
rect 4629 8925 4663 8959
rect 6469 8925 6503 8959
rect 7297 8925 7331 8959
rect 7941 8925 7975 8959
rect 8677 8925 8711 8959
rect 10241 8925 10275 8959
rect 17693 8925 17727 8959
rect 20913 8925 20947 8959
rect 24961 8925 24995 8959
rect 5917 8857 5951 8891
rect 8125 8857 8159 8891
rect 16681 8857 16715 8891
rect 24409 8857 24443 8891
rect 1869 8789 1903 8823
rect 4169 8789 4203 8823
rect 9413 8789 9447 8823
rect 9873 8789 9907 8823
rect 11621 8789 11655 8823
rect 12449 8789 12483 8823
rect 15393 8789 15427 8823
rect 17049 8789 17083 8823
rect 17601 8789 17635 8823
rect 19717 8789 19751 8823
rect 20361 8789 20395 8823
rect 22293 8789 22327 8823
rect 2421 8585 2455 8619
rect 2881 8585 2915 8619
rect 4997 8585 5031 8619
rect 6285 8585 6319 8619
rect 8217 8585 8251 8619
rect 9505 8585 9539 8619
rect 10885 8585 10919 8619
rect 11805 8585 11839 8619
rect 12265 8585 12299 8619
rect 15761 8585 15795 8619
rect 16129 8585 16163 8619
rect 19901 8585 19935 8619
rect 23489 8585 23523 8619
rect 24501 8585 24535 8619
rect 24869 8585 24903 8619
rect 25145 8585 25179 8619
rect 1501 8517 1535 8551
rect 6561 8517 6595 8551
rect 9873 8517 9907 8551
rect 12633 8517 12667 8551
rect 16405 8517 16439 8551
rect 18153 8517 18187 8551
rect 20085 8517 20119 8551
rect 21649 8517 21683 8551
rect 1961 8449 1995 8483
rect 2973 8449 3007 8483
rect 8769 8449 8803 8483
rect 10333 8449 10367 8483
rect 11345 8449 11379 8483
rect 11437 8449 11471 8483
rect 16957 8449 16991 8483
rect 17417 8449 17451 8483
rect 18705 8449 18739 8483
rect 19533 8449 19567 8483
rect 20637 8449 20671 8483
rect 21465 8449 21499 8483
rect 23949 8449 23983 8483
rect 5273 8381 5307 8415
rect 5457 8381 5491 8415
rect 6837 8381 6871 8415
rect 7665 8381 7699 8415
rect 8493 8381 8527 8415
rect 9689 8381 9723 8415
rect 10701 8381 10735 8415
rect 12449 8381 12483 8415
rect 13829 8381 13863 8415
rect 14096 8381 14130 8415
rect 19073 8381 19107 8415
rect 20361 8381 20395 8415
rect 21925 8381 21959 8415
rect 22569 8381 22603 8415
rect 23673 8381 23707 8415
rect 24961 8381 24995 8415
rect 25513 8381 25547 8415
rect 1961 8313 1995 8347
rect 2053 8313 2087 8347
rect 3218 8313 3252 8347
rect 5733 8313 5767 8347
rect 7113 8313 7147 8347
rect 8033 8313 8067 8347
rect 8677 8313 8711 8347
rect 9137 8313 9171 8347
rect 11345 8313 11379 8347
rect 16681 8313 16715 8347
rect 16865 8313 16899 8347
rect 18429 8313 18463 8347
rect 18613 8313 18647 8347
rect 20545 8313 20579 8347
rect 22201 8313 22235 8347
rect 4353 8245 4387 8279
rect 13093 8245 13127 8279
rect 13645 8245 13679 8279
rect 15209 8245 15243 8279
rect 17693 8245 17727 8279
rect 21005 8245 21039 8279
rect 22109 8245 22143 8279
rect 1409 8041 1443 8075
rect 2145 8041 2179 8075
rect 2973 8041 3007 8075
rect 4629 8041 4663 8075
rect 7113 8041 7147 8075
rect 7665 8041 7699 8075
rect 8125 8041 8159 8075
rect 8953 8041 8987 8075
rect 11345 8041 11379 8075
rect 12725 8041 12759 8075
rect 13645 8041 13679 8075
rect 14105 8041 14139 8075
rect 15025 8041 15059 8075
rect 15853 8041 15887 8075
rect 17417 8041 17451 8075
rect 18521 8041 18555 8075
rect 21557 8041 21591 8075
rect 23673 8041 23707 8075
rect 4721 7973 4755 8007
rect 6000 7973 6034 8007
rect 9321 7973 9355 8007
rect 13461 7973 13495 8007
rect 15945 7973 15979 8007
rect 18061 7973 18095 8007
rect 18153 7973 18187 8007
rect 19441 7973 19475 8007
rect 19625 7973 19659 8007
rect 21189 7973 21223 8007
rect 22008 7973 22042 8007
rect 24593 7973 24627 8007
rect 5733 7905 5767 7939
rect 8217 7905 8251 7939
rect 8493 7905 8527 7939
rect 10232 7905 10266 7939
rect 13737 7905 13771 7939
rect 14473 7905 14507 7939
rect 15669 7905 15703 7939
rect 24317 7905 24351 7939
rect 2973 7837 3007 7871
rect 3065 7837 3099 7871
rect 4629 7837 4663 7871
rect 9965 7837 9999 7871
rect 16313 7837 16347 7871
rect 17969 7837 18003 7871
rect 19717 7837 19751 7871
rect 21741 7837 21775 7871
rect 4169 7769 4203 7803
rect 13185 7769 13219 7803
rect 15393 7769 15427 7803
rect 17601 7769 17635 7803
rect 18981 7769 19015 7803
rect 2513 7701 2547 7735
rect 3709 7701 3743 7735
rect 5181 7701 5215 7735
rect 5457 7701 5491 7735
rect 11897 7701 11931 7735
rect 12265 7701 12299 7735
rect 16681 7701 16715 7735
rect 19165 7701 19199 7735
rect 20085 7701 20119 7735
rect 20453 7701 20487 7735
rect 23121 7701 23155 7735
rect 2145 7497 2179 7531
rect 3709 7497 3743 7531
rect 4629 7497 4663 7531
rect 5273 7497 5307 7531
rect 6285 7497 6319 7531
rect 7665 7497 7699 7531
rect 10425 7497 10459 7531
rect 13001 7497 13035 7531
rect 15577 7497 15611 7531
rect 16129 7497 16163 7531
rect 17509 7497 17543 7531
rect 18705 7497 18739 7531
rect 21465 7497 21499 7531
rect 21925 7497 21959 7531
rect 24685 7497 24719 7531
rect 25421 7497 25455 7531
rect 3433 7429 3467 7463
rect 4997 7429 5031 7463
rect 12633 7429 12667 7463
rect 22109 7429 22143 7463
rect 23765 7429 23799 7463
rect 2513 7361 2547 7395
rect 2697 7361 2731 7395
rect 4261 7361 4295 7395
rect 5733 7361 5767 7395
rect 7849 7361 7883 7395
rect 10885 7361 10919 7395
rect 12081 7361 12115 7395
rect 24317 7361 24351 7395
rect 1961 7293 1995 7327
rect 5825 7293 5859 7327
rect 10977 7293 11011 7327
rect 12449 7293 12483 7327
rect 13553 7293 13587 7327
rect 13820 7293 13854 7327
rect 16405 7293 16439 7327
rect 17049 7293 17083 7327
rect 18061 7293 18095 7327
rect 19257 7293 19291 7327
rect 22385 7293 22419 7327
rect 24041 7293 24075 7327
rect 25237 7293 25271 7327
rect 2605 7225 2639 7259
rect 3985 7225 4019 7259
rect 5733 7225 5767 7259
rect 7389 7225 7423 7259
rect 8094 7225 8128 7259
rect 11713 7225 11747 7259
rect 16681 7225 16715 7259
rect 19165 7225 19199 7259
rect 19524 7225 19558 7259
rect 22569 7225 22603 7259
rect 22661 7225 22695 7259
rect 23489 7225 23523 7259
rect 25789 7225 25823 7259
rect 3065 7157 3099 7191
rect 4169 7157 4203 7191
rect 6561 7157 6595 7191
rect 6837 7157 6871 7191
rect 9229 7157 9263 7191
rect 10057 7157 10091 7191
rect 10885 7157 10919 7191
rect 11345 7157 11379 7191
rect 13461 7157 13495 7191
rect 14933 7157 14967 7191
rect 15945 7157 15979 7191
rect 16589 7157 16623 7191
rect 18245 7157 18279 7191
rect 20637 7157 20671 7191
rect 23029 7157 23063 7191
rect 24225 7157 24259 7191
rect 6285 6953 6319 6987
rect 6653 6953 6687 6987
rect 7941 6953 7975 6987
rect 10425 6953 10459 6987
rect 13185 6953 13219 6987
rect 13553 6953 13587 6987
rect 15577 6953 15611 6987
rect 18245 6953 18279 6987
rect 22109 6953 22143 6987
rect 4528 6885 4562 6919
rect 14197 6885 14231 6919
rect 19809 6885 19843 6919
rect 1768 6817 1802 6851
rect 3709 6817 3743 6851
rect 4261 6817 4295 6851
rect 6929 6817 6963 6851
rect 9689 6817 9723 6851
rect 11233 6817 11267 6851
rect 14289 6817 14323 6851
rect 14657 6817 14691 6851
rect 15025 6817 15059 6851
rect 16120 6817 16154 6851
rect 17877 6817 17911 6851
rect 18797 6817 18831 6851
rect 19165 6817 19199 6851
rect 20729 6817 20763 6851
rect 20913 6817 20947 6851
rect 22385 6817 22419 6851
rect 22917 6817 22951 6851
rect 25145 6817 25179 6851
rect 1501 6749 1535 6783
rect 7849 6749 7883 6783
rect 8033 6749 8067 6783
rect 10977 6749 11011 6783
rect 14105 6749 14139 6783
rect 15853 6749 15887 6783
rect 19717 6749 19751 6783
rect 19901 6749 19935 6783
rect 21741 6749 21775 6783
rect 22668 6749 22702 6783
rect 5641 6681 5675 6715
rect 7481 6681 7515 6715
rect 13737 6681 13771 6715
rect 25329 6681 25363 6715
rect 2881 6613 2915 6647
rect 8401 6613 8435 6647
rect 8769 6613 8803 6647
rect 9413 6613 9447 6647
rect 9873 6613 9907 6647
rect 10701 6613 10735 6647
rect 12357 6613 12391 6647
rect 17233 6613 17267 6647
rect 19349 6613 19383 6647
rect 20269 6613 20303 6647
rect 21097 6613 21131 6647
rect 24041 6613 24075 6647
rect 1685 6409 1719 6443
rect 2053 6409 2087 6443
rect 3525 6409 3559 6443
rect 4261 6409 4295 6443
rect 5273 6409 5307 6443
rect 6285 6409 6319 6443
rect 6561 6409 6595 6443
rect 7205 6409 7239 6443
rect 9045 6409 9079 6443
rect 10793 6409 10827 6443
rect 13645 6409 13679 6443
rect 18889 6409 18923 6443
rect 19349 6409 19383 6443
rect 20821 6409 20855 6443
rect 23029 6409 23063 6443
rect 23397 6409 23431 6443
rect 7573 6341 7607 6375
rect 12541 6341 12575 6375
rect 22109 6341 22143 6375
rect 2145 6273 2179 6307
rect 5825 6273 5859 6307
rect 7665 6273 7699 6307
rect 16865 6273 16899 6307
rect 18337 6273 18371 6307
rect 22569 6273 22603 6307
rect 23673 6273 23707 6307
rect 2412 6205 2446 6239
rect 4721 6205 4755 6239
rect 7932 6205 7966 6239
rect 11345 6205 11379 6239
rect 11897 6205 11931 6239
rect 14105 6205 14139 6239
rect 16589 6205 16623 6239
rect 17693 6205 17727 6239
rect 18061 6205 18095 6239
rect 19441 6205 19475 6239
rect 19708 6205 19742 6239
rect 21925 6205 21959 6239
rect 25605 6205 25639 6239
rect 4997 6137 5031 6171
rect 5549 6137 5583 6171
rect 5733 6137 5767 6171
rect 11069 6137 11103 6171
rect 11253 6137 11287 6171
rect 12817 6137 12851 6171
rect 13093 6137 13127 6171
rect 14350 6137 14384 6171
rect 16405 6137 16439 6171
rect 22569 6137 22603 6171
rect 22661 6137 22695 6171
rect 23940 6137 23974 6171
rect 9781 6069 9815 6103
rect 10149 6069 10183 6103
rect 10609 6069 10643 6103
rect 12265 6069 12299 6103
rect 13001 6069 13035 6103
rect 15485 6069 15519 6103
rect 16037 6069 16071 6103
rect 17325 6069 17359 6103
rect 21373 6069 21407 6103
rect 25053 6069 25087 6103
rect 1409 5865 1443 5899
rect 2237 5865 2271 5899
rect 4353 5865 4387 5899
rect 4997 5865 5031 5899
rect 5549 5865 5583 5899
rect 6561 5865 6595 5899
rect 7389 5865 7423 5899
rect 8953 5865 8987 5899
rect 9689 5865 9723 5899
rect 10609 5865 10643 5899
rect 12081 5865 12115 5899
rect 12725 5865 12759 5899
rect 15025 5865 15059 5899
rect 15485 5865 15519 5899
rect 18613 5865 18647 5899
rect 19625 5865 19659 5899
rect 20085 5865 20119 5899
rect 22017 5865 22051 5899
rect 23029 5865 23063 5899
rect 23765 5865 23799 5899
rect 25513 5865 25547 5899
rect 2973 5797 3007 5831
rect 5089 5797 5123 5831
rect 7941 5797 7975 5831
rect 8125 5797 8159 5831
rect 8217 5797 8251 5831
rect 13185 5797 13219 5831
rect 14013 5797 14047 5831
rect 14197 5797 14231 5831
rect 14289 5797 14323 5831
rect 15945 5797 15979 5831
rect 16764 5797 16798 5831
rect 21189 5797 21223 5831
rect 22293 5797 22327 5831
rect 22845 5797 22879 5831
rect 2789 5729 2823 5763
rect 7113 5729 7147 5763
rect 10701 5729 10735 5763
rect 10968 5729 11002 5763
rect 15301 5729 15335 5763
rect 19441 5729 19475 5763
rect 20913 5729 20947 5763
rect 24041 5729 24075 5763
rect 25329 5729 25363 5763
rect 3065 5661 3099 5695
rect 4997 5661 5031 5695
rect 6469 5661 6503 5695
rect 6653 5661 6687 5695
rect 16497 5661 16531 5695
rect 19717 5661 19751 5695
rect 23121 5661 23155 5695
rect 24317 5661 24351 5695
rect 4537 5593 4571 5627
rect 6101 5593 6135 5627
rect 7665 5593 7699 5627
rect 8585 5593 8619 5627
rect 9505 5593 9539 5627
rect 13737 5593 13771 5627
rect 14749 5593 14783 5627
rect 20729 5593 20763 5627
rect 2513 5525 2547 5559
rect 3709 5525 3743 5559
rect 5917 5525 5951 5559
rect 10241 5525 10275 5559
rect 13553 5525 13587 5559
rect 16221 5525 16255 5559
rect 17877 5525 17911 5559
rect 18981 5525 19015 5559
rect 19165 5525 19199 5559
rect 22569 5525 22603 5559
rect 1961 5321 1995 5355
rect 3157 5321 3191 5355
rect 4721 5321 4755 5355
rect 6561 5321 6595 5355
rect 7297 5321 7331 5355
rect 8861 5321 8895 5355
rect 9781 5321 9815 5355
rect 10333 5321 10367 5355
rect 11253 5321 11287 5355
rect 12725 5321 12759 5355
rect 15393 5321 15427 5355
rect 15853 5321 15887 5355
rect 16773 5321 16807 5355
rect 17233 5321 17267 5355
rect 19073 5321 19107 5355
rect 20637 5321 20671 5355
rect 23489 5321 23523 5355
rect 24225 5321 24259 5355
rect 24777 5321 24811 5355
rect 25421 5321 25455 5355
rect 2145 5253 2179 5287
rect 3709 5253 3743 5287
rect 5273 5253 5307 5287
rect 6285 5253 6319 5287
rect 14289 5253 14323 5287
rect 22109 5253 22143 5287
rect 23949 5253 23983 5287
rect 2697 5185 2731 5219
rect 10793 5185 10827 5219
rect 10885 5185 10919 5219
rect 11897 5185 11931 5219
rect 13277 5185 13311 5219
rect 13645 5185 13679 5219
rect 16221 5185 16255 5219
rect 16405 5185 16439 5219
rect 19257 5185 19291 5219
rect 21557 5185 21591 5219
rect 22661 5185 22695 5219
rect 23029 5185 23063 5219
rect 2421 5117 2455 5151
rect 5549 5117 5583 5151
rect 7481 5117 7515 5151
rect 12173 5117 12207 5151
rect 13001 5117 13035 5151
rect 14105 5117 14139 5151
rect 14565 5117 14599 5151
rect 17509 5117 17543 5151
rect 18061 5117 18095 5151
rect 18613 5117 18647 5151
rect 21925 5117 21959 5151
rect 22385 5117 22419 5151
rect 24593 5117 24627 5151
rect 2605 5049 2639 5083
rect 3525 5049 3559 5083
rect 3985 5049 4019 5083
rect 4261 5049 4295 5083
rect 5825 5049 5859 5083
rect 7748 5049 7782 5083
rect 10793 5049 10827 5083
rect 13185 5049 13219 5083
rect 14749 5049 14783 5083
rect 14841 5049 14875 5083
rect 16313 5049 16347 5083
rect 19524 5049 19558 5083
rect 22569 5049 22603 5083
rect 4169 4981 4203 5015
rect 5089 4981 5123 5015
rect 5733 4981 5767 5015
rect 10149 4981 10183 5015
rect 18245 4981 18279 5015
rect 1869 4777 1903 4811
rect 2329 4777 2363 4811
rect 2973 4777 3007 4811
rect 4629 4777 4663 4811
rect 5549 4777 5583 4811
rect 6193 4777 6227 4811
rect 7757 4777 7791 4811
rect 8217 4777 8251 4811
rect 9413 4777 9447 4811
rect 12081 4777 12115 4811
rect 12725 4777 12759 4811
rect 12817 4777 12851 4811
rect 13461 4777 13495 4811
rect 17785 4777 17819 4811
rect 18429 4777 18463 4811
rect 22109 4777 22143 4811
rect 25237 4777 25271 4811
rect 25605 4777 25639 4811
rect 2789 4709 2823 4743
rect 3065 4709 3099 4743
rect 4445 4709 4479 4743
rect 5181 4709 5215 4743
rect 7849 4709 7883 4743
rect 8585 4709 8619 4743
rect 3709 4641 3743 4675
rect 6285 4641 6319 4675
rect 7113 4641 7147 4675
rect 10037 4641 10071 4675
rect 1409 4573 1443 4607
rect 4721 4573 4755 4607
rect 6193 4573 6227 4607
rect 7757 4573 7791 4607
rect 9781 4573 9815 4607
rect 2513 4505 2547 4539
rect 4169 4505 4203 4539
rect 5733 4505 5767 4539
rect 13277 4709 13311 4743
rect 14197 4709 14231 4743
rect 18797 4709 18831 4743
rect 19625 4709 19659 4743
rect 19809 4709 19843 4743
rect 21465 4709 21499 4743
rect 22836 4709 22870 4743
rect 14657 4641 14691 4675
rect 16120 4641 16154 4675
rect 19165 4641 19199 4675
rect 19901 4641 19935 4675
rect 21557 4641 21591 4675
rect 22569 4641 22603 4675
rect 25053 4641 25087 4675
rect 13553 4573 13587 4607
rect 15853 4573 15887 4607
rect 21373 4573 21407 4607
rect 24593 4573 24627 4607
rect 19349 4505 19383 4539
rect 20361 4505 20395 4539
rect 21005 4505 21039 4539
rect 6745 4437 6779 4471
rect 7297 4437 7331 4471
rect 9137 4437 9171 4471
rect 11161 4437 11195 4471
rect 11713 4437 11747 4471
rect 12817 4437 12851 4471
rect 13001 4437 13035 4471
rect 14933 4437 14967 4471
rect 15577 4437 15611 4471
rect 17233 4437 17267 4471
rect 20729 4437 20763 4471
rect 22385 4437 22419 4471
rect 23949 4437 23983 4471
rect 2881 4233 2915 4267
rect 4997 4233 5031 4267
rect 6193 4233 6227 4267
rect 6653 4233 6687 4267
rect 7573 4233 7607 4267
rect 8493 4233 8527 4267
rect 9137 4233 9171 4267
rect 10701 4233 10735 4267
rect 13645 4233 13679 4267
rect 19349 4233 19383 4267
rect 20913 4233 20947 4267
rect 22937 4233 22971 4267
rect 23305 4233 23339 4267
rect 25513 4233 25547 4267
rect 19533 4165 19567 4199
rect 1869 4097 1903 4131
rect 2513 4097 2547 4131
rect 5365 4097 5399 4131
rect 7389 4097 7423 4131
rect 7941 4097 7975 4131
rect 8125 4097 8159 4131
rect 10425 4097 10459 4131
rect 12173 4097 12207 4131
rect 14105 4097 14139 4131
rect 14841 4097 14875 4131
rect 16681 4097 16715 4131
rect 18889 4097 18923 4131
rect 20085 4097 20119 4131
rect 21465 4097 21499 4131
rect 22477 4097 22511 4131
rect 23857 4097 23891 4131
rect 24869 4097 24903 4131
rect 2053 4029 2087 4063
rect 2973 4029 3007 4063
rect 3240 4029 3274 4063
rect 5457 4029 5491 4063
rect 9689 4029 9723 4063
rect 10977 4029 11011 4063
rect 11253 4029 11287 4063
rect 11621 4029 11655 4063
rect 15577 4029 15611 4063
rect 16773 4029 16807 4063
rect 17877 4029 17911 4063
rect 18061 4029 18095 4063
rect 18337 4029 18371 4063
rect 23673 4029 23707 4063
rect 24409 4029 24443 4063
rect 24961 4029 24995 4063
rect 5733 3961 5767 3995
rect 8033 3961 8067 3995
rect 9413 3961 9447 3995
rect 9597 3961 9631 3995
rect 10149 3961 10183 3995
rect 11161 3961 11195 3995
rect 13001 3961 13035 3995
rect 13277 3961 13311 3995
rect 14565 3961 14599 3995
rect 16681 3961 16715 3995
rect 19809 3961 19843 3995
rect 21999 3961 22033 3995
rect 22569 3961 22603 3995
rect 25881 3961 25915 3995
rect 1491 3893 1525 3927
rect 1961 3893 1995 3927
rect 4353 3893 4387 3927
rect 8953 3893 8987 3927
rect 12715 3893 12749 3927
rect 13185 3893 13219 3927
rect 14279 3893 14313 3927
rect 14749 3893 14783 3927
rect 15853 3893 15887 3927
rect 16211 3893 16245 3927
rect 17141 3893 17175 3927
rect 19993 3893 20027 3927
rect 20453 3893 20487 3927
rect 21833 3893 21867 3927
rect 22477 3893 22511 3927
rect 25145 3893 25179 3927
rect 26249 3893 26283 3927
rect 1409 3689 1443 3723
rect 2329 3689 2363 3723
rect 2973 3689 3007 3723
rect 3433 3689 3467 3723
rect 3801 3689 3835 3723
rect 4905 3689 4939 3723
rect 5457 3689 5491 3723
rect 7481 3689 7515 3723
rect 8585 3689 8619 3723
rect 9505 3689 9539 3723
rect 11529 3689 11563 3723
rect 14105 3689 14139 3723
rect 15025 3689 15059 3723
rect 15853 3689 15887 3723
rect 18889 3689 18923 3723
rect 20269 3689 20303 3723
rect 20729 3689 20763 3723
rect 22293 3689 22327 3723
rect 23949 3689 23983 3723
rect 25237 3689 25271 3723
rect 25605 3689 25639 3723
rect 2789 3621 2823 3655
rect 5816 3621 5850 3655
rect 12265 3621 12299 3655
rect 12992 3621 13026 3655
rect 15669 3621 15703 3655
rect 17202 3621 17236 3655
rect 19717 3621 19751 3655
rect 21189 3621 21223 3655
rect 22836 3621 22870 3655
rect 4077 3553 4111 3587
rect 4353 3553 4387 3587
rect 7941 3553 7975 3587
rect 8677 3553 8711 3587
rect 10416 3553 10450 3587
rect 12633 3553 12667 3587
rect 16957 3553 16991 3587
rect 19441 3553 19475 3587
rect 20913 3553 20947 3587
rect 22017 3553 22051 3587
rect 22569 3553 22603 3587
rect 25053 3553 25087 3587
rect 3065 3485 3099 3519
rect 5549 3485 5583 3519
rect 8585 3485 8619 3519
rect 9965 3485 9999 3519
rect 10149 3485 10183 3519
rect 12725 3485 12759 3519
rect 15945 3485 15979 3519
rect 19349 3485 19383 3519
rect 2513 3417 2547 3451
rect 6929 3417 6963 3451
rect 9137 3417 9171 3451
rect 15393 3417 15427 3451
rect 24869 3417 24903 3451
rect 1961 3349 1995 3383
rect 8125 3349 8159 3383
rect 14749 3349 14783 3383
rect 16313 3349 16347 3383
rect 16773 3349 16807 3383
rect 18337 3349 18371 3383
rect 24501 3349 24535 3383
rect 25973 3349 26007 3383
rect 5273 3145 5307 3179
rect 6285 3145 6319 3179
rect 6561 3145 6595 3179
rect 9137 3145 9171 3179
rect 14289 3145 14323 3179
rect 15393 3145 15427 3179
rect 16865 3145 16899 3179
rect 17417 3145 17451 3179
rect 17785 3145 17819 3179
rect 18153 3145 18187 3179
rect 19349 3145 19383 3179
rect 20729 3145 20763 3179
rect 21005 3145 21039 3179
rect 22385 3145 22419 3179
rect 23397 3145 23431 3179
rect 24961 3145 24995 3179
rect 25789 3145 25823 3179
rect 19073 3077 19107 3111
rect 5733 3009 5767 3043
rect 9321 3009 9355 3043
rect 18521 3009 18555 3043
rect 1409 2941 1443 2975
rect 2605 2941 2639 2975
rect 2697 2941 2731 2975
rect 5089 2941 5123 2975
rect 5825 2941 5859 2975
rect 6837 2941 6871 2975
rect 7104 2941 7138 2975
rect 11253 2941 11287 2975
rect 12173 2941 12207 2975
rect 12725 2941 12759 2975
rect 12909 2941 12943 2975
rect 13176 2941 13210 2975
rect 15209 2941 15243 2975
rect 15485 2941 15519 2975
rect 1685 2873 1719 2907
rect 2964 2873 2998 2907
rect 5733 2873 5767 2907
rect 9566 2873 9600 2907
rect 15730 2873 15764 2907
rect 18705 2873 18739 2907
rect 19717 3077 19751 3111
rect 23029 3077 23063 3111
rect 24501 3077 24535 3111
rect 19533 3009 19567 3043
rect 20177 3009 20211 3043
rect 21465 3009 21499 3043
rect 23949 3009 23983 3043
rect 25329 3009 25363 3043
rect 20269 2941 20303 2975
rect 21189 2941 21223 2975
rect 21925 2941 21959 2975
rect 22477 2941 22511 2975
rect 23765 2941 23799 2975
rect 25053 2941 25087 2975
rect 26249 2941 26283 2975
rect 2237 2805 2271 2839
rect 4077 2805 4111 2839
rect 4629 2805 4663 2839
rect 8217 2805 8251 2839
rect 8769 2805 8803 2839
rect 10701 2805 10735 2839
rect 11621 2805 11655 2839
rect 14933 2805 14967 2839
rect 15209 2805 15243 2839
rect 18613 2805 18647 2839
rect 19349 2805 19383 2839
rect 20177 2805 20211 2839
rect 22661 2805 22695 2839
rect 1869 2601 1903 2635
rect 3893 2601 3927 2635
rect 5457 2601 5491 2635
rect 6009 2601 6043 2635
rect 7481 2601 7515 2635
rect 7941 2601 7975 2635
rect 8309 2601 8343 2635
rect 9137 2601 9171 2635
rect 9505 2601 9539 2635
rect 11161 2601 11195 2635
rect 15209 2601 15243 2635
rect 17601 2601 17635 2635
rect 20085 2601 20119 2635
rect 22201 2601 22235 2635
rect 1409 2533 1443 2567
rect 2329 2533 2363 2567
rect 2973 2533 3007 2567
rect 3065 2533 3099 2567
rect 3433 2533 3467 2567
rect 4322 2533 4356 2567
rect 7573 2533 7607 2567
rect 14381 2533 14415 2567
rect 15853 2533 15887 2567
rect 16037 2533 16071 2567
rect 16129 2533 16163 2567
rect 16957 2533 16991 2567
rect 18061 2533 18095 2567
rect 18889 2533 18923 2567
rect 21263 2533 21297 2567
rect 21741 2533 21775 2567
rect 21833 2533 21867 2567
rect 24317 2533 24351 2567
rect 4077 2465 4111 2499
rect 6653 2465 6687 2499
rect 7297 2465 7331 2499
rect 8493 2465 8527 2499
rect 9781 2465 9815 2499
rect 10037 2465 10071 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 14197 2465 14231 2499
rect 14841 2465 14875 2499
rect 16497 2465 16531 2499
rect 17049 2465 17083 2499
rect 18981 2465 19015 2499
rect 19901 2465 19935 2499
rect 20637 2465 20671 2499
rect 22569 2465 22603 2499
rect 22753 2465 22787 2499
rect 23305 2465 23339 2499
rect 24041 2465 24075 2499
rect 24777 2465 24811 2499
rect 25145 2465 25179 2499
rect 25329 2465 25363 2499
rect 25881 2465 25915 2499
rect 2881 2397 2915 2431
rect 12449 2397 12483 2431
rect 14473 2397 14507 2431
rect 18797 2397 18831 2431
rect 19717 2397 19751 2431
rect 21649 2397 21683 2431
rect 23673 2397 23707 2431
rect 7021 2329 7055 2363
rect 12817 2329 12851 2363
rect 13921 2329 13955 2363
rect 15577 2329 15611 2363
rect 18429 2329 18463 2363
rect 2513 2261 2547 2295
rect 8677 2261 8711 2295
rect 11713 2261 11747 2295
rect 13645 2261 13679 2295
rect 17233 2261 17267 2295
rect 20913 2261 20947 2295
rect 22937 2261 22971 2295
rect 25513 2261 25547 2295
<< metal1 >>
rect 22002 26596 22008 26648
rect 22060 26636 22066 26648
rect 23566 26636 23572 26648
rect 22060 26608 23572 26636
rect 22060 26596 22066 26608
rect 23566 26596 23572 26608
rect 23624 26596 23630 26648
rect 14642 26392 14648 26444
rect 14700 26432 14706 26444
rect 23474 26432 23480 26444
rect 14700 26404 23480 26432
rect 14700 26392 14706 26404
rect 23474 26392 23480 26404
rect 23532 26392 23538 26444
rect 3418 26256 3424 26308
rect 3476 26296 3482 26308
rect 11238 26296 11244 26308
rect 3476 26268 11244 26296
rect 3476 26256 3482 26268
rect 11238 26256 11244 26268
rect 11296 26256 11302 26308
rect 22186 26256 22192 26308
rect 22244 26296 22250 26308
rect 23474 26296 23480 26308
rect 22244 26268 23480 26296
rect 22244 26256 22250 26268
rect 23474 26256 23480 26268
rect 23532 26256 23538 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 3050 24828 3056 24880
rect 3108 24868 3114 24880
rect 15930 24868 15936 24880
rect 3108 24840 15936 24868
rect 3108 24828 3114 24840
rect 15930 24828 15936 24840
rect 15988 24828 15994 24880
rect 21174 24828 21180 24880
rect 21232 24868 21238 24880
rect 23474 24868 23480 24880
rect 21232 24840 23480 24868
rect 21232 24828 21238 24840
rect 23474 24828 23480 24840
rect 23532 24828 23538 24880
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 23842 19796 23848 19848
rect 23900 19836 23906 19848
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 23900 19808 24593 19836
rect 23900 19796 23906 19808
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 23750 19252 23756 19304
rect 23808 19292 23814 19304
rect 24581 19295 24639 19301
rect 24581 19292 24593 19295
rect 23808 19264 24593 19292
rect 23808 19252 23814 19264
rect 24581 19261 24593 19264
rect 24627 19292 24639 19295
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 24627 19264 25145 19292
rect 24627 19261 24639 19264
rect 24581 19255 24639 19261
rect 25133 19261 25145 19264
rect 25179 19261 25191 19295
rect 25133 19255 25191 19261
rect 24765 19159 24823 19165
rect 24765 19125 24777 19159
rect 24811 19156 24823 19159
rect 26878 19156 26884 19168
rect 24811 19128 26884 19156
rect 24811 19125 24823 19128
rect 24765 19119 24823 19125
rect 26878 19116 26884 19128
rect 26936 19116 26942 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 23474 18816 23480 18828
rect 23435 18788 23480 18816
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 24578 18816 24584 18828
rect 24539 18788 24584 18816
rect 24578 18776 24584 18788
rect 24636 18776 24642 18828
rect 22465 18751 22523 18757
rect 22465 18717 22477 18751
rect 22511 18748 22523 18751
rect 22830 18748 22836 18760
rect 22511 18720 22836 18748
rect 22511 18717 22523 18720
rect 22465 18711 22523 18717
rect 22830 18708 22836 18720
rect 22888 18708 22894 18760
rect 23661 18615 23719 18621
rect 23661 18581 23673 18615
rect 23707 18612 23719 18615
rect 24118 18612 24124 18624
rect 23707 18584 24124 18612
rect 23707 18581 23719 18584
rect 23661 18575 23719 18581
rect 24118 18572 24124 18584
rect 24176 18572 24182 18624
rect 24210 18572 24216 18624
rect 24268 18612 24274 18624
rect 24765 18615 24823 18621
rect 24765 18612 24777 18615
rect 24268 18584 24777 18612
rect 24268 18572 24274 18584
rect 24765 18581 24777 18584
rect 24811 18581 24823 18615
rect 24765 18575 24823 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 24670 18368 24676 18420
rect 24728 18408 24734 18420
rect 25133 18411 25191 18417
rect 25133 18408 25145 18411
rect 24728 18380 25145 18408
rect 24728 18368 24734 18380
rect 25133 18377 25145 18380
rect 25179 18377 25191 18411
rect 25133 18371 25191 18377
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 1443 18176 2084 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 2056 18080 2084 18176
rect 24412 18176 24593 18204
rect 750 18028 756 18080
rect 808 18068 814 18080
rect 1581 18071 1639 18077
rect 1581 18068 1593 18071
rect 808 18040 1593 18068
rect 808 18028 814 18040
rect 1581 18037 1593 18040
rect 1627 18037 1639 18071
rect 2038 18068 2044 18080
rect 1999 18040 2044 18068
rect 1581 18031 1639 18037
rect 2038 18028 2044 18040
rect 2096 18028 2102 18080
rect 20162 18068 20168 18080
rect 20123 18040 20168 18068
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 22370 18028 22376 18080
rect 22428 18068 22434 18080
rect 22557 18071 22615 18077
rect 22557 18068 22569 18071
rect 22428 18040 22569 18068
rect 22428 18028 22434 18040
rect 22557 18037 22569 18040
rect 22603 18037 22615 18071
rect 22557 18031 22615 18037
rect 23290 18028 23296 18080
rect 23348 18068 23354 18080
rect 23474 18068 23480 18080
rect 23348 18040 23480 18068
rect 23348 18028 23354 18040
rect 23474 18028 23480 18040
rect 23532 18068 23538 18080
rect 23845 18071 23903 18077
rect 23845 18068 23857 18071
rect 23532 18040 23857 18068
rect 23532 18028 23538 18040
rect 23845 18037 23857 18040
rect 23891 18037 23903 18071
rect 23845 18031 23903 18037
rect 24026 18028 24032 18080
rect 24084 18068 24090 18080
rect 24412 18077 24440 18176
rect 24581 18173 24593 18176
rect 24627 18173 24639 18207
rect 24581 18167 24639 18173
rect 24397 18071 24455 18077
rect 24397 18068 24409 18071
rect 24084 18040 24409 18068
rect 24084 18028 24090 18040
rect 24397 18037 24409 18040
rect 24443 18037 24455 18071
rect 24397 18031 24455 18037
rect 24765 18071 24823 18077
rect 24765 18037 24777 18071
rect 24811 18068 24823 18071
rect 25406 18068 25412 18080
rect 24811 18040 25412 18068
rect 24811 18037 24823 18040
rect 24765 18031 24823 18037
rect 25406 18028 25412 18040
rect 25464 18028 25470 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 22925 17867 22983 17873
rect 22925 17833 22937 17867
rect 22971 17864 22983 17867
rect 23382 17864 23388 17876
rect 22971 17836 23388 17864
rect 22971 17833 22983 17836
rect 22925 17827 22983 17833
rect 23382 17824 23388 17836
rect 23440 17824 23446 17876
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17697 1455 17731
rect 2498 17728 2504 17740
rect 2459 17700 2504 17728
rect 1397 17691 1455 17697
rect 1412 17660 1440 17691
rect 2498 17688 2504 17700
rect 2556 17688 2562 17740
rect 22462 17688 22468 17740
rect 22520 17728 22526 17740
rect 22741 17731 22799 17737
rect 22741 17728 22753 17731
rect 22520 17700 22753 17728
rect 22520 17688 22526 17700
rect 22741 17697 22753 17700
rect 22787 17697 22799 17731
rect 22741 17691 22799 17697
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24670 17728 24676 17740
rect 24627 17700 24676 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 2038 17660 2044 17672
rect 1412 17632 2044 17660
rect 2038 17620 2044 17632
rect 2096 17620 2102 17672
rect 19518 17660 19524 17672
rect 19479 17632 19524 17660
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 21361 17663 21419 17669
rect 21361 17629 21373 17663
rect 21407 17660 21419 17663
rect 21726 17660 21732 17672
rect 21407 17632 21732 17660
rect 21407 17629 21419 17632
rect 21361 17623 21419 17629
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 23014 17660 23020 17672
rect 22975 17632 23020 17660
rect 23014 17620 23020 17632
rect 23072 17620 23078 17672
rect 658 17484 664 17536
rect 716 17524 722 17536
rect 1581 17527 1639 17533
rect 1581 17524 1593 17527
rect 716 17496 1593 17524
rect 716 17484 722 17496
rect 1581 17493 1593 17496
rect 1627 17493 1639 17527
rect 1581 17487 1639 17493
rect 2590 17484 2596 17536
rect 2648 17524 2654 17536
rect 2685 17527 2743 17533
rect 2685 17524 2697 17527
rect 2648 17496 2697 17524
rect 2648 17484 2654 17496
rect 2685 17493 2697 17496
rect 2731 17493 2743 17527
rect 2685 17487 2743 17493
rect 22097 17527 22155 17533
rect 22097 17493 22109 17527
rect 22143 17524 22155 17527
rect 22465 17527 22523 17533
rect 22465 17524 22477 17527
rect 22143 17496 22477 17524
rect 22143 17493 22155 17496
rect 22097 17487 22155 17493
rect 22465 17493 22477 17496
rect 22511 17524 22523 17527
rect 22554 17524 22560 17536
rect 22511 17496 22560 17524
rect 22511 17493 22523 17496
rect 22465 17487 22523 17493
rect 22554 17484 22560 17496
rect 22612 17484 22618 17536
rect 23566 17484 23572 17536
rect 23624 17524 23630 17536
rect 24765 17527 24823 17533
rect 24765 17524 24777 17527
rect 23624 17496 24777 17524
rect 23624 17484 23630 17496
rect 24765 17493 24777 17496
rect 24811 17493 24823 17527
rect 24765 17487 24823 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2409 17323 2467 17329
rect 2409 17289 2421 17323
rect 2455 17320 2467 17323
rect 2498 17320 2504 17332
rect 2455 17292 2504 17320
rect 2455 17289 2467 17292
rect 2409 17283 2467 17289
rect 2498 17280 2504 17292
rect 2556 17280 2562 17332
rect 22462 17280 22468 17332
rect 22520 17320 22526 17332
rect 23017 17323 23075 17329
rect 23017 17320 23029 17323
rect 22520 17292 23029 17320
rect 22520 17280 22526 17292
rect 23017 17289 23029 17292
rect 23063 17289 23075 17323
rect 23017 17283 23075 17289
rect 2314 17212 2320 17264
rect 2372 17252 2378 17264
rect 2685 17255 2743 17261
rect 2685 17252 2697 17255
rect 2372 17224 2697 17252
rect 2372 17212 2378 17224
rect 2685 17221 2697 17224
rect 2731 17221 2743 17255
rect 2685 17215 2743 17221
rect 22097 17255 22155 17261
rect 22097 17221 22109 17255
rect 22143 17252 22155 17255
rect 23385 17255 23443 17261
rect 23385 17252 23397 17255
rect 22143 17224 23397 17252
rect 22143 17221 22155 17224
rect 22097 17215 22155 17221
rect 23385 17221 23397 17224
rect 23431 17221 23443 17255
rect 23385 17215 23443 17221
rect 25133 17255 25191 17261
rect 25133 17221 25145 17255
rect 25179 17252 25191 17255
rect 25774 17252 25780 17264
rect 25179 17224 25780 17252
rect 25179 17221 25191 17224
rect 25133 17215 25191 17221
rect 21545 17187 21603 17193
rect 21545 17153 21557 17187
rect 21591 17184 21603 17187
rect 23014 17184 23020 17196
rect 21591 17156 23020 17184
rect 21591 17153 21603 17156
rect 21545 17147 21603 17153
rect 23014 17144 23020 17156
rect 23072 17144 23078 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2501 17119 2559 17125
rect 1443 17088 2084 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 1581 16983 1639 16989
rect 1581 16949 1593 16983
rect 1627 16980 1639 16983
rect 1854 16980 1860 16992
rect 1627 16952 1860 16980
rect 1627 16949 1639 16952
rect 1581 16943 1639 16949
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 2056 16989 2084 17088
rect 2501 17085 2513 17119
rect 2547 17116 2559 17119
rect 20901 17119 20959 17125
rect 20901 17116 20913 17119
rect 2547 17088 3188 17116
rect 2547 17085 2559 17088
rect 2501 17079 2559 17085
rect 3160 16992 3188 17088
rect 20824 17088 20913 17116
rect 20824 16992 20852 17088
rect 20901 17085 20913 17088
rect 20947 17085 20959 17119
rect 23400 17116 23428 17215
rect 25774 17212 25780 17224
rect 25832 17212 25838 17264
rect 23661 17119 23719 17125
rect 23661 17116 23673 17119
rect 23400 17088 23673 17116
rect 20901 17079 20959 17085
rect 23661 17085 23673 17088
rect 23707 17085 23719 17119
rect 23661 17079 23719 17085
rect 24118 17076 24124 17128
rect 24176 17116 24182 17128
rect 24949 17119 25007 17125
rect 24949 17116 24961 17119
rect 24176 17088 24961 17116
rect 24176 17076 24182 17088
rect 24949 17085 24961 17088
rect 24995 17116 25007 17119
rect 25501 17119 25559 17125
rect 25501 17116 25513 17119
rect 24995 17088 25513 17116
rect 24995 17085 25007 17088
rect 24949 17079 25007 17085
rect 25501 17085 25513 17088
rect 25547 17085 25559 17119
rect 25501 17079 25559 17085
rect 22373 17051 22431 17057
rect 22373 17017 22385 17051
rect 22419 17017 22431 17051
rect 22646 17048 22652 17060
rect 22607 17020 22652 17048
rect 22373 17011 22431 17017
rect 2041 16983 2099 16989
rect 2041 16949 2053 16983
rect 2087 16980 2099 16983
rect 2682 16980 2688 16992
rect 2087 16952 2688 16980
rect 2087 16949 2099 16952
rect 2041 16943 2099 16949
rect 2682 16940 2688 16952
rect 2740 16940 2746 16992
rect 3142 16980 3148 16992
rect 3103 16952 3148 16980
rect 3142 16940 3148 16952
rect 3200 16940 3206 16992
rect 19889 16983 19947 16989
rect 19889 16949 19901 16983
rect 19935 16980 19947 16983
rect 20530 16980 20536 16992
rect 19935 16952 20536 16980
rect 19935 16949 19947 16952
rect 19889 16943 19947 16949
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 20806 16980 20812 16992
rect 20767 16952 20812 16980
rect 20806 16940 20812 16952
rect 20864 16940 20870 16992
rect 21082 16980 21088 16992
rect 21043 16952 21088 16980
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 21818 16980 21824 16992
rect 21779 16952 21824 16980
rect 21818 16940 21824 16952
rect 21876 16980 21882 16992
rect 22388 16980 22416 17011
rect 22646 17008 22652 17020
rect 22704 17008 22710 17060
rect 23474 17008 23480 17060
rect 23532 17048 23538 17060
rect 23937 17051 23995 17057
rect 23937 17048 23949 17051
rect 23532 17020 23949 17048
rect 23532 17008 23538 17020
rect 23937 17017 23949 17020
rect 23983 17017 23995 17051
rect 23937 17011 23995 17017
rect 22554 16980 22560 16992
rect 21876 16952 22416 16980
rect 22515 16952 22560 16980
rect 21876 16940 21882 16952
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 23658 16940 23664 16992
rect 23716 16980 23722 16992
rect 24581 16983 24639 16989
rect 24581 16980 24593 16983
rect 23716 16952 24593 16980
rect 23716 16940 23722 16952
rect 24581 16949 24593 16952
rect 24627 16980 24639 16983
rect 24670 16980 24676 16992
rect 24627 16952 24676 16980
rect 24627 16949 24639 16952
rect 24581 16943 24639 16949
rect 24670 16940 24676 16952
rect 24728 16940 24734 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2038 16776 2044 16788
rect 1999 16748 2044 16776
rect 2038 16736 2044 16748
rect 2096 16736 2102 16788
rect 2130 16736 2136 16788
rect 2188 16776 2194 16788
rect 2685 16779 2743 16785
rect 2685 16776 2697 16779
rect 2188 16748 2697 16776
rect 2188 16736 2194 16748
rect 2685 16745 2697 16748
rect 2731 16745 2743 16779
rect 2685 16739 2743 16745
rect 19797 16779 19855 16785
rect 19797 16745 19809 16779
rect 19843 16776 19855 16779
rect 21818 16776 21824 16788
rect 19843 16748 21824 16776
rect 19843 16745 19855 16748
rect 19797 16739 19855 16745
rect 21818 16736 21824 16748
rect 21876 16736 21882 16788
rect 22097 16779 22155 16785
rect 22097 16745 22109 16779
rect 22143 16776 22155 16779
rect 22646 16776 22652 16788
rect 22143 16748 22652 16776
rect 22143 16745 22155 16748
rect 22097 16739 22155 16745
rect 22646 16736 22652 16748
rect 22704 16776 22710 16788
rect 23934 16776 23940 16788
rect 22704 16748 23940 16776
rect 22704 16736 22710 16748
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 25225 16779 25283 16785
rect 25225 16745 25237 16779
rect 25271 16776 25283 16779
rect 25958 16776 25964 16788
rect 25271 16748 25964 16776
rect 25271 16745 25283 16748
rect 25225 16739 25283 16745
rect 25958 16736 25964 16748
rect 26016 16736 26022 16788
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2056 16640 2084 16736
rect 4617 16711 4675 16717
rect 4617 16677 4629 16711
rect 4663 16708 4675 16711
rect 4890 16708 4896 16720
rect 4663 16680 4896 16708
rect 4663 16677 4675 16680
rect 4617 16671 4675 16677
rect 4890 16668 4896 16680
rect 4948 16668 4954 16720
rect 22824 16711 22882 16717
rect 22824 16677 22836 16711
rect 22870 16708 22882 16711
rect 23014 16708 23020 16720
rect 22870 16680 23020 16708
rect 22870 16677 22882 16680
rect 22824 16671 22882 16677
rect 23014 16668 23020 16680
rect 23072 16668 23078 16720
rect 1443 16612 2084 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 2498 16600 2504 16652
rect 2556 16640 2562 16652
rect 2556 16612 2601 16640
rect 2556 16600 2562 16612
rect 2682 16600 2688 16652
rect 2740 16600 2746 16652
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4430 16640 4436 16652
rect 4120 16612 4436 16640
rect 4120 16600 4126 16612
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 10134 16640 10140 16652
rect 9999 16612 10140 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 15804 16612 16313 16640
rect 15804 16600 15810 16612
rect 16301 16609 16313 16612
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 17589 16643 17647 16649
rect 17589 16609 17601 16643
rect 17635 16640 17647 16643
rect 17862 16640 17868 16652
rect 17635 16612 17868 16640
rect 17635 16609 17647 16612
rect 17589 16603 17647 16609
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 18782 16640 18788 16652
rect 18743 16612 18788 16640
rect 18782 16600 18788 16612
rect 18840 16600 18846 16652
rect 21453 16643 21511 16649
rect 21453 16609 21465 16643
rect 21499 16640 21511 16643
rect 21818 16640 21824 16652
rect 21499 16612 21824 16640
rect 21499 16609 21511 16612
rect 21453 16603 21511 16609
rect 21818 16600 21824 16612
rect 21876 16600 21882 16652
rect 22465 16643 22523 16649
rect 22465 16609 22477 16643
rect 22511 16640 22523 16643
rect 23382 16640 23388 16652
rect 22511 16612 23388 16640
rect 22511 16609 22523 16612
rect 22465 16603 22523 16609
rect 23382 16600 23388 16612
rect 23440 16600 23446 16652
rect 25041 16643 25099 16649
rect 25041 16609 25053 16643
rect 25087 16640 25099 16643
rect 25314 16640 25320 16652
rect 25087 16612 25320 16640
rect 25087 16609 25099 16612
rect 25041 16603 25099 16609
rect 25314 16600 25320 16612
rect 25372 16600 25378 16652
rect 2700 16572 2728 16600
rect 4080 16572 4108 16600
rect 2700 16544 4108 16572
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 5258 16572 5264 16584
rect 4755 16544 5264 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 22554 16572 22560 16584
rect 22515 16544 22560 16572
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 21177 16507 21235 16513
rect 21177 16473 21189 16507
rect 21223 16504 21235 16507
rect 21542 16504 21548 16516
rect 21223 16476 21548 16504
rect 21223 16473 21235 16476
rect 21177 16467 21235 16473
rect 21542 16464 21548 16476
rect 21600 16464 21606 16516
rect 1210 16396 1216 16448
rect 1268 16436 1274 16448
rect 1581 16439 1639 16445
rect 1581 16436 1593 16439
rect 1268 16408 1593 16436
rect 1268 16396 1274 16408
rect 1581 16405 1593 16408
rect 1627 16405 1639 16439
rect 1581 16399 1639 16405
rect 2409 16439 2467 16445
rect 2409 16405 2421 16439
rect 2455 16436 2467 16439
rect 2866 16436 2872 16448
rect 2455 16408 2872 16436
rect 2455 16405 2467 16408
rect 2409 16399 2467 16405
rect 2866 16396 2872 16408
rect 2924 16396 2930 16448
rect 2958 16396 2964 16448
rect 3016 16436 3022 16448
rect 3145 16439 3203 16445
rect 3145 16436 3157 16439
rect 3016 16408 3157 16436
rect 3016 16396 3022 16408
rect 3145 16405 3157 16408
rect 3191 16436 3203 16439
rect 4157 16439 4215 16445
rect 4157 16436 4169 16439
rect 3191 16408 4169 16436
rect 3191 16405 3203 16408
rect 3145 16399 3203 16405
rect 4157 16405 4169 16408
rect 4203 16405 4215 16439
rect 4157 16399 4215 16405
rect 10505 16439 10563 16445
rect 10505 16405 10517 16439
rect 10551 16436 10563 16439
rect 10962 16436 10968 16448
rect 10551 16408 10968 16436
rect 10551 16405 10563 16408
rect 10505 16399 10563 16405
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 14277 16439 14335 16445
rect 14277 16405 14289 16439
rect 14323 16436 14335 16439
rect 14826 16436 14832 16448
rect 14323 16408 14832 16436
rect 14323 16405 14335 16408
rect 14277 16399 14335 16405
rect 14826 16396 14832 16408
rect 14884 16396 14890 16448
rect 21266 16396 21272 16448
rect 21324 16436 21330 16448
rect 21637 16439 21695 16445
rect 21637 16436 21649 16439
rect 21324 16408 21649 16436
rect 21324 16396 21330 16408
rect 21637 16405 21649 16408
rect 21683 16405 21695 16439
rect 21637 16399 21695 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 3973 16235 4031 16241
rect 3973 16201 3985 16235
rect 4019 16232 4031 16235
rect 4062 16232 4068 16244
rect 4019 16204 4068 16232
rect 4019 16201 4031 16204
rect 3973 16195 4031 16201
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 22465 16235 22523 16241
rect 22465 16201 22477 16235
rect 22511 16232 22523 16235
rect 23014 16232 23020 16244
rect 22511 16204 23020 16232
rect 22511 16201 22523 16204
rect 22465 16195 22523 16201
rect 23014 16192 23020 16204
rect 23072 16192 23078 16244
rect 2222 16124 2228 16176
rect 2280 16164 2286 16176
rect 2685 16167 2743 16173
rect 2685 16164 2697 16167
rect 2280 16136 2697 16164
rect 2280 16124 2286 16136
rect 2685 16133 2697 16136
rect 2731 16133 2743 16167
rect 2685 16127 2743 16133
rect 4157 16167 4215 16173
rect 4157 16133 4169 16167
rect 4203 16164 4215 16167
rect 4798 16164 4804 16176
rect 4203 16136 4804 16164
rect 4203 16133 4215 16136
rect 4157 16127 4215 16133
rect 4798 16124 4804 16136
rect 4856 16124 4862 16176
rect 10505 16167 10563 16173
rect 10505 16133 10517 16167
rect 10551 16164 10563 16167
rect 11790 16164 11796 16176
rect 10551 16136 11796 16164
rect 10551 16133 10563 16136
rect 10505 16127 10563 16133
rect 11790 16124 11796 16136
rect 11848 16124 11854 16176
rect 14277 16167 14335 16173
rect 14277 16133 14289 16167
rect 14323 16164 14335 16167
rect 15654 16164 15660 16176
rect 14323 16136 15660 16164
rect 14323 16133 14335 16136
rect 14277 16127 14335 16133
rect 15654 16124 15660 16136
rect 15712 16124 15718 16176
rect 2038 16096 2044 16108
rect 1412 16068 2044 16096
rect 1412 16037 1440 16068
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 14826 16096 14832 16108
rect 14787 16068 14832 16096
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 15997 2559 16031
rect 5813 16031 5871 16037
rect 5813 16028 5825 16031
rect 2501 15991 2559 15997
rect 4632 16000 5825 16028
rect 2516 15960 2544 15991
rect 4632 15972 4660 16000
rect 5813 15997 5825 16000
rect 5859 15997 5871 16031
rect 5813 15991 5871 15997
rect 10321 16031 10379 16037
rect 10321 15997 10333 16031
rect 10367 16028 10379 16031
rect 10686 16028 10692 16040
rect 10367 16000 10692 16028
rect 10367 15997 10379 16000
rect 10321 15991 10379 15997
rect 10686 15988 10692 16000
rect 10744 16028 10750 16040
rect 11057 16031 11115 16037
rect 11057 16028 11069 16031
rect 10744 16000 11069 16028
rect 10744 15988 10750 16000
rect 11057 15997 11069 16000
rect 11103 16028 11115 16031
rect 11882 16028 11888 16040
rect 11103 16000 11888 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 23934 16037 23940 16040
rect 14093 16031 14151 16037
rect 14093 15997 14105 16031
rect 14139 16028 14151 16031
rect 19981 16031 20039 16037
rect 14139 16000 14780 16028
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 14752 15972 14780 16000
rect 19981 15997 19993 16031
rect 20027 16028 20039 16031
rect 21085 16031 21143 16037
rect 21085 16028 21097 16031
rect 20027 16000 20668 16028
rect 20027 15997 20039 16000
rect 19981 15991 20039 15997
rect 3145 15963 3203 15969
rect 3145 15960 3157 15963
rect 2516 15932 3157 15960
rect 3145 15929 3157 15932
rect 3191 15960 3203 15963
rect 4062 15960 4068 15972
rect 3191 15932 4068 15960
rect 3191 15929 3203 15932
rect 3145 15923 3203 15929
rect 4062 15920 4068 15932
rect 4120 15920 4126 15972
rect 4338 15920 4344 15972
rect 4396 15960 4402 15972
rect 4433 15963 4491 15969
rect 4433 15960 4445 15963
rect 4396 15932 4445 15960
rect 4396 15920 4402 15932
rect 4433 15929 4445 15932
rect 4479 15929 4491 15963
rect 4614 15960 4620 15972
rect 4527 15932 4620 15960
rect 4433 15923 4491 15929
rect 4614 15920 4620 15932
rect 4672 15920 4678 15972
rect 4706 15920 4712 15972
rect 4764 15960 4770 15972
rect 5077 15963 5135 15969
rect 5077 15960 5089 15963
rect 4764 15932 5089 15960
rect 4764 15920 4770 15932
rect 5077 15929 5089 15932
rect 5123 15929 5135 15963
rect 9950 15960 9956 15972
rect 9863 15932 9956 15960
rect 5077 15923 5135 15929
rect 9950 15920 9956 15932
rect 10008 15960 10014 15972
rect 10781 15963 10839 15969
rect 10781 15960 10793 15963
rect 10008 15932 10793 15960
rect 10008 15920 10014 15932
rect 10781 15929 10793 15932
rect 10827 15929 10839 15963
rect 10962 15960 10968 15972
rect 10923 15932 10968 15960
rect 10781 15923 10839 15929
rect 10962 15920 10968 15932
rect 11020 15920 11026 15972
rect 14550 15960 14556 15972
rect 14511 15932 14556 15960
rect 14550 15920 14556 15932
rect 14608 15920 14614 15972
rect 14734 15960 14740 15972
rect 14695 15932 14740 15960
rect 14734 15920 14740 15932
rect 14792 15920 14798 15972
rect 20640 15904 20668 16000
rect 20916 16000 21097 16028
rect 20916 15904 20944 16000
rect 21085 15997 21097 16000
rect 21131 15997 21143 16031
rect 23661 16031 23719 16037
rect 23661 16028 23673 16031
rect 21085 15991 21143 15997
rect 23400 16000 23673 16028
rect 21352 15963 21410 15969
rect 21352 15929 21364 15963
rect 21398 15960 21410 15963
rect 21542 15960 21548 15972
rect 21398 15932 21548 15960
rect 21398 15929 21410 15932
rect 21352 15923 21410 15929
rect 21542 15920 21548 15932
rect 21600 15920 21606 15972
rect 937 15895 995 15901
rect 937 15861 949 15895
rect 983 15892 995 15895
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 983 15864 1593 15892
rect 983 15861 995 15864
rect 937 15855 995 15861
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 2409 15895 2467 15901
rect 2409 15861 2421 15895
rect 2455 15892 2467 15895
rect 2498 15892 2504 15904
rect 2455 15864 2504 15892
rect 2455 15861 2467 15864
rect 2409 15855 2467 15861
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 3605 15895 3663 15901
rect 3605 15861 3617 15895
rect 3651 15892 3663 15895
rect 4890 15892 4896 15904
rect 3651 15864 4896 15892
rect 3651 15861 3663 15864
rect 3605 15855 3663 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 5258 15852 5264 15904
rect 5316 15892 5322 15904
rect 5445 15895 5503 15901
rect 5445 15892 5457 15895
rect 5316 15864 5457 15892
rect 5316 15852 5322 15864
rect 5445 15861 5457 15864
rect 5491 15861 5503 15895
rect 5445 15855 5503 15861
rect 6273 15895 6331 15901
rect 6273 15861 6285 15895
rect 6319 15892 6331 15895
rect 6546 15892 6552 15904
rect 6319 15864 6552 15892
rect 6319 15861 6331 15864
rect 6273 15855 6331 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 6822 15892 6828 15904
rect 6687 15864 6828 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 16301 15895 16359 15901
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 16482 15892 16488 15904
rect 16347 15864 16488 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 18966 15892 18972 15904
rect 18927 15864 18972 15892
rect 18966 15852 18972 15864
rect 19024 15852 19030 15904
rect 20165 15895 20223 15901
rect 20165 15861 20177 15895
rect 20211 15892 20223 15895
rect 20438 15892 20444 15904
rect 20211 15864 20444 15892
rect 20211 15861 20223 15864
rect 20165 15855 20223 15861
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 20622 15892 20628 15904
rect 20583 15864 20628 15892
rect 20622 15852 20628 15864
rect 20680 15852 20686 15904
rect 20898 15892 20904 15904
rect 20859 15864 20904 15892
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 23106 15892 23112 15904
rect 22612 15864 23112 15892
rect 22612 15852 22618 15864
rect 23106 15852 23112 15864
rect 23164 15892 23170 15904
rect 23400 15901 23428 16000
rect 23661 15997 23673 16000
rect 23707 15997 23719 16031
rect 23928 16028 23940 16037
rect 23895 16000 23940 16028
rect 23661 15991 23719 15997
rect 23928 15991 23940 16000
rect 23934 15988 23940 15991
rect 23992 15988 23998 16040
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 23164 15864 23397 15892
rect 23164 15852 23170 15864
rect 23385 15861 23397 15864
rect 23431 15861 23443 15895
rect 25038 15892 25044 15904
rect 24999 15864 25044 15892
rect 23385 15855 23443 15861
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 25314 15852 25320 15904
rect 25372 15892 25378 15904
rect 25593 15895 25651 15901
rect 25593 15892 25605 15895
rect 25372 15864 25605 15892
rect 25372 15852 25378 15864
rect 25593 15861 25605 15864
rect 25639 15861 25651 15895
rect 25593 15855 25651 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2958 15688 2964 15700
rect 2919 15660 2964 15688
rect 2958 15648 2964 15660
rect 3016 15648 3022 15700
rect 11882 15688 11888 15700
rect 11843 15660 11888 15688
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 14277 15691 14335 15697
rect 14277 15657 14289 15691
rect 14323 15688 14335 15691
rect 14550 15688 14556 15700
rect 14323 15660 14556 15688
rect 14323 15657 14335 15660
rect 14277 15651 14335 15657
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 19797 15691 19855 15697
rect 19797 15657 19809 15691
rect 19843 15688 19855 15691
rect 19978 15688 19984 15700
rect 19843 15660 19984 15688
rect 19843 15657 19855 15660
rect 19797 15651 19855 15657
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 22925 15691 22983 15697
rect 22925 15657 22937 15691
rect 22971 15688 22983 15691
rect 23014 15688 23020 15700
rect 22971 15660 23020 15688
rect 22971 15657 22983 15660
rect 22925 15651 22983 15657
rect 23014 15648 23020 15660
rect 23072 15648 23078 15700
rect 23753 15691 23811 15697
rect 23753 15657 23765 15691
rect 23799 15688 23811 15691
rect 23934 15688 23940 15700
rect 23799 15660 23940 15688
rect 23799 15657 23811 15660
rect 23753 15651 23811 15657
rect 23934 15648 23940 15660
rect 23992 15648 23998 15700
rect 4890 15620 4896 15632
rect 4803 15592 4896 15620
rect 4890 15580 4896 15592
rect 4948 15620 4954 15632
rect 5442 15620 5448 15632
rect 4948 15592 5448 15620
rect 4948 15580 4954 15592
rect 5442 15580 5448 15592
rect 5500 15580 5506 15632
rect 9953 15623 10011 15629
rect 9953 15589 9965 15623
rect 9999 15620 10011 15623
rect 10594 15620 10600 15632
rect 9999 15592 10600 15620
rect 9999 15589 10011 15592
rect 9953 15583 10011 15589
rect 10594 15580 10600 15592
rect 10652 15620 10658 15632
rect 10750 15623 10808 15629
rect 10750 15620 10762 15623
rect 10652 15592 10762 15620
rect 10652 15580 10658 15592
rect 10750 15589 10762 15592
rect 10796 15589 10808 15623
rect 15654 15620 15660 15632
rect 15615 15592 15660 15620
rect 10750 15583 10808 15589
rect 15654 15580 15660 15592
rect 15712 15580 15718 15632
rect 15838 15620 15844 15632
rect 15799 15592 15844 15620
rect 15838 15580 15844 15592
rect 15896 15580 15902 15632
rect 20717 15623 20775 15629
rect 20717 15589 20729 15623
rect 20763 15620 20775 15623
rect 21818 15620 21824 15632
rect 20763 15592 21824 15620
rect 20763 15589 20775 15592
rect 20717 15583 20775 15589
rect 21818 15580 21824 15592
rect 21876 15580 21882 15632
rect 15672 15552 15700 15580
rect 16574 15552 16580 15564
rect 15672 15524 16580 15552
rect 16574 15512 16580 15524
rect 16632 15512 16638 15564
rect 18138 15552 18144 15564
rect 18099 15524 18144 15552
rect 18138 15512 18144 15524
rect 18196 15512 18202 15564
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19889 15555 19947 15561
rect 19889 15552 19901 15555
rect 19392 15524 19901 15552
rect 19392 15512 19398 15524
rect 19889 15521 19901 15524
rect 19935 15552 19947 15555
rect 20990 15552 20996 15564
rect 19935 15524 20996 15552
rect 19935 15521 19947 15524
rect 19889 15515 19947 15521
rect 20990 15512 20996 15524
rect 21048 15552 21054 15564
rect 21157 15555 21215 15561
rect 21157 15552 21169 15555
rect 21048 15524 21169 15552
rect 21048 15512 21054 15524
rect 21157 15521 21169 15524
rect 21203 15521 21215 15555
rect 21157 15515 21215 15521
rect 24204 15555 24262 15561
rect 24204 15521 24216 15555
rect 24250 15552 24262 15555
rect 25038 15552 25044 15564
rect 24250 15524 25044 15552
rect 24250 15521 24262 15524
rect 24204 15515 24262 15521
rect 25038 15512 25044 15524
rect 25096 15512 25102 15564
rect 1854 15444 1860 15496
rect 1912 15484 1918 15496
rect 2498 15484 2504 15496
rect 1912 15456 2504 15484
rect 1912 15444 1918 15456
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 2958 15484 2964 15496
rect 2919 15456 2964 15484
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 4890 15484 4896 15496
rect 3099 15456 3133 15484
rect 4851 15456 4896 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 2317 15419 2375 15425
rect 2317 15385 2329 15419
rect 2363 15416 2375 15419
rect 3068 15416 3096 15447
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15484 5043 15487
rect 5074 15484 5080 15496
rect 5031 15456 5080 15484
rect 5031 15453 5043 15456
rect 4985 15447 5043 15453
rect 5074 15444 5080 15456
rect 5132 15444 5138 15496
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 5905 15487 5963 15493
rect 5905 15484 5917 15487
rect 5592 15456 5917 15484
rect 5592 15444 5598 15456
rect 5905 15453 5917 15456
rect 5951 15453 5963 15487
rect 7006 15484 7012 15496
rect 6967 15456 7012 15484
rect 5905 15447 5963 15453
rect 7006 15444 7012 15456
rect 7064 15444 7070 15496
rect 8478 15484 8484 15496
rect 8439 15456 8484 15484
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 10502 15484 10508 15496
rect 10463 15456 10508 15484
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15484 13047 15487
rect 13078 15484 13084 15496
rect 13035 15456 13084 15484
rect 13035 15453 13047 15456
rect 12989 15447 13047 15453
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 15470 15444 15476 15496
rect 15528 15484 15534 15496
rect 15933 15487 15991 15493
rect 15933 15484 15945 15487
rect 15528 15456 15945 15484
rect 15528 15444 15534 15456
rect 15933 15453 15945 15456
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 17129 15487 17187 15493
rect 17129 15453 17141 15487
rect 17175 15484 17187 15487
rect 17586 15484 17592 15496
rect 17175 15456 17592 15484
rect 17175 15453 17187 15456
rect 17129 15447 17187 15453
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19484 15456 19717 15484
rect 19484 15444 19490 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 20898 15484 20904 15496
rect 20859 15456 20904 15484
rect 19705 15447 19763 15453
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 23934 15484 23940 15496
rect 23895 15456 23940 15484
rect 23934 15444 23940 15456
rect 23992 15444 23998 15496
rect 3418 15416 3424 15428
rect 2363 15388 3424 15416
rect 2363 15385 2375 15388
rect 2317 15379 2375 15385
rect 3418 15376 3424 15388
rect 3476 15376 3482 15428
rect 3513 15419 3571 15425
rect 3513 15385 3525 15419
rect 3559 15416 3571 15419
rect 4062 15416 4068 15428
rect 3559 15388 4068 15416
rect 3559 15385 3571 15388
rect 3513 15379 3571 15385
rect 4062 15376 4068 15388
rect 4120 15376 4126 15428
rect 4433 15419 4491 15425
rect 4433 15385 4445 15419
rect 4479 15416 4491 15419
rect 4614 15416 4620 15428
rect 4479 15388 4620 15416
rect 4479 15385 4491 15388
rect 4433 15379 4491 15385
rect 4614 15376 4620 15388
rect 4672 15376 4678 15428
rect 6270 15376 6276 15428
rect 6328 15416 6334 15428
rect 6733 15419 6791 15425
rect 6733 15416 6745 15419
rect 6328 15388 6745 15416
rect 6328 15376 6334 15388
rect 6733 15385 6745 15388
rect 6779 15385 6791 15419
rect 6733 15379 6791 15385
rect 19337 15419 19395 15425
rect 19337 15385 19349 15419
rect 19383 15416 19395 15419
rect 20714 15416 20720 15428
rect 19383 15388 20720 15416
rect 19383 15385 19395 15388
rect 19337 15379 19395 15385
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 1854 15348 1860 15360
rect 1815 15320 1860 15348
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 2501 15351 2559 15357
rect 2501 15317 2513 15351
rect 2547 15348 2559 15351
rect 2590 15348 2596 15360
rect 2547 15320 2596 15348
rect 2547 15317 2559 15320
rect 2501 15311 2559 15317
rect 2590 15308 2596 15320
rect 2648 15308 2654 15360
rect 3881 15351 3939 15357
rect 3881 15317 3893 15351
rect 3927 15348 3939 15351
rect 4338 15348 4344 15360
rect 3927 15320 4344 15348
rect 3927 15317 3939 15320
rect 3881 15311 3939 15317
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 5350 15348 5356 15360
rect 5311 15320 5356 15348
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 5813 15351 5871 15357
rect 5813 15317 5825 15351
rect 5859 15348 5871 15351
rect 5994 15348 6000 15360
rect 5859 15320 6000 15348
rect 5859 15317 5871 15320
rect 5813 15311 5871 15317
rect 5994 15308 6000 15320
rect 6052 15308 6058 15360
rect 6454 15348 6460 15360
rect 6415 15320 6460 15348
rect 6454 15308 6460 15320
rect 6512 15308 6518 15360
rect 12529 15351 12587 15357
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 12986 15348 12992 15360
rect 12575 15320 12992 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 15378 15348 15384 15360
rect 15339 15320 15384 15348
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 18322 15348 18328 15360
rect 18283 15320 18328 15348
rect 18322 15308 18328 15320
rect 18380 15308 18386 15360
rect 20346 15348 20352 15360
rect 20307 15320 20352 15348
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 21542 15308 21548 15360
rect 21600 15348 21606 15360
rect 22281 15351 22339 15357
rect 22281 15348 22293 15351
rect 21600 15320 22293 15348
rect 21600 15308 21606 15320
rect 22281 15317 22293 15320
rect 22327 15317 22339 15351
rect 22281 15311 22339 15317
rect 22554 15308 22560 15360
rect 22612 15348 22618 15360
rect 23201 15351 23259 15357
rect 23201 15348 23213 15351
rect 22612 15320 23213 15348
rect 22612 15308 22618 15320
rect 23201 15317 23213 15320
rect 23247 15317 23259 15351
rect 23201 15311 23259 15317
rect 24946 15308 24952 15360
rect 25004 15348 25010 15360
rect 25317 15351 25375 15357
rect 25317 15348 25329 15351
rect 25004 15320 25329 15348
rect 25004 15308 25010 15320
rect 25317 15317 25329 15320
rect 25363 15317 25375 15351
rect 25317 15311 25375 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2866 15144 2872 15156
rect 2827 15116 2872 15144
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 4341 15147 4399 15153
rect 4341 15113 4353 15147
rect 4387 15144 4399 15147
rect 4706 15144 4712 15156
rect 4387 15116 4712 15144
rect 4387 15113 4399 15116
rect 4341 15107 4399 15113
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 5353 15147 5411 15153
rect 5353 15113 5365 15147
rect 5399 15144 5411 15147
rect 5442 15144 5448 15156
rect 5399 15116 5448 15144
rect 5399 15113 5411 15116
rect 5353 15107 5411 15113
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 9674 15144 9680 15156
rect 9635 15116 9680 15144
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 9950 15144 9956 15156
rect 9911 15116 9956 15144
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 11790 15144 11796 15156
rect 11751 15116 11796 15144
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 14645 15147 14703 15153
rect 14645 15113 14657 15147
rect 14691 15144 14703 15147
rect 15470 15144 15476 15156
rect 14691 15116 15476 15144
rect 14691 15113 14703 15116
rect 14645 15107 14703 15113
rect 15470 15104 15476 15116
rect 15528 15144 15534 15156
rect 16390 15144 16396 15156
rect 15528 15116 16396 15144
rect 15528 15104 15534 15116
rect 16390 15104 16396 15116
rect 16448 15144 16454 15156
rect 16485 15147 16543 15153
rect 16485 15144 16497 15147
rect 16448 15116 16497 15144
rect 16448 15104 16454 15116
rect 16485 15113 16497 15116
rect 16531 15113 16543 15147
rect 16485 15107 16543 15113
rect 16574 15104 16580 15156
rect 16632 15144 16638 15156
rect 17037 15147 17095 15153
rect 17037 15144 17049 15147
rect 16632 15116 17049 15144
rect 16632 15104 16638 15116
rect 17037 15113 17049 15116
rect 17083 15113 17095 15147
rect 17037 15107 17095 15113
rect 18417 15147 18475 15153
rect 18417 15113 18429 15147
rect 18463 15144 18475 15147
rect 19242 15144 19248 15156
rect 18463 15116 19248 15144
rect 18463 15113 18475 15116
rect 18417 15107 18475 15113
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 19337 15147 19395 15153
rect 19337 15113 19349 15147
rect 19383 15144 19395 15147
rect 19426 15144 19432 15156
rect 19383 15116 19432 15144
rect 19383 15113 19395 15116
rect 19337 15107 19395 15113
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 20990 15144 20996 15156
rect 20951 15116 20996 15144
rect 20990 15104 20996 15116
rect 21048 15144 21054 15156
rect 21913 15147 21971 15153
rect 21913 15144 21925 15147
rect 21048 15116 21925 15144
rect 21048 15104 21054 15116
rect 21913 15113 21925 15116
rect 21959 15113 21971 15147
rect 21913 15107 21971 15113
rect 1762 14968 1768 15020
rect 1820 15008 1826 15020
rect 2884 15008 2912 15104
rect 12529 15079 12587 15085
rect 12529 15045 12541 15079
rect 12575 15076 12587 15079
rect 13906 15076 13912 15088
rect 12575 15048 13912 15076
rect 12575 15045 12587 15048
rect 12529 15039 12587 15045
rect 13906 15036 13912 15048
rect 13964 15036 13970 15088
rect 24489 15079 24547 15085
rect 24489 15045 24501 15079
rect 24535 15076 24547 15079
rect 24670 15076 24676 15088
rect 24535 15048 24676 15076
rect 24535 15045 24547 15048
rect 24489 15039 24547 15045
rect 24670 15036 24676 15048
rect 24728 15036 24734 15088
rect 2961 15011 3019 15017
rect 2961 15008 2973 15011
rect 1820 14980 2973 15008
rect 1820 14968 1826 14980
rect 2961 14977 2973 14980
rect 3007 14977 3019 15011
rect 2961 14971 3019 14977
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 15008 10563 15011
rect 10594 15008 10600 15020
rect 10551 14980 10600 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 10594 14968 10600 14980
rect 10652 15008 10658 15020
rect 11146 15008 11152 15020
rect 10652 14980 11152 15008
rect 10652 14968 10658 14980
rect 11146 14968 11152 14980
rect 11204 15008 11210 15020
rect 11241 15011 11299 15017
rect 11241 15008 11253 15011
rect 11204 14980 11253 15008
rect 11204 14968 11210 14980
rect 11241 14977 11253 14980
rect 11287 14977 11299 15011
rect 11241 14971 11299 14977
rect 12989 15011 13047 15017
rect 12989 14977 13001 15011
rect 13035 15008 13047 15011
rect 14093 15011 14151 15017
rect 13035 14980 13216 15008
rect 13035 14977 13047 14980
rect 12989 14971 13047 14977
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14909 1455 14943
rect 1397 14903 1455 14909
rect 1412 14872 1440 14903
rect 5258 14900 5264 14952
rect 5316 14940 5322 14952
rect 5445 14943 5503 14949
rect 5445 14940 5457 14943
rect 5316 14912 5457 14940
rect 5316 14900 5322 14912
rect 5445 14909 5457 14912
rect 5491 14940 5503 14943
rect 6181 14943 6239 14949
rect 6181 14940 6193 14943
rect 5491 14912 6193 14940
rect 5491 14909 5503 14912
rect 5445 14903 5503 14909
rect 6181 14909 6193 14912
rect 6227 14909 6239 14943
rect 6181 14903 6239 14909
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 2038 14872 2044 14884
rect 1412 14844 2044 14872
rect 2038 14832 2044 14844
rect 2096 14832 2102 14884
rect 2501 14875 2559 14881
rect 2501 14841 2513 14875
rect 2547 14872 2559 14875
rect 3142 14872 3148 14884
rect 2547 14844 3148 14872
rect 2547 14841 2559 14844
rect 2501 14835 2559 14841
rect 3142 14832 3148 14844
rect 3200 14881 3206 14884
rect 3200 14875 3264 14881
rect 3200 14841 3218 14875
rect 3252 14841 3264 14875
rect 3200 14835 3264 14841
rect 5721 14875 5779 14881
rect 5721 14841 5733 14875
rect 5767 14872 5779 14875
rect 6730 14872 6736 14884
rect 5767 14844 6736 14872
rect 5767 14841 5779 14844
rect 5721 14835 5779 14841
rect 3200 14832 3206 14835
rect 6730 14832 6736 14844
rect 6788 14832 6794 14884
rect 1578 14804 1584 14816
rect 1539 14776 1584 14804
rect 1578 14764 1584 14776
rect 1636 14764 1642 14816
rect 4982 14804 4988 14816
rect 4943 14776 4988 14804
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 6638 14804 6644 14816
rect 6599 14776 6644 14804
rect 6638 14764 6644 14776
rect 6696 14804 6702 14816
rect 6840 14804 6868 14903
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10229 14943 10287 14949
rect 10229 14940 10241 14943
rect 10192 14912 10241 14940
rect 10192 14900 10198 14912
rect 10229 14909 10241 14912
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12802 14940 12808 14952
rect 12299 14912 12808 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12802 14900 12808 14912
rect 12860 14940 12866 14952
rect 13081 14943 13139 14949
rect 13081 14940 13093 14943
rect 12860 14912 13093 14940
rect 12860 14900 12866 14912
rect 13081 14909 13093 14912
rect 13127 14909 13139 14943
rect 13081 14903 13139 14909
rect 6914 14832 6920 14884
rect 6972 14872 6978 14884
rect 7070 14875 7128 14881
rect 7070 14872 7082 14875
rect 6972 14844 7082 14872
rect 6972 14832 6978 14844
rect 7070 14841 7082 14844
rect 7116 14841 7128 14875
rect 7070 14835 7128 14841
rect 9674 14832 9680 14884
rect 9732 14872 9738 14884
rect 10413 14875 10471 14881
rect 10413 14872 10425 14875
rect 9732 14844 10425 14872
rect 9732 14832 9738 14844
rect 10413 14841 10425 14844
rect 10459 14841 10471 14875
rect 10413 14835 10471 14841
rect 10502 14832 10508 14884
rect 10560 14872 10566 14884
rect 10965 14875 11023 14881
rect 10965 14872 10977 14875
rect 10560 14844 10977 14872
rect 10560 14832 10566 14844
rect 10965 14841 10977 14844
rect 11011 14872 11023 14875
rect 12342 14872 12348 14884
rect 11011 14844 12348 14872
rect 11011 14841 11023 14844
rect 10965 14835 11023 14841
rect 12342 14832 12348 14844
rect 12400 14832 12406 14884
rect 12986 14872 12992 14884
rect 12947 14844 12992 14872
rect 12986 14832 12992 14844
rect 13044 14832 13050 14884
rect 6696 14776 6868 14804
rect 6696 14764 6702 14776
rect 7834 14764 7840 14816
rect 7892 14804 7898 14816
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 7892 14776 8217 14804
rect 7892 14764 7898 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 9122 14764 9128 14816
rect 9180 14804 9186 14816
rect 9309 14807 9367 14813
rect 9309 14804 9321 14807
rect 9180 14776 9321 14804
rect 9180 14764 9186 14776
rect 9309 14773 9321 14776
rect 9355 14773 9367 14807
rect 9309 14767 9367 14773
rect 11882 14764 11888 14816
rect 11940 14804 11946 14816
rect 13188 14804 13216 14980
rect 14093 14977 14105 15011
rect 14139 15008 14151 15011
rect 14550 15008 14556 15020
rect 14139 14980 14556 15008
rect 14139 14977 14151 14980
rect 14093 14971 14151 14977
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 15008 23167 15011
rect 25038 15008 25044 15020
rect 23155 14980 25044 15008
rect 23155 14977 23167 14980
rect 23109 14971 23167 14977
rect 25038 14968 25044 14980
rect 25096 14968 25102 15020
rect 15102 14940 15108 14952
rect 15063 14912 15108 14940
rect 15102 14900 15108 14912
rect 15160 14900 15166 14952
rect 18230 14900 18236 14952
rect 18288 14940 18294 14952
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18288 14912 18521 14940
rect 18288 14900 18294 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 19613 14943 19671 14949
rect 19613 14940 19625 14943
rect 19484 14912 19625 14940
rect 19484 14900 19490 14912
rect 19613 14909 19625 14912
rect 19659 14940 19671 14943
rect 20898 14940 20904 14952
rect 19659 14912 20904 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 20898 14900 20904 14912
rect 20956 14900 20962 14952
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 23937 14943 23995 14949
rect 22152 14912 22197 14940
rect 22152 14900 22158 14912
rect 23937 14909 23949 14943
rect 23983 14940 23995 14943
rect 23983 14912 24900 14940
rect 23983 14909 23995 14912
rect 23937 14903 23995 14909
rect 24872 14884 24900 14912
rect 14826 14832 14832 14884
rect 14884 14872 14890 14884
rect 15350 14875 15408 14881
rect 15350 14872 15362 14875
rect 14884 14844 15362 14872
rect 14884 14832 14890 14844
rect 15350 14841 15362 14844
rect 15396 14872 15408 14875
rect 15654 14872 15660 14884
rect 15396 14844 15660 14872
rect 15396 14841 15408 14844
rect 15350 14835 15408 14841
rect 15654 14832 15660 14844
rect 15712 14832 15718 14884
rect 17865 14875 17923 14881
rect 17865 14841 17877 14875
rect 17911 14872 17923 14875
rect 18138 14872 18144 14884
rect 17911 14844 18144 14872
rect 17911 14841 17923 14844
rect 17865 14835 17923 14841
rect 18138 14832 18144 14844
rect 18196 14872 18202 14884
rect 19242 14872 19248 14884
rect 18196 14844 19248 14872
rect 18196 14832 18202 14844
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 19880 14875 19938 14881
rect 19880 14841 19892 14875
rect 19926 14872 19938 14875
rect 20346 14872 20352 14884
rect 19926 14844 20352 14872
rect 19926 14841 19938 14844
rect 19880 14835 19938 14841
rect 20346 14832 20352 14844
rect 20404 14872 20410 14884
rect 22373 14875 22431 14881
rect 20404 14844 20668 14872
rect 20404 14832 20410 14844
rect 20640 14816 20668 14844
rect 22373 14841 22385 14875
rect 22419 14872 22431 14875
rect 23290 14872 23296 14884
rect 22419 14844 23296 14872
rect 22419 14841 22431 14844
rect 22373 14835 22431 14841
rect 23290 14832 23296 14844
rect 23348 14832 23354 14884
rect 24302 14872 24308 14884
rect 24215 14844 24308 14872
rect 24302 14832 24308 14844
rect 24360 14872 24366 14884
rect 24765 14875 24823 14881
rect 24765 14872 24777 14875
rect 24360 14844 24777 14872
rect 24360 14832 24366 14844
rect 24765 14841 24777 14844
rect 24811 14841 24823 14875
rect 24765 14835 24823 14841
rect 24854 14832 24860 14884
rect 24912 14872 24918 14884
rect 24949 14875 25007 14881
rect 24949 14872 24961 14875
rect 24912 14844 24961 14872
rect 24912 14832 24918 14844
rect 24949 14841 24961 14844
rect 24995 14841 25007 14875
rect 24949 14835 25007 14841
rect 11940 14776 13216 14804
rect 15013 14807 15071 14813
rect 11940 14764 11946 14776
rect 15013 14773 15025 14807
rect 15059 14804 15071 14807
rect 15102 14804 15108 14816
rect 15059 14776 15108 14804
rect 15059 14773 15071 14776
rect 15013 14767 15071 14773
rect 15102 14764 15108 14776
rect 15160 14804 15166 14816
rect 15562 14804 15568 14816
rect 15160 14776 15568 14804
rect 15160 14764 15166 14776
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 18690 14804 18696 14816
rect 18651 14776 18696 14804
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 20622 14764 20628 14816
rect 20680 14764 20686 14816
rect 21637 14807 21695 14813
rect 21637 14773 21649 14807
rect 21683 14804 21695 14807
rect 22646 14804 22652 14816
rect 21683 14776 22652 14804
rect 21683 14773 21695 14776
rect 21637 14767 21695 14773
rect 22646 14764 22652 14776
rect 22704 14804 22710 14816
rect 23106 14804 23112 14816
rect 22704 14776 23112 14804
rect 22704 14764 22710 14776
rect 23106 14764 23112 14776
rect 23164 14804 23170 14816
rect 23385 14807 23443 14813
rect 23385 14804 23397 14807
rect 23164 14776 23397 14804
rect 23164 14764 23170 14776
rect 23385 14773 23397 14776
rect 23431 14804 23443 14807
rect 23934 14804 23940 14816
rect 23431 14776 23940 14804
rect 23431 14773 23443 14776
rect 23385 14767 23443 14773
rect 23934 14764 23940 14776
rect 23992 14764 23998 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 3142 14600 3148 14612
rect 3055 14572 3148 14600
rect 2774 14492 2780 14544
rect 2832 14532 2838 14544
rect 3068 14541 3096 14572
rect 3142 14560 3148 14572
rect 3200 14600 3206 14612
rect 3881 14603 3939 14609
rect 3881 14600 3893 14603
rect 3200 14572 3893 14600
rect 3200 14560 3206 14572
rect 3881 14569 3893 14572
rect 3927 14600 3939 14603
rect 5074 14600 5080 14612
rect 3927 14572 5080 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 5074 14560 5080 14572
rect 5132 14560 5138 14612
rect 7190 14560 7196 14612
rect 7248 14600 7254 14612
rect 7745 14603 7803 14609
rect 7745 14600 7757 14603
rect 7248 14572 7757 14600
rect 7248 14560 7254 14572
rect 7745 14569 7757 14572
rect 7791 14569 7803 14603
rect 7745 14563 7803 14569
rect 9953 14603 10011 14609
rect 9953 14569 9965 14603
rect 9999 14600 10011 14603
rect 10134 14600 10140 14612
rect 9999 14572 10140 14600
rect 9999 14569 10011 14572
rect 9953 14563 10011 14569
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 10505 14603 10563 14609
rect 10505 14569 10517 14603
rect 10551 14600 10563 14603
rect 10686 14600 10692 14612
rect 10551 14572 10692 14600
rect 10551 14569 10563 14572
rect 10505 14563 10563 14569
rect 10686 14560 10692 14572
rect 10744 14600 10750 14612
rect 11330 14600 11336 14612
rect 10744 14572 11336 14600
rect 10744 14560 10750 14572
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 15654 14560 15660 14612
rect 15712 14600 15718 14612
rect 15749 14603 15807 14609
rect 15749 14600 15761 14603
rect 15712 14572 15761 14600
rect 15712 14560 15718 14572
rect 15749 14569 15761 14572
rect 15795 14569 15807 14603
rect 15749 14563 15807 14569
rect 19337 14603 19395 14609
rect 19337 14569 19349 14603
rect 19383 14600 19395 14603
rect 19978 14600 19984 14612
rect 19383 14572 19984 14600
rect 19383 14569 19395 14572
rect 19337 14563 19395 14569
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20714 14600 20720 14612
rect 20675 14572 20720 14600
rect 20714 14560 20720 14572
rect 20772 14600 20778 14612
rect 21453 14603 21511 14609
rect 21453 14600 21465 14603
rect 20772 14572 21465 14600
rect 20772 14560 20778 14572
rect 21453 14569 21465 14572
rect 21499 14569 21511 14603
rect 21453 14563 21511 14569
rect 22094 14560 22100 14612
rect 22152 14600 22158 14612
rect 24581 14603 24639 14609
rect 22152 14572 22197 14600
rect 22152 14560 22158 14572
rect 24581 14569 24593 14603
rect 24627 14600 24639 14603
rect 25038 14600 25044 14612
rect 24627 14572 25044 14600
rect 24627 14569 24639 14572
rect 24581 14563 24639 14569
rect 25038 14560 25044 14572
rect 25096 14560 25102 14612
rect 2961 14535 3019 14541
rect 2832 14504 2877 14532
rect 2832 14492 2838 14504
rect 2961 14501 2973 14535
rect 3007 14501 3019 14535
rect 2961 14495 3019 14501
rect 3053 14535 3111 14541
rect 3053 14501 3065 14535
rect 3099 14501 3111 14535
rect 3053 14495 3111 14501
rect 2976 14464 3004 14495
rect 4706 14492 4712 14544
rect 4764 14532 4770 14544
rect 4954 14535 5012 14541
rect 4954 14532 4966 14535
rect 4764 14504 4966 14532
rect 4764 14492 4770 14504
rect 4954 14501 4966 14504
rect 5000 14501 5012 14535
rect 4954 14495 5012 14501
rect 7006 14492 7012 14544
rect 7064 14532 7070 14544
rect 7561 14535 7619 14541
rect 7561 14532 7573 14535
rect 7064 14504 7573 14532
rect 7064 14492 7070 14504
rect 7561 14501 7573 14504
rect 7607 14501 7619 14535
rect 7561 14495 7619 14501
rect 7834 14492 7840 14544
rect 7892 14532 7898 14544
rect 10965 14535 11023 14541
rect 7892 14504 7937 14532
rect 7892 14492 7898 14504
rect 10965 14501 10977 14535
rect 11011 14532 11023 14535
rect 11054 14532 11060 14544
rect 11011 14504 11060 14532
rect 11011 14501 11023 14504
rect 10965 14495 11023 14501
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 11149 14535 11207 14541
rect 11149 14501 11161 14535
rect 11195 14501 11207 14535
rect 11149 14495 11207 14501
rect 3326 14464 3332 14476
rect 2976 14436 3332 14464
rect 3326 14424 3332 14436
rect 3384 14424 3390 14476
rect 10870 14424 10876 14476
rect 10928 14464 10934 14476
rect 11164 14464 11192 14495
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 12710 14532 12716 14544
rect 11848 14504 12716 14532
rect 11848 14492 11854 14504
rect 12710 14492 12716 14504
rect 12768 14492 12774 14544
rect 16390 14492 16396 14544
rect 16448 14532 16454 14544
rect 16574 14541 16580 14544
rect 16546 14535 16580 14541
rect 16546 14532 16558 14535
rect 16448 14504 16558 14532
rect 16448 14492 16454 14504
rect 16546 14501 16558 14504
rect 16632 14532 16638 14544
rect 16632 14504 16694 14532
rect 16546 14495 16580 14501
rect 16574 14492 16580 14495
rect 16632 14492 16638 14504
rect 20530 14492 20536 14544
rect 20588 14532 20594 14544
rect 21269 14535 21327 14541
rect 21269 14532 21281 14535
rect 20588 14504 21281 14532
rect 20588 14492 20594 14504
rect 21269 14501 21281 14504
rect 21315 14532 21327 14535
rect 21358 14532 21364 14544
rect 21315 14504 21364 14532
rect 21315 14501 21327 14504
rect 21269 14495 21327 14501
rect 21358 14492 21364 14504
rect 21416 14492 21422 14544
rect 24302 14532 24308 14544
rect 21458 14504 24308 14532
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 10928 14436 11192 14464
rect 11256 14436 12817 14464
rect 10928 14424 10934 14436
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 2590 14396 2596 14408
rect 1443 14368 2596 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 2866 14356 2872 14408
rect 2924 14396 2930 14408
rect 4614 14396 4620 14408
rect 2924 14368 4620 14396
rect 2924 14356 2930 14368
rect 4614 14356 4620 14368
rect 4672 14396 4678 14408
rect 4709 14399 4767 14405
rect 4709 14396 4721 14399
rect 4672 14368 4721 14396
rect 4672 14356 4678 14368
rect 4709 14365 4721 14368
rect 4755 14365 4767 14399
rect 4709 14359 4767 14365
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 11256 14405 11284 14436
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 15562 14424 15568 14476
rect 15620 14464 15626 14476
rect 16301 14467 16359 14473
rect 16301 14464 16313 14467
rect 15620 14436 16313 14464
rect 15620 14424 15626 14436
rect 16301 14433 16313 14436
rect 16347 14464 16359 14467
rect 16942 14464 16948 14476
rect 16347 14436 16948 14464
rect 16347 14433 16359 14436
rect 16301 14427 16359 14433
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 19705 14467 19763 14473
rect 19705 14433 19717 14467
rect 19751 14464 19763 14467
rect 20070 14464 20076 14476
rect 19751 14436 20076 14464
rect 19751 14433 19763 14436
rect 19705 14427 19763 14433
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 21458 14464 21486 14504
rect 24302 14492 24308 14504
rect 24360 14492 24366 14544
rect 25314 14532 25320 14544
rect 25275 14504 25320 14532
rect 25314 14492 25320 14504
rect 25372 14492 25378 14544
rect 20171 14436 21486 14464
rect 22557 14467 22615 14473
rect 11241 14399 11299 14405
rect 11241 14396 11253 14399
rect 11204 14368 11253 14396
rect 11204 14356 11210 14368
rect 11241 14365 11253 14368
rect 11287 14365 11299 14399
rect 12710 14396 12716 14408
rect 12671 14368 12716 14396
rect 11241 14359 11299 14365
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 12986 14356 12992 14408
rect 13044 14396 13050 14408
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13044 14368 13737 14396
rect 13044 14356 13050 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 13725 14359 13783 14365
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 18414 14356 18420 14408
rect 18472 14396 18478 14408
rect 20171 14396 20199 14436
rect 22557 14433 22569 14467
rect 22603 14464 22615 14467
rect 22646 14464 22652 14476
rect 22603 14436 22652 14464
rect 22603 14433 22615 14436
rect 22557 14427 22615 14433
rect 22646 14424 22652 14436
rect 22704 14424 22710 14476
rect 22824 14467 22882 14473
rect 22824 14433 22836 14467
rect 22870 14464 22882 14467
rect 23106 14464 23112 14476
rect 22870 14436 23112 14464
rect 22870 14433 22882 14436
rect 22824 14427 22882 14433
rect 23106 14424 23112 14436
rect 23164 14424 23170 14476
rect 25038 14464 25044 14476
rect 24999 14436 25044 14464
rect 25038 14424 25044 14436
rect 25096 14424 25102 14476
rect 18472 14368 20199 14396
rect 18472 14356 18478 14368
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 21542 14396 21548 14408
rect 20772 14368 21548 14396
rect 20772 14356 20778 14368
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 2317 14331 2375 14337
rect 1412 14300 2176 14328
rect 1412 14272 1440 14300
rect 1394 14220 1400 14272
rect 1452 14220 1458 14272
rect 1949 14263 2007 14269
rect 1949 14229 1961 14263
rect 1995 14260 2007 14263
rect 2038 14260 2044 14272
rect 1995 14232 2044 14260
rect 1995 14229 2007 14232
rect 1949 14223 2007 14229
rect 2038 14220 2044 14232
rect 2096 14220 2102 14272
rect 2148 14260 2176 14300
rect 2317 14297 2329 14331
rect 2363 14328 2375 14331
rect 3142 14328 3148 14340
rect 2363 14300 3148 14328
rect 2363 14297 2375 14300
rect 2317 14291 2375 14297
rect 3142 14288 3148 14300
rect 3200 14288 3206 14340
rect 7282 14328 7288 14340
rect 7243 14300 7288 14328
rect 7282 14288 7288 14300
rect 7340 14288 7346 14340
rect 10689 14331 10747 14337
rect 10689 14297 10701 14331
rect 10735 14328 10747 14331
rect 10962 14328 10968 14340
rect 10735 14300 10968 14328
rect 10735 14297 10747 14300
rect 10689 14291 10747 14297
rect 10962 14288 10968 14300
rect 11020 14288 11026 14340
rect 14734 14288 14740 14340
rect 14792 14328 14798 14340
rect 15838 14328 15844 14340
rect 14792 14300 15844 14328
rect 14792 14288 14798 14300
rect 15838 14288 15844 14300
rect 15896 14328 15902 14340
rect 16117 14331 16175 14337
rect 16117 14328 16129 14331
rect 15896 14300 16129 14328
rect 15896 14288 15902 14300
rect 16117 14297 16129 14300
rect 16163 14297 16175 14331
rect 16117 14291 16175 14297
rect 20993 14331 21051 14337
rect 20993 14297 21005 14331
rect 21039 14328 21051 14331
rect 22094 14328 22100 14340
rect 21039 14300 22100 14328
rect 21039 14297 21051 14300
rect 20993 14291 21051 14297
rect 22094 14288 22100 14300
rect 22152 14288 22158 14340
rect 2501 14263 2559 14269
rect 2501 14260 2513 14263
rect 2148 14232 2513 14260
rect 2501 14229 2513 14232
rect 2547 14229 2559 14263
rect 2501 14223 2559 14229
rect 2682 14220 2688 14272
rect 2740 14260 2746 14272
rect 3421 14263 3479 14269
rect 3421 14260 3433 14263
rect 2740 14232 3433 14260
rect 2740 14220 2746 14232
rect 3421 14229 3433 14232
rect 3467 14229 3479 14263
rect 4246 14260 4252 14272
rect 4207 14232 4252 14260
rect 3421 14223 3479 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 6086 14260 6092 14272
rect 6047 14232 6092 14260
rect 6086 14220 6092 14232
rect 6144 14260 6150 14272
rect 6825 14263 6883 14269
rect 6825 14260 6837 14263
rect 6144 14232 6837 14260
rect 6144 14220 6150 14232
rect 6825 14229 6837 14232
rect 6871 14260 6883 14263
rect 6914 14260 6920 14272
rect 6871 14232 6920 14260
rect 6871 14229 6883 14232
rect 6825 14223 6883 14229
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 8297 14263 8355 14269
rect 8297 14229 8309 14263
rect 8343 14260 8355 14263
rect 8386 14260 8392 14272
rect 8343 14232 8392 14260
rect 8343 14229 8355 14232
rect 8297 14223 8355 14229
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 8570 14260 8576 14272
rect 8531 14232 8576 14260
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 8938 14260 8944 14272
rect 8899 14232 8944 14260
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 9401 14263 9459 14269
rect 9401 14260 9413 14263
rect 9272 14232 9413 14260
rect 9272 14220 9278 14232
rect 9401 14229 9413 14232
rect 9447 14229 9459 14263
rect 11606 14260 11612 14272
rect 11567 14232 11612 14260
rect 9401 14223 9459 14229
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 11974 14260 11980 14272
rect 11935 14232 11980 14260
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12250 14260 12256 14272
rect 12211 14232 12256 14260
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12434 14220 12440 14272
rect 12492 14260 12498 14272
rect 13170 14260 13176 14272
rect 12492 14232 13176 14260
rect 12492 14220 12498 14232
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 17678 14260 17684 14272
rect 17639 14232 17684 14260
rect 17678 14220 17684 14232
rect 17736 14220 17742 14272
rect 18230 14220 18236 14272
rect 18288 14260 18294 14272
rect 18509 14263 18567 14269
rect 18509 14260 18521 14263
rect 18288 14232 18521 14260
rect 18288 14220 18294 14232
rect 18509 14229 18521 14232
rect 18555 14229 18567 14263
rect 19886 14260 19892 14272
rect 19847 14232 19892 14260
rect 18509 14223 18567 14229
rect 19886 14220 19892 14232
rect 19944 14220 19950 14272
rect 19978 14220 19984 14272
rect 20036 14260 20042 14272
rect 20257 14263 20315 14269
rect 20257 14260 20269 14263
rect 20036 14232 20269 14260
rect 20036 14220 20042 14232
rect 20257 14229 20269 14232
rect 20303 14229 20315 14263
rect 20257 14223 20315 14229
rect 20898 14220 20904 14272
rect 20956 14260 20962 14272
rect 23658 14260 23664 14272
rect 20956 14232 23664 14260
rect 20956 14220 20962 14232
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 23934 14260 23940 14272
rect 23895 14232 23940 14260
rect 23934 14220 23940 14232
rect 23992 14220 23998 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1673 14059 1731 14065
rect 1673 14025 1685 14059
rect 1719 14056 1731 14059
rect 1719 14028 2728 14056
rect 1719 14025 1731 14028
rect 1673 14019 1731 14025
rect 2700 13988 2728 14028
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 3697 14059 3755 14065
rect 3697 14056 3709 14059
rect 2832 14028 3709 14056
rect 2832 14016 2838 14028
rect 3697 14025 3709 14028
rect 3743 14025 3755 14059
rect 4338 14056 4344 14068
rect 4299 14028 4344 14056
rect 3697 14019 3755 14025
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 4706 14016 4712 14068
rect 4764 14056 4770 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 4764 14028 5641 14056
rect 4764 14016 4770 14028
rect 5629 14025 5641 14028
rect 5675 14025 5687 14059
rect 5629 14019 5687 14025
rect 6638 14016 6644 14068
rect 6696 14016 6702 14068
rect 7190 14056 7196 14068
rect 7151 14028 7196 14056
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 10778 14056 10784 14068
rect 10739 14028 10784 14056
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11790 14056 11796 14068
rect 11751 14028 11796 14056
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 12710 14056 12716 14068
rect 12299 14028 12716 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 13817 14059 13875 14065
rect 13817 14056 13829 14059
rect 12860 14028 13829 14056
rect 12860 14016 12866 14028
rect 13817 14025 13829 14028
rect 13863 14025 13875 14059
rect 13817 14019 13875 14025
rect 14829 14059 14887 14065
rect 14829 14025 14841 14059
rect 14875 14056 14887 14059
rect 15562 14056 15568 14068
rect 14875 14028 15568 14056
rect 14875 14025 14887 14028
rect 14829 14019 14887 14025
rect 3142 13988 3148 14000
rect 2700 13960 3004 13988
rect 3103 13960 3148 13988
rect 1762 13920 1768 13932
rect 1723 13892 1768 13920
rect 1762 13880 1768 13892
rect 1820 13880 1826 13932
rect 2976 13920 3004 13960
rect 3142 13948 3148 13960
rect 3200 13948 3206 14000
rect 4614 13948 4620 14000
rect 4672 13988 4678 14000
rect 5261 13991 5319 13997
rect 5261 13988 5273 13991
rect 4672 13960 5273 13988
rect 4672 13948 4678 13960
rect 5261 13957 5273 13960
rect 5307 13988 5319 13991
rect 6457 13991 6515 13997
rect 6457 13988 6469 13991
rect 5307 13960 6469 13988
rect 5307 13957 5319 13960
rect 5261 13951 5319 13957
rect 6457 13957 6469 13960
rect 6503 13988 6515 13991
rect 6549 13991 6607 13997
rect 6549 13988 6561 13991
rect 6503 13960 6561 13988
rect 6503 13957 6515 13960
rect 6457 13951 6515 13957
rect 6549 13957 6561 13960
rect 6595 13988 6607 13991
rect 6656 13988 6684 14016
rect 6595 13960 6684 13988
rect 9861 13991 9919 13997
rect 6595 13957 6607 13960
rect 6549 13951 6607 13957
rect 9861 13957 9873 13991
rect 9907 13988 9919 13991
rect 11146 13988 11152 14000
rect 9907 13960 11152 13988
rect 9907 13957 9919 13960
rect 9861 13951 9919 13957
rect 11146 13948 11152 13960
rect 11204 13948 11210 14000
rect 11330 13948 11336 14000
rect 11388 13988 11394 14000
rect 12434 13988 12440 14000
rect 11388 13960 12440 13988
rect 11388 13948 11394 13960
rect 12434 13948 12440 13960
rect 12492 13948 12498 14000
rect 3326 13920 3332 13932
rect 2976 13892 3332 13920
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13920 4951 13923
rect 5074 13920 5080 13932
rect 4939 13892 5080 13920
rect 4939 13889 4951 13892
rect 4893 13883 4951 13889
rect 5074 13880 5080 13892
rect 5132 13880 5138 13932
rect 6273 13923 6331 13929
rect 6273 13889 6285 13923
rect 6319 13920 6331 13923
rect 6638 13920 6644 13932
rect 6319 13892 6644 13920
rect 6319 13889 6331 13892
rect 6273 13883 6331 13889
rect 6638 13880 6644 13892
rect 6696 13920 6702 13932
rect 6696 13892 7420 13920
rect 6696 13880 6702 13892
rect 2038 13861 2044 13864
rect 2032 13852 2044 13861
rect 1999 13824 2044 13852
rect 2032 13815 2044 13824
rect 2038 13812 2044 13815
rect 2096 13812 2102 13864
rect 4338 13812 4344 13864
rect 4396 13852 4402 13864
rect 4617 13855 4675 13861
rect 4617 13852 4629 13855
rect 4396 13824 4629 13852
rect 4396 13812 4402 13824
rect 4617 13821 4629 13824
rect 4663 13821 4675 13855
rect 4617 13815 4675 13821
rect 6457 13855 6515 13861
rect 6457 13821 6469 13855
rect 6503 13852 6515 13855
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 6503 13824 7297 13852
rect 6503 13821 6515 13824
rect 6457 13815 6515 13821
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 7392 13852 7420 13892
rect 10962 13880 10968 13932
rect 11020 13920 11026 13932
rect 11241 13923 11299 13929
rect 11241 13920 11253 13923
rect 11020 13892 11253 13920
rect 11020 13880 11026 13892
rect 11241 13889 11253 13892
rect 11287 13920 11299 13923
rect 11606 13920 11612 13932
rect 11287 13892 11612 13920
rect 11287 13889 11299 13892
rect 11241 13883 11299 13889
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 13538 13880 13544 13932
rect 13596 13920 13602 13932
rect 14936 13929 14964 14028
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 15654 14016 15660 14068
rect 15712 14056 15718 14068
rect 16301 14059 16359 14065
rect 16301 14056 16313 14059
rect 15712 14028 16313 14056
rect 15712 14016 15718 14028
rect 16301 14025 16313 14028
rect 16347 14025 16359 14059
rect 21358 14056 21364 14068
rect 21319 14028 21364 14056
rect 16301 14019 16359 14025
rect 21358 14016 21364 14028
rect 21416 14016 21422 14068
rect 21726 14016 21732 14068
rect 21784 14056 21790 14068
rect 21821 14059 21879 14065
rect 21821 14056 21833 14059
rect 21784 14028 21833 14056
rect 21784 14016 21790 14028
rect 21821 14025 21833 14028
rect 21867 14025 21879 14059
rect 21821 14019 21879 14025
rect 18509 13991 18567 13997
rect 18509 13957 18521 13991
rect 18555 13988 18567 13991
rect 19334 13988 19340 14000
rect 18555 13960 19340 13988
rect 18555 13957 18567 13960
rect 18509 13951 18567 13957
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 20622 13948 20628 14000
rect 20680 13988 20686 14000
rect 20809 13991 20867 13997
rect 20809 13988 20821 13991
rect 20680 13960 20821 13988
rect 20680 13948 20686 13960
rect 20809 13957 20821 13960
rect 20855 13957 20867 13991
rect 20809 13951 20867 13957
rect 14921 13923 14979 13929
rect 14921 13920 14933 13923
rect 13596 13892 14933 13920
rect 13596 13880 13602 13892
rect 14921 13889 14933 13892
rect 14967 13889 14979 13923
rect 21836 13920 21864 14019
rect 23382 14016 23388 14068
rect 23440 14056 23446 14068
rect 23842 14056 23848 14068
rect 23440 14028 23848 14056
rect 23440 14016 23446 14028
rect 23842 14016 23848 14028
rect 23900 14016 23906 14068
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25501 14059 25559 14065
rect 25501 14056 25513 14059
rect 24912 14028 25513 14056
rect 24912 14016 24918 14028
rect 25501 14025 25513 14028
rect 25547 14025 25559 14059
rect 25501 14019 25559 14025
rect 22094 13948 22100 14000
rect 22152 13988 22158 14000
rect 22152 13960 22197 13988
rect 22152 13948 22158 13960
rect 22465 13923 22523 13929
rect 22465 13920 22477 13923
rect 21836 13892 22477 13920
rect 14921 13883 14979 13889
rect 22465 13889 22477 13892
rect 22511 13889 22523 13923
rect 22465 13883 22523 13889
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 23014 13920 23020 13932
rect 22695 13892 23020 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 23014 13880 23020 13892
rect 23072 13920 23078 13932
rect 23934 13920 23940 13932
rect 23072 13892 23940 13920
rect 23072 13880 23078 13892
rect 23934 13880 23940 13892
rect 23992 13880 23998 13932
rect 7552 13855 7610 13861
rect 7552 13852 7564 13855
rect 7392 13824 7564 13852
rect 7285 13815 7343 13821
rect 7552 13821 7564 13824
rect 7598 13852 7610 13855
rect 7834 13852 7840 13864
rect 7598 13824 7840 13852
rect 7598 13821 7610 13824
rect 7552 13815 7610 13821
rect 7300 13784 7328 13815
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13852 9551 13855
rect 12250 13852 12256 13864
rect 9539 13824 12256 13852
rect 9539 13821 9551 13824
rect 9493 13815 9551 13821
rect 7650 13784 7656 13796
rect 7300 13756 7656 13784
rect 7650 13744 7656 13756
rect 7708 13744 7714 13796
rect 10229 13787 10287 13793
rect 10229 13753 10241 13787
rect 10275 13784 10287 13787
rect 11054 13784 11060 13796
rect 10275 13756 11060 13784
rect 10275 13753 10287 13756
rect 10229 13747 10287 13753
rect 11054 13744 11060 13756
rect 11112 13744 11118 13796
rect 11256 13793 11284 13824
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 12434 13852 12440 13864
rect 12395 13824 12440 13852
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12704 13855 12762 13861
rect 12704 13821 12716 13855
rect 12750 13852 12762 13855
rect 13170 13852 13176 13864
rect 12750 13824 13176 13852
rect 12750 13821 12762 13824
rect 12704 13815 12762 13821
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 15177 13855 15235 13861
rect 15177 13852 15189 13855
rect 15120 13824 15189 13852
rect 11241 13787 11299 13793
rect 11241 13753 11253 13787
rect 11287 13753 11299 13787
rect 11241 13747 11299 13753
rect 11330 13744 11336 13796
rect 11388 13784 11394 13796
rect 11388 13756 11433 13784
rect 11388 13744 11394 13756
rect 14826 13744 14832 13796
rect 14884 13784 14890 13796
rect 15120 13784 15148 13824
rect 15177 13821 15189 13824
rect 15223 13821 15235 13855
rect 18322 13852 18328 13864
rect 18235 13824 18328 13852
rect 15177 13815 15235 13821
rect 18322 13812 18328 13824
rect 18380 13852 18386 13864
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 18380 13824 18889 13852
rect 18380 13812 18386 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 19426 13852 19432 13864
rect 19339 13824 19432 13852
rect 18877 13815 18935 13821
rect 19426 13812 19432 13824
rect 19484 13852 19490 13864
rect 24118 13852 24124 13864
rect 19484 13824 19840 13852
rect 24079 13824 24124 13852
rect 19484 13812 19490 13824
rect 14884 13756 15148 13784
rect 14884 13744 14890 13756
rect 19150 13744 19156 13796
rect 19208 13784 19214 13796
rect 19674 13787 19732 13793
rect 19674 13784 19686 13787
rect 19208 13756 19686 13784
rect 19208 13744 19214 13756
rect 19674 13753 19686 13756
rect 19720 13753 19732 13787
rect 19674 13747 19732 13753
rect 1210 13676 1216 13728
rect 1268 13716 1274 13728
rect 1486 13716 1492 13728
rect 1268 13688 1492 13716
rect 1268 13676 1274 13688
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 4154 13716 4160 13728
rect 4067 13688 4160 13716
rect 4154 13676 4160 13688
rect 4212 13716 4218 13728
rect 4801 13719 4859 13725
rect 4801 13716 4813 13719
rect 4212 13688 4813 13716
rect 4212 13676 4218 13688
rect 4801 13685 4813 13688
rect 4847 13716 4859 13719
rect 4982 13716 4988 13728
rect 4847 13688 4988 13716
rect 4847 13685 4859 13688
rect 4801 13679 4859 13685
rect 4982 13676 4988 13688
rect 5040 13676 5046 13728
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 7466 13716 7472 13728
rect 6972 13688 7472 13716
rect 6972 13676 6978 13688
rect 7466 13676 7472 13688
rect 7524 13676 7530 13728
rect 7834 13676 7840 13728
rect 7892 13716 7898 13728
rect 8665 13719 8723 13725
rect 8665 13716 8677 13719
rect 7892 13688 8677 13716
rect 7892 13676 7898 13688
rect 8665 13685 8677 13688
rect 8711 13685 8723 13719
rect 8665 13679 8723 13685
rect 10597 13719 10655 13725
rect 10597 13685 10609 13719
rect 10643 13716 10655 13719
rect 10778 13716 10784 13728
rect 10643 13688 10784 13716
rect 10643 13685 10655 13688
rect 10597 13679 10655 13685
rect 10778 13676 10784 13688
rect 10836 13676 10842 13728
rect 14366 13716 14372 13728
rect 14327 13688 14372 13716
rect 14366 13676 14372 13688
rect 14424 13676 14430 13728
rect 16206 13676 16212 13728
rect 16264 13716 16270 13728
rect 16390 13716 16396 13728
rect 16264 13688 16396 13716
rect 16264 13676 16270 13688
rect 16390 13676 16396 13688
rect 16448 13676 16454 13728
rect 16942 13716 16948 13728
rect 16855 13688 16948 13716
rect 16942 13676 16948 13688
rect 17000 13716 17006 13728
rect 17218 13716 17224 13728
rect 17000 13688 17224 13716
rect 17000 13676 17006 13688
rect 17218 13676 17224 13688
rect 17276 13676 17282 13728
rect 19337 13719 19395 13725
rect 19337 13685 19349 13719
rect 19383 13716 19395 13719
rect 19812 13716 19840 13824
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 24388 13855 24446 13861
rect 24388 13821 24400 13855
rect 24434 13852 24446 13855
rect 24946 13852 24952 13864
rect 24434 13824 24952 13852
rect 24434 13821 24446 13824
rect 24388 13815 24446 13821
rect 22094 13744 22100 13796
rect 22152 13784 22158 13796
rect 22554 13784 22560 13796
rect 22152 13756 22560 13784
rect 22152 13744 22158 13756
rect 22554 13744 22560 13756
rect 22612 13744 22618 13796
rect 23477 13787 23535 13793
rect 23477 13753 23489 13787
rect 23523 13784 23535 13787
rect 24403 13784 24431 13815
rect 24946 13812 24952 13824
rect 25004 13812 25010 13864
rect 23523 13756 24431 13784
rect 23523 13753 23535 13756
rect 23477 13747 23535 13753
rect 19978 13716 19984 13728
rect 19383 13688 19984 13716
rect 19383 13685 19395 13688
rect 19337 13679 19395 13685
rect 19978 13676 19984 13688
rect 20036 13676 20042 13728
rect 22738 13676 22744 13728
rect 22796 13716 22802 13728
rect 23017 13719 23075 13725
rect 23017 13716 23029 13719
rect 22796 13688 23029 13716
rect 22796 13676 22802 13688
rect 23017 13685 23029 13688
rect 23063 13716 23075 13719
rect 23937 13719 23995 13725
rect 23937 13716 23949 13719
rect 23063 13688 23949 13716
rect 23063 13685 23075 13688
rect 23017 13679 23075 13685
rect 23937 13685 23949 13688
rect 23983 13716 23995 13719
rect 24118 13716 24124 13728
rect 23983 13688 24124 13716
rect 23983 13685 23995 13688
rect 23937 13679 23995 13685
rect 24118 13676 24124 13688
rect 24176 13676 24182 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1394 13472 1400 13524
rect 1452 13512 1458 13524
rect 1762 13512 1768 13524
rect 1452 13484 1768 13512
rect 1452 13472 1458 13484
rect 1762 13472 1768 13484
rect 1820 13472 1826 13524
rect 3697 13515 3755 13521
rect 3697 13481 3709 13515
rect 3743 13512 3755 13515
rect 4706 13512 4712 13524
rect 3743 13484 4712 13512
rect 3743 13481 3755 13484
rect 3697 13475 3755 13481
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 5074 13512 5080 13524
rect 5035 13484 5080 13512
rect 5074 13472 5080 13484
rect 5132 13472 5138 13524
rect 5442 13472 5448 13524
rect 5500 13472 5506 13524
rect 6638 13512 6644 13524
rect 6599 13484 6644 13512
rect 6638 13472 6644 13484
rect 6696 13472 6702 13524
rect 7006 13512 7012 13524
rect 6967 13484 7012 13512
rect 7006 13472 7012 13484
rect 7064 13472 7070 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 7484 13484 8953 13512
rect 2774 13404 2780 13456
rect 2832 13444 2838 13456
rect 4614 13444 4620 13456
rect 2832 13416 2877 13444
rect 4527 13416 4620 13444
rect 2832 13404 2838 13416
rect 4614 13404 4620 13416
rect 4672 13444 4678 13456
rect 5460 13444 5488 13472
rect 5994 13444 6000 13456
rect 4672 13416 5488 13444
rect 5955 13416 6000 13444
rect 4672 13404 4678 13416
rect 5994 13404 6000 13416
rect 6052 13404 6058 13456
rect 6181 13447 6239 13453
rect 6181 13413 6193 13447
rect 6227 13444 6239 13447
rect 7190 13444 7196 13456
rect 6227 13416 7196 13444
rect 6227 13413 6239 13416
rect 6181 13407 6239 13413
rect 7190 13404 7196 13416
rect 7248 13444 7254 13456
rect 7484 13444 7512 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 8941 13475 8999 13481
rect 11057 13515 11115 13521
rect 11057 13481 11069 13515
rect 11103 13512 11115 13515
rect 11146 13512 11152 13524
rect 11103 13484 11152 13512
rect 11103 13481 11115 13484
rect 11057 13475 11115 13481
rect 11146 13472 11152 13484
rect 11204 13512 11210 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 11204 13484 11621 13512
rect 11204 13472 11210 13484
rect 11609 13481 11621 13484
rect 11655 13512 11667 13515
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11655 13484 12081 13512
rect 11655 13481 11667 13484
rect 11609 13475 11667 13481
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 15654 13472 15660 13524
rect 15712 13512 15718 13524
rect 16117 13515 16175 13521
rect 16117 13512 16129 13515
rect 15712 13484 16129 13512
rect 15712 13472 15718 13484
rect 16117 13481 16129 13484
rect 16163 13512 16175 13515
rect 16390 13512 16396 13524
rect 16163 13484 16396 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 16574 13512 16580 13524
rect 16535 13484 16580 13512
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 20070 13472 20076 13524
rect 20128 13512 20134 13524
rect 20257 13515 20315 13521
rect 20257 13512 20269 13515
rect 20128 13484 20269 13512
rect 20128 13472 20134 13484
rect 20257 13481 20269 13484
rect 20303 13481 20315 13515
rect 20714 13512 20720 13524
rect 20675 13484 20720 13512
rect 20257 13475 20315 13481
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 21174 13472 21180 13524
rect 21232 13512 21238 13524
rect 21453 13515 21511 13521
rect 21453 13512 21465 13515
rect 21232 13484 21465 13512
rect 21232 13472 21238 13484
rect 21453 13481 21465 13484
rect 21499 13481 21511 13515
rect 24670 13512 24676 13524
rect 24631 13484 24676 13512
rect 21453 13475 21511 13481
rect 24670 13472 24676 13484
rect 24728 13472 24734 13524
rect 7742 13444 7748 13456
rect 7248 13416 7512 13444
rect 7655 13416 7748 13444
rect 7248 13404 7254 13416
rect 7742 13404 7748 13416
rect 7800 13444 7806 13456
rect 8573 13447 8631 13453
rect 8573 13444 8585 13447
rect 7800 13416 8585 13444
rect 7800 13404 7806 13416
rect 8573 13413 8585 13416
rect 8619 13413 8631 13447
rect 13538 13444 13544 13456
rect 8573 13407 8631 13413
rect 12728 13416 13544 13444
rect 1670 13336 1676 13388
rect 1728 13376 1734 13388
rect 2593 13379 2651 13385
rect 2593 13376 2605 13379
rect 1728 13348 2605 13376
rect 1728 13336 1734 13348
rect 2593 13345 2605 13348
rect 2639 13345 2651 13379
rect 2593 13339 2651 13345
rect 3510 13336 3516 13388
rect 3568 13376 3574 13388
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 3568 13348 4445 13376
rect 3568 13336 3574 13348
rect 4433 13345 4445 13348
rect 4479 13376 4491 13379
rect 5442 13376 5448 13388
rect 4479 13348 5448 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 7558 13376 7564 13388
rect 7519 13348 7564 13376
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 7834 13376 7840 13388
rect 7795 13348 7840 13376
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 9933 13379 9991 13385
rect 9933 13376 9945 13379
rect 9456 13348 9945 13376
rect 9456 13336 9462 13348
rect 9933 13345 9945 13348
rect 9979 13345 9991 13379
rect 9933 13339 9991 13345
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 12728 13385 12756 13416
rect 13538 13404 13544 13416
rect 13596 13404 13602 13456
rect 16206 13404 16212 13456
rect 16264 13444 16270 13456
rect 17037 13447 17095 13453
rect 17037 13444 17049 13447
rect 16264 13416 17049 13444
rect 16264 13404 16270 13416
rect 17037 13413 17049 13416
rect 17083 13444 17095 13447
rect 17396 13447 17454 13453
rect 17396 13444 17408 13447
rect 17083 13416 17408 13444
rect 17083 13413 17095 13416
rect 17037 13407 17095 13413
rect 17396 13413 17408 13416
rect 17442 13444 17454 13447
rect 17678 13444 17684 13456
rect 17442 13416 17684 13444
rect 17442 13413 17454 13416
rect 17396 13407 17454 13413
rect 17678 13404 17684 13416
rect 17736 13404 17742 13456
rect 22186 13444 22192 13456
rect 21744 13416 22192 13444
rect 12529 13379 12587 13385
rect 12529 13376 12541 13379
rect 12492 13348 12541 13376
rect 12492 13336 12498 13348
rect 12529 13345 12541 13348
rect 12575 13376 12587 13379
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12575 13348 12725 13376
rect 12575 13345 12587 13348
rect 12529 13339 12587 13345
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 12969 13379 13027 13385
rect 12969 13376 12981 13379
rect 12860 13348 12981 13376
rect 12860 13336 12866 13348
rect 12969 13345 12981 13348
rect 13015 13345 13027 13379
rect 12969 13339 13027 13345
rect 17129 13379 17187 13385
rect 17129 13345 17141 13379
rect 17175 13376 17187 13379
rect 17218 13376 17224 13388
rect 17175 13348 17224 13376
rect 17175 13345 17187 13348
rect 17129 13339 17187 13345
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13376 19763 13379
rect 20346 13376 20352 13388
rect 19751 13348 20352 13376
rect 19751 13345 19763 13348
rect 19705 13339 19763 13345
rect 20346 13336 20352 13348
rect 20404 13336 20410 13388
rect 21269 13379 21327 13385
rect 21269 13345 21281 13379
rect 21315 13376 21327 13379
rect 21744 13376 21772 13416
rect 22186 13404 22192 13416
rect 22244 13404 22250 13456
rect 23014 13453 23020 13456
rect 23008 13444 23020 13453
rect 22940 13416 23020 13444
rect 21315 13348 21772 13376
rect 22097 13379 22155 13385
rect 21315 13345 21327 13348
rect 21269 13339 21327 13345
rect 22097 13345 22109 13379
rect 22143 13376 22155 13379
rect 22940 13376 22968 13416
rect 23008 13407 23020 13416
rect 23014 13404 23020 13407
rect 23072 13404 23078 13456
rect 25222 13376 25228 13388
rect 22143 13348 22968 13376
rect 25183 13348 25228 13376
rect 22143 13345 22155 13348
rect 22097 13339 22155 13345
rect 25222 13336 25228 13348
rect 25280 13336 25286 13388
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13277 2927 13311
rect 2869 13271 2927 13277
rect 2317 13175 2375 13181
rect 2317 13141 2329 13175
rect 2363 13172 2375 13175
rect 2682 13172 2688 13184
rect 2363 13144 2688 13172
rect 2363 13141 2375 13144
rect 2317 13135 2375 13141
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 2884 13172 2912 13271
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4709 13311 4767 13317
rect 4709 13308 4721 13311
rect 4120 13280 4721 13308
rect 4120 13268 4126 13280
rect 4709 13277 4721 13280
rect 4755 13308 4767 13311
rect 5074 13308 5080 13320
rect 4755 13280 5080 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 6236 13280 6285 13308
rect 6236 13268 6242 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 9732 13280 9777 13308
rect 9732 13268 9738 13280
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15896 13280 16129 13308
rect 15896 13268 15902 13280
rect 16117 13277 16129 13280
rect 16163 13308 16175 13311
rect 16298 13308 16304 13320
rect 16163 13280 16304 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 21542 13308 21548 13320
rect 21503 13280 21548 13308
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 22554 13268 22560 13320
rect 22612 13308 22618 13320
rect 22738 13308 22744 13320
rect 22612 13280 22744 13308
rect 22612 13268 22618 13280
rect 22738 13268 22744 13280
rect 22796 13268 22802 13320
rect 4154 13240 4160 13252
rect 4067 13212 4160 13240
rect 4154 13200 4160 13212
rect 4212 13240 4218 13252
rect 5350 13240 5356 13252
rect 4212 13212 5356 13240
rect 4212 13200 4218 13212
rect 5350 13200 5356 13212
rect 5408 13200 5414 13252
rect 5718 13240 5724 13252
rect 5679 13212 5724 13240
rect 5718 13200 5724 13212
rect 5776 13200 5782 13252
rect 7285 13243 7343 13249
rect 7285 13209 7297 13243
rect 7331 13240 7343 13243
rect 8202 13240 8208 13252
rect 7331 13212 8208 13240
rect 7331 13209 7343 13212
rect 7285 13203 7343 13209
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 15657 13243 15715 13249
rect 15657 13209 15669 13243
rect 15703 13240 15715 13243
rect 16666 13240 16672 13252
rect 15703 13212 16672 13240
rect 15703 13209 15715 13212
rect 15657 13203 15715 13209
rect 16666 13200 16672 13212
rect 16724 13200 16730 13252
rect 3142 13172 3148 13184
rect 2884 13144 3148 13172
rect 3142 13132 3148 13144
rect 3200 13172 3206 13184
rect 3237 13175 3295 13181
rect 3237 13172 3249 13175
rect 3200 13144 3249 13172
rect 3200 13132 3206 13144
rect 3237 13141 3249 13144
rect 3283 13141 3295 13175
rect 3237 13135 3295 13141
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 5445 13175 5503 13181
rect 5445 13172 5457 13175
rect 3384 13144 5457 13172
rect 3384 13132 3390 13144
rect 5445 13141 5457 13144
rect 5491 13141 5503 13175
rect 8294 13172 8300 13184
rect 8255 13144 8300 13172
rect 5445 13135 5503 13141
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 9493 13175 9551 13181
rect 9493 13141 9505 13175
rect 9539 13172 9551 13175
rect 9674 13172 9680 13184
rect 9539 13144 9680 13172
rect 9539 13141 9551 13144
rect 9493 13135 9551 13141
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 14093 13175 14151 13181
rect 14093 13141 14105 13175
rect 14139 13172 14151 13175
rect 14182 13172 14188 13184
rect 14139 13144 14188 13172
rect 14139 13141 14151 13144
rect 14093 13135 14151 13141
rect 14182 13132 14188 13144
rect 14240 13172 14246 13184
rect 14826 13172 14832 13184
rect 14240 13144 14832 13172
rect 14240 13132 14246 13144
rect 14826 13132 14832 13144
rect 14884 13172 14890 13184
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 14884 13144 14933 13172
rect 14884 13132 14890 13144
rect 14921 13141 14933 13144
rect 14967 13141 14979 13175
rect 18506 13172 18512 13184
rect 18467 13144 18512 13172
rect 14921 13135 14979 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 19150 13132 19156 13184
rect 19208 13172 19214 13184
rect 19429 13175 19487 13181
rect 19429 13172 19441 13175
rect 19208 13144 19441 13172
rect 19208 13132 19214 13144
rect 19429 13141 19441 13144
rect 19475 13141 19487 13175
rect 19429 13135 19487 13141
rect 19889 13175 19947 13181
rect 19889 13141 19901 13175
rect 19935 13172 19947 13175
rect 20070 13172 20076 13184
rect 19935 13144 20076 13172
rect 19935 13141 19947 13144
rect 19889 13135 19947 13141
rect 20070 13132 20076 13144
rect 20128 13132 20134 13184
rect 20990 13172 20996 13184
rect 20951 13144 20996 13172
rect 20990 13132 20996 13144
rect 21048 13132 21054 13184
rect 22649 13175 22707 13181
rect 22649 13141 22661 13175
rect 22695 13172 22707 13175
rect 23106 13172 23112 13184
rect 22695 13144 23112 13172
rect 22695 13141 22707 13144
rect 22649 13135 22707 13141
rect 23106 13132 23112 13144
rect 23164 13132 23170 13184
rect 24118 13172 24124 13184
rect 24079 13144 24124 13172
rect 24118 13132 24124 13144
rect 24176 13132 24182 13184
rect 25038 13172 25044 13184
rect 24999 13144 25044 13172
rect 25038 13132 25044 13144
rect 25096 13132 25102 13184
rect 25409 13175 25467 13181
rect 25409 13141 25421 13175
rect 25455 13172 25467 13175
rect 26142 13172 26148 13184
rect 25455 13144 26148 13172
rect 25455 13141 25467 13144
rect 25409 13135 25467 13141
rect 26142 13132 26148 13144
rect 26200 13132 26206 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1670 12968 1676 12980
rect 1631 12940 1676 12968
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 1949 12971 2007 12977
rect 1949 12968 1961 12971
rect 1912 12940 1961 12968
rect 1912 12928 1918 12940
rect 1949 12937 1961 12940
rect 1995 12937 2007 12971
rect 3510 12968 3516 12980
rect 3471 12940 3516 12968
rect 1949 12931 2007 12937
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 4614 12968 4620 12980
rect 4575 12940 4620 12968
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 5258 12968 5264 12980
rect 5219 12940 5264 12968
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 7469 12971 7527 12977
rect 7469 12937 7481 12971
rect 7515 12968 7527 12971
rect 7834 12968 7840 12980
rect 7515 12940 7840 12968
rect 7515 12937 7527 12940
rect 7469 12931 7527 12937
rect 3326 12900 3332 12912
rect 2424 12872 3332 12900
rect 1946 12792 1952 12844
rect 2004 12832 2010 12844
rect 2424 12841 2452 12872
rect 3326 12860 3332 12872
rect 3384 12860 3390 12912
rect 3697 12903 3755 12909
rect 3697 12869 3709 12903
rect 3743 12900 3755 12903
rect 3743 12872 5672 12900
rect 3743 12869 3755 12872
rect 3697 12863 3755 12869
rect 2409 12835 2467 12841
rect 2409 12832 2421 12835
rect 2004 12804 2421 12832
rect 2004 12792 2010 12804
rect 2409 12801 2421 12804
rect 2455 12801 2467 12835
rect 2409 12795 2467 12801
rect 2498 12792 2504 12844
rect 2556 12832 2562 12844
rect 2866 12832 2872 12844
rect 2556 12804 2872 12832
rect 2556 12792 2562 12804
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 4154 12832 4160 12844
rect 4115 12804 4160 12832
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12832 4307 12835
rect 4706 12832 4712 12844
rect 4295 12804 4712 12832
rect 4295 12801 4307 12804
rect 4249 12795 4307 12801
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 5644 12841 5672 12872
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12832 5687 12835
rect 5718 12832 5724 12844
rect 5675 12804 5724 12832
rect 5675 12801 5687 12804
rect 5629 12795 5687 12801
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 4430 12724 4436 12776
rect 4488 12764 4494 12776
rect 4614 12764 4620 12776
rect 4488 12736 4620 12764
rect 4488 12724 4494 12736
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5813 12767 5871 12773
rect 5813 12764 5825 12767
rect 5123 12736 5825 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5813 12733 5825 12736
rect 5859 12764 5871 12767
rect 6086 12764 6092 12776
rect 5859 12736 6092 12764
rect 5859 12733 5871 12736
rect 5813 12727 5871 12733
rect 6086 12724 6092 12736
rect 6144 12724 6150 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 7484 12764 7512 12931
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 9398 12968 9404 12980
rect 9359 12940 9404 12968
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 10873 12971 10931 12977
rect 10873 12937 10885 12971
rect 10919 12968 10931 12971
rect 10962 12968 10968 12980
rect 10919 12940 10968 12968
rect 10919 12937 10931 12940
rect 10873 12931 10931 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 13538 12968 13544 12980
rect 13499 12940 13544 12968
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 14369 12971 14427 12977
rect 14369 12937 14381 12971
rect 14415 12968 14427 12971
rect 14734 12968 14740 12980
rect 14415 12940 14740 12968
rect 14415 12937 14427 12940
rect 14369 12931 14427 12937
rect 14734 12928 14740 12940
rect 14792 12928 14798 12980
rect 15930 12968 15936 12980
rect 15891 12940 15936 12968
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 21821 12971 21879 12977
rect 21821 12968 21833 12971
rect 21232 12940 21833 12968
rect 21232 12928 21238 12940
rect 21821 12937 21833 12940
rect 21867 12937 21879 12971
rect 22186 12968 22192 12980
rect 22147 12940 22192 12968
rect 21821 12931 21879 12937
rect 22186 12928 22192 12940
rect 22244 12928 22250 12980
rect 23382 12968 23388 12980
rect 23343 12940 23388 12968
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 24029 12971 24087 12977
rect 24029 12937 24041 12971
rect 24075 12968 24087 12971
rect 25038 12968 25044 12980
rect 24075 12940 25044 12968
rect 24075 12937 24087 12940
rect 24029 12931 24087 12937
rect 25038 12928 25044 12940
rect 25096 12928 25102 12980
rect 25222 12968 25228 12980
rect 25183 12940 25228 12968
rect 25222 12928 25228 12940
rect 25280 12928 25286 12980
rect 25682 12968 25688 12980
rect 25643 12940 25688 12968
rect 25682 12928 25688 12940
rect 25740 12928 25746 12980
rect 12434 12860 12440 12912
rect 12492 12900 12498 12912
rect 12529 12903 12587 12909
rect 12529 12900 12541 12903
rect 12492 12872 12541 12900
rect 12492 12860 12498 12872
rect 12529 12869 12541 12872
rect 12575 12869 12587 12903
rect 12529 12863 12587 12869
rect 14550 12860 14556 12912
rect 14608 12900 14614 12912
rect 14826 12900 14832 12912
rect 14608 12872 14832 12900
rect 14608 12860 14614 12872
rect 14826 12860 14832 12872
rect 14884 12860 14890 12912
rect 15657 12903 15715 12909
rect 15657 12869 15669 12903
rect 15703 12900 15715 12903
rect 15838 12900 15844 12912
rect 15703 12872 15844 12900
rect 15703 12869 15715 12872
rect 15657 12863 15715 12869
rect 15838 12860 15844 12872
rect 15896 12860 15902 12912
rect 16209 12903 16267 12909
rect 16209 12869 16221 12903
rect 16255 12900 16267 12903
rect 16390 12900 16396 12912
rect 16255 12872 16396 12900
rect 16255 12869 16267 12872
rect 16209 12863 16267 12869
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 18417 12903 18475 12909
rect 18417 12869 18429 12903
rect 18463 12900 18475 12903
rect 19426 12900 19432 12912
rect 18463 12872 19432 12900
rect 18463 12869 18475 12872
rect 18417 12863 18475 12869
rect 19426 12860 19432 12872
rect 19484 12860 19490 12912
rect 7650 12792 7656 12844
rect 7708 12832 7714 12844
rect 7837 12835 7895 12841
rect 7837 12832 7849 12835
rect 7708 12804 7849 12832
rect 7708 12792 7714 12804
rect 7837 12801 7849 12804
rect 7883 12832 7895 12835
rect 8021 12835 8079 12841
rect 8021 12832 8033 12835
rect 7883 12804 8033 12832
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 8021 12801 8033 12804
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 11146 12792 11152 12844
rect 11204 12832 11210 12844
rect 11425 12835 11483 12841
rect 11425 12832 11437 12835
rect 11204 12804 11437 12832
rect 11204 12792 11210 12804
rect 11425 12801 11437 12804
rect 11471 12801 11483 12835
rect 11425 12795 11483 12801
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 12986 12832 12992 12844
rect 11931 12804 12992 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12832 14243 12835
rect 14734 12832 14740 12844
rect 14231 12804 14740 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 16574 12832 16580 12844
rect 16535 12804 16580 12832
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 16761 12835 16819 12841
rect 16761 12801 16773 12835
rect 16807 12832 16819 12835
rect 17678 12832 17684 12844
rect 16807 12804 17684 12832
rect 16807 12801 16819 12804
rect 16761 12795 16819 12801
rect 17678 12792 17684 12804
rect 17736 12832 17742 12844
rect 18506 12832 18512 12844
rect 17736 12804 18512 12832
rect 17736 12792 17742 12804
rect 18506 12792 18512 12804
rect 18564 12792 18570 12844
rect 18782 12832 18788 12844
rect 18743 12804 18788 12832
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 22554 12792 22560 12844
rect 22612 12832 22618 12844
rect 22925 12835 22983 12841
rect 22925 12832 22937 12835
rect 22612 12804 22937 12832
rect 22612 12792 22618 12804
rect 22925 12801 22937 12804
rect 22971 12801 22983 12835
rect 22925 12795 22983 12801
rect 24486 12792 24492 12844
rect 24544 12832 24550 12844
rect 24581 12835 24639 12841
rect 24581 12832 24593 12835
rect 24544 12804 24593 12832
rect 24544 12792 24550 12804
rect 24581 12801 24593 12804
rect 24627 12832 24639 12835
rect 24946 12832 24952 12844
rect 24627 12804 24952 12832
rect 24627 12801 24639 12804
rect 24581 12795 24639 12801
rect 24946 12792 24952 12804
rect 25004 12792 25010 12844
rect 6871 12736 7512 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 14642 12724 14648 12776
rect 14700 12764 14706 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14700 12736 14933 12764
rect 14700 12724 14706 12736
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 14921 12727 14979 12733
rect 15654 12724 15660 12776
rect 15712 12764 15718 12776
rect 15838 12764 15844 12776
rect 15712 12736 15844 12764
rect 15712 12724 15718 12736
rect 15838 12724 15844 12736
rect 15896 12724 15902 12776
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 19889 12767 19947 12773
rect 19889 12764 19901 12767
rect 19843 12736 19901 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 19889 12733 19901 12736
rect 19935 12764 19947 12767
rect 19978 12764 19984 12776
rect 19935 12736 19984 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 20156 12767 20214 12773
rect 20156 12764 20168 12767
rect 20088 12736 20168 12764
rect 2498 12696 2504 12708
rect 2459 12668 2504 12696
rect 2498 12656 2504 12668
rect 2556 12656 2562 12708
rect 4154 12696 4160 12708
rect 4115 12668 4160 12696
rect 4154 12656 4160 12668
rect 4212 12656 4218 12708
rect 4798 12656 4804 12708
rect 4856 12696 4862 12708
rect 5721 12699 5779 12705
rect 5721 12696 5733 12699
rect 4856 12668 5733 12696
rect 4856 12656 4862 12668
rect 5721 12665 5733 12668
rect 5767 12696 5779 12699
rect 5994 12696 6000 12708
rect 5767 12668 6000 12696
rect 5767 12665 5779 12668
rect 5721 12659 5779 12665
rect 5994 12656 6000 12668
rect 6052 12656 6058 12708
rect 6178 12656 6184 12708
rect 6236 12696 6242 12708
rect 6273 12699 6331 12705
rect 6273 12696 6285 12699
rect 6236 12668 6285 12696
rect 6236 12656 6242 12668
rect 6273 12665 6285 12668
rect 6319 12696 6331 12699
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 6319 12668 6653 12696
rect 6319 12665 6331 12668
rect 6273 12659 6331 12665
rect 6641 12665 6653 12668
rect 6687 12696 6699 12699
rect 7926 12696 7932 12708
rect 6687 12668 7932 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 7926 12656 7932 12668
rect 7984 12696 7990 12708
rect 8294 12705 8300 12708
rect 8266 12699 8300 12705
rect 8266 12696 8278 12699
rect 7984 12668 8278 12696
rect 7984 12656 7990 12668
rect 8266 12665 8278 12668
rect 8352 12696 8358 12708
rect 8352 12668 8414 12696
rect 8266 12659 8300 12665
rect 8294 12656 8300 12659
rect 8352 12656 8358 12668
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 10045 12699 10103 12705
rect 10045 12696 10057 12699
rect 9824 12668 10057 12696
rect 9824 12656 9830 12668
rect 10045 12665 10057 12668
rect 10091 12696 10103 12699
rect 10962 12696 10968 12708
rect 10091 12668 10968 12696
rect 10091 12665 10103 12668
rect 10045 12659 10103 12665
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 11054 12656 11060 12708
rect 11112 12696 11118 12708
rect 11149 12699 11207 12705
rect 11149 12696 11161 12699
rect 11112 12668 11161 12696
rect 11112 12656 11118 12668
rect 11149 12665 11161 12668
rect 11195 12665 11207 12699
rect 11149 12659 11207 12665
rect 13081 12699 13139 12705
rect 13081 12665 13093 12699
rect 13127 12696 13139 12699
rect 13630 12696 13636 12708
rect 13127 12668 13636 12696
rect 13127 12665 13139 12668
rect 13081 12659 13139 12665
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 13814 12656 13820 12708
rect 13872 12696 13878 12708
rect 14366 12696 14372 12708
rect 13872 12668 14372 12696
rect 13872 12656 13878 12668
rect 14366 12656 14372 12668
rect 14424 12696 14430 12708
rect 14829 12699 14887 12705
rect 14829 12696 14841 12699
rect 14424 12668 14841 12696
rect 14424 12656 14430 12668
rect 14829 12665 14841 12668
rect 14875 12665 14887 12699
rect 14829 12659 14887 12665
rect 15930 12656 15936 12708
rect 15988 12696 15994 12708
rect 16669 12699 16727 12705
rect 16669 12696 16681 12699
rect 15988 12668 16681 12696
rect 15988 12656 15994 12668
rect 16669 12665 16681 12668
rect 16715 12665 16727 12699
rect 17770 12696 17776 12708
rect 17731 12668 17776 12696
rect 16669 12659 16727 12665
rect 17770 12656 17776 12668
rect 17828 12696 17834 12708
rect 18874 12696 18880 12708
rect 17828 12668 18880 12696
rect 17828 12656 17834 12668
rect 18874 12656 18880 12668
rect 18932 12656 18938 12708
rect 18969 12699 19027 12705
rect 18969 12665 18981 12699
rect 19015 12696 19027 12699
rect 19429 12699 19487 12705
rect 19015 12668 19196 12696
rect 19015 12665 19027 12668
rect 18969 12659 19027 12665
rect 19168 12640 19196 12668
rect 19429 12665 19441 12699
rect 19475 12696 19487 12699
rect 20088 12696 20116 12736
rect 20156 12733 20168 12736
rect 20202 12764 20214 12767
rect 20714 12764 20720 12776
rect 20202 12736 20720 12764
rect 20202 12733 20214 12736
rect 20156 12727 20214 12733
rect 20714 12724 20720 12736
rect 20772 12764 20778 12776
rect 21542 12764 21548 12776
rect 20772 12736 21548 12764
rect 20772 12724 20778 12736
rect 21542 12724 21548 12736
rect 21600 12724 21606 12776
rect 22373 12767 22431 12773
rect 22373 12733 22385 12767
rect 22419 12764 22431 12767
rect 22646 12764 22652 12776
rect 22419 12736 22652 12764
rect 22419 12733 22431 12736
rect 22373 12727 22431 12733
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 23382 12724 23388 12776
rect 23440 12764 23446 12776
rect 24305 12767 24363 12773
rect 24305 12764 24317 12767
rect 23440 12736 24317 12764
rect 23440 12724 23446 12736
rect 24305 12733 24317 12736
rect 24351 12733 24363 12767
rect 25498 12764 25504 12776
rect 25459 12736 25504 12764
rect 24305 12727 24363 12733
rect 25498 12724 25504 12736
rect 25556 12764 25562 12776
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 25556 12736 26065 12764
rect 25556 12724 25562 12736
rect 26053 12733 26065 12736
rect 26099 12733 26111 12767
rect 26053 12727 26111 12733
rect 19475 12668 20116 12696
rect 19475 12665 19487 12668
rect 19429 12659 19487 12665
rect 2409 12631 2467 12637
rect 2409 12597 2421 12631
rect 2455 12628 2467 12631
rect 2682 12628 2688 12640
rect 2455 12600 2688 12628
rect 2455 12597 2467 12600
rect 2409 12591 2467 12597
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 2961 12631 3019 12637
rect 2961 12628 2973 12631
rect 2832 12600 2973 12628
rect 2832 12588 2838 12600
rect 2961 12597 2973 12600
rect 3007 12628 3019 12631
rect 3326 12628 3332 12640
rect 3007 12600 3332 12628
rect 3007 12597 3019 12600
rect 2961 12591 3019 12597
rect 3326 12588 3332 12600
rect 3384 12588 3390 12640
rect 7006 12628 7012 12640
rect 6967 12600 7012 12628
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 10686 12628 10692 12640
rect 10599 12600 10692 12628
rect 10686 12588 10692 12600
rect 10744 12628 10750 12640
rect 11330 12628 11336 12640
rect 10744 12600 11336 12628
rect 10744 12588 10750 12600
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 11698 12588 11704 12640
rect 11756 12628 11762 12640
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 11756 12600 12265 12628
rect 11756 12588 11762 12600
rect 12253 12597 12265 12600
rect 12299 12628 12311 12631
rect 12989 12631 13047 12637
rect 12989 12628 13001 12631
rect 12299 12600 13001 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 12989 12597 13001 12600
rect 13035 12597 13047 12631
rect 17218 12628 17224 12640
rect 17179 12600 17224 12628
rect 12989 12591 13047 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 19150 12588 19156 12640
rect 19208 12628 19214 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 19208 12600 21281 12628
rect 19208 12588 19214 12600
rect 21269 12597 21281 12600
rect 21315 12628 21327 12631
rect 21542 12628 21548 12640
rect 21315 12600 21548 12628
rect 21315 12597 21327 12600
rect 21269 12591 21327 12597
rect 21542 12588 21548 12600
rect 21600 12588 21606 12640
rect 22557 12631 22615 12637
rect 22557 12597 22569 12631
rect 22603 12628 22615 12631
rect 22738 12628 22744 12640
rect 22603 12600 22744 12628
rect 22603 12597 22615 12600
rect 22557 12591 22615 12597
rect 22738 12588 22744 12600
rect 22796 12588 22802 12640
rect 24489 12631 24547 12637
rect 24489 12597 24501 12631
rect 24535 12628 24547 12631
rect 24670 12628 24676 12640
rect 24535 12600 24676 12628
rect 24535 12597 24547 12600
rect 24489 12591 24547 12597
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2038 12384 2044 12436
rect 2096 12424 2102 12436
rect 2777 12427 2835 12433
rect 2777 12424 2789 12427
rect 2096 12396 2789 12424
rect 2096 12384 2102 12396
rect 2777 12393 2789 12396
rect 2823 12393 2835 12427
rect 2777 12387 2835 12393
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 4062 12424 4068 12436
rect 3927 12396 4068 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6454 12424 6460 12436
rect 6144 12396 6460 12424
rect 6144 12384 6150 12396
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 7009 12427 7067 12433
rect 7009 12424 7021 12427
rect 6696 12396 7021 12424
rect 6696 12384 6702 12396
rect 7009 12393 7021 12396
rect 7055 12424 7067 12427
rect 8294 12424 8300 12436
rect 7055 12396 7880 12424
rect 8255 12396 8300 12424
rect 7055 12393 7067 12396
rect 7009 12387 7067 12393
rect 4617 12359 4675 12365
rect 4617 12325 4629 12359
rect 4663 12356 4675 12359
rect 4798 12356 4804 12368
rect 4663 12328 4804 12356
rect 4663 12325 4675 12328
rect 4617 12319 4675 12325
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 6178 12356 6184 12368
rect 6139 12328 6184 12356
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 7098 12316 7104 12368
rect 7156 12356 7162 12368
rect 7282 12356 7288 12368
rect 7156 12328 7288 12356
rect 7156 12316 7162 12328
rect 7282 12316 7288 12328
rect 7340 12316 7346 12368
rect 7650 12316 7656 12368
rect 7708 12356 7714 12368
rect 7852 12365 7880 12396
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 9306 12424 9312 12436
rect 9267 12396 9312 12424
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 12897 12427 12955 12433
rect 12897 12424 12909 12427
rect 12860 12396 12909 12424
rect 12860 12384 12866 12396
rect 12897 12393 12909 12396
rect 12943 12393 12955 12427
rect 12897 12387 12955 12393
rect 13449 12427 13507 12433
rect 13449 12393 13461 12427
rect 13495 12424 13507 12427
rect 13538 12424 13544 12436
rect 13495 12396 13544 12424
rect 13495 12393 13507 12396
rect 13449 12387 13507 12393
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14366 12424 14372 12436
rect 14148 12396 14372 12424
rect 14148 12384 14154 12396
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 14734 12424 14740 12436
rect 14695 12396 14740 12424
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 16356 12396 16405 12424
rect 16356 12384 16362 12396
rect 16393 12393 16405 12396
rect 16439 12393 16451 12427
rect 18782 12424 18788 12436
rect 18743 12396 18788 12424
rect 16393 12387 16451 12393
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 19150 12424 19156 12436
rect 19111 12396 19156 12424
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 20254 12384 20260 12436
rect 20312 12424 20318 12436
rect 20530 12424 20536 12436
rect 20312 12396 20536 12424
rect 20312 12384 20318 12396
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 20622 12384 20628 12436
rect 20680 12384 20686 12436
rect 20990 12384 20996 12436
rect 21048 12424 21054 12436
rect 21453 12427 21511 12433
rect 21453 12424 21465 12427
rect 21048 12396 21465 12424
rect 21048 12384 21054 12396
rect 21453 12393 21465 12396
rect 21499 12424 21511 12427
rect 21634 12424 21640 12436
rect 21499 12396 21640 12424
rect 21499 12393 21511 12396
rect 21453 12387 21511 12393
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 22646 12384 22652 12436
rect 22704 12424 22710 12436
rect 22833 12427 22891 12433
rect 22704 12396 22784 12424
rect 22704 12384 22710 12396
rect 7745 12359 7803 12365
rect 7745 12356 7757 12359
rect 7708 12328 7757 12356
rect 7708 12316 7714 12328
rect 7745 12325 7757 12328
rect 7791 12325 7803 12359
rect 7745 12319 7803 12325
rect 7837 12359 7895 12365
rect 7837 12325 7849 12359
rect 7883 12356 7895 12359
rect 7926 12356 7932 12368
rect 7883 12328 7932 12356
rect 7883 12325 7895 12328
rect 7837 12319 7895 12325
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 9858 12316 9864 12368
rect 9916 12356 9922 12368
rect 9953 12359 10011 12365
rect 9953 12356 9965 12359
rect 9916 12328 9965 12356
rect 9916 12316 9922 12328
rect 9953 12325 9965 12328
rect 9999 12325 10011 12359
rect 9953 12319 10011 12325
rect 10689 12359 10747 12365
rect 10689 12325 10701 12359
rect 10735 12356 10747 12359
rect 11054 12356 11060 12368
rect 10735 12328 11060 12356
rect 10735 12325 10747 12328
rect 10689 12319 10747 12325
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 14185 12359 14243 12365
rect 14185 12325 14197 12359
rect 14231 12356 14243 12359
rect 14274 12356 14280 12368
rect 14231 12328 14280 12356
rect 14231 12325 14243 12328
rect 14185 12319 14243 12325
rect 14274 12316 14280 12328
rect 14332 12356 14338 12368
rect 14458 12356 14464 12368
rect 14332 12328 14464 12356
rect 14332 12316 14338 12328
rect 14458 12316 14464 12328
rect 14516 12316 14522 12368
rect 17028 12359 17086 12365
rect 17028 12325 17040 12359
rect 17074 12356 17086 12359
rect 17678 12356 17684 12368
rect 17074 12328 17684 12356
rect 17074 12325 17086 12328
rect 17028 12319 17086 12325
rect 17678 12316 17684 12328
rect 17736 12316 17742 12368
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 19797 12359 19855 12365
rect 19797 12356 19809 12359
rect 19392 12328 19809 12356
rect 19392 12316 19398 12328
rect 19797 12325 19809 12328
rect 19843 12356 19855 12359
rect 20441 12359 20499 12365
rect 20441 12356 20453 12359
rect 19843 12328 20453 12356
rect 19843 12325 19855 12328
rect 19797 12319 19855 12325
rect 20441 12325 20453 12328
rect 20487 12325 20499 12359
rect 20441 12319 20499 12325
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 1664 12291 1722 12297
rect 1664 12257 1676 12291
rect 1710 12288 1722 12291
rect 4433 12291 4491 12297
rect 1710 12260 2452 12288
rect 1710 12257 1722 12260
rect 1664 12251 1722 12257
rect 2424 12220 2452 12260
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 4982 12288 4988 12300
rect 4479 12260 4988 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 5537 12291 5595 12297
rect 5537 12257 5549 12291
rect 5583 12288 5595 12291
rect 5994 12288 6000 12300
rect 5583 12260 6000 12288
rect 5583 12257 5595 12260
rect 5537 12251 5595 12257
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 9674 12288 9680 12300
rect 9587 12260 9680 12288
rect 9674 12248 9680 12260
rect 9732 12288 9738 12300
rect 10870 12288 10876 12300
rect 9732 12260 10876 12288
rect 9732 12248 9738 12260
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 11238 12297 11244 12300
rect 11232 12288 11244 12297
rect 11199 12260 11244 12288
rect 11232 12251 11244 12260
rect 11238 12248 11244 12251
rect 11296 12248 11302 12300
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 15013 12291 15071 12297
rect 15013 12288 15025 12291
rect 13872 12260 15025 12288
rect 13872 12248 13878 12260
rect 15013 12257 15025 12260
rect 15059 12288 15071 12291
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 15059 12260 15301 12288
rect 15059 12257 15071 12260
rect 15013 12251 15071 12257
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 16761 12291 16819 12297
rect 16761 12257 16773 12291
rect 16807 12288 16819 12291
rect 17310 12288 17316 12300
rect 16807 12260 17316 12288
rect 16807 12257 16819 12260
rect 16761 12251 16819 12257
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 18966 12248 18972 12300
rect 19024 12288 19030 12300
rect 19889 12291 19947 12297
rect 19889 12288 19901 12291
rect 19024 12260 19901 12288
rect 19024 12248 19030 12260
rect 19889 12257 19901 12260
rect 19935 12288 19947 12291
rect 20640 12288 20668 12384
rect 21542 12356 21548 12368
rect 21503 12328 21548 12356
rect 21542 12316 21548 12328
rect 21600 12316 21606 12368
rect 21266 12288 21272 12300
rect 19935 12260 20668 12288
rect 21227 12260 21272 12288
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 21266 12248 21272 12260
rect 21324 12248 21330 12300
rect 2498 12220 2504 12232
rect 2411 12192 2504 12220
rect 2498 12180 2504 12192
rect 2556 12220 2562 12232
rect 4706 12220 4712 12232
rect 2556 12192 3464 12220
rect 4667 12192 4712 12220
rect 2556 12180 2562 12192
rect 3436 12096 3464 12192
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 4890 12180 4896 12232
rect 4948 12220 4954 12232
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 4948 12192 5181 12220
rect 4948 12180 4954 12192
rect 5169 12189 5181 12192
rect 5215 12220 5227 12223
rect 6178 12220 6184 12232
rect 5215 12192 6184 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 6178 12180 6184 12192
rect 6236 12220 6242 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 6236 12192 6285 12220
rect 6236 12180 6242 12192
rect 6273 12189 6285 12192
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 7374 12180 7380 12232
rect 7432 12220 7438 12232
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 7432 12192 7757 12220
rect 7432 12180 7438 12192
rect 7745 12189 7757 12192
rect 7791 12220 7803 12223
rect 8386 12220 8392 12232
rect 7791 12192 8392 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 10962 12220 10968 12232
rect 10923 12192 10968 12220
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 14090 12220 14096 12232
rect 14051 12192 14096 12220
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14274 12220 14280 12232
rect 14235 12192 14280 12220
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 15565 12223 15623 12229
rect 15565 12189 15577 12223
rect 15611 12220 15623 12223
rect 15930 12220 15936 12232
rect 15611 12192 15936 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 19426 12180 19432 12232
rect 19484 12220 19490 12232
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 19484 12192 19809 12220
rect 19484 12180 19490 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 3510 12112 3516 12164
rect 3568 12152 3574 12164
rect 4157 12155 4215 12161
rect 4157 12152 4169 12155
rect 3568 12124 4169 12152
rect 3568 12112 3574 12124
rect 4157 12121 4169 12124
rect 4203 12152 4215 12155
rect 5534 12152 5540 12164
rect 4203 12124 5540 12152
rect 4203 12121 4215 12124
rect 4157 12115 4215 12121
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 5721 12155 5779 12161
rect 5721 12121 5733 12155
rect 5767 12152 5779 12155
rect 5767 12124 6776 12152
rect 5767 12121 5779 12124
rect 5721 12115 5779 12121
rect 937 12087 995 12093
rect 937 12053 949 12087
rect 983 12084 995 12087
rect 1578 12084 1584 12096
rect 983 12056 1584 12084
rect 983 12053 995 12056
rect 937 12047 995 12053
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 3418 12084 3424 12096
rect 3379 12056 3424 12084
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 6638 12084 6644 12096
rect 6599 12056 6644 12084
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 6748 12084 6776 12124
rect 7190 12112 7196 12164
rect 7248 12152 7254 12164
rect 7285 12155 7343 12161
rect 7285 12152 7297 12155
rect 7248 12124 7297 12152
rect 7248 12112 7254 12124
rect 7285 12121 7297 12124
rect 7331 12121 7343 12155
rect 8570 12152 8576 12164
rect 8531 12124 8576 12152
rect 7285 12115 7343 12121
rect 8570 12112 8576 12124
rect 8628 12112 8634 12164
rect 10134 12112 10140 12164
rect 10192 12152 10198 12164
rect 10689 12155 10747 12161
rect 10689 12152 10701 12155
rect 10192 12124 10701 12152
rect 10192 12112 10198 12124
rect 10689 12121 10701 12124
rect 10735 12152 10747 12155
rect 10781 12155 10839 12161
rect 10781 12152 10793 12155
rect 10735 12124 10793 12152
rect 10735 12121 10747 12124
rect 10689 12115 10747 12121
rect 10781 12121 10793 12124
rect 10827 12121 10839 12155
rect 13722 12152 13728 12164
rect 13683 12124 13728 12152
rect 10781 12115 10839 12121
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 19812 12152 19840 12183
rect 20162 12180 20168 12232
rect 20220 12220 20226 12232
rect 20530 12220 20536 12232
rect 20220 12192 20536 12220
rect 20220 12180 20226 12192
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 21560 12220 21588 12316
rect 22278 12248 22284 12300
rect 22336 12288 22342 12300
rect 22646 12288 22652 12300
rect 22336 12260 22652 12288
rect 22336 12248 22342 12260
rect 22646 12248 22652 12260
rect 22704 12248 22710 12300
rect 22094 12220 22100 12232
rect 21560 12192 22100 12220
rect 22094 12180 22100 12192
rect 22152 12180 22158 12232
rect 22756 12220 22784 12396
rect 22833 12393 22845 12427
rect 22879 12424 22891 12427
rect 23014 12424 23020 12436
rect 22879 12396 23020 12424
rect 22879 12393 22891 12396
rect 22833 12387 22891 12393
rect 23014 12384 23020 12396
rect 23072 12384 23078 12436
rect 24486 12424 24492 12436
rect 24447 12396 24492 12424
rect 24486 12384 24492 12396
rect 24544 12384 24550 12436
rect 23842 12316 23848 12368
rect 23900 12356 23906 12368
rect 23937 12359 23995 12365
rect 23937 12356 23949 12359
rect 23900 12328 23949 12356
rect 23900 12316 23906 12328
rect 23937 12325 23949 12328
rect 23983 12325 23995 12359
rect 25222 12356 25228 12368
rect 25183 12328 25228 12356
rect 23937 12319 23995 12325
rect 25222 12316 25228 12328
rect 25280 12316 25286 12368
rect 23106 12248 23112 12300
rect 23164 12288 23170 12300
rect 23293 12291 23351 12297
rect 23293 12288 23305 12291
rect 23164 12260 23305 12288
rect 23164 12248 23170 12260
rect 23293 12257 23305 12260
rect 23339 12288 23351 12291
rect 24949 12291 25007 12297
rect 23339 12260 24072 12288
rect 23339 12257 23351 12260
rect 23293 12251 23351 12257
rect 22388 12192 22784 12220
rect 20254 12152 20260 12164
rect 19812 12124 20260 12152
rect 20254 12112 20260 12124
rect 20312 12112 20318 12164
rect 20441 12155 20499 12161
rect 20441 12121 20453 12155
rect 20487 12152 20499 12155
rect 20993 12155 21051 12161
rect 20993 12152 21005 12155
rect 20487 12124 21005 12152
rect 20487 12121 20499 12124
rect 20441 12115 20499 12121
rect 20993 12121 21005 12124
rect 21039 12121 21051 12155
rect 20993 12115 21051 12121
rect 22005 12155 22063 12161
rect 22005 12121 22017 12155
rect 22051 12152 22063 12155
rect 22388 12152 22416 12192
rect 23566 12180 23572 12232
rect 23624 12220 23630 12232
rect 24044 12229 24072 12260
rect 24949 12257 24961 12291
rect 24995 12288 25007 12291
rect 25038 12288 25044 12300
rect 24995 12260 25044 12288
rect 24995 12257 25007 12260
rect 24949 12251 25007 12257
rect 25038 12248 25044 12260
rect 25096 12288 25102 12300
rect 25314 12288 25320 12300
rect 25096 12260 25320 12288
rect 25096 12248 25102 12260
rect 25314 12248 25320 12260
rect 25372 12248 25378 12300
rect 23845 12223 23903 12229
rect 23845 12220 23857 12223
rect 23624 12192 23857 12220
rect 23624 12180 23630 12192
rect 23845 12189 23857 12192
rect 23891 12189 23903 12223
rect 23845 12183 23903 12189
rect 24029 12223 24087 12229
rect 24029 12189 24041 12223
rect 24075 12220 24087 12223
rect 24854 12220 24860 12232
rect 24075 12192 24860 12220
rect 24075 12189 24087 12192
rect 24029 12183 24087 12189
rect 24854 12180 24860 12192
rect 24912 12180 24918 12232
rect 22051 12124 22416 12152
rect 22051 12121 22063 12124
rect 22005 12115 22063 12121
rect 22388 12096 22416 12124
rect 23382 12112 23388 12164
rect 23440 12152 23446 12164
rect 23477 12155 23535 12161
rect 23477 12152 23489 12155
rect 23440 12124 23489 12152
rect 23440 12112 23446 12124
rect 23477 12121 23489 12124
rect 23523 12121 23535 12155
rect 23477 12115 23535 12121
rect 7006 12084 7012 12096
rect 6748 12056 7012 12084
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8720 12056 8953 12084
rect 8720 12044 8726 12056
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 8941 12047 8999 12053
rect 9490 12044 9496 12096
rect 9548 12084 9554 12096
rect 10413 12087 10471 12093
rect 10413 12084 10425 12087
rect 9548 12056 10425 12084
rect 9548 12044 9554 12056
rect 10413 12053 10425 12056
rect 10459 12053 10471 12087
rect 10413 12047 10471 12053
rect 12250 12044 12256 12096
rect 12308 12084 12314 12096
rect 12345 12087 12403 12093
rect 12345 12084 12357 12087
rect 12308 12056 12357 12084
rect 12308 12044 12314 12056
rect 12345 12053 12357 12056
rect 12391 12053 12403 12087
rect 12345 12047 12403 12053
rect 15838 12044 15844 12096
rect 15896 12084 15902 12096
rect 16025 12087 16083 12093
rect 16025 12084 16037 12087
rect 15896 12056 16037 12084
rect 15896 12044 15902 12056
rect 16025 12053 16037 12056
rect 16071 12053 16083 12087
rect 18138 12084 18144 12096
rect 18099 12056 18144 12084
rect 16025 12047 16083 12053
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 19337 12087 19395 12093
rect 19337 12053 19349 12087
rect 19383 12084 19395 12087
rect 20162 12084 20168 12096
rect 19383 12056 20168 12084
rect 19383 12053 19395 12056
rect 19337 12047 19395 12053
rect 20162 12044 20168 12056
rect 20220 12044 20226 12096
rect 20346 12084 20352 12096
rect 20307 12056 20352 12084
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 20714 12084 20720 12096
rect 20675 12056 20720 12084
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 22278 12084 22284 12096
rect 22239 12056 22284 12084
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 22370 12044 22376 12096
rect 22428 12044 22434 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 1452 11852 1593 11880
rect 1452 11840 1458 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 1581 11843 1639 11849
rect 1596 11608 1624 11843
rect 1670 11840 1676 11892
rect 1728 11880 1734 11892
rect 2222 11880 2228 11892
rect 1728 11852 2228 11880
rect 1728 11840 1734 11852
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 3142 11880 3148 11892
rect 3103 11852 3148 11880
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 3237 11883 3295 11889
rect 3237 11849 3249 11883
rect 3283 11880 3295 11883
rect 3513 11883 3571 11889
rect 3513 11880 3525 11883
rect 3283 11852 3525 11880
rect 3283 11849 3295 11852
rect 3237 11843 3295 11849
rect 3513 11849 3525 11852
rect 3559 11880 3571 11883
rect 4982 11880 4988 11892
rect 3559 11852 4988 11880
rect 3559 11849 3571 11852
rect 3513 11843 3571 11849
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 7377 11883 7435 11889
rect 7377 11849 7389 11883
rect 7423 11880 7435 11883
rect 7558 11880 7564 11892
rect 7423 11852 7564 11880
rect 7423 11849 7435 11852
rect 7377 11843 7435 11849
rect 7558 11840 7564 11852
rect 7616 11880 7622 11892
rect 8662 11880 8668 11892
rect 7616 11852 8668 11880
rect 7616 11840 7622 11852
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 10870 11880 10876 11892
rect 10831 11852 10876 11880
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11296 11852 11805 11880
rect 11296 11840 11302 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 12897 11883 12955 11889
rect 12897 11849 12909 11883
rect 12943 11880 12955 11883
rect 14274 11880 14280 11892
rect 12943 11852 14280 11880
rect 12943 11849 12955 11852
rect 12897 11843 12955 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 14737 11883 14795 11889
rect 14737 11849 14749 11883
rect 14783 11880 14795 11883
rect 14826 11880 14832 11892
rect 14783 11852 14832 11880
rect 14783 11849 14795 11852
rect 14737 11843 14795 11849
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 15657 11883 15715 11889
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 16206 11880 16212 11892
rect 15703 11852 16212 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 17678 11840 17684 11892
rect 17736 11880 17742 11892
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 17736 11852 17785 11880
rect 17736 11840 17742 11852
rect 17773 11849 17785 11852
rect 17819 11849 17831 11883
rect 18966 11880 18972 11892
rect 18927 11852 18972 11880
rect 17773 11843 17831 11849
rect 18966 11840 18972 11852
rect 19024 11840 19030 11892
rect 19978 11880 19984 11892
rect 19812 11852 19984 11880
rect 1857 11815 1915 11821
rect 1857 11781 1869 11815
rect 1903 11812 1915 11815
rect 2406 11812 2412 11824
rect 1903 11784 2412 11812
rect 1903 11781 1915 11784
rect 1857 11775 1915 11781
rect 2406 11772 2412 11784
rect 2464 11772 2470 11824
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 1872 11716 2237 11744
rect 1872 11688 1900 11716
rect 2225 11713 2237 11716
rect 2271 11713 2283 11747
rect 3160 11744 3188 11840
rect 8018 11812 8024 11824
rect 7760 11784 8024 11812
rect 3160 11716 4108 11744
rect 2225 11707 2283 11713
rect 1854 11636 1860 11688
rect 1912 11636 1918 11688
rect 3973 11679 4031 11685
rect 3973 11676 3985 11679
rect 2148 11648 3985 11676
rect 2148 11608 2176 11648
rect 2314 11608 2320 11620
rect 1596 11580 2176 11608
rect 2275 11580 2320 11608
rect 1872 11552 1900 11580
rect 2314 11568 2320 11580
rect 2372 11568 2378 11620
rect 2409 11611 2467 11617
rect 2409 11577 2421 11611
rect 2455 11577 2467 11611
rect 2409 11571 2467 11577
rect 1854 11500 1860 11552
rect 1912 11500 1918 11552
rect 1946 11500 1952 11552
rect 2004 11540 2010 11552
rect 2424 11540 2452 11571
rect 2004 11512 2452 11540
rect 2004 11500 2010 11512
rect 2682 11500 2688 11552
rect 2740 11540 2746 11552
rect 3237 11543 3295 11549
rect 3237 11540 3249 11543
rect 2740 11512 3249 11540
rect 2740 11500 2746 11512
rect 3237 11509 3249 11512
rect 3283 11509 3295 11543
rect 3712 11540 3740 11648
rect 3973 11645 3985 11648
rect 4019 11645 4031 11679
rect 4080 11676 4108 11716
rect 4982 11704 4988 11756
rect 5040 11744 5046 11756
rect 7374 11744 7380 11756
rect 5040 11716 7380 11744
rect 5040 11704 5046 11716
rect 7374 11704 7380 11716
rect 7432 11744 7438 11756
rect 7760 11753 7788 11784
rect 8018 11772 8024 11784
rect 8076 11772 8082 11824
rect 8110 11772 8116 11824
rect 8168 11812 8174 11824
rect 8941 11815 8999 11821
rect 8941 11812 8953 11815
rect 8168 11784 8953 11812
rect 8168 11772 8174 11784
rect 8941 11781 8953 11784
rect 8987 11781 8999 11815
rect 8941 11775 8999 11781
rect 16485 11815 16543 11821
rect 16485 11781 16497 11815
rect 16531 11812 16543 11815
rect 16574 11812 16580 11824
rect 16531 11784 16580 11812
rect 16531 11781 16543 11784
rect 16485 11775 16543 11781
rect 16574 11772 16580 11784
rect 16632 11772 16638 11824
rect 7745 11747 7803 11753
rect 7745 11744 7757 11747
rect 7432 11716 7757 11744
rect 7432 11704 7438 11716
rect 7745 11713 7757 11716
rect 7791 11713 7803 11747
rect 7926 11744 7932 11756
rect 7887 11716 7932 11744
rect 7745 11707 7803 11713
rect 7926 11704 7932 11716
rect 7984 11704 7990 11756
rect 9306 11744 9312 11756
rect 9267 11716 9312 11744
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 9490 11744 9496 11756
rect 9451 11716 9496 11744
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 11333 11747 11391 11753
rect 11333 11744 11345 11747
rect 9999 11716 11345 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 11333 11713 11345 11716
rect 11379 11744 11391 11747
rect 12342 11744 12348 11756
rect 11379 11716 12348 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 16390 11704 16396 11756
rect 16448 11744 16454 11756
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 16448 11716 16957 11744
rect 16448 11704 16454 11716
rect 16945 11713 16957 11716
rect 16991 11744 17003 11747
rect 17954 11744 17960 11756
rect 16991 11716 17960 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 4229 11679 4287 11685
rect 4229 11676 4241 11679
rect 4080 11648 4241 11676
rect 3973 11639 4031 11645
rect 4229 11645 4241 11648
rect 4275 11676 4287 11679
rect 4706 11676 4712 11688
rect 4275 11648 4712 11676
rect 4275 11645 4287 11648
rect 4229 11639 4287 11645
rect 4706 11636 4712 11648
rect 4764 11636 4770 11688
rect 7193 11679 7251 11685
rect 7193 11645 7205 11679
rect 7239 11676 7251 11679
rect 8386 11676 8392 11688
rect 7239 11648 7880 11676
rect 8347 11648 8392 11676
rect 7239 11645 7251 11648
rect 7193 11639 7251 11645
rect 7852 11620 7880 11648
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 9508 11676 9536 11704
rect 8803 11648 9536 11676
rect 13357 11679 13415 11685
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 13357 11645 13369 11679
rect 13403 11676 13415 11679
rect 13446 11676 13452 11688
rect 13403 11648 13452 11676
rect 13403 11645 13415 11648
rect 13357 11639 13415 11645
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 13630 11685 13636 11688
rect 13624 11676 13636 11685
rect 13591 11648 13636 11676
rect 13624 11639 13636 11648
rect 13630 11636 13636 11639
rect 13688 11636 13694 11688
rect 18046 11676 18052 11688
rect 18007 11648 18052 11676
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 18966 11636 18972 11688
rect 19024 11676 19030 11688
rect 19812 11685 19840 11852
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 21177 11883 21235 11889
rect 21177 11880 21189 11883
rect 20772 11852 21189 11880
rect 20772 11840 20778 11852
rect 21177 11849 21189 11852
rect 21223 11849 21235 11883
rect 21177 11843 21235 11849
rect 21266 11840 21272 11892
rect 21324 11880 21330 11892
rect 21729 11883 21787 11889
rect 21729 11880 21741 11883
rect 21324 11852 21741 11880
rect 21324 11840 21330 11852
rect 21729 11849 21741 11852
rect 21775 11849 21787 11883
rect 21729 11843 21787 11849
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 24762 11880 24768 11892
rect 22152 11852 22197 11880
rect 24723 11852 24768 11880
rect 22152 11840 22158 11852
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 25406 11880 25412 11892
rect 25367 11852 25412 11880
rect 25406 11840 25412 11852
rect 25464 11840 25470 11892
rect 23382 11772 23388 11824
rect 23440 11812 23446 11824
rect 23753 11815 23811 11821
rect 23753 11812 23765 11815
rect 23440 11784 23765 11812
rect 23440 11772 23446 11784
rect 23753 11781 23765 11784
rect 23799 11781 23811 11815
rect 23753 11775 23811 11781
rect 23842 11772 23848 11824
rect 23900 11812 23906 11824
rect 25133 11815 25191 11821
rect 25133 11812 25145 11815
rect 23900 11784 25145 11812
rect 23900 11772 23906 11784
rect 25133 11781 25145 11784
rect 25179 11812 25191 11815
rect 25590 11812 25596 11824
rect 25179 11784 25596 11812
rect 25179 11781 25191 11784
rect 25133 11775 25191 11781
rect 25590 11772 25596 11784
rect 25648 11772 25654 11824
rect 24118 11704 24124 11756
rect 24176 11744 24182 11756
rect 24305 11747 24363 11753
rect 24305 11744 24317 11747
rect 24176 11716 24317 11744
rect 24176 11704 24182 11716
rect 24305 11713 24317 11716
rect 24351 11713 24363 11747
rect 24305 11707 24363 11713
rect 19613 11679 19671 11685
rect 19613 11676 19625 11679
rect 19024 11648 19625 11676
rect 19024 11636 19030 11648
rect 19613 11645 19625 11648
rect 19659 11676 19671 11679
rect 19797 11679 19855 11685
rect 19797 11676 19809 11679
rect 19659 11648 19809 11676
rect 19659 11645 19671 11648
rect 19613 11639 19671 11645
rect 19797 11645 19809 11648
rect 19843 11645 19855 11679
rect 22278 11676 22284 11688
rect 22239 11648 22284 11676
rect 19797 11639 19855 11645
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 23477 11679 23535 11685
rect 23477 11645 23489 11679
rect 23523 11676 23535 11679
rect 23566 11676 23572 11688
rect 23523 11648 23572 11676
rect 23523 11645 23535 11648
rect 23477 11639 23535 11645
rect 23566 11636 23572 11648
rect 23624 11636 23630 11688
rect 25222 11676 25228 11688
rect 25183 11648 25228 11676
rect 25222 11636 25228 11648
rect 25280 11676 25286 11688
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 25280 11648 25789 11676
rect 25280 11636 25286 11648
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 3878 11608 3884 11620
rect 3791 11580 3884 11608
rect 3878 11568 3884 11580
rect 3936 11608 3942 11620
rect 4798 11608 4804 11620
rect 3936 11580 4804 11608
rect 3936 11568 3942 11580
rect 4798 11568 4804 11580
rect 4856 11568 4862 11620
rect 5810 11568 5816 11620
rect 5868 11608 5874 11620
rect 6549 11611 6607 11617
rect 6549 11608 6561 11611
rect 5868 11580 6561 11608
rect 5868 11568 5874 11580
rect 6549 11577 6561 11580
rect 6595 11608 6607 11611
rect 7650 11608 7656 11620
rect 6595 11580 7656 11608
rect 6595 11577 6607 11580
rect 6549 11571 6607 11577
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 7834 11608 7840 11620
rect 7795 11580 7840 11608
rect 7834 11568 7840 11580
rect 7892 11568 7898 11620
rect 10689 11611 10747 11617
rect 10689 11577 10701 11611
rect 10735 11608 10747 11611
rect 11425 11611 11483 11617
rect 11425 11608 11437 11611
rect 10735 11580 11437 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 11425 11577 11437 11580
rect 11471 11608 11483 11611
rect 13262 11608 13268 11620
rect 11471 11580 12848 11608
rect 13175 11580 13268 11608
rect 11471 11577 11483 11580
rect 11425 11571 11483 11577
rect 4246 11540 4252 11552
rect 3712 11512 4252 11540
rect 3237 11503 3295 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 5350 11540 5356 11552
rect 5311 11512 5356 11540
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 5902 11540 5908 11552
rect 5863 11512 5908 11540
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 6822 11540 6828 11552
rect 6696 11512 6828 11540
rect 6696 11500 6702 11512
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 9398 11540 9404 11552
rect 9359 11512 9404 11540
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 10321 11543 10379 11549
rect 10321 11509 10333 11543
rect 10367 11540 10379 11543
rect 10870 11540 10876 11552
rect 10367 11512 10876 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 10870 11500 10876 11512
rect 10928 11540 10934 11552
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 10928 11512 11345 11540
rect 10928 11500 10934 11512
rect 11333 11509 11345 11512
rect 11379 11509 11391 11543
rect 12250 11540 12256 11552
rect 12211 11512 12256 11540
rect 11333 11503 11391 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 12820 11540 12848 11580
rect 13262 11568 13268 11580
rect 13320 11608 13326 11620
rect 14090 11608 14096 11620
rect 13320 11580 14096 11608
rect 13320 11568 13326 11580
rect 14090 11568 14096 11580
rect 14148 11568 14154 11620
rect 16301 11611 16359 11617
rect 16301 11577 16313 11611
rect 16347 11608 16359 11611
rect 17037 11611 17095 11617
rect 17037 11608 17049 11611
rect 16347 11580 17049 11608
rect 16347 11577 16359 11580
rect 16301 11571 16359 11577
rect 17037 11577 17049 11580
rect 17083 11608 17095 11611
rect 18138 11608 18144 11620
rect 17083 11580 18144 11608
rect 17083 11577 17095 11580
rect 17037 11571 17095 11577
rect 18138 11568 18144 11580
rect 18196 11568 18202 11620
rect 20042 11611 20100 11617
rect 20042 11608 20054 11611
rect 19444 11580 20054 11608
rect 19444 11552 19472 11580
rect 20042 11577 20054 11580
rect 20088 11577 20100 11611
rect 23106 11608 23112 11620
rect 23019 11580 23112 11608
rect 20042 11571 20100 11577
rect 23106 11568 23112 11580
rect 23164 11608 23170 11620
rect 24029 11611 24087 11617
rect 24029 11608 24041 11611
rect 23164 11580 24041 11608
rect 23164 11568 23170 11580
rect 24029 11577 24041 11580
rect 24075 11577 24087 11611
rect 24029 11571 24087 11577
rect 14826 11540 14832 11552
rect 12820 11512 14832 11540
rect 14826 11500 14832 11512
rect 14884 11500 14890 11552
rect 16942 11540 16948 11552
rect 16903 11512 16948 11540
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 17497 11543 17555 11549
rect 17497 11540 17509 11543
rect 17276 11512 17509 11540
rect 17276 11500 17282 11512
rect 17497 11509 17509 11512
rect 17543 11540 17555 11543
rect 17770 11540 17776 11552
rect 17543 11512 17776 11540
rect 17543 11509 17555 11512
rect 17497 11503 17555 11509
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 18233 11543 18291 11549
rect 18233 11509 18245 11543
rect 18279 11540 18291 11543
rect 18414 11540 18420 11552
rect 18279 11512 18420 11540
rect 18279 11509 18291 11512
rect 18233 11503 18291 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 19337 11543 19395 11549
rect 19337 11509 19349 11543
rect 19383 11540 19395 11543
rect 19426 11540 19432 11552
rect 19383 11512 19432 11540
rect 19383 11509 19395 11512
rect 19337 11503 19395 11509
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 22462 11540 22468 11552
rect 22423 11512 22468 11540
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 24213 11543 24271 11549
rect 24213 11509 24225 11543
rect 24259 11540 24271 11543
rect 24762 11540 24768 11552
rect 24259 11512 24768 11540
rect 24259 11509 24271 11512
rect 24213 11503 24271 11509
rect 24762 11500 24768 11512
rect 24820 11500 24826 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1946 11336 1952 11348
rect 1907 11308 1952 11336
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 3513 11339 3571 11345
rect 3513 11336 3525 11339
rect 3476 11308 3525 11336
rect 3476 11296 3482 11308
rect 3513 11305 3525 11308
rect 3559 11336 3571 11339
rect 5350 11336 5356 11348
rect 3559 11308 5356 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 7009 11339 7067 11345
rect 7009 11336 7021 11339
rect 6880 11308 7021 11336
rect 6880 11296 6886 11308
rect 7009 11305 7021 11308
rect 7055 11336 7067 11339
rect 7926 11336 7932 11348
rect 7055 11308 7932 11336
rect 7055 11305 7067 11308
rect 7009 11299 7067 11305
rect 7926 11296 7932 11308
rect 7984 11336 7990 11348
rect 7984 11308 8156 11336
rect 7984 11296 7990 11308
rect 2961 11271 3019 11277
rect 2961 11237 2973 11271
rect 3007 11268 3019 11271
rect 3789 11271 3847 11277
rect 3789 11268 3801 11271
rect 3007 11240 3801 11268
rect 3007 11237 3019 11240
rect 2961 11231 3019 11237
rect 3789 11237 3801 11240
rect 3835 11268 3847 11271
rect 3970 11268 3976 11280
rect 3835 11240 3976 11268
rect 3835 11237 3847 11240
rect 3789 11231 3847 11237
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 4246 11268 4252 11280
rect 4207 11240 4252 11268
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 4706 11268 4712 11280
rect 4667 11240 4712 11268
rect 4706 11228 4712 11240
rect 4764 11228 4770 11280
rect 5252 11271 5310 11277
rect 5252 11237 5264 11271
rect 5298 11268 5310 11271
rect 5442 11268 5448 11280
rect 5298 11240 5448 11268
rect 5298 11237 5310 11240
rect 5252 11231 5310 11237
rect 5442 11228 5448 11240
rect 5500 11228 5506 11280
rect 7374 11268 7380 11280
rect 7335 11240 7380 11268
rect 7374 11228 7380 11240
rect 7432 11228 7438 11280
rect 8128 11277 8156 11308
rect 8294 11296 8300 11348
rect 8352 11336 8358 11348
rect 8849 11339 8907 11345
rect 8849 11336 8861 11339
rect 8352 11308 8861 11336
rect 8352 11296 8358 11308
rect 8849 11305 8861 11308
rect 8895 11336 8907 11339
rect 9398 11336 9404 11348
rect 8895 11308 9404 11336
rect 8895 11305 8907 11308
rect 8849 11299 8907 11305
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 11422 11336 11428 11348
rect 11335 11308 11428 11336
rect 11422 11296 11428 11308
rect 11480 11336 11486 11348
rect 12250 11336 12256 11348
rect 11480 11308 12256 11336
rect 11480 11296 11486 11308
rect 12250 11296 12256 11308
rect 12308 11336 12314 11348
rect 13173 11339 13231 11345
rect 13173 11336 13185 11339
rect 12308 11308 13185 11336
rect 12308 11296 12314 11308
rect 13173 11305 13185 11308
rect 13219 11336 13231 11339
rect 13630 11336 13636 11348
rect 13219 11308 13636 11336
rect 13219 11305 13231 11308
rect 13173 11299 13231 11305
rect 13630 11296 13636 11308
rect 13688 11336 13694 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 13688 11308 14105 11336
rect 13688 11296 13694 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14093 11299 14151 11305
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 17129 11339 17187 11345
rect 17129 11336 17141 11339
rect 16724 11308 17141 11336
rect 16724 11296 16730 11308
rect 17129 11305 17141 11308
rect 17175 11336 17187 11339
rect 17310 11336 17316 11348
rect 17175 11308 17316 11336
rect 17175 11305 17187 11308
rect 17129 11299 17187 11305
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 17954 11336 17960 11348
rect 17915 11308 17960 11336
rect 17954 11296 17960 11308
rect 18012 11296 18018 11348
rect 18138 11296 18144 11348
rect 18196 11336 18202 11348
rect 18877 11339 18935 11345
rect 18877 11336 18889 11339
rect 18196 11308 18889 11336
rect 18196 11296 18202 11308
rect 18877 11305 18889 11308
rect 18923 11305 18935 11339
rect 19334 11336 19340 11348
rect 19295 11308 19340 11336
rect 18877 11299 18935 11305
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 20254 11336 20260 11348
rect 20215 11308 20260 11336
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 20714 11336 20720 11348
rect 20675 11308 20720 11336
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 21634 11336 21640 11348
rect 21595 11308 21640 11336
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 24118 11296 24124 11348
rect 24176 11336 24182 11348
rect 24673 11339 24731 11345
rect 24673 11336 24685 11339
rect 24176 11308 24685 11336
rect 24176 11296 24182 11308
rect 24673 11305 24685 11308
rect 24719 11305 24731 11339
rect 25038 11336 25044 11348
rect 24999 11308 25044 11336
rect 24673 11299 24731 11305
rect 25038 11296 25044 11308
rect 25096 11296 25102 11348
rect 25406 11336 25412 11348
rect 25367 11308 25412 11336
rect 25406 11296 25412 11308
rect 25464 11296 25470 11348
rect 8021 11271 8079 11277
rect 8021 11268 8033 11271
rect 7944 11240 8033 11268
rect 2317 11203 2375 11209
rect 2317 11169 2329 11203
rect 2363 11200 2375 11203
rect 3053 11203 3111 11209
rect 3053 11200 3065 11203
rect 2363 11172 3065 11200
rect 2363 11169 2375 11172
rect 2317 11163 2375 11169
rect 3053 11169 3065 11172
rect 3099 11200 3111 11203
rect 3418 11200 3424 11212
rect 3099 11172 3424 11200
rect 3099 11169 3111 11172
rect 3053 11163 3111 11169
rect 3418 11160 3424 11172
rect 3476 11160 3482 11212
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3510 11132 3516 11144
rect 3007 11104 3516 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 4264 11132 4292 11228
rect 4724 11200 4752 11228
rect 7944 11212 7972 11240
rect 8021 11237 8033 11240
rect 8067 11237 8079 11271
rect 8021 11231 8079 11237
rect 8113 11271 8171 11277
rect 8113 11237 8125 11271
rect 8159 11237 8171 11271
rect 8113 11231 8171 11237
rect 9306 11228 9312 11280
rect 9364 11268 9370 11280
rect 10229 11271 10287 11277
rect 10229 11268 10241 11271
rect 9364 11240 10241 11268
rect 9364 11228 9370 11240
rect 10229 11237 10241 11240
rect 10275 11237 10287 11271
rect 10229 11231 10287 11237
rect 10778 11228 10784 11280
rect 10836 11268 10842 11280
rect 13722 11268 13728 11280
rect 10836 11240 13728 11268
rect 10836 11228 10842 11240
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 15562 11268 15568 11280
rect 15523 11240 15568 11268
rect 15562 11228 15568 11240
rect 15620 11228 15626 11280
rect 16209 11271 16267 11277
rect 16209 11237 16221 11271
rect 16255 11268 16267 11271
rect 16482 11268 16488 11280
rect 16255 11240 16488 11268
rect 16255 11237 16267 11240
rect 16209 11231 16267 11237
rect 16482 11228 16488 11240
rect 16540 11268 16546 11280
rect 17221 11271 17279 11277
rect 17221 11268 17233 11271
rect 16540 11240 17233 11268
rect 16540 11228 16546 11240
rect 17221 11237 17233 11240
rect 17267 11268 17279 11271
rect 17678 11268 17684 11280
rect 17267 11240 17684 11268
rect 17267 11237 17279 11240
rect 17221 11231 17279 11237
rect 17678 11228 17684 11240
rect 17736 11228 17742 11280
rect 18506 11228 18512 11280
rect 18564 11268 18570 11280
rect 19978 11268 19984 11280
rect 18564 11240 19984 11268
rect 18564 11228 18570 11240
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 20346 11228 20352 11280
rect 20404 11268 20410 11280
rect 21177 11271 21235 11277
rect 21177 11268 21189 11271
rect 20404 11240 21189 11268
rect 20404 11228 20410 11240
rect 21177 11237 21189 11240
rect 21223 11237 21235 11271
rect 21177 11231 21235 11237
rect 22649 11271 22707 11277
rect 22649 11237 22661 11271
rect 22695 11268 22707 11271
rect 23008 11271 23066 11277
rect 23008 11268 23020 11271
rect 22695 11240 23020 11268
rect 22695 11237 22707 11240
rect 22649 11231 22707 11237
rect 23008 11237 23020 11240
rect 23054 11268 23066 11271
rect 24136 11268 24164 11296
rect 23054 11240 24164 11268
rect 23054 11237 23066 11240
rect 23008 11231 23066 11237
rect 4724 11172 6408 11200
rect 4982 11132 4988 11144
rect 4264 11104 4988 11132
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 2314 11024 2320 11076
rect 2372 11064 2378 11076
rect 6380 11073 6408 11172
rect 7926 11160 7932 11212
rect 7984 11160 7990 11212
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9916 11172 10057 11200
rect 9916 11160 9922 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 12049 11203 12107 11209
rect 12049 11200 12061 11203
rect 11664 11172 12061 11200
rect 11664 11160 11670 11172
rect 12049 11169 12061 11172
rect 12095 11169 12107 11203
rect 12049 11163 12107 11169
rect 14458 11160 14464 11212
rect 14516 11160 14522 11212
rect 14826 11160 14832 11212
rect 14884 11200 14890 11212
rect 15289 11203 15347 11209
rect 15289 11200 15301 11203
rect 14884 11172 15301 11200
rect 14884 11160 14890 11172
rect 15289 11169 15301 11172
rect 15335 11200 15347 11203
rect 15378 11200 15384 11212
rect 15335 11172 15384 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 18141 11203 18199 11209
rect 18141 11169 18153 11203
rect 18187 11169 18199 11203
rect 19702 11200 19708 11212
rect 19663 11172 19708 11200
rect 18141 11163 18199 11169
rect 8018 11132 8024 11144
rect 7979 11104 8024 11132
rect 8018 11092 8024 11104
rect 8076 11092 8082 11144
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9950 11132 9956 11144
rect 9539 11104 9956 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9950 11092 9956 11104
rect 10008 11132 10014 11144
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 10008 11104 10333 11132
rect 10008 11092 10014 11104
rect 10321 11101 10333 11104
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11057 11135 11115 11141
rect 11057 11132 11069 11135
rect 11020 11104 11069 11132
rect 11020 11092 11026 11104
rect 11057 11101 11069 11104
rect 11103 11132 11115 11135
rect 11790 11132 11796 11144
rect 11103 11104 11796 11132
rect 11103 11101 11115 11104
rect 11057 11095 11115 11101
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 13817 11135 13875 11141
rect 13817 11101 13829 11135
rect 13863 11132 13875 11135
rect 14274 11132 14280 11144
rect 13863 11104 14280 11132
rect 13863 11101 13875 11104
rect 13817 11095 13875 11101
rect 14274 11092 14280 11104
rect 14332 11132 14338 11144
rect 14476 11132 14504 11160
rect 14332 11104 14504 11132
rect 17129 11135 17187 11141
rect 14332 11092 14338 11104
rect 17129 11101 17141 11135
rect 17175 11132 17187 11135
rect 17218 11132 17224 11144
rect 17175 11104 17224 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 2501 11067 2559 11073
rect 2501 11064 2513 11067
rect 2372 11036 2513 11064
rect 2372 11024 2378 11036
rect 2501 11033 2513 11036
rect 2547 11033 2559 11067
rect 2501 11027 2559 11033
rect 6365 11067 6423 11073
rect 6365 11033 6377 11067
rect 6411 11033 6423 11067
rect 6365 11027 6423 11033
rect 7561 11067 7619 11073
rect 7561 11033 7573 11067
rect 7607 11064 7619 11067
rect 7742 11064 7748 11076
rect 7607 11036 7748 11064
rect 7607 11033 7619 11036
rect 7561 11027 7619 11033
rect 7742 11024 7748 11036
rect 7800 11024 7806 11076
rect 9766 11064 9772 11076
rect 9727 11036 9772 11064
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 14461 11067 14519 11073
rect 14461 11064 14473 11067
rect 13648 11036 14473 11064
rect 8570 10996 8576 11008
rect 8531 10968 8576 10996
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 13538 10956 13544 11008
rect 13596 10996 13602 11008
rect 13648 10996 13676 11036
rect 14461 11033 14473 11036
rect 14507 11033 14519 11067
rect 14461 11027 14519 11033
rect 15105 11067 15163 11073
rect 15105 11033 15117 11067
rect 15151 11033 15163 11067
rect 15105 11027 15163 11033
rect 16669 11067 16727 11073
rect 16669 11033 16681 11067
rect 16715 11064 16727 11067
rect 16942 11064 16948 11076
rect 16715 11036 16948 11064
rect 16715 11033 16727 11036
rect 16669 11027 16727 11033
rect 13596 10968 13676 10996
rect 15120 10996 15148 11027
rect 16942 11024 16948 11036
rect 17000 11064 17006 11076
rect 17589 11067 17647 11073
rect 17589 11064 17601 11067
rect 17000 11036 17601 11064
rect 17000 11024 17006 11036
rect 17589 11033 17601 11036
rect 17635 11033 17647 11067
rect 18156 11064 18184 11163
rect 19702 11160 19708 11172
rect 19760 11160 19766 11212
rect 20162 11160 20168 11212
rect 20220 11200 20226 11212
rect 20714 11200 20720 11212
rect 20220 11172 20720 11200
rect 20220 11160 20226 11172
rect 20714 11160 20720 11172
rect 20772 11200 20778 11212
rect 20901 11203 20959 11209
rect 20901 11200 20913 11203
rect 20772 11172 20913 11200
rect 20772 11160 20778 11172
rect 20901 11169 20913 11172
rect 20947 11169 20959 11203
rect 20901 11163 20959 11169
rect 25225 11203 25283 11209
rect 25225 11169 25237 11203
rect 25271 11200 25283 11203
rect 25590 11200 25596 11212
rect 25271 11172 25596 11200
rect 25271 11169 25283 11172
rect 25225 11163 25283 11169
rect 25590 11160 25596 11172
rect 25648 11160 25654 11212
rect 18322 11132 18328 11144
rect 18283 11104 18328 11132
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 19426 11092 19432 11144
rect 19484 11132 19490 11144
rect 20254 11132 20260 11144
rect 19484 11104 20260 11132
rect 19484 11092 19490 11104
rect 20254 11092 20260 11104
rect 20312 11092 20318 11144
rect 22554 11092 22560 11144
rect 22612 11132 22618 11144
rect 22741 11135 22799 11141
rect 22741 11132 22753 11135
rect 22612 11104 22753 11132
rect 22612 11092 22618 11104
rect 22741 11101 22753 11104
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 17589 11027 17647 11033
rect 17880 11036 18184 11064
rect 19889 11067 19947 11073
rect 15654 10996 15660 11008
rect 15120 10968 15660 10996
rect 13596 10956 13602 10968
rect 15654 10956 15660 10968
rect 15712 10956 15718 11008
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 17678 10996 17684 11008
rect 16632 10968 17684 10996
rect 16632 10956 16638 10968
rect 17678 10956 17684 10968
rect 17736 10996 17742 11008
rect 17880 10996 17908 11036
rect 19889 11033 19901 11067
rect 19935 11064 19947 11067
rect 20346 11064 20352 11076
rect 19935 11036 20352 11064
rect 19935 11033 19947 11036
rect 19889 11027 19947 11033
rect 20346 11024 20352 11036
rect 20404 11024 20410 11076
rect 17736 10968 17908 10996
rect 17736 10956 17742 10968
rect 18230 10956 18236 11008
rect 18288 10996 18294 11008
rect 18690 10996 18696 11008
rect 18288 10968 18696 10996
rect 18288 10956 18294 10968
rect 18690 10956 18696 10968
rect 18748 10956 18754 11008
rect 22097 10999 22155 11005
rect 22097 10965 22109 10999
rect 22143 10996 22155 10999
rect 22370 10996 22376 11008
rect 22143 10968 22376 10996
rect 22143 10965 22155 10968
rect 22097 10959 22155 10965
rect 22370 10956 22376 10968
rect 22428 10956 22434 11008
rect 22756 10996 22784 11095
rect 23658 10996 23664 11008
rect 22756 10968 23664 10996
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 23750 10956 23756 11008
rect 23808 10996 23814 11008
rect 24121 10999 24179 11005
rect 24121 10996 24133 10999
rect 23808 10968 24133 10996
rect 23808 10956 23814 10968
rect 24121 10965 24133 10968
rect 24167 10965 24179 10999
rect 24121 10959 24179 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2225 10795 2283 10801
rect 2225 10761 2237 10795
rect 2271 10792 2283 10795
rect 2958 10792 2964 10804
rect 2271 10764 2964 10792
rect 2271 10761 2283 10764
rect 2225 10755 2283 10761
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 3970 10792 3976 10804
rect 3931 10764 3976 10792
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 4982 10792 4988 10804
rect 4943 10764 4988 10792
rect 4982 10752 4988 10764
rect 5040 10792 5046 10804
rect 5258 10792 5264 10804
rect 5040 10764 5264 10792
rect 5040 10752 5046 10764
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 6181 10795 6239 10801
rect 6181 10792 6193 10795
rect 5592 10764 6193 10792
rect 5592 10752 5598 10764
rect 6181 10761 6193 10764
rect 6227 10761 6239 10795
rect 6181 10755 6239 10761
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 6822 10792 6828 10804
rect 6687 10764 6828 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 7837 10795 7895 10801
rect 7837 10761 7849 10795
rect 7883 10792 7895 10795
rect 8018 10792 8024 10804
rect 7883 10764 8024 10792
rect 7883 10761 7895 10764
rect 7837 10755 7895 10761
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 10870 10792 10876 10804
rect 10831 10764 10876 10792
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 12526 10752 12532 10804
rect 12584 10792 12590 10804
rect 12805 10795 12863 10801
rect 12805 10792 12817 10795
rect 12584 10764 12817 10792
rect 12584 10752 12590 10764
rect 12805 10761 12817 10764
rect 12851 10792 12863 10795
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12851 10764 12909 10792
rect 12851 10761 12863 10764
rect 12805 10755 12863 10761
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 13446 10792 13452 10804
rect 12897 10755 12955 10761
rect 13096 10764 13452 10792
rect 1762 10684 1768 10736
rect 1820 10724 1826 10736
rect 2409 10727 2467 10733
rect 2409 10724 2421 10727
rect 1820 10696 2421 10724
rect 1820 10684 1826 10696
rect 2409 10693 2421 10696
rect 2455 10693 2467 10727
rect 2409 10687 2467 10693
rect 5166 10684 5172 10736
rect 5224 10724 5230 10736
rect 7926 10724 7932 10736
rect 5224 10696 7932 10724
rect 5224 10684 5230 10696
rect 7926 10684 7932 10696
rect 7984 10724 7990 10736
rect 8113 10727 8171 10733
rect 8113 10724 8125 10727
rect 7984 10696 8125 10724
rect 7984 10684 7990 10696
rect 8113 10693 8125 10696
rect 8159 10724 8171 10727
rect 8202 10724 8208 10736
rect 8159 10696 8208 10724
rect 8159 10693 8171 10696
rect 8113 10687 8171 10693
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 11790 10684 11796 10736
rect 11848 10724 11854 10736
rect 11885 10727 11943 10733
rect 11885 10724 11897 10727
rect 11848 10696 11897 10724
rect 11848 10684 11854 10696
rect 11885 10693 11897 10696
rect 11931 10724 11943 10727
rect 13096 10724 13124 10764
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 14826 10792 14832 10804
rect 14599 10764 14832 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 16482 10792 16488 10804
rect 16443 10764 16488 10792
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 20714 10792 20720 10804
rect 20675 10764 20720 10792
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 11931 10696 13124 10724
rect 13173 10727 13231 10733
rect 11931 10693 11943 10696
rect 11885 10687 11943 10693
rect 13173 10693 13185 10727
rect 13219 10724 13231 10727
rect 13998 10724 14004 10736
rect 13219 10696 14004 10724
rect 13219 10693 13231 10696
rect 13173 10687 13231 10693
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 14734 10684 14740 10736
rect 14792 10724 14798 10736
rect 15105 10727 15163 10733
rect 15105 10724 15117 10727
rect 14792 10696 15117 10724
rect 14792 10684 14798 10696
rect 15105 10693 15117 10696
rect 15151 10693 15163 10727
rect 15105 10687 15163 10693
rect 22097 10727 22155 10733
rect 22097 10693 22109 10727
rect 22143 10724 22155 10727
rect 23474 10724 23480 10736
rect 22143 10696 23480 10724
rect 22143 10693 22155 10696
rect 22097 10687 22155 10693
rect 23474 10684 23480 10696
rect 23532 10684 23538 10736
rect 2590 10616 2596 10668
rect 2648 10656 2654 10668
rect 2774 10656 2780 10668
rect 2648 10628 2780 10656
rect 2648 10616 2654 10628
rect 2774 10616 2780 10628
rect 2832 10656 2838 10668
rect 2961 10659 3019 10665
rect 2832 10628 2877 10656
rect 2832 10616 2838 10628
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3234 10656 3240 10668
rect 3007 10628 3240 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3234 10616 3240 10628
rect 3292 10656 3298 10668
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 3292 10628 4537 10656
rect 3292 10616 3298 10628
rect 4525 10625 4537 10628
rect 4571 10656 4583 10659
rect 4706 10656 4712 10668
rect 4571 10628 4712 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 6362 10656 6368 10668
rect 5767 10628 6368 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 11422 10656 11428 10668
rect 11383 10628 11428 10656
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 13725 10659 13783 10665
rect 13725 10656 13737 10659
rect 12492 10628 13737 10656
rect 12492 10616 12498 10628
rect 13725 10625 13737 10628
rect 13771 10656 13783 10659
rect 14093 10659 14151 10665
rect 14093 10656 14105 10659
rect 13771 10628 14105 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 14093 10625 14105 10628
rect 14139 10625 14151 10659
rect 15654 10656 15660 10668
rect 15615 10628 15660 10656
rect 14093 10619 14151 10625
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 20714 10616 20720 10668
rect 20772 10656 20778 10668
rect 20772 10628 22324 10656
rect 20772 10616 20778 10628
rect 3786 10588 3792 10600
rect 3699 10560 3792 10588
rect 3786 10548 3792 10560
rect 3844 10588 3850 10600
rect 4246 10588 4252 10600
rect 3844 10560 4252 10588
rect 3844 10548 3850 10560
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 5350 10548 5356 10600
rect 5408 10588 5414 10600
rect 5445 10591 5503 10597
rect 5445 10588 5457 10591
rect 5408 10560 5457 10588
rect 5408 10548 5414 10560
rect 5445 10557 5457 10560
rect 5491 10557 5503 10591
rect 5445 10551 5503 10557
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10588 7067 10591
rect 8110 10588 8116 10600
rect 7055 10560 8116 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8294 10588 8300 10600
rect 8255 10560 8300 10588
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 8570 10597 8576 10600
rect 8564 10588 8576 10597
rect 8531 10560 8576 10588
rect 8564 10551 8576 10560
rect 8570 10548 8576 10551
rect 8628 10548 8634 10600
rect 12805 10591 12863 10597
rect 12805 10557 12817 10591
rect 12851 10588 12863 10591
rect 13446 10588 13452 10600
rect 12851 10560 13452 10588
rect 12851 10557 12863 10560
rect 12805 10551 12863 10557
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 14642 10548 14648 10600
rect 14700 10588 14706 10600
rect 15381 10591 15439 10597
rect 15381 10588 15393 10591
rect 14700 10560 15393 10588
rect 14700 10548 14706 10560
rect 15381 10557 15393 10560
rect 15427 10557 15439 10591
rect 15381 10551 15439 10557
rect 16577 10591 16635 10597
rect 16577 10557 16589 10591
rect 16623 10557 16635 10591
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 16577 10551 16635 10557
rect 17788 10560 18061 10588
rect 2869 10523 2927 10529
rect 2869 10489 2881 10523
rect 2915 10520 2927 10523
rect 2958 10520 2964 10532
rect 2915 10492 2964 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 2958 10480 2964 10492
rect 3016 10480 3022 10532
rect 7282 10520 7288 10532
rect 7243 10492 7288 10520
rect 7282 10480 7288 10492
rect 7340 10480 7346 10532
rect 11149 10523 11207 10529
rect 11149 10489 11161 10523
rect 11195 10489 11207 10523
rect 12526 10520 12532 10532
rect 11149 10483 11207 10489
rect 11716 10492 12532 10520
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 3421 10455 3479 10461
rect 3421 10421 3433 10455
rect 3467 10452 3479 10455
rect 4430 10452 4436 10464
rect 3467 10424 4436 10452
rect 3467 10421 3479 10424
rect 3421 10415 3479 10421
rect 4430 10412 4436 10424
rect 4488 10452 4494 10464
rect 7374 10452 7380 10464
rect 4488 10424 7380 10452
rect 4488 10412 4494 10424
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 9674 10452 9680 10464
rect 9635 10424 9680 10452
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 9916 10424 10241 10452
rect 9916 10412 9922 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 10686 10452 10692 10464
rect 10647 10424 10692 10452
rect 10229 10415 10287 10421
rect 10686 10412 10692 10424
rect 10744 10452 10750 10464
rect 11164 10452 11192 10483
rect 10744 10424 11192 10452
rect 11333 10455 11391 10461
rect 10744 10412 10750 10424
rect 11333 10421 11345 10455
rect 11379 10452 11391 10455
rect 11716 10452 11744 10492
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 13354 10480 13360 10532
rect 13412 10520 13418 10532
rect 13633 10523 13691 10529
rect 13633 10520 13645 10523
rect 13412 10492 13645 10520
rect 13412 10480 13418 10492
rect 13633 10489 13645 10492
rect 13679 10489 13691 10523
rect 16022 10520 16028 10532
rect 15983 10492 16028 10520
rect 13633 10483 13691 10489
rect 16022 10480 16028 10492
rect 16080 10520 16086 10532
rect 16592 10520 16620 10551
rect 16080 10492 16620 10520
rect 16853 10523 16911 10529
rect 16080 10480 16086 10492
rect 16853 10489 16865 10523
rect 16899 10520 16911 10523
rect 17126 10520 17132 10532
rect 16899 10492 17132 10520
rect 16899 10489 16911 10492
rect 16853 10483 16911 10489
rect 17126 10480 17132 10492
rect 17184 10480 17190 10532
rect 12250 10452 12256 10464
rect 11379 10424 11744 10452
rect 12163 10424 12256 10452
rect 11379 10421 11391 10424
rect 11333 10415 11391 10421
rect 12250 10412 12256 10424
rect 12308 10452 12314 10464
rect 13372 10452 13400 10480
rect 17788 10464 17816 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 18138 10548 18144 10600
rect 18196 10588 18202 10600
rect 18305 10591 18363 10597
rect 18305 10588 18317 10591
rect 18196 10560 18317 10588
rect 18196 10548 18202 10560
rect 18305 10557 18317 10560
rect 18351 10557 18363 10591
rect 18305 10551 18363 10557
rect 19702 10548 19708 10600
rect 19760 10588 19766 10600
rect 20070 10588 20076 10600
rect 19760 10560 20076 10588
rect 19760 10548 19766 10560
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10588 20867 10591
rect 21542 10588 21548 10600
rect 20855 10560 21548 10588
rect 20855 10557 20867 10560
rect 20809 10551 20867 10557
rect 21542 10548 21548 10560
rect 21600 10548 21606 10600
rect 21913 10591 21971 10597
rect 21913 10557 21925 10591
rect 21959 10588 21971 10591
rect 22296 10588 22324 10628
rect 22370 10616 22376 10668
rect 22428 10656 22434 10668
rect 22649 10659 22707 10665
rect 22649 10656 22661 10659
rect 22428 10628 22661 10656
rect 22428 10616 22434 10628
rect 22649 10625 22661 10628
rect 22695 10656 22707 10659
rect 22695 10628 23796 10656
rect 22695 10625 22707 10628
rect 22649 10619 22707 10625
rect 23768 10600 23796 10628
rect 23658 10588 23664 10600
rect 21959 10560 22232 10588
rect 22296 10560 22600 10588
rect 21959 10557 21971 10560
rect 21913 10551 21971 10557
rect 22204 10532 22232 10560
rect 20898 10480 20904 10532
rect 20956 10520 20962 10532
rect 20956 10492 22140 10520
rect 20956 10480 20962 10492
rect 12308 10424 13400 10452
rect 12308 10412 12314 10424
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 13780 10424 14933 10452
rect 13780 10412 13786 10424
rect 14921 10421 14933 10424
rect 14967 10452 14979 10455
rect 15565 10455 15623 10461
rect 15565 10452 15577 10455
rect 14967 10424 15577 10452
rect 14967 10421 14979 10424
rect 14921 10415 14979 10421
rect 15565 10421 15577 10424
rect 15611 10452 15623 10455
rect 16390 10452 16396 10464
rect 15611 10424 16396 10452
rect 15611 10421 15623 10424
rect 15565 10415 15623 10421
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 17313 10455 17371 10461
rect 17313 10452 17325 10455
rect 17276 10424 17325 10452
rect 17276 10412 17282 10424
rect 17313 10421 17325 10424
rect 17359 10421 17371 10455
rect 17770 10452 17776 10464
rect 17731 10424 17776 10452
rect 17313 10415 17371 10421
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 18506 10412 18512 10464
rect 18564 10452 18570 10464
rect 19429 10455 19487 10461
rect 19429 10452 19441 10455
rect 18564 10424 19441 10452
rect 18564 10412 18570 10424
rect 19429 10421 19441 10424
rect 19475 10421 19487 10455
rect 19429 10415 19487 10421
rect 20993 10455 21051 10461
rect 20993 10421 21005 10455
rect 21039 10452 21051 10455
rect 21266 10452 21272 10464
rect 21039 10424 21272 10452
rect 21039 10421 21051 10424
rect 20993 10415 21051 10421
rect 21266 10412 21272 10424
rect 21324 10412 21330 10464
rect 21453 10455 21511 10461
rect 21453 10421 21465 10455
rect 21499 10452 21511 10455
rect 21542 10452 21548 10464
rect 21499 10424 21548 10452
rect 21499 10421 21511 10424
rect 21453 10415 21511 10421
rect 21542 10412 21548 10424
rect 21600 10412 21606 10464
rect 22112 10452 22140 10492
rect 22186 10480 22192 10532
rect 22244 10520 22250 10532
rect 22572 10529 22600 10560
rect 23492 10560 23664 10588
rect 22373 10523 22431 10529
rect 22373 10520 22385 10523
rect 22244 10492 22385 10520
rect 22244 10480 22250 10492
rect 22373 10489 22385 10492
rect 22419 10489 22431 10523
rect 22373 10483 22431 10489
rect 22557 10523 22615 10529
rect 22557 10489 22569 10523
rect 22603 10520 22615 10523
rect 23382 10520 23388 10532
rect 22603 10492 23388 10520
rect 22603 10489 22615 10492
rect 22557 10483 22615 10489
rect 23382 10480 23388 10492
rect 23440 10480 23446 10532
rect 23492 10461 23520 10560
rect 23658 10548 23664 10560
rect 23716 10548 23722 10600
rect 23750 10548 23756 10600
rect 23808 10588 23814 10600
rect 23917 10591 23975 10597
rect 23917 10588 23929 10591
rect 23808 10560 23929 10588
rect 23808 10548 23814 10560
rect 23917 10557 23929 10560
rect 23963 10557 23975 10591
rect 23917 10551 23975 10557
rect 23017 10455 23075 10461
rect 23017 10452 23029 10455
rect 22112 10424 23029 10452
rect 23017 10421 23029 10424
rect 23063 10452 23075 10455
rect 23477 10455 23535 10461
rect 23477 10452 23489 10455
rect 23063 10424 23489 10452
rect 23063 10421 23075 10424
rect 23017 10415 23075 10421
rect 23477 10421 23489 10424
rect 23523 10421 23535 10455
rect 25038 10452 25044 10464
rect 24999 10424 25044 10452
rect 23477 10415 23535 10421
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 25590 10452 25596 10464
rect 25551 10424 25596 10452
rect 25590 10412 25596 10424
rect 25648 10412 25654 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 1854 10248 1860 10260
rect 1719 10220 1860 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 3234 10248 3240 10260
rect 2832 10220 2877 10248
rect 3195 10220 3240 10248
rect 2832 10208 2838 10220
rect 3234 10208 3240 10220
rect 3292 10248 3298 10260
rect 4249 10251 4307 10257
rect 4249 10248 4261 10251
rect 3292 10220 4261 10248
rect 3292 10208 3298 10220
rect 4249 10217 4261 10220
rect 4295 10217 4307 10251
rect 4249 10211 4307 10217
rect 4522 10208 4528 10260
rect 4580 10248 4586 10260
rect 4985 10251 5043 10257
rect 4985 10248 4997 10251
rect 4580 10220 4997 10248
rect 4580 10208 4586 10220
rect 4985 10217 4997 10220
rect 5031 10217 5043 10251
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 4985 10211 5043 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 8021 10251 8079 10257
rect 8021 10217 8033 10251
rect 8067 10248 8079 10251
rect 8110 10248 8116 10260
rect 8067 10220 8116 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 8294 10248 8300 10260
rect 8255 10220 8300 10248
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 8938 10248 8944 10260
rect 8496 10220 8944 10248
rect 1394 10140 1400 10192
rect 1452 10180 1458 10192
rect 2332 10180 2360 10208
rect 4798 10180 4804 10192
rect 1452 10152 2360 10180
rect 4759 10152 4804 10180
rect 1452 10140 1458 10152
rect 4798 10140 4804 10152
rect 4856 10140 4862 10192
rect 5077 10183 5135 10189
rect 5077 10149 5089 10183
rect 5123 10180 5135 10183
rect 5534 10180 5540 10192
rect 5123 10152 5540 10180
rect 5123 10149 5135 10152
rect 5077 10143 5135 10149
rect 5534 10140 5540 10152
rect 5592 10180 5598 10192
rect 6242 10183 6300 10189
rect 6242 10180 6254 10183
rect 5592 10152 6254 10180
rect 5592 10140 5598 10152
rect 6242 10149 6254 10152
rect 6288 10180 6300 10183
rect 6454 10180 6460 10192
rect 6288 10152 6460 10180
rect 6288 10149 6300 10152
rect 6242 10143 6300 10149
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 1762 10072 1768 10124
rect 1820 10112 1826 10124
rect 2133 10115 2191 10121
rect 2133 10112 2145 10115
rect 1820 10084 2145 10112
rect 1820 10072 1826 10084
rect 2133 10081 2145 10084
rect 2179 10081 2191 10115
rect 2133 10075 2191 10081
rect 2774 10072 2780 10124
rect 2832 10112 2838 10124
rect 5166 10112 5172 10124
rect 2832 10084 5172 10112
rect 2832 10072 2838 10084
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 5997 10115 6055 10121
rect 5997 10112 6009 10115
rect 5500 10084 6009 10112
rect 5500 10072 5506 10084
rect 5997 10081 6009 10084
rect 6043 10081 6055 10115
rect 5997 10075 6055 10081
rect 2406 10044 2412 10056
rect 2367 10016 2412 10044
rect 2406 10004 2412 10016
rect 2464 10044 2470 10056
rect 3418 10044 3424 10056
rect 2464 10016 3424 10044
rect 2464 10004 2470 10016
rect 3418 10004 3424 10016
rect 3476 10044 3482 10056
rect 3513 10047 3571 10053
rect 3513 10044 3525 10047
rect 3476 10016 3525 10044
rect 3476 10004 3482 10016
rect 3513 10013 3525 10016
rect 3559 10013 3571 10047
rect 3513 10007 3571 10013
rect 4525 9979 4583 9985
rect 4525 9945 4537 9979
rect 4571 9976 4583 9979
rect 4706 9976 4712 9988
rect 4571 9948 4712 9976
rect 4571 9945 4583 9948
rect 4525 9939 4583 9945
rect 4706 9936 4712 9948
rect 4764 9936 4770 9988
rect 8312 9920 8340 10208
rect 8496 10121 8524 10220
rect 8938 10208 8944 10220
rect 8996 10248 9002 10260
rect 8996 10220 11560 10248
rect 8996 10208 9002 10220
rect 10226 10180 10232 10192
rect 10187 10152 10232 10180
rect 10226 10140 10232 10152
rect 10284 10140 10290 10192
rect 11532 10189 11560 10220
rect 13722 10208 13728 10260
rect 13780 10248 13786 10260
rect 13998 10248 14004 10260
rect 13780 10220 14004 10248
rect 13780 10208 13786 10220
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 14642 10208 14648 10260
rect 14700 10248 14706 10260
rect 15013 10251 15071 10257
rect 15013 10248 15025 10251
rect 14700 10220 15025 10248
rect 14700 10208 14706 10220
rect 15013 10217 15025 10220
rect 15059 10217 15071 10251
rect 17310 10248 17316 10260
rect 15013 10211 15071 10217
rect 15488 10220 15976 10248
rect 17271 10220 17316 10248
rect 11517 10183 11575 10189
rect 11517 10149 11529 10183
rect 11563 10149 11575 10183
rect 13170 10180 13176 10192
rect 13131 10152 13176 10180
rect 11517 10143 11575 10149
rect 13170 10140 13176 10152
rect 13228 10140 13234 10192
rect 13354 10140 13360 10192
rect 13412 10180 13418 10192
rect 15488 10180 15516 10220
rect 15654 10189 15660 10192
rect 15648 10180 15660 10189
rect 13412 10152 15516 10180
rect 15615 10152 15660 10180
rect 13412 10140 13418 10152
rect 15648 10143 15660 10152
rect 15654 10140 15660 10143
rect 15712 10140 15718 10192
rect 15838 10140 15844 10192
rect 15896 10140 15902 10192
rect 15948 10180 15976 10220
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 17678 10248 17684 10260
rect 17639 10220 17684 10248
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 18230 10208 18236 10260
rect 18288 10248 18294 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 18288 10220 18429 10248
rect 18288 10208 18294 10220
rect 18417 10217 18429 10220
rect 18463 10248 18475 10251
rect 18598 10248 18604 10260
rect 18463 10220 18604 10248
rect 18463 10217 18475 10220
rect 18417 10211 18475 10217
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 20714 10248 20720 10260
rect 20675 10220 20720 10248
rect 20714 10208 20720 10220
rect 20772 10208 20778 10260
rect 22830 10248 22836 10260
rect 22791 10220 22836 10248
rect 22830 10208 22836 10220
rect 22888 10208 22894 10260
rect 23750 10248 23756 10260
rect 23711 10220 23756 10248
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 17402 10180 17408 10192
rect 15948 10152 17408 10180
rect 17402 10140 17408 10152
rect 17460 10140 17466 10192
rect 18506 10140 18512 10192
rect 18564 10180 18570 10192
rect 18564 10152 18609 10180
rect 18564 10140 18570 10152
rect 21910 10140 21916 10192
rect 21968 10180 21974 10192
rect 21968 10152 22876 10180
rect 21968 10140 21974 10152
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10081 8539 10115
rect 8481 10075 8539 10081
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 10318 10112 10324 10124
rect 9732 10084 10324 10112
rect 9732 10072 9738 10084
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 11241 10115 11299 10121
rect 11241 10081 11253 10115
rect 11287 10112 11299 10115
rect 11974 10112 11980 10124
rect 11287 10084 11980 10112
rect 11287 10081 11299 10084
rect 11241 10075 11299 10081
rect 10134 10044 10140 10056
rect 10095 10016 10140 10044
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 8662 9976 8668 9988
rect 8623 9948 8668 9976
rect 8662 9936 8668 9948
rect 8720 9936 8726 9988
rect 9125 9979 9183 9985
rect 9125 9945 9137 9979
rect 9171 9976 9183 9979
rect 9490 9976 9496 9988
rect 9171 9948 9496 9976
rect 9171 9945 9183 9948
rect 9125 9939 9183 9945
rect 9490 9936 9496 9948
rect 9548 9936 9554 9988
rect 9769 9979 9827 9985
rect 9769 9945 9781 9979
rect 9815 9976 9827 9979
rect 11256 9976 11284 10075
rect 11974 10072 11980 10084
rect 12032 10072 12038 10124
rect 12986 10112 12992 10124
rect 12947 10084 12992 10112
rect 12986 10072 12992 10084
rect 13044 10112 13050 10124
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13044 10084 13645 10112
rect 13044 10072 13050 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 14185 10115 14243 10121
rect 14185 10081 14197 10115
rect 14231 10112 14243 10115
rect 14642 10112 14648 10124
rect 14231 10084 14648 10112
rect 14231 10081 14243 10084
rect 14185 10075 14243 10081
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 15381 10115 15439 10121
rect 15381 10081 15393 10115
rect 15427 10112 15439 10115
rect 15856 10112 15884 10140
rect 22848 10124 22876 10152
rect 15427 10084 15884 10112
rect 15427 10081 15439 10084
rect 15381 10075 15439 10081
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 18233 10115 18291 10121
rect 18233 10112 18245 10115
rect 18104 10084 18245 10112
rect 18104 10072 18110 10084
rect 18233 10081 18245 10084
rect 18279 10081 18291 10115
rect 18233 10075 18291 10081
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 21726 10121 21732 10124
rect 19521 10115 19579 10121
rect 19521 10112 19533 10115
rect 19484 10084 19533 10112
rect 19484 10072 19490 10084
rect 19521 10081 19533 10084
rect 19567 10081 19579 10115
rect 19521 10075 19579 10081
rect 21361 10115 21419 10121
rect 21361 10081 21373 10115
rect 21407 10112 21419 10115
rect 21720 10112 21732 10121
rect 21407 10084 21732 10112
rect 21407 10081 21419 10084
rect 21361 10075 21419 10081
rect 21720 10075 21732 10084
rect 21726 10072 21732 10075
rect 21784 10072 21790 10124
rect 22830 10072 22836 10124
rect 22888 10072 22894 10124
rect 23658 10072 23664 10124
rect 23716 10112 23722 10124
rect 23937 10115 23995 10121
rect 23937 10112 23949 10115
rect 23716 10084 23949 10112
rect 23716 10072 23722 10084
rect 23937 10081 23949 10084
rect 23983 10081 23995 10115
rect 23937 10075 23995 10081
rect 24204 10115 24262 10121
rect 24204 10081 24216 10115
rect 24250 10112 24262 10115
rect 25038 10112 25044 10124
rect 24250 10084 25044 10112
rect 24250 10081 24262 10084
rect 24204 10075 24262 10081
rect 25038 10072 25044 10084
rect 25096 10072 25102 10124
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 12492 10016 13277 10044
rect 12492 10004 12498 10016
rect 13265 10013 13277 10016
rect 13311 10044 13323 10047
rect 13446 10044 13452 10056
rect 13311 10016 13452 10044
rect 13311 10013 13323 10016
rect 13265 10007 13323 10013
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 16390 10004 16396 10056
rect 16448 10044 16454 10056
rect 19150 10044 19156 10056
rect 16448 10016 19156 10044
rect 16448 10004 16454 10016
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 20898 10004 20904 10056
rect 20956 10044 20962 10056
rect 21453 10047 21511 10053
rect 21453 10044 21465 10047
rect 20956 10016 21465 10044
rect 20956 10004 20962 10016
rect 21453 10013 21465 10016
rect 21499 10013 21511 10047
rect 21453 10007 21511 10013
rect 9815 9948 11284 9976
rect 9815 9945 9827 9948
rect 9769 9939 9827 9945
rect 12158 9936 12164 9988
rect 12216 9976 12222 9988
rect 12713 9979 12771 9985
rect 12216 9948 12664 9976
rect 12216 9936 12222 9948
rect 1857 9911 1915 9917
rect 1857 9877 1869 9911
rect 1903 9908 1915 9911
rect 2314 9908 2320 9920
rect 1903 9880 2320 9908
rect 1903 9877 1915 9880
rect 1857 9871 1915 9877
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 5350 9868 5356 9920
rect 5408 9908 5414 9920
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 5408 9880 5825 9908
rect 5408 9868 5414 9880
rect 5813 9877 5825 9880
rect 5859 9877 5871 9911
rect 5813 9871 5871 9877
rect 7377 9911 7435 9917
rect 7377 9877 7389 9911
rect 7423 9908 7435 9911
rect 7466 9908 7472 9920
rect 7423 9880 7472 9908
rect 7423 9877 7435 9880
rect 7377 9871 7435 9877
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 8294 9868 8300 9920
rect 8352 9868 8358 9920
rect 9306 9868 9312 9920
rect 9364 9908 9370 9920
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 9364 9880 9413 9908
rect 9364 9868 9370 9880
rect 9401 9877 9413 9880
rect 9447 9877 9459 9911
rect 9401 9871 9459 9877
rect 10873 9911 10931 9917
rect 10873 9877 10885 9911
rect 10919 9908 10931 9911
rect 10962 9908 10968 9920
rect 10919 9880 10968 9908
rect 10919 9877 10931 9880
rect 10873 9871 10931 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11664 9880 11989 9908
rect 11664 9868 11670 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 11977 9871 12035 9877
rect 12437 9911 12495 9917
rect 12437 9877 12449 9911
rect 12483 9908 12495 9911
rect 12526 9908 12532 9920
rect 12483 9880 12532 9908
rect 12483 9877 12495 9880
rect 12437 9871 12495 9877
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 12636 9908 12664 9948
rect 12713 9945 12725 9979
rect 12759 9976 12771 9979
rect 13630 9976 13636 9988
rect 12759 9948 13636 9976
rect 12759 9945 12771 9948
rect 12713 9939 12771 9945
rect 13630 9936 13636 9948
rect 13688 9976 13694 9988
rect 14645 9979 14703 9985
rect 14645 9976 14657 9979
rect 13688 9948 14657 9976
rect 13688 9936 13694 9948
rect 14645 9945 14657 9948
rect 14691 9945 14703 9979
rect 16850 9976 16856 9988
rect 14645 9939 14703 9945
rect 16316 9948 16856 9976
rect 15378 9908 15384 9920
rect 12636 9880 15384 9908
rect 15378 9868 15384 9880
rect 15436 9908 15442 9920
rect 16316 9908 16344 9948
rect 16850 9936 16856 9948
rect 16908 9936 16914 9988
rect 18138 9936 18144 9988
rect 18196 9976 18202 9988
rect 18877 9979 18935 9985
rect 18877 9976 18889 9979
rect 18196 9948 18889 9976
rect 18196 9936 18202 9948
rect 18877 9945 18889 9948
rect 18923 9976 18935 9979
rect 18966 9976 18972 9988
rect 18923 9948 18972 9976
rect 18923 9945 18935 9948
rect 18877 9939 18935 9945
rect 18966 9936 18972 9948
rect 19024 9936 19030 9988
rect 15436 9880 16344 9908
rect 15436 9868 15442 9880
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 16761 9911 16819 9917
rect 16761 9908 16773 9911
rect 16632 9880 16773 9908
rect 16632 9868 16638 9880
rect 16761 9877 16773 9880
rect 16807 9877 16819 9911
rect 16761 9871 16819 9877
rect 17957 9911 18015 9917
rect 17957 9877 17969 9911
rect 18003 9908 18015 9911
rect 18598 9908 18604 9920
rect 18003 9880 18604 9908
rect 18003 9877 18015 9880
rect 17957 9871 18015 9877
rect 18598 9868 18604 9880
rect 18656 9868 18662 9920
rect 19337 9911 19395 9917
rect 19337 9877 19349 9911
rect 19383 9908 19395 9911
rect 19610 9908 19616 9920
rect 19383 9880 19616 9908
rect 19383 9877 19395 9880
rect 19337 9871 19395 9877
rect 19610 9868 19616 9880
rect 19668 9868 19674 9920
rect 19705 9911 19763 9917
rect 19705 9877 19717 9911
rect 19751 9908 19763 9911
rect 20530 9908 20536 9920
rect 19751 9880 20536 9908
rect 19751 9877 19763 9880
rect 19705 9871 19763 9877
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 24946 9868 24952 9920
rect 25004 9908 25010 9920
rect 25317 9911 25375 9917
rect 25317 9908 25329 9911
rect 25004 9880 25329 9908
rect 25004 9868 25010 9880
rect 25317 9877 25329 9880
rect 25363 9877 25375 9911
rect 25317 9871 25375 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1854 9704 1860 9716
rect 1688 9676 1860 9704
rect 1688 9577 1716 9676
rect 1854 9664 1860 9676
rect 1912 9664 1918 9716
rect 4522 9704 4528 9716
rect 4080 9676 4528 9704
rect 4080 9645 4108 9676
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 5442 9664 5448 9716
rect 5500 9704 5506 9716
rect 6089 9707 6147 9713
rect 6089 9704 6101 9707
rect 5500 9676 6101 9704
rect 5500 9664 5506 9676
rect 6089 9673 6101 9676
rect 6135 9673 6147 9707
rect 6454 9704 6460 9716
rect 6415 9676 6460 9704
rect 6089 9667 6147 9673
rect 4065 9639 4123 9645
rect 4065 9605 4077 9639
rect 4111 9605 4123 9639
rect 6104 9636 6132 9667
rect 6454 9664 6460 9676
rect 6512 9704 6518 9716
rect 6822 9704 6828 9716
rect 6512 9676 6828 9704
rect 6512 9664 6518 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 8665 9707 8723 9713
rect 8665 9704 8677 9707
rect 8628 9676 8677 9704
rect 8628 9664 8634 9676
rect 8665 9673 8677 9676
rect 8711 9673 8723 9707
rect 10318 9704 10324 9716
rect 10279 9676 10324 9704
rect 8665 9667 8723 9673
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 15654 9704 15660 9716
rect 13320 9676 13768 9704
rect 13320 9664 13326 9676
rect 7101 9639 7159 9645
rect 7101 9636 7113 9639
rect 6104 9608 7113 9636
rect 4065 9599 4123 9605
rect 7101 9605 7113 9608
rect 7147 9636 7159 9639
rect 10870 9636 10876 9648
rect 7147 9608 7328 9636
rect 10831 9608 10876 9636
rect 7147 9605 7159 9608
rect 7101 9599 7159 9605
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 2958 9528 2964 9580
rect 3016 9568 3022 9580
rect 3697 9571 3755 9577
rect 3697 9568 3709 9571
rect 3016 9540 3709 9568
rect 3016 9528 3022 9540
rect 3697 9537 3709 9540
rect 3743 9568 3755 9571
rect 4154 9568 4160 9580
rect 3743 9540 4160 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 7300 9577 7328 9608
rect 10870 9596 10876 9608
rect 10928 9596 10934 9648
rect 12253 9639 12311 9645
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 12434 9636 12440 9648
rect 12299 9608 12440 9636
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 13173 9639 13231 9645
rect 13173 9605 13185 9639
rect 13219 9636 13231 9639
rect 13354 9636 13360 9648
rect 13219 9608 13360 9636
rect 13219 9605 13231 9608
rect 13173 9599 13231 9605
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 13740 9636 13768 9676
rect 15120 9676 15660 9704
rect 15120 9648 15148 9676
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 18230 9664 18236 9716
rect 18288 9704 18294 9716
rect 18601 9707 18659 9713
rect 18601 9704 18613 9707
rect 18288 9676 18613 9704
rect 18288 9664 18294 9676
rect 18601 9673 18613 9676
rect 18647 9673 18659 9707
rect 18601 9667 18659 9673
rect 18782 9664 18788 9716
rect 18840 9704 18846 9716
rect 23382 9704 23388 9716
rect 18840 9676 23388 9704
rect 18840 9664 18846 9676
rect 23382 9664 23388 9676
rect 23440 9664 23446 9716
rect 23658 9664 23664 9716
rect 23716 9704 23722 9716
rect 23845 9707 23903 9713
rect 23845 9704 23857 9707
rect 23716 9676 23857 9704
rect 23716 9664 23722 9676
rect 23845 9673 23857 9676
rect 23891 9673 23903 9707
rect 23845 9667 23903 9673
rect 14093 9639 14151 9645
rect 14093 9636 14105 9639
rect 13740 9608 14105 9636
rect 14093 9605 14105 9608
rect 14139 9605 14151 9639
rect 14093 9599 14151 9605
rect 15102 9596 15108 9648
rect 15160 9596 15166 9648
rect 17865 9639 17923 9645
rect 17865 9605 17877 9639
rect 17911 9636 17923 9639
rect 17954 9636 17960 9648
rect 17911 9608 17960 9636
rect 17911 9605 17923 9608
rect 17865 9599 17923 9605
rect 17954 9596 17960 9608
rect 18012 9636 18018 9648
rect 18506 9636 18512 9648
rect 18012 9608 18512 9636
rect 18012 9596 18018 9608
rect 18506 9596 18512 9608
rect 18564 9596 18570 9648
rect 20257 9639 20315 9645
rect 20257 9605 20269 9639
rect 20303 9636 20315 9639
rect 21174 9636 21180 9648
rect 20303 9608 21180 9636
rect 20303 9605 20315 9608
rect 20257 9599 20315 9605
rect 21174 9596 21180 9608
rect 21232 9596 21238 9648
rect 23477 9639 23535 9645
rect 23477 9605 23489 9639
rect 23523 9636 23535 9639
rect 23566 9636 23572 9648
rect 23523 9608 23572 9636
rect 23523 9605 23535 9608
rect 23477 9599 23535 9605
rect 23566 9596 23572 9608
rect 23624 9596 23630 9648
rect 24118 9636 24124 9648
rect 24079 9608 24124 9636
rect 24118 9596 24124 9608
rect 24176 9596 24182 9648
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 11425 9571 11483 9577
rect 11425 9537 11437 9571
rect 11471 9568 11483 9571
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 11471 9540 11897 9568
rect 11471 9537 11483 9540
rect 11425 9531 11483 9537
rect 11885 9537 11897 9540
rect 11931 9568 11943 9571
rect 12342 9568 12348 9580
rect 11931 9540 12348 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 1940 9503 1998 9509
rect 1940 9469 1952 9503
rect 1986 9500 1998 9503
rect 2406 9500 2412 9512
rect 1986 9472 2412 9500
rect 1986 9469 1998 9472
rect 1940 9463 1998 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 7300 9500 7328 9531
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 13538 9568 13544 9580
rect 13499 9540 13544 9568
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 18046 9528 18052 9580
rect 18104 9568 18110 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 18104 9540 18245 9568
rect 18104 9528 18110 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 21082 9528 21088 9580
rect 21140 9568 21146 9580
rect 21269 9571 21327 9577
rect 21269 9568 21281 9571
rect 21140 9540 21281 9568
rect 21140 9528 21146 9540
rect 21269 9537 21281 9540
rect 21315 9537 21327 9571
rect 21269 9531 21327 9537
rect 22005 9571 22063 9577
rect 22005 9537 22017 9571
rect 22051 9568 22063 9571
rect 22094 9568 22100 9580
rect 22051 9540 22100 9568
rect 22051 9537 22063 9540
rect 22005 9531 22063 9537
rect 22094 9528 22100 9540
rect 22152 9568 22158 9580
rect 22741 9571 22799 9577
rect 22741 9568 22753 9571
rect 22152 9540 22753 9568
rect 22152 9528 22158 9540
rect 22741 9537 22753 9540
rect 22787 9537 22799 9571
rect 22741 9531 22799 9537
rect 24486 9528 24492 9580
rect 24544 9568 24550 9580
rect 24581 9571 24639 9577
rect 24581 9568 24593 9571
rect 24544 9540 24593 9568
rect 24544 9528 24550 9540
rect 24581 9537 24593 9540
rect 24627 9568 24639 9571
rect 25593 9571 25651 9577
rect 25593 9568 25605 9571
rect 24627 9540 25605 9568
rect 24627 9537 24639 9540
rect 24581 9531 24639 9537
rect 25593 9537 25605 9540
rect 25639 9537 25651 9571
rect 25593 9531 25651 9537
rect 8294 9500 8300 9512
rect 7300 9472 8300 9500
rect 8294 9460 8300 9472
rect 8352 9500 8358 9512
rect 8938 9500 8944 9512
rect 8352 9472 8944 9500
rect 8352 9460 8358 9472
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 12989 9503 13047 9509
rect 12989 9469 13001 9503
rect 13035 9500 13047 9503
rect 13725 9503 13783 9509
rect 13725 9500 13737 9503
rect 13035 9472 13737 9500
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 13725 9469 13737 9472
rect 13771 9500 13783 9503
rect 13814 9500 13820 9512
rect 13771 9472 13820 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15243 9472 15485 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15740 9503 15798 9509
rect 15740 9500 15752 9503
rect 15473 9463 15531 9469
rect 15580 9472 15752 9500
rect 4424 9435 4482 9441
rect 4424 9401 4436 9435
rect 4470 9432 4482 9435
rect 4522 9432 4528 9444
rect 4470 9404 4528 9432
rect 4470 9401 4482 9404
rect 4424 9395 4482 9401
rect 4522 9392 4528 9404
rect 4580 9392 4586 9444
rect 7466 9392 7472 9444
rect 7524 9441 7530 9444
rect 7524 9435 7588 9441
rect 7524 9401 7542 9435
rect 7576 9401 7588 9435
rect 9674 9432 9680 9444
rect 9635 9404 9680 9432
rect 7524 9395 7588 9401
rect 7524 9392 7530 9395
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 10689 9435 10747 9441
rect 10689 9401 10701 9435
rect 10735 9432 10747 9435
rect 11146 9432 11152 9444
rect 10735 9404 11152 9432
rect 10735 9401 10747 9404
rect 10689 9395 10747 9401
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 13630 9432 13636 9444
rect 13591 9404 13636 9432
rect 13630 9392 13636 9404
rect 13688 9392 13694 9444
rect 14645 9435 14703 9441
rect 14645 9401 14657 9435
rect 14691 9432 14703 9435
rect 14826 9432 14832 9444
rect 14691 9404 14832 9432
rect 14691 9401 14703 9404
rect 14645 9395 14703 9401
rect 14826 9392 14832 9404
rect 14884 9432 14890 9444
rect 15580 9432 15608 9472
rect 15740 9469 15752 9472
rect 15786 9500 15798 9503
rect 16022 9500 16028 9512
rect 15786 9472 16028 9500
rect 15786 9469 15798 9472
rect 15740 9463 15798 9469
rect 16022 9460 16028 9472
rect 16080 9500 16086 9512
rect 16482 9500 16488 9512
rect 16080 9472 16488 9500
rect 16080 9460 16086 9472
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 18877 9503 18935 9509
rect 18877 9469 18889 9503
rect 18923 9469 18935 9503
rect 19144 9503 19202 9509
rect 19144 9500 19156 9503
rect 18877 9463 18935 9469
rect 18984 9472 19156 9500
rect 17405 9435 17463 9441
rect 17405 9432 17417 9435
rect 14884 9404 15608 9432
rect 16592 9404 17417 9432
rect 14884 9392 14890 9404
rect 16592 9376 16620 9404
rect 17405 9401 17417 9404
rect 17451 9401 17463 9435
rect 17405 9395 17463 9401
rect 17770 9392 17776 9444
rect 17828 9432 17834 9444
rect 18138 9432 18144 9444
rect 17828 9404 18144 9432
rect 17828 9392 17834 9404
rect 18138 9392 18144 9404
rect 18196 9432 18202 9444
rect 18892 9432 18920 9463
rect 18984 9444 19012 9472
rect 19144 9469 19156 9472
rect 19190 9500 19202 9503
rect 19610 9500 19616 9512
rect 19190 9472 19616 9500
rect 19190 9469 19202 9472
rect 19144 9463 19202 9469
rect 19610 9460 19616 9472
rect 19668 9460 19674 9512
rect 20714 9460 20720 9512
rect 20772 9500 20778 9512
rect 21729 9503 21787 9509
rect 21729 9500 21741 9503
rect 20772 9472 21741 9500
rect 20772 9460 20778 9472
rect 21729 9469 21741 9472
rect 21775 9500 21787 9503
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 21775 9472 22385 9500
rect 21775 9469 21787 9472
rect 21729 9463 21787 9469
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 25409 9503 25467 9509
rect 25409 9500 25421 9503
rect 22373 9463 22431 9469
rect 24596 9472 25421 9500
rect 24596 9444 24624 9472
rect 25409 9469 25421 9472
rect 25455 9469 25467 9503
rect 25409 9463 25467 9469
rect 18196 9404 18920 9432
rect 18196 9392 18202 9404
rect 18966 9392 18972 9444
rect 19024 9392 19030 9444
rect 21082 9392 21088 9444
rect 21140 9432 21146 9444
rect 21634 9432 21640 9444
rect 21140 9404 21640 9432
rect 21140 9392 21146 9404
rect 21634 9392 21640 9404
rect 21692 9432 21698 9444
rect 21913 9435 21971 9441
rect 21913 9432 21925 9435
rect 21692 9404 21925 9432
rect 21692 9392 21698 9404
rect 21913 9401 21925 9404
rect 21959 9401 21971 9435
rect 21913 9395 21971 9401
rect 23566 9392 23572 9444
rect 23624 9432 23630 9444
rect 24578 9432 24584 9444
rect 23624 9404 24440 9432
rect 24491 9404 24584 9432
rect 23624 9392 23630 9404
rect 3050 9364 3056 9376
rect 3011 9336 3056 9364
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 4982 9324 4988 9376
rect 5040 9364 5046 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5040 9336 5549 9364
rect 5040 9324 5046 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 9214 9364 9220 9376
rect 9175 9336 9220 9364
rect 5537 9327 5595 9333
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 9766 9364 9772 9376
rect 9727 9336 9772 9364
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11330 9364 11336 9376
rect 11020 9336 11336 9364
rect 11020 9324 11026 9336
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 13170 9324 13176 9376
rect 13228 9364 13234 9376
rect 14921 9367 14979 9373
rect 14921 9364 14933 9367
rect 13228 9336 14933 9364
rect 13228 9324 13234 9336
rect 14921 9333 14933 9336
rect 14967 9364 14979 9367
rect 15197 9367 15255 9373
rect 15197 9364 15209 9367
rect 14967 9336 15209 9364
rect 14967 9333 14979 9336
rect 14921 9327 14979 9333
rect 15197 9333 15209 9336
rect 15243 9364 15255 9367
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 15243 9336 15301 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15289 9333 15301 9336
rect 15335 9364 15347 9367
rect 15838 9364 15844 9376
rect 15335 9336 15844 9364
rect 15335 9333 15347 9336
rect 15289 9327 15347 9333
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 16574 9324 16580 9376
rect 16632 9324 16638 9376
rect 16850 9364 16856 9376
rect 16811 9336 16856 9364
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 20898 9364 20904 9376
rect 20859 9336 20904 9364
rect 20898 9324 20904 9336
rect 20956 9324 20962 9376
rect 21443 9367 21501 9373
rect 21443 9333 21455 9367
rect 21489 9364 21501 9367
rect 21818 9364 21824 9376
rect 21489 9336 21824 9364
rect 21489 9333 21501 9336
rect 21443 9327 21501 9333
rect 21818 9324 21824 9336
rect 21876 9324 21882 9376
rect 24412 9364 24440 9404
rect 24578 9392 24584 9404
rect 24636 9392 24642 9444
rect 24673 9435 24731 9441
rect 24673 9401 24685 9435
rect 24719 9432 24731 9435
rect 24946 9432 24952 9444
rect 24719 9404 24952 9432
rect 24719 9401 24731 9404
rect 24673 9395 24731 9401
rect 24688 9364 24716 9395
rect 24946 9392 24952 9404
rect 25004 9392 25010 9444
rect 25038 9364 25044 9376
rect 24412 9336 24716 9364
rect 24999 9336 25044 9364
rect 25038 9324 25044 9336
rect 25096 9324 25102 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1452 9132 1593 9160
rect 1452 9120 1458 9132
rect 1581 9129 1593 9132
rect 1627 9160 1639 9163
rect 2130 9160 2136 9172
rect 1627 9132 2136 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 3050 9160 3056 9172
rect 2424 9132 3056 9160
rect 2424 9104 2452 9132
rect 3050 9120 3056 9132
rect 3108 9120 3114 9172
rect 3418 9160 3424 9172
rect 3379 9132 3424 9160
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 3881 9163 3939 9169
rect 3881 9129 3893 9163
rect 3927 9160 3939 9163
rect 4522 9160 4528 9172
rect 3927 9132 4528 9160
rect 3927 9129 3939 9132
rect 3881 9123 3939 9129
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 5077 9163 5135 9169
rect 5077 9160 5089 9163
rect 4856 9132 5089 9160
rect 4856 9120 4862 9132
rect 5077 9129 5089 9132
rect 5123 9129 5135 9163
rect 5534 9160 5540 9172
rect 5495 9132 5540 9160
rect 5077 9123 5135 9129
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 5626 9120 5632 9172
rect 5684 9160 5690 9172
rect 6362 9160 6368 9172
rect 5684 9132 6368 9160
rect 5684 9120 5690 9132
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 6914 9160 6920 9172
rect 6875 9132 6920 9160
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7156 9132 8616 9160
rect 7156 9120 7162 9132
rect 2271 9095 2329 9101
rect 2271 9092 2283 9095
rect 2148 9064 2283 9092
rect 1854 8820 1860 8832
rect 1815 8792 1860 8820
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 2148 8820 2176 9064
rect 2271 9061 2283 9064
rect 2317 9061 2329 9095
rect 2271 9055 2329 9061
rect 2406 9052 2412 9104
rect 2464 9092 2470 9104
rect 2464 9064 2557 9092
rect 2464 9052 2470 9064
rect 3436 9024 3464 9120
rect 4617 9095 4675 9101
rect 4617 9061 4629 9095
rect 4663 9092 4675 9095
rect 4890 9092 4896 9104
rect 4663 9064 4896 9092
rect 4663 9061 4675 9064
rect 4617 9055 4675 9061
rect 4890 9052 4896 9064
rect 4948 9052 4954 9104
rect 6181 9095 6239 9101
rect 6181 9061 6193 9095
rect 6227 9092 6239 9095
rect 6638 9092 6644 9104
rect 6227 9064 6644 9092
rect 6227 9061 6239 9064
rect 6181 9055 6239 9061
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 8294 9052 8300 9104
rect 8352 9092 8358 9104
rect 8389 9095 8447 9101
rect 8389 9092 8401 9095
rect 8352 9064 8401 9092
rect 8352 9052 8358 9064
rect 8389 9061 8401 9064
rect 8435 9092 8447 9095
rect 8478 9092 8484 9104
rect 8435 9064 8484 9092
rect 8435 9061 8447 9064
rect 8389 9055 8447 9061
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 8588 9101 8616 9132
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 14090 9160 14096 9172
rect 13504 9132 14096 9160
rect 13504 9120 13510 9132
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 14734 9160 14740 9172
rect 14695 9132 14740 9160
rect 14734 9120 14740 9132
rect 14792 9160 14798 9172
rect 15841 9163 15899 9169
rect 15841 9160 15853 9163
rect 14792 9132 15853 9160
rect 14792 9120 14798 9132
rect 15841 9129 15853 9132
rect 15887 9129 15899 9163
rect 15841 9123 15899 9129
rect 18966 9120 18972 9172
rect 19024 9160 19030 9172
rect 19061 9163 19119 9169
rect 19061 9160 19073 9163
rect 19024 9132 19073 9160
rect 19024 9120 19030 9132
rect 19061 9129 19073 9132
rect 19107 9129 19119 9163
rect 19061 9123 19119 9129
rect 20073 9163 20131 9169
rect 20073 9129 20085 9163
rect 20119 9160 20131 9163
rect 20438 9160 20444 9172
rect 20119 9132 20444 9160
rect 20119 9129 20131 9132
rect 20073 9123 20131 9129
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 23474 9120 23480 9172
rect 23532 9160 23538 9172
rect 23661 9163 23719 9169
rect 23661 9160 23673 9163
rect 23532 9132 23673 9160
rect 23532 9120 23538 9132
rect 23661 9129 23673 9132
rect 23707 9129 23719 9163
rect 23661 9123 23719 9129
rect 24121 9163 24179 9169
rect 24121 9129 24133 9163
rect 24167 9160 24179 9163
rect 24486 9160 24492 9172
rect 24167 9132 24492 9160
rect 24167 9129 24179 9132
rect 24121 9123 24179 9129
rect 24486 9120 24492 9132
rect 24544 9120 24550 9172
rect 24854 9160 24860 9172
rect 24767 9132 24860 9160
rect 24854 9120 24860 9132
rect 24912 9160 24918 9172
rect 26234 9160 26240 9172
rect 24912 9132 26240 9160
rect 24912 9120 24918 9132
rect 26234 9120 26240 9132
rect 26292 9120 26298 9172
rect 8573 9095 8631 9101
rect 8573 9061 8585 9095
rect 8619 9092 8631 9095
rect 9030 9092 9036 9104
rect 8619 9064 8800 9092
rect 8991 9064 9036 9092
rect 8619 9061 8631 9064
rect 8573 9055 8631 9061
rect 4709 9027 4767 9033
rect 4709 9024 4721 9027
rect 3436 8996 4721 9024
rect 4709 8993 4721 8996
rect 4755 9024 4767 9027
rect 4982 9024 4988 9036
rect 4755 8996 4988 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 2314 8956 2320 8968
rect 2275 8928 2320 8956
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8956 4675 8959
rect 5074 8956 5080 8968
rect 4663 8928 5080 8956
rect 4663 8925 4675 8928
rect 4617 8919 4675 8925
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 6454 8956 6460 8968
rect 6415 8928 6460 8956
rect 6454 8916 6460 8928
rect 6512 8956 6518 8968
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 6512 8928 7297 8956
rect 6512 8916 6518 8928
rect 7285 8925 7297 8928
rect 7331 8956 7343 8959
rect 7466 8956 7472 8968
rect 7331 8928 7472 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8570 8956 8576 8968
rect 7975 8928 8576 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 8570 8916 8576 8928
rect 8628 8956 8634 8968
rect 8665 8959 8723 8965
rect 8665 8956 8677 8959
rect 8628 8928 8677 8956
rect 8628 8916 8634 8928
rect 8665 8925 8677 8928
rect 8711 8925 8723 8959
rect 8665 8919 8723 8925
rect 5350 8848 5356 8900
rect 5408 8848 5414 8900
rect 5905 8891 5963 8897
rect 5905 8857 5917 8891
rect 5951 8888 5963 8891
rect 6730 8888 6736 8900
rect 5951 8860 6736 8888
rect 5951 8857 5963 8860
rect 5905 8851 5963 8857
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 8110 8888 8116 8900
rect 8071 8860 8116 8888
rect 8110 8848 8116 8860
rect 8168 8848 8174 8900
rect 8386 8848 8392 8900
rect 8444 8888 8450 8900
rect 8772 8888 8800 9064
rect 9030 9052 9036 9064
rect 9088 9052 9094 9104
rect 12342 9052 12348 9104
rect 12400 9092 12406 9104
rect 12958 9095 13016 9101
rect 12958 9092 12970 9095
rect 12400 9064 12970 9092
rect 12400 9052 12406 9064
rect 12958 9061 12970 9064
rect 13004 9061 13016 9095
rect 12958 9055 13016 9061
rect 13170 9052 13176 9104
rect 13228 9052 13234 9104
rect 15102 9092 15108 9104
rect 15063 9064 15108 9092
rect 15102 9052 15108 9064
rect 15160 9052 15166 9104
rect 15286 9052 15292 9104
rect 15344 9092 15350 9104
rect 15657 9095 15715 9101
rect 15657 9092 15669 9095
rect 15344 9064 15669 9092
rect 15344 9052 15350 9064
rect 15657 9061 15669 9064
rect 15703 9092 15715 9095
rect 15746 9092 15752 9104
rect 15703 9064 15752 9092
rect 15703 9061 15715 9064
rect 15657 9055 15715 9061
rect 15746 9052 15752 9064
rect 15804 9052 15810 9104
rect 15933 9095 15991 9101
rect 15933 9061 15945 9095
rect 15979 9092 15991 9095
rect 16022 9092 16028 9104
rect 15979 9064 16028 9092
rect 15979 9061 15991 9064
rect 15933 9055 15991 9061
rect 16022 9052 16028 9064
rect 16080 9052 16086 9104
rect 17954 9101 17960 9104
rect 17948 9092 17960 9101
rect 17915 9064 17960 9092
rect 17948 9055 17960 9064
rect 17954 9052 17960 9055
rect 18012 9052 18018 9104
rect 21174 9101 21180 9104
rect 21168 9092 21180 9101
rect 21087 9064 21180 9092
rect 21168 9055 21180 9064
rect 21232 9092 21238 9104
rect 22094 9092 22100 9104
rect 21232 9064 22100 9092
rect 21174 9052 21180 9055
rect 21232 9052 21238 9064
rect 22094 9052 22100 9064
rect 22152 9052 22158 9104
rect 25498 9052 25504 9104
rect 25556 9092 25562 9104
rect 26418 9092 26424 9104
rect 25556 9064 26424 9092
rect 25556 9052 25562 9064
rect 26418 9052 26424 9064
rect 26476 9052 26482 9104
rect 10496 9027 10554 9033
rect 10496 8993 10508 9027
rect 10542 9024 10554 9027
rect 11790 9024 11796 9036
rect 10542 8996 11796 9024
rect 10542 8993 10554 8996
rect 10496 8987 10554 8993
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 9024 12771 9027
rect 13188 9024 13216 9052
rect 16298 9024 16304 9036
rect 12759 8996 13216 9024
rect 16259 8996 16304 9024
rect 12759 8993 12771 8996
rect 12713 8987 12771 8993
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 17770 8984 17776 9036
rect 17828 8984 17834 9036
rect 20162 8984 20168 9036
rect 20220 9024 20226 9036
rect 22462 9024 22468 9036
rect 20220 8996 22468 9024
rect 20220 8984 20226 8996
rect 22462 8984 22468 8996
rect 22520 8984 22526 9036
rect 24670 9024 24676 9036
rect 24631 8996 24676 9024
rect 24670 8984 24676 8996
rect 24728 8984 24734 9036
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 10192 8928 10241 8956
rect 10192 8916 10198 8928
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 15470 8916 15476 8968
rect 15528 8956 15534 8968
rect 16390 8956 16396 8968
rect 15528 8928 16396 8956
rect 15528 8916 15534 8928
rect 16390 8916 16396 8928
rect 16448 8916 16454 8968
rect 17402 8916 17408 8968
rect 17460 8956 17466 8968
rect 17681 8959 17739 8965
rect 17681 8956 17693 8959
rect 17460 8928 17693 8956
rect 17460 8916 17466 8928
rect 17681 8925 17693 8928
rect 17727 8956 17739 8959
rect 17788 8956 17816 8984
rect 20898 8956 20904 8968
rect 17727 8928 17816 8956
rect 20859 8928 20904 8956
rect 17727 8925 17739 8928
rect 17681 8919 17739 8925
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 23658 8916 23664 8968
rect 23716 8956 23722 8968
rect 24949 8959 25007 8965
rect 24949 8956 24961 8959
rect 23716 8928 24961 8956
rect 23716 8916 23722 8928
rect 24949 8925 24961 8928
rect 24995 8956 25007 8959
rect 25038 8956 25044 8968
rect 24995 8928 25044 8956
rect 24995 8925 25007 8928
rect 24949 8919 25007 8925
rect 25038 8916 25044 8928
rect 25096 8916 25102 8968
rect 16666 8888 16672 8900
rect 8444 8860 8800 8888
rect 16627 8860 16672 8888
rect 8444 8848 8450 8860
rect 16666 8848 16672 8860
rect 16724 8848 16730 8900
rect 24397 8891 24455 8897
rect 24397 8857 24409 8891
rect 24443 8888 24455 8891
rect 24578 8888 24584 8900
rect 24443 8860 24584 8888
rect 24443 8857 24455 8860
rect 24397 8851 24455 8857
rect 24578 8848 24584 8860
rect 24636 8848 24642 8900
rect 4157 8823 4215 8829
rect 4157 8820 4169 8823
rect 2148 8792 4169 8820
rect 4157 8789 4169 8792
rect 4203 8820 4215 8823
rect 5368 8820 5396 8848
rect 9398 8820 9404 8832
rect 4203 8792 5396 8820
rect 9359 8792 9404 8820
rect 4203 8789 4215 8792
rect 4157 8783 4215 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 9861 8823 9919 8829
rect 9861 8820 9873 8823
rect 9732 8792 9873 8820
rect 9732 8780 9738 8792
rect 9861 8789 9873 8792
rect 9907 8789 9919 8823
rect 11606 8820 11612 8832
rect 11567 8792 11612 8820
rect 9861 8783 9919 8789
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 15381 8823 15439 8829
rect 12492 8792 12537 8820
rect 12492 8780 12498 8792
rect 15381 8789 15393 8823
rect 15427 8820 15439 8823
rect 16482 8820 16488 8832
rect 15427 8792 16488 8820
rect 15427 8789 15439 8792
rect 15381 8783 15439 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 17034 8820 17040 8832
rect 16995 8792 17040 8820
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 17586 8820 17592 8832
rect 17547 8792 17592 8820
rect 17586 8780 17592 8792
rect 17644 8780 17650 8832
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 19702 8820 19708 8832
rect 19484 8792 19708 8820
rect 19484 8780 19490 8792
rect 19702 8780 19708 8792
rect 19760 8780 19766 8832
rect 20162 8780 20168 8832
rect 20220 8820 20226 8832
rect 20349 8823 20407 8829
rect 20349 8820 20361 8823
rect 20220 8792 20361 8820
rect 20220 8780 20226 8792
rect 20349 8789 20361 8792
rect 20395 8789 20407 8823
rect 20349 8783 20407 8789
rect 22281 8823 22339 8829
rect 22281 8789 22293 8823
rect 22327 8820 22339 8823
rect 22370 8820 22376 8832
rect 22327 8792 22376 8820
rect 22327 8789 22339 8792
rect 22281 8783 22339 8789
rect 22370 8780 22376 8792
rect 22428 8780 22434 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 1946 8616 1952 8628
rect 1728 8588 1952 8616
rect 1728 8576 1734 8588
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 2406 8616 2412 8628
rect 2367 8588 2412 8616
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 2958 8616 2964 8628
rect 2915 8588 2964 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 4982 8616 4988 8628
rect 4943 8588 4988 8616
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6454 8616 6460 8628
rect 6319 8588 6460 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 8202 8616 8208 8628
rect 8163 8588 8208 8616
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 8996 8588 9505 8616
rect 8996 8576 9002 8588
rect 9493 8585 9505 8588
rect 9539 8616 9551 8619
rect 10134 8616 10140 8628
rect 9539 8588 10140 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10778 8576 10784 8628
rect 10836 8616 10842 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 10836 8588 10885 8616
rect 10836 8576 10842 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 11790 8616 11796 8628
rect 11751 8588 11796 8616
rect 10873 8579 10931 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12342 8616 12348 8628
rect 12299 8588 12348 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 1489 8551 1547 8557
rect 1489 8517 1501 8551
rect 1535 8548 1547 8551
rect 2130 8548 2136 8560
rect 1535 8520 2136 8548
rect 1535 8517 1547 8520
rect 1489 8511 1547 8517
rect 2130 8508 2136 8520
rect 2188 8508 2194 8560
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2976 8489 3004 8576
rect 4890 8508 4896 8560
rect 4948 8548 4954 8560
rect 6549 8551 6607 8557
rect 6549 8548 6561 8551
rect 4948 8520 6561 8548
rect 4948 8508 4954 8520
rect 6549 8517 6561 8520
rect 6595 8517 6607 8551
rect 6549 8511 6607 8517
rect 9861 8551 9919 8557
rect 9861 8517 9873 8551
rect 9907 8548 9919 8551
rect 9950 8548 9956 8560
rect 9907 8520 9956 8548
rect 9907 8517 9919 8520
rect 9861 8511 9919 8517
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 11698 8548 11704 8560
rect 11348 8520 11704 8548
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 5626 8480 5632 8492
rect 5408 8452 5632 8480
rect 5408 8440 5414 8452
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6178 8480 6184 8492
rect 5960 8452 6184 8480
rect 5960 8440 5966 8452
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 6638 8480 6644 8492
rect 6512 8452 6644 8480
rect 6512 8440 6518 8452
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 8570 8440 8576 8492
rect 8628 8480 8634 8492
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8628 8452 8769 8480
rect 8628 8440 8634 8452
rect 8757 8449 8769 8452
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8480 10379 8483
rect 11238 8480 11244 8492
rect 10367 8452 11244 8480
rect 10367 8449 10379 8452
rect 10321 8443 10379 8449
rect 11238 8440 11244 8452
rect 11296 8480 11302 8492
rect 11348 8489 11376 8520
rect 11698 8508 11704 8520
rect 11756 8508 11762 8560
rect 11333 8483 11391 8489
rect 11333 8480 11345 8483
rect 11296 8452 11345 8480
rect 11296 8440 11302 8452
rect 11333 8449 11345 8452
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 11425 8483 11483 8489
rect 11425 8449 11437 8483
rect 11471 8480 11483 8483
rect 12268 8480 12296 8579
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 15746 8616 15752 8628
rect 15707 8588 15752 8616
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 16114 8616 16120 8628
rect 16075 8588 16120 8616
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 19889 8619 19947 8625
rect 19889 8585 19901 8619
rect 19935 8616 19947 8619
rect 19978 8616 19984 8628
rect 19935 8588 19984 8616
rect 19935 8585 19947 8588
rect 19889 8579 19947 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 21358 8576 21364 8628
rect 21416 8616 21422 8628
rect 23477 8619 23535 8625
rect 21416 8588 21772 8616
rect 21416 8576 21422 8588
rect 12618 8548 12624 8560
rect 12579 8520 12624 8548
rect 12618 8508 12624 8520
rect 12676 8508 12682 8560
rect 16390 8548 16396 8560
rect 16351 8520 16396 8548
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 18138 8548 18144 8560
rect 18099 8520 18144 8548
rect 18138 8508 18144 8520
rect 18196 8508 18202 8560
rect 20073 8551 20131 8557
rect 20073 8517 20085 8551
rect 20119 8548 20131 8551
rect 20714 8548 20720 8560
rect 20119 8520 20720 8548
rect 20119 8517 20131 8520
rect 20073 8511 20131 8517
rect 20714 8508 20720 8520
rect 20772 8508 20778 8560
rect 21634 8548 21640 8560
rect 21595 8520 21640 8548
rect 21634 8508 21640 8520
rect 21692 8508 21698 8560
rect 21744 8548 21772 8588
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 23658 8616 23664 8628
rect 23523 8588 23664 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 24489 8619 24547 8625
rect 24489 8585 24501 8619
rect 24535 8616 24547 8619
rect 24670 8616 24676 8628
rect 24535 8588 24676 8616
rect 24535 8585 24547 8588
rect 24489 8579 24547 8585
rect 24504 8548 24532 8579
rect 24670 8576 24676 8588
rect 24728 8576 24734 8628
rect 24854 8616 24860 8628
rect 24815 8588 24860 8616
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 25130 8616 25136 8628
rect 25091 8588 25136 8616
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 21744 8520 24532 8548
rect 12710 8480 12716 8492
rect 11471 8452 12716 8480
rect 11471 8449 11483 8452
rect 11425 8443 11483 8449
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16356 8452 16957 8480
rect 16356 8440 16362 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 18693 8483 18751 8489
rect 18693 8480 18705 8483
rect 17451 8452 18705 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 18693 8449 18705 8452
rect 18739 8480 18751 8483
rect 18966 8480 18972 8492
rect 18739 8452 18972 8480
rect 18739 8449 18751 8452
rect 18693 8443 18751 8449
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8480 19579 8483
rect 20625 8483 20683 8489
rect 20625 8480 20637 8483
rect 19567 8452 20637 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 20625 8449 20637 8452
rect 20671 8480 20683 8483
rect 21174 8480 21180 8492
rect 20671 8452 21180 8480
rect 20671 8449 20683 8452
rect 20625 8443 20683 8449
rect 21174 8440 21180 8452
rect 21232 8440 21238 8492
rect 21453 8483 21511 8489
rect 21453 8449 21465 8483
rect 21499 8480 21511 8483
rect 22370 8480 22376 8492
rect 21499 8452 22376 8480
rect 21499 8449 21511 8452
rect 21453 8443 21511 8449
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 23934 8480 23940 8492
rect 23895 8452 23940 8480
rect 23934 8440 23940 8452
rect 23992 8440 23998 8492
rect 2498 8412 2504 8424
rect 1964 8384 2504 8412
rect 1964 8353 1992 8384
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 5261 8415 5319 8421
rect 5261 8412 5273 8415
rect 3068 8384 5273 8412
rect 1949 8347 2007 8353
rect 1949 8313 1961 8347
rect 1995 8313 2007 8347
rect 1949 8307 2007 8313
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8344 2099 8347
rect 2682 8344 2688 8356
rect 2087 8316 2688 8344
rect 2087 8313 2099 8316
rect 2041 8307 2099 8313
rect 2682 8304 2688 8316
rect 2740 8344 2746 8356
rect 3068 8344 3096 8384
rect 5261 8381 5273 8384
rect 5307 8381 5319 8415
rect 5442 8412 5448 8424
rect 5403 8384 5448 8412
rect 5261 8375 5319 8381
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6788 8384 6837 8412
rect 6788 8372 6794 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 8481 8415 8539 8421
rect 8481 8412 8493 8415
rect 7699 8384 8493 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 8481 8381 8493 8384
rect 8527 8412 8539 8415
rect 9674 8412 9680 8424
rect 8527 8384 9536 8412
rect 9635 8384 9680 8412
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 2740 8316 3096 8344
rect 2740 8304 2746 8316
rect 3142 8304 3148 8356
rect 3200 8353 3206 8356
rect 3200 8347 3264 8353
rect 3200 8313 3218 8347
rect 3252 8313 3264 8347
rect 5718 8344 5724 8356
rect 5679 8316 5724 8344
rect 3200 8307 3264 8313
rect 3200 8304 3206 8307
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 7098 8344 7104 8356
rect 7059 8316 7104 8344
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 8021 8347 8079 8353
rect 8021 8313 8033 8347
rect 8067 8344 8079 8347
rect 8386 8344 8392 8356
rect 8067 8316 8392 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 8662 8344 8668 8356
rect 8623 8316 8668 8344
rect 8662 8304 8668 8316
rect 8720 8344 8726 8356
rect 9125 8347 9183 8353
rect 9125 8344 9137 8347
rect 8720 8316 9137 8344
rect 8720 8304 8726 8316
rect 9125 8313 9137 8316
rect 9171 8344 9183 8347
rect 9306 8344 9312 8356
rect 9171 8316 9312 8344
rect 9171 8313 9183 8316
rect 9125 8307 9183 8313
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 9508 8344 9536 8384
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 10686 8412 10692 8424
rect 10599 8384 10692 8412
rect 10686 8372 10692 8384
rect 10744 8412 10750 8424
rect 10744 8384 11376 8412
rect 10744 8372 10750 8384
rect 9582 8344 9588 8356
rect 9508 8316 9588 8344
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 11348 8353 11376 8384
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 14090 8421 14096 8424
rect 13817 8415 13875 8421
rect 13817 8412 13829 8415
rect 12492 8384 12537 8412
rect 13648 8384 13829 8412
rect 12492 8372 12498 8384
rect 11333 8347 11391 8353
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 11882 8344 11888 8356
rect 11379 8316 11888 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 4341 8279 4399 8285
rect 4341 8245 4353 8279
rect 4387 8276 4399 8279
rect 4706 8276 4712 8288
rect 4387 8248 4712 8276
rect 4387 8245 4399 8248
rect 4341 8239 4399 8245
rect 4706 8236 4712 8248
rect 4764 8276 4770 8288
rect 5258 8276 5264 8288
rect 4764 8248 5264 8276
rect 4764 8236 4770 8248
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 9674 8236 9680 8288
rect 9732 8276 9738 8288
rect 9858 8276 9864 8288
rect 9732 8248 9864 8276
rect 9732 8236 9738 8248
rect 9858 8236 9864 8248
rect 9916 8276 9922 8288
rect 12158 8276 12164 8288
rect 9916 8248 12164 8276
rect 9916 8236 9922 8248
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 13081 8279 13139 8285
rect 13081 8245 13093 8279
rect 13127 8276 13139 8279
rect 13170 8276 13176 8288
rect 13127 8248 13176 8276
rect 13127 8245 13139 8248
rect 13081 8239 13139 8245
rect 13170 8236 13176 8248
rect 13228 8276 13234 8288
rect 13648 8285 13676 8384
rect 13817 8381 13829 8384
rect 13863 8381 13875 8415
rect 14084 8412 14096 8421
rect 14051 8384 14096 8412
rect 13817 8375 13875 8381
rect 14084 8375 14096 8384
rect 14090 8372 14096 8375
rect 14148 8372 14154 8424
rect 16114 8372 16120 8424
rect 16172 8412 16178 8424
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 16172 8384 16896 8412
rect 16172 8372 16178 8384
rect 16868 8353 16896 8384
rect 18616 8384 19073 8412
rect 18616 8356 18644 8384
rect 19061 8381 19073 8384
rect 19107 8381 19119 8415
rect 19061 8375 19119 8381
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 20349 8415 20407 8421
rect 20349 8412 20361 8415
rect 20036 8384 20361 8412
rect 20036 8372 20042 8384
rect 20349 8381 20361 8384
rect 20395 8381 20407 8415
rect 21910 8412 21916 8424
rect 21871 8384 21916 8412
rect 20349 8375 20407 8381
rect 21910 8372 21916 8384
rect 21968 8412 21974 8424
rect 22557 8415 22615 8421
rect 22557 8412 22569 8415
rect 21968 8384 22569 8412
rect 21968 8372 21974 8384
rect 22557 8381 22569 8384
rect 22603 8381 22615 8415
rect 22557 8375 22615 8381
rect 23474 8372 23480 8424
rect 23532 8412 23538 8424
rect 23661 8415 23719 8421
rect 23661 8412 23673 8415
rect 23532 8384 23673 8412
rect 23532 8372 23538 8384
rect 23661 8381 23673 8384
rect 23707 8381 23719 8415
rect 24946 8412 24952 8424
rect 24907 8384 24952 8412
rect 23661 8375 23719 8381
rect 24946 8372 24952 8384
rect 25004 8412 25010 8424
rect 25501 8415 25559 8421
rect 25501 8412 25513 8415
rect 25004 8384 25513 8412
rect 25004 8372 25010 8384
rect 25501 8381 25513 8384
rect 25547 8381 25559 8415
rect 25501 8375 25559 8381
rect 16669 8347 16727 8353
rect 16669 8344 16681 8347
rect 16500 8316 16681 8344
rect 13633 8279 13691 8285
rect 13633 8276 13645 8279
rect 13228 8248 13645 8276
rect 13228 8236 13234 8248
rect 13633 8245 13645 8248
rect 13679 8245 13691 8279
rect 13633 8239 13691 8245
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 15197 8279 15255 8285
rect 15197 8276 15209 8279
rect 13872 8248 15209 8276
rect 13872 8236 13878 8248
rect 15197 8245 15209 8248
rect 15243 8245 15255 8279
rect 15197 8239 15255 8245
rect 16298 8236 16304 8288
rect 16356 8276 16362 8288
rect 16500 8276 16528 8316
rect 16669 8313 16681 8316
rect 16715 8313 16727 8347
rect 16669 8307 16727 8313
rect 16853 8347 16911 8353
rect 16853 8313 16865 8347
rect 16899 8313 16911 8347
rect 16853 8307 16911 8313
rect 17586 8304 17592 8356
rect 17644 8344 17650 8356
rect 18417 8347 18475 8353
rect 18417 8344 18429 8347
rect 17644 8316 18429 8344
rect 17644 8304 17650 8316
rect 18417 8313 18429 8316
rect 18463 8313 18475 8347
rect 18598 8344 18604 8356
rect 18559 8316 18604 8344
rect 18417 8307 18475 8313
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 20438 8304 20444 8356
rect 20496 8344 20502 8356
rect 20533 8347 20591 8353
rect 20533 8344 20545 8347
rect 20496 8316 20545 8344
rect 20496 8304 20502 8316
rect 20533 8313 20545 8316
rect 20579 8313 20591 8347
rect 20533 8307 20591 8313
rect 22189 8347 22247 8353
rect 22189 8313 22201 8347
rect 22235 8344 22247 8347
rect 22370 8344 22376 8356
rect 22235 8316 22376 8344
rect 22235 8313 22247 8316
rect 22189 8307 22247 8313
rect 22370 8304 22376 8316
rect 22428 8304 22434 8356
rect 24210 8304 24216 8356
rect 24268 8344 24274 8356
rect 26786 8344 26792 8356
rect 24268 8316 26792 8344
rect 24268 8304 24274 8316
rect 26786 8304 26792 8316
rect 26844 8304 26850 8356
rect 16356 8248 16528 8276
rect 16356 8236 16362 8248
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 17681 8279 17739 8285
rect 17681 8276 17693 8279
rect 17460 8248 17693 8276
rect 17460 8236 17466 8248
rect 17681 8245 17693 8248
rect 17727 8245 17739 8279
rect 17681 8239 17739 8245
rect 20898 8236 20904 8288
rect 20956 8276 20962 8288
rect 20993 8279 21051 8285
rect 20993 8276 21005 8279
rect 20956 8248 21005 8276
rect 20956 8236 20962 8248
rect 20993 8245 21005 8248
rect 21039 8245 21051 8279
rect 20993 8239 21051 8245
rect 21542 8236 21548 8288
rect 21600 8276 21606 8288
rect 22097 8279 22155 8285
rect 22097 8276 22109 8279
rect 21600 8248 22109 8276
rect 21600 8236 21606 8248
rect 22097 8245 22109 8248
rect 22143 8245 22155 8279
rect 22097 8239 22155 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1397 8075 1455 8081
rect 1397 8041 1409 8075
rect 1443 8072 1455 8075
rect 1762 8072 1768 8084
rect 1443 8044 1768 8072
rect 1443 8041 1455 8044
rect 1397 8035 1455 8041
rect 1762 8032 1768 8044
rect 1820 8032 1826 8084
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 2222 8072 2228 8084
rect 2179 8044 2228 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2958 8072 2964 8084
rect 2919 8044 2964 8072
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 4617 8075 4675 8081
rect 4617 8072 4629 8075
rect 4488 8044 4629 8072
rect 4488 8032 4494 8044
rect 4617 8041 4629 8044
rect 4663 8041 4675 8075
rect 4617 8035 4675 8041
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 5408 8044 6316 8072
rect 5408 8032 5414 8044
rect 4522 7964 4528 8016
rect 4580 8004 4586 8016
rect 4709 8007 4767 8013
rect 4709 8004 4721 8007
rect 4580 7976 4721 8004
rect 4580 7964 4586 7976
rect 4709 7973 4721 7976
rect 4755 7973 4767 8007
rect 4709 7967 4767 7973
rect 5988 8007 6046 8013
rect 5988 7973 6000 8007
rect 6034 8004 6046 8007
rect 6178 8004 6184 8016
rect 6034 7976 6184 8004
rect 6034 7973 6046 7976
rect 5988 7967 6046 7973
rect 6178 7964 6184 7976
rect 6236 7964 6242 8016
rect 6288 8004 6316 8044
rect 6822 8032 6828 8084
rect 6880 8072 6886 8084
rect 7101 8075 7159 8081
rect 7101 8072 7113 8075
rect 6880 8044 7113 8072
rect 6880 8032 6886 8044
rect 7101 8041 7113 8044
rect 7147 8041 7159 8075
rect 7650 8072 7656 8084
rect 7611 8044 7656 8072
rect 7101 8035 7159 8041
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8202 8072 8208 8084
rect 8159 8044 8208 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8628 8044 8953 8072
rect 8628 8032 8634 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 10962 8032 10968 8084
rect 11020 8072 11026 8084
rect 11333 8075 11391 8081
rect 11333 8072 11345 8075
rect 11020 8044 11345 8072
rect 11020 8032 11026 8044
rect 11333 8041 11345 8044
rect 11379 8072 11391 8075
rect 11790 8072 11796 8084
rect 11379 8044 11796 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 12710 8072 12716 8084
rect 12671 8044 12716 8072
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13722 8072 13728 8084
rect 13679 8044 13728 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13872 8044 14105 8072
rect 13872 8032 13878 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14884 8044 15025 8072
rect 14884 8032 14890 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15838 8072 15844 8084
rect 15799 8044 15844 8072
rect 15013 8035 15071 8041
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 17405 8075 17463 8081
rect 17405 8041 17417 8075
rect 17451 8072 17463 8075
rect 18322 8072 18328 8084
rect 17451 8044 18328 8072
rect 17451 8041 17463 8044
rect 17405 8035 17463 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 18506 8072 18512 8084
rect 18467 8044 18512 8072
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 21542 8072 21548 8084
rect 20772 8044 21548 8072
rect 20772 8032 20778 8044
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 23658 8072 23664 8084
rect 23619 8044 23664 8072
rect 23658 8032 23664 8044
rect 23716 8032 23722 8084
rect 7006 8004 7012 8016
rect 6288 7976 7012 8004
rect 7006 7964 7012 7976
rect 7064 8004 7070 8016
rect 9309 8007 9367 8013
rect 9309 8004 9321 8007
rect 7064 7976 9321 8004
rect 7064 7964 7070 7976
rect 9309 7973 9321 7976
rect 9355 7973 9367 8007
rect 13446 8004 13452 8016
rect 13407 7976 13452 8004
rect 9309 7967 9367 7973
rect 13446 7964 13452 7976
rect 13504 7964 13510 8016
rect 15930 7964 15936 8016
rect 15988 8004 15994 8016
rect 15988 7976 16033 8004
rect 15988 7964 15994 7976
rect 17494 7964 17500 8016
rect 17552 8004 17558 8016
rect 18049 8007 18107 8013
rect 18049 8004 18061 8007
rect 17552 7976 18061 8004
rect 17552 7964 17558 7976
rect 18049 7973 18061 7976
rect 18095 7973 18107 8007
rect 18049 7967 18107 7973
rect 18141 8007 18199 8013
rect 18141 7973 18153 8007
rect 18187 8004 18199 8007
rect 18524 8004 18552 8032
rect 18187 7976 18552 8004
rect 18187 7973 18199 7976
rect 18141 7967 18199 7973
rect 19150 7964 19156 8016
rect 19208 8004 19214 8016
rect 19334 8004 19340 8016
rect 19208 7976 19340 8004
rect 19208 7964 19214 7976
rect 19334 7964 19340 7976
rect 19392 8004 19398 8016
rect 19429 8007 19487 8013
rect 19429 8004 19441 8007
rect 19392 7976 19441 8004
rect 19392 7964 19398 7976
rect 19429 7973 19441 7976
rect 19475 7973 19487 8007
rect 19429 7967 19487 7973
rect 19613 8007 19671 8013
rect 19613 7973 19625 8007
rect 19659 7973 19671 8007
rect 21174 8004 21180 8016
rect 21135 7976 21180 8004
rect 19613 7967 19671 7973
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 5684 7908 5733 7936
rect 5684 7896 5690 7908
rect 5721 7905 5733 7908
rect 5767 7936 5779 7939
rect 6362 7936 6368 7948
rect 5767 7908 6368 7936
rect 5767 7905 5779 7908
rect 5721 7899 5779 7905
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 8202 7936 8208 7948
rect 8163 7908 8208 7936
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8478 7936 8484 7948
rect 8439 7908 8484 7936
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 10220 7939 10278 7945
rect 10220 7905 10232 7939
rect 10266 7936 10278 7939
rect 11330 7936 11336 7948
rect 10266 7908 11336 7936
rect 10266 7905 10278 7908
rect 10220 7899 10278 7905
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 13725 7939 13783 7945
rect 13725 7905 13737 7939
rect 13771 7936 13783 7939
rect 14090 7936 14096 7948
rect 13771 7908 14096 7936
rect 13771 7905 13783 7908
rect 13725 7899 13783 7905
rect 14090 7896 14096 7908
rect 14148 7936 14154 7948
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 14148 7908 14473 7936
rect 14148 7896 14154 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 15654 7936 15660 7948
rect 15615 7908 15660 7936
rect 14461 7899 14519 7905
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 18230 7896 18236 7948
rect 18288 7936 18294 7948
rect 19628 7936 19656 7967
rect 21174 7964 21180 7976
rect 21232 7964 21238 8016
rect 21996 8007 22054 8013
rect 21996 7973 22008 8007
rect 22042 8004 22054 8007
rect 22370 8004 22376 8016
rect 22042 7976 22376 8004
rect 22042 7973 22054 7976
rect 21996 7967 22054 7973
rect 22370 7964 22376 7976
rect 22428 7964 22434 8016
rect 23842 7964 23848 8016
rect 23900 8004 23906 8016
rect 24581 8007 24639 8013
rect 24581 8004 24593 8007
rect 23900 7976 24593 8004
rect 23900 7964 23906 7976
rect 24581 7973 24593 7976
rect 24627 7973 24639 8007
rect 24581 7967 24639 7973
rect 18288 7908 19656 7936
rect 18288 7896 18294 7908
rect 21542 7896 21548 7948
rect 21600 7936 21606 7948
rect 23566 7936 23572 7948
rect 21600 7908 23572 7936
rect 21600 7896 21606 7908
rect 23566 7896 23572 7908
rect 23624 7896 23630 7948
rect 24118 7896 24124 7948
rect 24176 7936 24182 7948
rect 24305 7939 24363 7945
rect 24305 7936 24317 7939
rect 24176 7908 24317 7936
rect 24176 7896 24182 7908
rect 24305 7905 24317 7908
rect 24351 7905 24363 7939
rect 24305 7899 24363 7905
rect 2958 7868 2964 7880
rect 2919 7840 2964 7868
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3142 7868 3148 7880
rect 3099 7840 3148 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 4614 7868 4620 7880
rect 4575 7840 4620 7868
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7837 10011 7871
rect 9953 7831 10011 7837
rect 1854 7760 1860 7812
rect 1912 7800 1918 7812
rect 2590 7800 2596 7812
rect 1912 7772 2596 7800
rect 1912 7760 1918 7772
rect 2590 7760 2596 7772
rect 2648 7760 2654 7812
rect 4157 7803 4215 7809
rect 4157 7769 4169 7803
rect 4203 7800 4215 7803
rect 4890 7800 4896 7812
rect 4203 7772 4896 7800
rect 4203 7769 4215 7772
rect 4157 7763 4215 7769
rect 4890 7760 4896 7772
rect 4948 7760 4954 7812
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 2501 7735 2559 7741
rect 2501 7732 2513 7735
rect 2372 7704 2513 7732
rect 2372 7692 2378 7704
rect 2501 7701 2513 7704
rect 2547 7701 2559 7735
rect 2501 7695 2559 7701
rect 3697 7735 3755 7741
rect 3697 7701 3709 7735
rect 3743 7732 3755 7735
rect 3786 7732 3792 7744
rect 3743 7704 3792 7732
rect 3743 7701 3755 7704
rect 3697 7695 3755 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 5169 7735 5227 7741
rect 5169 7732 5181 7735
rect 4304 7704 5181 7732
rect 4304 7692 4310 7704
rect 5169 7701 5181 7704
rect 5215 7732 5227 7735
rect 5445 7735 5503 7741
rect 5445 7732 5457 7735
rect 5215 7704 5457 7732
rect 5215 7701 5227 7704
rect 5169 7695 5227 7701
rect 5445 7701 5457 7704
rect 5491 7701 5503 7735
rect 5445 7695 5503 7701
rect 9030 7692 9036 7744
rect 9088 7732 9094 7744
rect 9858 7732 9864 7744
rect 9088 7704 9864 7732
rect 9088 7692 9094 7704
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 9968 7732 9996 7831
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 15672 7868 15700 7896
rect 16298 7868 16304 7880
rect 11204 7840 15700 7868
rect 16259 7840 16304 7868
rect 11204 7828 11210 7840
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 17954 7868 17960 7880
rect 17915 7840 17960 7868
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 19705 7871 19763 7877
rect 19705 7868 19717 7871
rect 19536 7840 19717 7868
rect 13173 7803 13231 7809
rect 13173 7769 13185 7803
rect 13219 7800 13231 7803
rect 13538 7800 13544 7812
rect 13219 7772 13544 7800
rect 13219 7769 13231 7772
rect 13173 7763 13231 7769
rect 13538 7760 13544 7772
rect 13596 7760 13602 7812
rect 15378 7800 15384 7812
rect 15339 7772 15384 7800
rect 15378 7760 15384 7772
rect 15436 7760 15442 7812
rect 17586 7800 17592 7812
rect 17547 7772 17592 7800
rect 17586 7760 17592 7772
rect 17644 7760 17650 7812
rect 18969 7803 19027 7809
rect 18969 7769 18981 7803
rect 19015 7800 19027 7803
rect 19536 7800 19564 7840
rect 19705 7837 19717 7840
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 20898 7800 20904 7812
rect 19015 7772 19564 7800
rect 19015 7769 19027 7772
rect 18969 7763 19027 7769
rect 19536 7744 19564 7772
rect 20088 7772 20904 7800
rect 10134 7732 10140 7744
rect 9968 7704 10140 7732
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 11238 7692 11244 7744
rect 11296 7732 11302 7744
rect 11885 7735 11943 7741
rect 11885 7732 11897 7735
rect 11296 7704 11897 7732
rect 11296 7692 11302 7704
rect 11885 7701 11897 7704
rect 11931 7701 11943 7735
rect 12250 7732 12256 7744
rect 12211 7704 12256 7732
rect 11885 7695 11943 7701
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 16666 7732 16672 7744
rect 16627 7704 16672 7732
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 19150 7732 19156 7744
rect 19111 7704 19156 7732
rect 19150 7692 19156 7704
rect 19208 7692 19214 7744
rect 19518 7692 19524 7744
rect 19576 7692 19582 7744
rect 19886 7692 19892 7744
rect 19944 7732 19950 7744
rect 20088 7741 20116 7772
rect 20898 7760 20904 7772
rect 20956 7800 20962 7812
rect 21744 7800 21772 7831
rect 22738 7828 22744 7880
rect 22796 7868 22802 7880
rect 23106 7868 23112 7880
rect 22796 7840 23112 7868
rect 22796 7828 22802 7840
rect 23106 7828 23112 7840
rect 23164 7828 23170 7880
rect 20956 7772 21772 7800
rect 20956 7760 20962 7772
rect 20073 7735 20131 7741
rect 20073 7732 20085 7735
rect 19944 7704 20085 7732
rect 19944 7692 19950 7704
rect 20073 7701 20085 7704
rect 20119 7701 20131 7735
rect 20438 7732 20444 7744
rect 20399 7704 20444 7732
rect 20073 7695 20131 7701
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 23106 7732 23112 7744
rect 23067 7704 23112 7732
rect 23106 7692 23112 7704
rect 23164 7692 23170 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 2866 7528 2872 7540
rect 2179 7500 2872 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 3694 7528 3700 7540
rect 3655 7500 3700 7528
rect 3694 7488 3700 7500
rect 3752 7488 3758 7540
rect 4614 7528 4620 7540
rect 4575 7500 4620 7528
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 5261 7531 5319 7537
rect 5261 7497 5273 7531
rect 5307 7528 5319 7531
rect 5442 7528 5448 7540
rect 5307 7500 5448 7528
rect 5307 7497 5319 7500
rect 5261 7491 5319 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 6273 7531 6331 7537
rect 6273 7497 6285 7531
rect 6319 7528 6331 7531
rect 6362 7528 6368 7540
rect 6319 7500 6368 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 6362 7488 6368 7500
rect 6420 7528 6426 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 6420 7500 7665 7528
rect 6420 7488 6426 7500
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 3421 7463 3479 7469
rect 3421 7429 3433 7463
rect 3467 7460 3479 7463
rect 4430 7460 4436 7472
rect 3467 7432 4436 7460
rect 3467 7429 3479 7432
rect 3421 7423 3479 7429
rect 4430 7420 4436 7432
rect 4488 7420 4494 7472
rect 4522 7420 4528 7472
rect 4580 7460 4586 7472
rect 4985 7463 5043 7469
rect 4985 7460 4997 7463
rect 4580 7432 4997 7460
rect 4580 7420 4586 7432
rect 4985 7429 4997 7432
rect 5031 7429 5043 7463
rect 4985 7423 5043 7429
rect 2222 7352 2228 7404
rect 2280 7392 2286 7404
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 2280 7364 2513 7392
rect 2280 7352 2286 7364
rect 2501 7361 2513 7364
rect 2547 7361 2559 7395
rect 2501 7355 2559 7361
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7392 2743 7395
rect 3510 7392 3516 7404
rect 2731 7364 3516 7392
rect 2731 7361 2743 7364
rect 2685 7355 2743 7361
rect 3510 7352 3516 7364
rect 3568 7392 3574 7404
rect 4246 7392 4252 7404
rect 3568 7364 4252 7392
rect 3568 7352 3574 7364
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 5500 7364 5733 7392
rect 5500 7352 5506 7364
rect 5721 7361 5733 7364
rect 5767 7392 5779 7395
rect 6270 7392 6276 7404
rect 5767 7364 6276 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 7558 7352 7564 7404
rect 7616 7392 7622 7404
rect 7668 7392 7696 7491
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 9548 7500 10425 7528
rect 9548 7488 9554 7500
rect 10413 7497 10425 7500
rect 10459 7497 10471 7531
rect 10413 7491 10471 7497
rect 12894 7488 12900 7540
rect 12952 7528 12958 7540
rect 12989 7531 13047 7537
rect 12989 7528 13001 7531
rect 12952 7500 13001 7528
rect 12952 7488 12958 7500
rect 12989 7497 13001 7500
rect 13035 7497 13047 7531
rect 12989 7491 13047 7497
rect 15565 7531 15623 7537
rect 15565 7497 15577 7531
rect 15611 7528 15623 7531
rect 15838 7528 15844 7540
rect 15611 7500 15844 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 16114 7528 16120 7540
rect 16075 7500 16120 7528
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 17494 7528 17500 7540
rect 17455 7500 17500 7528
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 18230 7488 18236 7540
rect 18288 7528 18294 7540
rect 18693 7531 18751 7537
rect 18693 7528 18705 7531
rect 18288 7500 18705 7528
rect 18288 7488 18294 7500
rect 18693 7497 18705 7500
rect 18739 7497 18751 7531
rect 18693 7491 18751 7497
rect 20898 7488 20904 7540
rect 20956 7528 20962 7540
rect 21453 7531 21511 7537
rect 21453 7528 21465 7531
rect 20956 7500 21465 7528
rect 20956 7488 20962 7500
rect 21453 7497 21465 7500
rect 21499 7497 21511 7531
rect 21453 7491 21511 7497
rect 21913 7531 21971 7537
rect 21913 7497 21925 7531
rect 21959 7528 21971 7531
rect 22278 7528 22284 7540
rect 21959 7500 22284 7528
rect 21959 7497 21971 7500
rect 21913 7491 21971 7497
rect 12621 7463 12679 7469
rect 12621 7460 12633 7463
rect 10235 7432 12633 7460
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 7616 7364 7849 7392
rect 7616 7352 7622 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 10235 7392 10263 7432
rect 12621 7429 12633 7432
rect 12667 7429 12679 7463
rect 12621 7423 12679 7429
rect 9824 7364 10263 7392
rect 9824 7352 9830 7364
rect 10778 7352 10784 7404
rect 10836 7392 10842 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 10836 7364 10885 7392
rect 10836 7352 10842 7364
rect 10873 7361 10885 7364
rect 10919 7392 10931 7395
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 10919 7364 12081 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 5813 7327 5871 7333
rect 1995 7296 2636 7324
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 2608 7268 2636 7296
rect 5813 7293 5825 7327
rect 5859 7324 5871 7327
rect 6638 7324 6644 7336
rect 5859 7296 6644 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 6638 7284 6644 7296
rect 6696 7324 6702 7336
rect 6822 7324 6828 7336
rect 6696 7296 6828 7324
rect 6696 7284 6702 7296
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 10962 7324 10968 7336
rect 10923 7296 10968 7324
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 12894 7324 12900 7336
rect 12483 7296 12900 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 13170 7284 13176 7336
rect 13228 7324 13234 7336
rect 13814 7333 13820 7336
rect 13541 7327 13599 7333
rect 13541 7324 13553 7327
rect 13228 7296 13553 7324
rect 13228 7284 13234 7296
rect 13541 7293 13553 7296
rect 13587 7293 13599 7327
rect 13808 7324 13820 7333
rect 13775 7296 13820 7324
rect 13541 7287 13599 7293
rect 13808 7287 13820 7296
rect 2590 7256 2596 7268
rect 2551 7228 2596 7256
rect 2590 7216 2596 7228
rect 2648 7216 2654 7268
rect 3602 7216 3608 7268
rect 3660 7256 3666 7268
rect 3786 7256 3792 7268
rect 3660 7228 3792 7256
rect 3660 7216 3666 7228
rect 3786 7216 3792 7228
rect 3844 7256 3850 7268
rect 3973 7259 4031 7265
rect 3973 7256 3985 7259
rect 3844 7228 3985 7256
rect 3844 7216 3850 7228
rect 3973 7225 3985 7228
rect 4019 7225 4031 7259
rect 3973 7219 4031 7225
rect 5350 7216 5356 7268
rect 5408 7256 5414 7268
rect 5721 7259 5779 7265
rect 5721 7256 5733 7259
rect 5408 7228 5733 7256
rect 5408 7216 5414 7228
rect 5721 7225 5733 7228
rect 5767 7256 5779 7259
rect 6086 7256 6092 7268
rect 5767 7228 6092 7256
rect 5767 7225 5779 7228
rect 5721 7219 5779 7225
rect 6086 7216 6092 7228
rect 6144 7216 6150 7268
rect 7377 7259 7435 7265
rect 7377 7225 7389 7259
rect 7423 7256 7435 7259
rect 8018 7256 8024 7268
rect 7423 7228 8024 7256
rect 7423 7225 7435 7228
rect 7377 7219 7435 7225
rect 8018 7216 8024 7228
rect 8076 7265 8082 7268
rect 8076 7259 8140 7265
rect 8076 7225 8094 7259
rect 8128 7225 8140 7259
rect 11701 7259 11759 7265
rect 11701 7256 11713 7259
rect 8076 7219 8140 7225
rect 11072 7228 11713 7256
rect 8076 7216 8082 7219
rect 3050 7188 3056 7200
rect 3011 7160 3056 7188
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 4154 7188 4160 7200
rect 4115 7160 4160 7188
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6420 7160 6561 7188
rect 6420 7148 6426 7160
rect 6549 7157 6561 7160
rect 6595 7157 6607 7191
rect 6822 7188 6828 7200
rect 6783 7160 6828 7188
rect 6549 7151 6607 7157
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 9214 7188 9220 7200
rect 9175 7160 9220 7188
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 10045 7191 10103 7197
rect 10045 7157 10057 7191
rect 10091 7188 10103 7191
rect 10134 7188 10140 7200
rect 10091 7160 10140 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 10870 7188 10876 7200
rect 10831 7160 10876 7188
rect 10870 7148 10876 7160
rect 10928 7188 10934 7200
rect 11072 7188 11100 7228
rect 11701 7225 11713 7228
rect 11747 7225 11759 7259
rect 11701 7219 11759 7225
rect 11330 7188 11336 7200
rect 10928 7160 11100 7188
rect 11291 7160 11336 7188
rect 10928 7148 10934 7160
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 13449 7191 13507 7197
rect 13449 7157 13461 7191
rect 13495 7188 13507 7191
rect 13556 7188 13584 7287
rect 13814 7284 13820 7287
rect 13872 7284 13878 7336
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 16393 7327 16451 7333
rect 16393 7324 16405 7327
rect 14700 7296 16405 7324
rect 14700 7284 14706 7296
rect 16393 7293 16405 7296
rect 16439 7324 16451 7327
rect 17037 7327 17095 7333
rect 17037 7324 17049 7327
rect 16439 7296 17049 7324
rect 16439 7293 16451 7296
rect 16393 7287 16451 7293
rect 17037 7293 17049 7296
rect 17083 7293 17095 7327
rect 17037 7287 17095 7293
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7324 18107 7327
rect 18322 7324 18328 7336
rect 18095 7296 18328 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 19245 7327 19303 7333
rect 19245 7324 19257 7327
rect 18932 7296 19257 7324
rect 18932 7284 18938 7296
rect 19245 7293 19257 7296
rect 19291 7324 19303 7327
rect 19886 7324 19892 7336
rect 19291 7296 19892 7324
rect 19291 7293 19303 7296
rect 19245 7287 19303 7293
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 21468 7324 21496 7491
rect 22278 7488 22284 7500
rect 22336 7528 22342 7540
rect 23014 7528 23020 7540
rect 22336 7500 23020 7528
rect 22336 7488 22342 7500
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 24118 7488 24124 7540
rect 24176 7528 24182 7540
rect 24673 7531 24731 7537
rect 24673 7528 24685 7531
rect 24176 7500 24685 7528
rect 24176 7488 24182 7500
rect 24673 7497 24685 7500
rect 24719 7497 24731 7531
rect 25406 7528 25412 7540
rect 25367 7500 25412 7528
rect 24673 7491 24731 7497
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 22097 7463 22155 7469
rect 22097 7429 22109 7463
rect 22143 7460 22155 7463
rect 22554 7460 22560 7472
rect 22143 7432 22560 7460
rect 22143 7429 22155 7432
rect 22097 7423 22155 7429
rect 22554 7420 22560 7432
rect 22612 7420 22618 7472
rect 23753 7463 23811 7469
rect 23753 7429 23765 7463
rect 23799 7460 23811 7463
rect 23842 7460 23848 7472
rect 23799 7432 23848 7460
rect 23799 7429 23811 7432
rect 23753 7423 23811 7429
rect 23842 7420 23848 7432
rect 23900 7420 23906 7472
rect 22646 7352 22652 7404
rect 22704 7352 22710 7404
rect 23106 7352 23112 7404
rect 23164 7392 23170 7404
rect 24305 7395 24363 7401
rect 24305 7392 24317 7395
rect 23164 7364 24317 7392
rect 23164 7352 23170 7364
rect 24305 7361 24317 7364
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 22094 7324 22100 7336
rect 21468 7296 22100 7324
rect 22094 7284 22100 7296
rect 22152 7284 22158 7336
rect 22278 7284 22284 7336
rect 22336 7324 22342 7336
rect 22373 7327 22431 7333
rect 22373 7324 22385 7327
rect 22336 7296 22385 7324
rect 22336 7284 22342 7296
rect 22373 7293 22385 7296
rect 22419 7293 22431 7327
rect 22664 7324 22692 7352
rect 22373 7287 22431 7293
rect 22572 7296 22692 7324
rect 16666 7256 16672 7268
rect 16627 7228 16672 7256
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 19153 7259 19211 7265
rect 19153 7225 19165 7259
rect 19199 7256 19211 7259
rect 19334 7256 19340 7268
rect 19199 7228 19340 7256
rect 19199 7225 19211 7228
rect 19153 7219 19211 7225
rect 19334 7216 19340 7228
rect 19392 7216 19398 7268
rect 19518 7265 19524 7268
rect 19512 7256 19524 7265
rect 19479 7228 19524 7256
rect 19512 7219 19524 7228
rect 19518 7216 19524 7219
rect 19576 7216 19582 7268
rect 22572 7265 22600 7296
rect 23658 7284 23664 7336
rect 23716 7324 23722 7336
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 23716 7296 24041 7324
rect 23716 7284 23722 7296
rect 24029 7293 24041 7296
rect 24075 7293 24087 7327
rect 24029 7287 24087 7293
rect 25225 7327 25283 7333
rect 25225 7293 25237 7327
rect 25271 7293 25283 7327
rect 25225 7287 25283 7293
rect 22557 7259 22615 7265
rect 22557 7225 22569 7259
rect 22603 7225 22615 7259
rect 22557 7219 22615 7225
rect 22649 7259 22707 7265
rect 22649 7225 22661 7259
rect 22695 7225 22707 7259
rect 23474 7256 23480 7268
rect 23435 7228 23480 7256
rect 22649 7219 22707 7225
rect 13814 7188 13820 7200
rect 13495 7160 13820 7188
rect 13495 7157 13507 7160
rect 13449 7151 13507 7157
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 14642 7148 14648 7200
rect 14700 7188 14706 7200
rect 14921 7191 14979 7197
rect 14921 7188 14933 7191
rect 14700 7160 14933 7188
rect 14700 7148 14706 7160
rect 14921 7157 14933 7160
rect 14967 7157 14979 7191
rect 14921 7151 14979 7157
rect 15933 7191 15991 7197
rect 15933 7157 15945 7191
rect 15979 7188 15991 7191
rect 16298 7188 16304 7200
rect 15979 7160 16304 7188
rect 15979 7157 15991 7160
rect 15933 7151 15991 7157
rect 16298 7148 16304 7160
rect 16356 7188 16362 7200
rect 16577 7191 16635 7197
rect 16577 7188 16589 7191
rect 16356 7160 16589 7188
rect 16356 7148 16362 7160
rect 16577 7157 16589 7160
rect 16623 7188 16635 7191
rect 16758 7188 16764 7200
rect 16623 7160 16764 7188
rect 16623 7157 16635 7160
rect 16577 7151 16635 7157
rect 16758 7148 16764 7160
rect 16816 7148 16822 7200
rect 18233 7191 18291 7197
rect 18233 7157 18245 7191
rect 18279 7188 18291 7191
rect 18322 7188 18328 7200
rect 18279 7160 18328 7188
rect 18279 7157 18291 7160
rect 18233 7151 18291 7157
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 20254 7148 20260 7200
rect 20312 7188 20318 7200
rect 20622 7188 20628 7200
rect 20312 7160 20628 7188
rect 20312 7148 20318 7160
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 22186 7148 22192 7200
rect 22244 7188 22250 7200
rect 22664 7188 22692 7219
rect 23474 7216 23480 7228
rect 23532 7216 23538 7268
rect 25240 7256 25268 7287
rect 25777 7259 25835 7265
rect 25777 7256 25789 7259
rect 25240 7228 25789 7256
rect 23017 7191 23075 7197
rect 23017 7188 23029 7191
rect 22244 7160 23029 7188
rect 22244 7148 22250 7160
rect 23017 7157 23029 7160
rect 23063 7188 23075 7191
rect 23106 7188 23112 7200
rect 23063 7160 23112 7188
rect 23063 7157 23075 7160
rect 23017 7151 23075 7157
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 23492 7188 23520 7216
rect 24213 7191 24271 7197
rect 24213 7188 24225 7191
rect 23492 7160 24225 7188
rect 24213 7157 24225 7160
rect 24259 7188 24271 7191
rect 25240 7188 25268 7228
rect 25777 7225 25789 7228
rect 25823 7225 25835 7259
rect 25777 7219 25835 7225
rect 24259 7160 25268 7188
rect 24259 7157 24271 7160
rect 24213 7151 24271 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 6270 6984 6276 6996
rect 6231 6956 6276 6984
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 6638 6984 6644 6996
rect 6599 6956 6644 6984
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 7926 6984 7932 6996
rect 7887 6956 7932 6984
rect 7926 6944 7932 6956
rect 7984 6944 7990 6996
rect 10413 6987 10471 6993
rect 10413 6953 10425 6987
rect 10459 6984 10471 6987
rect 10962 6984 10968 6996
rect 10459 6956 10968 6984
rect 10459 6953 10471 6956
rect 10413 6947 10471 6953
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 13173 6987 13231 6993
rect 13173 6953 13185 6987
rect 13219 6984 13231 6987
rect 13446 6984 13452 6996
rect 13219 6956 13452 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 13541 6987 13599 6993
rect 13541 6953 13553 6987
rect 13587 6984 13599 6987
rect 14090 6984 14096 6996
rect 13587 6956 14096 6984
rect 13587 6953 13599 6956
rect 13541 6947 13599 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 15565 6987 15623 6993
rect 15565 6953 15577 6987
rect 15611 6984 15623 6987
rect 15654 6984 15660 6996
rect 15611 6956 15660 6984
rect 15611 6953 15623 6956
rect 15565 6947 15623 6953
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 18233 6987 18291 6993
rect 18233 6953 18245 6987
rect 18279 6984 18291 6987
rect 18506 6984 18512 6996
rect 18279 6956 18512 6984
rect 18279 6953 18291 6956
rect 18233 6947 18291 6953
rect 18506 6944 18512 6956
rect 18564 6944 18570 6996
rect 22097 6987 22155 6993
rect 22097 6953 22109 6987
rect 22143 6984 22155 6987
rect 22646 6984 22652 6996
rect 22143 6956 22652 6984
rect 22143 6953 22155 6956
rect 22097 6947 22155 6953
rect 22646 6944 22652 6956
rect 22704 6944 22710 6996
rect 4516 6919 4574 6925
rect 4516 6885 4528 6919
rect 4562 6916 4574 6919
rect 4706 6916 4712 6928
rect 4562 6888 4712 6916
rect 4562 6885 4574 6888
rect 4516 6879 4574 6885
rect 4706 6876 4712 6888
rect 4764 6876 4770 6928
rect 10686 6916 10692 6928
rect 8220 6888 10692 6916
rect 1762 6857 1768 6860
rect 1756 6848 1768 6857
rect 1723 6820 1768 6848
rect 1756 6811 1768 6820
rect 1762 6808 1768 6811
rect 1820 6808 1826 6860
rect 3697 6851 3755 6857
rect 3697 6817 3709 6851
rect 3743 6848 3755 6851
rect 4154 6848 4160 6860
rect 3743 6820 4160 6848
rect 3743 6817 3755 6820
rect 3697 6811 3755 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 6914 6848 6920 6860
rect 4304 6820 4349 6848
rect 6875 6820 6920 6848
rect 4304 6808 4310 6820
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7190 6808 7196 6860
rect 7248 6848 7254 6860
rect 8220 6848 8248 6888
rect 10686 6876 10692 6888
rect 10744 6876 10750 6928
rect 14185 6919 14243 6925
rect 14185 6916 14197 6919
rect 13556 6888 14197 6916
rect 13556 6860 13584 6888
rect 14185 6885 14197 6888
rect 14231 6885 14243 6919
rect 17402 6916 17408 6928
rect 14185 6879 14243 6885
rect 15856 6888 17408 6916
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 7248 6820 8248 6848
rect 9416 6820 9689 6848
rect 7248 6808 7254 6820
rect 1486 6780 1492 6792
rect 1447 6752 1492 6780
rect 1486 6740 1492 6752
rect 1544 6740 1550 6792
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8018 6780 8024 6792
rect 7979 6752 8024 6780
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 5626 6712 5632 6724
rect 5587 6684 5632 6712
rect 5626 6672 5632 6684
rect 5684 6712 5690 6724
rect 5994 6712 6000 6724
rect 5684 6684 6000 6712
rect 5684 6672 5690 6684
rect 5994 6672 6000 6684
rect 6052 6672 6058 6724
rect 7466 6712 7472 6724
rect 7427 6684 7472 6712
rect 7466 6672 7472 6684
rect 7524 6672 7530 6724
rect 8846 6712 8852 6724
rect 7576 6684 8852 6712
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 2869 6647 2927 6653
rect 2869 6644 2881 6647
rect 2740 6616 2881 6644
rect 2740 6604 2746 6616
rect 2869 6613 2881 6616
rect 2915 6613 2927 6647
rect 2869 6607 2927 6613
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 7576 6644 7604 6684
rect 8846 6672 8852 6684
rect 8904 6672 8910 6724
rect 8386 6644 8392 6656
rect 3476 6616 7604 6644
rect 8347 6616 8392 6644
rect 3476 6604 3482 6616
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8754 6644 8760 6656
rect 8715 6616 8760 6644
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 9416 6653 9444 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11221 6851 11279 6857
rect 11221 6848 11233 6851
rect 11112 6820 11233 6848
rect 11112 6808 11118 6820
rect 11221 6817 11233 6820
rect 11267 6817 11279 6851
rect 11221 6811 11279 6817
rect 13538 6808 13544 6860
rect 13596 6808 13602 6860
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 14056 6820 14289 6848
rect 14056 6808 14062 6820
rect 14277 6817 14289 6820
rect 14323 6848 14335 6851
rect 14642 6848 14648 6860
rect 14323 6820 14648 6848
rect 14323 6817 14335 6820
rect 14277 6811 14335 6817
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 14734 6808 14740 6860
rect 14792 6848 14798 6860
rect 15013 6851 15071 6857
rect 15013 6848 15025 6851
rect 14792 6820 15025 6848
rect 14792 6808 14798 6820
rect 15013 6817 15025 6820
rect 15059 6817 15071 6851
rect 15013 6811 15071 6817
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9364 6616 9413 6644
rect 9364 6604 9370 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9858 6644 9864 6656
rect 9819 6616 9864 6644
rect 9401 6607 9459 6613
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 10686 6644 10692 6656
rect 10647 6616 10692 6644
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 10980 6644 11008 6743
rect 12802 6740 12808 6792
rect 12860 6780 12866 6792
rect 13630 6780 13636 6792
rect 12860 6752 13636 6780
rect 12860 6740 12866 6752
rect 13630 6740 13636 6752
rect 13688 6780 13694 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13688 6752 14105 6780
rect 13688 6740 13694 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 15562 6740 15568 6792
rect 15620 6780 15626 6792
rect 15856 6789 15884 6888
rect 17402 6876 17408 6888
rect 17460 6876 17466 6928
rect 19058 6876 19064 6928
rect 19116 6916 19122 6928
rect 19610 6916 19616 6928
rect 19116 6888 19616 6916
rect 19116 6876 19122 6888
rect 19610 6876 19616 6888
rect 19668 6916 19674 6928
rect 19797 6919 19855 6925
rect 19797 6916 19809 6919
rect 19668 6888 19809 6916
rect 19668 6876 19674 6888
rect 19797 6885 19809 6888
rect 19843 6916 19855 6919
rect 20070 6916 20076 6928
rect 19843 6888 20076 6916
rect 19843 6885 19855 6888
rect 19797 6879 19855 6885
rect 20070 6876 20076 6888
rect 20128 6876 20134 6928
rect 23842 6916 23848 6928
rect 23400 6888 23848 6916
rect 23400 6860 23428 6888
rect 23842 6876 23848 6888
rect 23900 6876 23906 6928
rect 16114 6857 16120 6860
rect 16108 6848 16120 6857
rect 16075 6820 16120 6848
rect 16108 6811 16120 6820
rect 16172 6848 16178 6860
rect 16666 6848 16672 6860
rect 16172 6820 16672 6848
rect 16114 6808 16120 6811
rect 16172 6808 16178 6820
rect 16666 6808 16672 6820
rect 16724 6808 16730 6860
rect 17862 6848 17868 6860
rect 17823 6820 17868 6848
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 18785 6851 18843 6857
rect 18785 6817 18797 6851
rect 18831 6848 18843 6851
rect 19153 6851 19211 6857
rect 19153 6848 19165 6851
rect 18831 6820 19165 6848
rect 18831 6817 18843 6820
rect 18785 6811 18843 6817
rect 19153 6817 19165 6820
rect 19199 6848 19211 6851
rect 19518 6848 19524 6860
rect 19199 6820 19524 6848
rect 19199 6817 19211 6820
rect 19153 6811 19211 6817
rect 19518 6808 19524 6820
rect 19576 6848 19582 6860
rect 20714 6848 20720 6860
rect 19576 6820 19932 6848
rect 20675 6820 20720 6848
rect 19576 6808 19582 6820
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15620 6752 15853 6780
rect 15620 6740 15626 6752
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19904 6789 19932 6820
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 20901 6851 20959 6857
rect 20901 6817 20913 6851
rect 20947 6848 20959 6851
rect 21174 6848 21180 6860
rect 20947 6820 21180 6848
rect 20947 6817 20959 6820
rect 20901 6811 20959 6817
rect 21174 6808 21180 6820
rect 21232 6808 21238 6860
rect 22370 6848 22376 6860
rect 22331 6820 22376 6848
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 22905 6851 22963 6857
rect 22905 6848 22917 6851
rect 22572 6820 22917 6848
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 19392 6752 19717 6780
rect 19392 6740 19398 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 19889 6783 19947 6789
rect 19889 6749 19901 6783
rect 19935 6780 19947 6783
rect 21729 6783 21787 6789
rect 19935 6752 20852 6780
rect 19935 6749 19947 6752
rect 19889 6743 19947 6749
rect 13722 6712 13728 6724
rect 13683 6684 13728 6712
rect 13722 6672 13728 6684
rect 13780 6672 13786 6724
rect 13814 6672 13820 6724
rect 13872 6712 13878 6724
rect 19720 6712 19748 6743
rect 20070 6712 20076 6724
rect 13872 6684 14136 6712
rect 19720 6684 20076 6712
rect 13872 6672 13878 6684
rect 14108 6656 14136 6684
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 20824 6656 20852 6752
rect 21729 6749 21741 6783
rect 21775 6780 21787 6783
rect 22186 6780 22192 6792
rect 21775 6752 22192 6780
rect 21775 6749 21787 6752
rect 21729 6743 21787 6749
rect 22186 6740 22192 6752
rect 22244 6780 22250 6792
rect 22572 6780 22600 6820
rect 22905 6817 22917 6820
rect 22951 6817 22963 6851
rect 22905 6811 22963 6817
rect 23382 6808 23388 6860
rect 23440 6808 23446 6860
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6848 25191 6851
rect 25590 6848 25596 6860
rect 25179 6820 25596 6848
rect 25179 6817 25191 6820
rect 25133 6811 25191 6817
rect 25590 6808 25596 6820
rect 25648 6808 25654 6860
rect 22244 6752 22600 6780
rect 22244 6740 22250 6752
rect 22646 6740 22652 6792
rect 22704 6789 22710 6792
rect 22704 6780 22714 6789
rect 22704 6752 22749 6780
rect 22704 6743 22714 6752
rect 22704 6740 22710 6743
rect 25314 6712 25320 6724
rect 25275 6684 25320 6712
rect 25314 6672 25320 6684
rect 25372 6672 25378 6724
rect 11146 6644 11152 6656
rect 10980 6616 11152 6644
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 11330 6604 11336 6656
rect 11388 6644 11394 6656
rect 12345 6647 12403 6653
rect 12345 6644 12357 6647
rect 11388 6616 12357 6644
rect 11388 6604 11394 6616
rect 12345 6613 12357 6616
rect 12391 6613 12403 6647
rect 12345 6607 12403 6613
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 17218 6644 17224 6656
rect 17179 6616 17224 6644
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 19334 6644 19340 6656
rect 19295 6616 19340 6644
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 20254 6644 20260 6656
rect 20215 6616 20260 6644
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 20806 6604 20812 6656
rect 20864 6604 20870 6656
rect 21082 6644 21088 6656
rect 21043 6616 21088 6644
rect 21082 6604 21088 6616
rect 21140 6604 21146 6656
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 22646 6644 22652 6656
rect 22152 6616 22652 6644
rect 22152 6604 22158 6616
rect 22646 6604 22652 6616
rect 22704 6604 22710 6656
rect 24026 6644 24032 6656
rect 23987 6616 24032 6644
rect 24026 6604 24032 6616
rect 24084 6604 24090 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1486 6400 1492 6452
rect 1544 6440 1550 6452
rect 1673 6443 1731 6449
rect 1673 6440 1685 6443
rect 1544 6412 1685 6440
rect 1544 6400 1550 6412
rect 1673 6409 1685 6412
rect 1719 6440 1731 6443
rect 2041 6443 2099 6449
rect 2041 6440 2053 6443
rect 1719 6412 2053 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 2041 6409 2053 6412
rect 2087 6440 2099 6443
rect 3510 6440 3516 6452
rect 2087 6412 3188 6440
rect 3471 6412 3516 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 2148 6313 2176 6412
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6273 2191 6307
rect 3160 6304 3188 6412
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 4246 6440 4252 6452
rect 4207 6412 4252 6440
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 5261 6443 5319 6449
rect 5261 6409 5273 6443
rect 5307 6440 5319 6443
rect 5442 6440 5448 6452
rect 5307 6412 5448 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 6270 6440 6276 6452
rect 6231 6412 6276 6440
rect 6270 6400 6276 6412
rect 6328 6440 6334 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6328 6412 6561 6440
rect 6328 6400 6334 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 7193 6443 7251 6449
rect 7193 6409 7205 6443
rect 7239 6440 7251 6443
rect 8018 6440 8024 6452
rect 7239 6412 8024 6440
rect 7239 6409 7251 6412
rect 7193 6403 7251 6409
rect 8018 6400 8024 6412
rect 8076 6440 8082 6452
rect 9033 6443 9091 6449
rect 9033 6440 9045 6443
rect 8076 6412 9045 6440
rect 8076 6400 8082 6412
rect 9033 6409 9045 6412
rect 9079 6409 9091 6443
rect 10778 6440 10784 6452
rect 10739 6412 10784 6440
rect 9033 6403 9091 6409
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 13630 6440 13636 6452
rect 13591 6412 13636 6440
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 17402 6400 17408 6452
rect 17460 6440 17466 6452
rect 18874 6440 18880 6452
rect 17460 6412 18880 6440
rect 17460 6400 17466 6412
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 19337 6443 19395 6449
rect 19337 6409 19349 6443
rect 19383 6440 19395 6443
rect 19610 6440 19616 6452
rect 19383 6412 19616 6440
rect 19383 6409 19395 6412
rect 19337 6403 19395 6409
rect 19610 6400 19616 6412
rect 19668 6400 19674 6452
rect 20806 6440 20812 6452
rect 20767 6412 20812 6440
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 22646 6400 22652 6452
rect 22704 6440 22710 6452
rect 23017 6443 23075 6449
rect 23017 6440 23029 6443
rect 22704 6412 23029 6440
rect 22704 6400 22710 6412
rect 23017 6409 23029 6412
rect 23063 6440 23075 6443
rect 23385 6443 23443 6449
rect 23385 6440 23397 6443
rect 23063 6412 23397 6440
rect 23063 6409 23075 6412
rect 23017 6403 23075 6409
rect 23385 6409 23397 6412
rect 23431 6409 23443 6443
rect 23385 6403 23443 6409
rect 4264 6304 4292 6400
rect 3160 6276 4292 6304
rect 2133 6267 2191 6273
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5132 6276 5825 6304
rect 5132 6264 5138 6276
rect 5813 6273 5825 6276
rect 5859 6304 5871 6307
rect 6288 6304 6316 6400
rect 7558 6372 7564 6384
rect 7519 6344 7564 6372
rect 7558 6332 7564 6344
rect 7616 6372 7622 6384
rect 12526 6372 12532 6384
rect 7616 6344 7696 6372
rect 12487 6344 12532 6372
rect 7616 6332 7622 6344
rect 7668 6313 7696 6344
rect 12526 6332 12532 6344
rect 12584 6332 12590 6384
rect 22097 6375 22155 6381
rect 22097 6341 22109 6375
rect 22143 6372 22155 6375
rect 23290 6372 23296 6384
rect 22143 6344 23296 6372
rect 22143 6341 22155 6344
rect 22097 6335 22155 6341
rect 23290 6332 23296 6344
rect 23348 6332 23354 6384
rect 23400 6372 23428 6403
rect 23400 6344 23704 6372
rect 5859 6276 6316 6304
rect 7653 6307 7711 6313
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 7653 6273 7665 6307
rect 7699 6273 7711 6307
rect 13538 6304 13544 6316
rect 7653 6267 7711 6273
rect 11808 6276 13544 6304
rect 2222 6196 2228 6248
rect 2280 6236 2286 6248
rect 2400 6239 2458 6245
rect 2400 6236 2412 6239
rect 2280 6208 2412 6236
rect 2280 6196 2286 6208
rect 2400 6205 2412 6208
rect 2446 6236 2458 6239
rect 2682 6236 2688 6248
rect 2446 6208 2688 6236
rect 2446 6205 2458 6208
rect 2400 6199 2458 6205
rect 2682 6196 2688 6208
rect 2740 6196 2746 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 7920 6239 7978 6245
rect 4755 6208 5764 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 5736 6180 5764 6208
rect 7920 6205 7932 6239
rect 7966 6236 7978 6239
rect 8386 6236 8392 6248
rect 7966 6208 8392 6236
rect 7966 6205 7978 6208
rect 7920 6199 7978 6205
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 11330 6236 11336 6248
rect 9824 6208 11336 6236
rect 9824 6196 9830 6208
rect 11330 6196 11336 6208
rect 11388 6196 11394 6248
rect 3234 6128 3240 6180
rect 3292 6168 3298 6180
rect 4985 6171 5043 6177
rect 4985 6168 4997 6171
rect 3292 6140 4997 6168
rect 3292 6128 3298 6140
rect 4985 6137 4997 6140
rect 5031 6168 5043 6171
rect 5537 6171 5595 6177
rect 5537 6168 5549 6171
rect 5031 6140 5549 6168
rect 5031 6137 5043 6140
rect 4985 6131 5043 6137
rect 5537 6137 5549 6140
rect 5583 6137 5595 6171
rect 5718 6168 5724 6180
rect 5679 6140 5724 6168
rect 5537 6131 5595 6137
rect 5552 6100 5580 6131
rect 5718 6128 5724 6140
rect 5776 6128 5782 6180
rect 9674 6128 9680 6180
rect 9732 6168 9738 6180
rect 10686 6168 10692 6180
rect 9732 6140 10692 6168
rect 9732 6128 9738 6140
rect 10686 6128 10692 6140
rect 10744 6168 10750 6180
rect 11057 6171 11115 6177
rect 11057 6168 11069 6171
rect 10744 6140 11069 6168
rect 10744 6128 10750 6140
rect 11057 6137 11069 6140
rect 11103 6137 11115 6171
rect 11057 6131 11115 6137
rect 11241 6171 11299 6177
rect 11241 6137 11253 6171
rect 11287 6168 11299 6171
rect 11808 6168 11836 6276
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 16850 6304 16856 6316
rect 16811 6276 16856 6304
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 18325 6307 18383 6313
rect 18325 6273 18337 6307
rect 18371 6304 18383 6307
rect 19242 6304 19248 6316
rect 18371 6276 19248 6304
rect 18371 6273 18383 6276
rect 18325 6267 18383 6273
rect 19242 6264 19248 6276
rect 19300 6264 19306 6316
rect 22370 6264 22376 6316
rect 22428 6304 22434 6316
rect 22557 6307 22615 6313
rect 22557 6304 22569 6307
rect 22428 6276 22569 6304
rect 22428 6264 22434 6276
rect 22557 6273 22569 6276
rect 22603 6304 22615 6307
rect 23382 6304 23388 6316
rect 22603 6276 23388 6304
rect 22603 6273 22615 6276
rect 22557 6267 22615 6273
rect 23382 6264 23388 6276
rect 23440 6264 23446 6316
rect 23676 6313 23704 6344
rect 23661 6307 23719 6313
rect 23661 6273 23673 6307
rect 23707 6273 23719 6307
rect 23661 6267 23719 6273
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 14090 6236 14096 6248
rect 11931 6208 12940 6236
rect 14051 6208 14096 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 11287 6140 11836 6168
rect 12268 6140 12817 6168
rect 11287 6137 11299 6140
rect 11241 6131 11299 6137
rect 5994 6100 6000 6112
rect 5552 6072 6000 6100
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10134 6100 10140 6112
rect 10095 6072 10140 6100
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10597 6103 10655 6109
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 11256 6100 11284 6131
rect 12268 6112 12296 6140
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 12805 6131 12863 6137
rect 12250 6100 12256 6112
rect 10643 6072 11284 6100
rect 12211 6072 12256 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12912 6100 12940 6208
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 16574 6236 16580 6248
rect 16535 6208 16580 6236
rect 16574 6196 16580 6208
rect 16632 6236 16638 6248
rect 17681 6239 17739 6245
rect 17681 6236 17693 6239
rect 16632 6208 17693 6236
rect 16632 6196 16638 6208
rect 17681 6205 17693 6208
rect 17727 6205 17739 6239
rect 18046 6236 18052 6248
rect 18007 6208 18052 6236
rect 17681 6199 17739 6205
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 18874 6196 18880 6248
rect 18932 6236 18938 6248
rect 19429 6239 19487 6245
rect 19429 6236 19441 6239
rect 18932 6208 19441 6236
rect 18932 6196 18938 6208
rect 19429 6205 19441 6208
rect 19475 6205 19487 6239
rect 19429 6199 19487 6205
rect 19696 6239 19754 6245
rect 19696 6205 19708 6239
rect 19742 6236 19754 6239
rect 20254 6236 20260 6248
rect 19742 6208 20260 6236
rect 19742 6205 19754 6208
rect 19696 6199 19754 6205
rect 20254 6196 20260 6208
rect 20312 6196 20318 6248
rect 21913 6239 21971 6245
rect 21913 6205 21925 6239
rect 21959 6236 21971 6239
rect 25590 6236 25596 6248
rect 21959 6208 22692 6236
rect 25551 6208 25596 6236
rect 21959 6205 21971 6208
rect 21913 6199 21971 6205
rect 13078 6168 13084 6180
rect 13039 6140 13084 6168
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 13998 6128 14004 6180
rect 14056 6168 14062 6180
rect 14338 6171 14396 6177
rect 14338 6168 14350 6171
rect 14056 6140 14350 6168
rect 14056 6128 14062 6140
rect 14338 6137 14350 6140
rect 14384 6137 14396 6171
rect 16114 6168 16120 6180
rect 14338 6131 14396 6137
rect 15488 6140 16120 6168
rect 12989 6103 13047 6109
rect 12989 6100 13001 6103
rect 12912 6072 13001 6100
rect 12989 6069 13001 6072
rect 13035 6100 13047 6103
rect 13170 6100 13176 6112
rect 13035 6072 13176 6100
rect 13035 6069 13047 6072
rect 12989 6063 13047 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 15378 6060 15384 6112
rect 15436 6100 15442 6112
rect 15488 6109 15516 6140
rect 16114 6128 16120 6140
rect 16172 6168 16178 6180
rect 16393 6171 16451 6177
rect 16393 6168 16405 6171
rect 16172 6140 16405 6168
rect 16172 6128 16178 6140
rect 16393 6137 16405 6140
rect 16439 6137 16451 6171
rect 22554 6168 22560 6180
rect 22515 6140 22560 6168
rect 16393 6131 16451 6137
rect 22554 6128 22560 6140
rect 22612 6128 22618 6180
rect 22664 6177 22692 6208
rect 25590 6196 25596 6208
rect 25648 6196 25654 6248
rect 22649 6171 22707 6177
rect 22649 6137 22661 6171
rect 22695 6168 22707 6171
rect 23928 6171 23986 6177
rect 23928 6168 23940 6171
rect 22695 6140 23940 6168
rect 22695 6137 22707 6140
rect 22649 6131 22707 6137
rect 23928 6137 23940 6140
rect 23974 6168 23986 6171
rect 24026 6168 24032 6180
rect 23974 6140 24032 6168
rect 23974 6137 23986 6140
rect 23928 6131 23986 6137
rect 24026 6128 24032 6140
rect 24084 6128 24090 6180
rect 15473 6103 15531 6109
rect 15473 6100 15485 6103
rect 15436 6072 15485 6100
rect 15436 6060 15442 6072
rect 15473 6069 15485 6072
rect 15519 6069 15531 6103
rect 15473 6063 15531 6069
rect 15562 6060 15568 6112
rect 15620 6100 15626 6112
rect 16025 6103 16083 6109
rect 16025 6100 16037 6103
rect 15620 6072 16037 6100
rect 15620 6060 15626 6072
rect 16025 6069 16037 6072
rect 16071 6069 16083 6103
rect 17310 6100 17316 6112
rect 17271 6072 17316 6100
rect 16025 6063 16083 6069
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 21174 6060 21180 6112
rect 21232 6100 21238 6112
rect 21361 6103 21419 6109
rect 21361 6100 21373 6103
rect 21232 6072 21373 6100
rect 21232 6060 21238 6072
rect 21361 6069 21373 6072
rect 21407 6069 21419 6103
rect 21361 6063 21419 6069
rect 24118 6060 24124 6112
rect 24176 6100 24182 6112
rect 25041 6103 25099 6109
rect 25041 6100 25053 6103
rect 24176 6072 25053 6100
rect 24176 6060 24182 6072
rect 25041 6069 25053 6072
rect 25087 6069 25099 6103
rect 25041 6063 25099 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1394 5896 1400 5908
rect 1355 5868 1400 5896
rect 1394 5856 1400 5868
rect 1452 5856 1458 5908
rect 2222 5896 2228 5908
rect 2183 5868 2228 5896
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 4341 5899 4399 5905
rect 4341 5865 4353 5899
rect 4387 5896 4399 5899
rect 4706 5896 4712 5908
rect 4387 5868 4712 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 4982 5896 4988 5908
rect 4943 5868 4988 5896
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5537 5899 5595 5905
rect 5537 5896 5549 5899
rect 5224 5868 5549 5896
rect 5224 5856 5230 5868
rect 5537 5865 5549 5868
rect 5583 5896 5595 5899
rect 6362 5896 6368 5908
rect 5583 5868 6368 5896
rect 5583 5865 5595 5868
rect 5537 5859 5595 5865
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 6546 5896 6552 5908
rect 6507 5868 6552 5896
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7377 5899 7435 5905
rect 7377 5896 7389 5899
rect 6972 5868 7389 5896
rect 6972 5856 6978 5868
rect 7377 5865 7389 5868
rect 7423 5896 7435 5899
rect 8938 5896 8944 5908
rect 7423 5868 7972 5896
rect 8899 5868 8944 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 2866 5788 2872 5840
rect 2924 5828 2930 5840
rect 2961 5831 3019 5837
rect 2961 5828 2973 5831
rect 2924 5800 2973 5828
rect 2924 5788 2930 5800
rect 2961 5797 2973 5800
rect 3007 5797 3019 5831
rect 2961 5791 3019 5797
rect 5074 5788 5080 5840
rect 5132 5828 5138 5840
rect 7944 5837 7972 5868
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 9674 5896 9680 5908
rect 9635 5868 9680 5896
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 10597 5899 10655 5905
rect 10597 5865 10609 5899
rect 10643 5896 10655 5899
rect 11054 5896 11060 5908
rect 10643 5868 11060 5896
rect 10643 5865 10655 5868
rect 10597 5859 10655 5865
rect 11054 5856 11060 5868
rect 11112 5896 11118 5908
rect 11606 5896 11612 5908
rect 11112 5868 11612 5896
rect 11112 5856 11118 5868
rect 11606 5856 11612 5868
rect 11664 5896 11670 5908
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 11664 5868 12081 5896
rect 11664 5856 11670 5868
rect 12069 5865 12081 5868
rect 12115 5896 12127 5899
rect 12713 5899 12771 5905
rect 12713 5896 12725 5899
rect 12115 5868 12725 5896
rect 12115 5865 12127 5868
rect 12069 5859 12127 5865
rect 12713 5865 12725 5868
rect 12759 5896 12771 5899
rect 13078 5896 13084 5908
rect 12759 5868 13084 5896
rect 12759 5865 12771 5868
rect 12713 5859 12771 5865
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 15013 5899 15071 5905
rect 15013 5896 15025 5899
rect 13872 5868 15025 5896
rect 13872 5856 13878 5868
rect 15013 5865 15025 5868
rect 15059 5865 15071 5899
rect 15470 5896 15476 5908
rect 15431 5868 15476 5896
rect 15013 5859 15071 5865
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 18601 5899 18659 5905
rect 18601 5865 18613 5899
rect 18647 5896 18659 5899
rect 19150 5896 19156 5908
rect 18647 5868 19156 5896
rect 18647 5865 18659 5868
rect 18601 5859 18659 5865
rect 19150 5856 19156 5868
rect 19208 5896 19214 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 19208 5868 19625 5896
rect 19208 5856 19214 5868
rect 19613 5865 19625 5868
rect 19659 5865 19671 5899
rect 20070 5896 20076 5908
rect 20031 5868 20076 5896
rect 19613 5859 19671 5865
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 22005 5899 22063 5905
rect 22005 5865 22017 5899
rect 22051 5896 22063 5899
rect 22554 5896 22560 5908
rect 22051 5868 22560 5896
rect 22051 5865 22063 5868
rect 22005 5859 22063 5865
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 23017 5899 23075 5905
rect 23017 5896 23029 5899
rect 22756 5868 23029 5896
rect 7929 5831 7987 5837
rect 5132 5800 5177 5828
rect 5132 5788 5138 5800
rect 7929 5797 7941 5831
rect 7975 5797 7987 5831
rect 8110 5828 8116 5840
rect 8071 5800 8116 5828
rect 7929 5791 7987 5797
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 8205 5831 8263 5837
rect 8205 5797 8217 5831
rect 8251 5828 8263 5831
rect 8386 5828 8392 5840
rect 8251 5800 8392 5828
rect 8251 5797 8263 5800
rect 8205 5791 8263 5797
rect 2777 5763 2835 5769
rect 2777 5729 2789 5763
rect 2823 5760 2835 5763
rect 3326 5760 3332 5772
rect 2823 5732 3332 5760
rect 2823 5729 2835 5732
rect 2777 5723 2835 5729
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 4522 5760 4528 5772
rect 4120 5732 4528 5760
rect 4120 5720 4126 5732
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 7101 5763 7159 5769
rect 7101 5729 7113 5763
rect 7147 5760 7159 5763
rect 8220 5760 8248 5791
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 10134 5788 10140 5840
rect 10192 5828 10198 5840
rect 11146 5828 11152 5840
rect 10192 5800 11152 5828
rect 10192 5788 10198 5800
rect 10704 5769 10732 5800
rect 11146 5788 11152 5800
rect 11204 5788 11210 5840
rect 13173 5831 13231 5837
rect 13173 5797 13185 5831
rect 13219 5828 13231 5831
rect 13219 5800 13676 5828
rect 13219 5797 13231 5800
rect 13173 5791 13231 5797
rect 10962 5769 10968 5772
rect 7147 5732 8248 5760
rect 10689 5763 10747 5769
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 10689 5729 10701 5763
rect 10735 5729 10747 5763
rect 10956 5760 10968 5769
rect 10923 5732 10968 5760
rect 10689 5723 10747 5729
rect 10956 5723 10968 5732
rect 10962 5720 10968 5723
rect 11020 5720 11026 5772
rect 13648 5760 13676 5800
rect 13722 5788 13728 5840
rect 13780 5828 13786 5840
rect 14001 5831 14059 5837
rect 14001 5828 14013 5831
rect 13780 5800 14013 5828
rect 13780 5788 13786 5800
rect 14001 5797 14013 5800
rect 14047 5797 14059 5831
rect 14182 5828 14188 5840
rect 14143 5800 14188 5828
rect 14001 5791 14059 5797
rect 14182 5788 14188 5800
rect 14240 5788 14246 5840
rect 14277 5831 14335 5837
rect 14277 5797 14289 5831
rect 14323 5828 14335 5831
rect 15378 5828 15384 5840
rect 14323 5800 15384 5828
rect 14323 5797 14335 5800
rect 14277 5791 14335 5797
rect 14292 5760 14320 5791
rect 15378 5788 15384 5800
rect 15436 5788 15442 5840
rect 15933 5831 15991 5837
rect 15933 5797 15945 5831
rect 15979 5828 15991 5831
rect 16752 5831 16810 5837
rect 16752 5828 16764 5831
rect 15979 5800 16764 5828
rect 15979 5797 15991 5800
rect 15933 5791 15991 5797
rect 16752 5797 16764 5800
rect 16798 5828 16810 5831
rect 17218 5828 17224 5840
rect 16798 5800 17224 5828
rect 16798 5797 16810 5800
rect 16752 5791 16810 5797
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 21177 5831 21235 5837
rect 21177 5797 21189 5831
rect 21223 5828 21235 5831
rect 21726 5828 21732 5840
rect 21223 5800 21732 5828
rect 21223 5797 21235 5800
rect 21177 5791 21235 5797
rect 21726 5788 21732 5800
rect 21784 5788 21790 5840
rect 22186 5788 22192 5840
rect 22244 5828 22250 5840
rect 22281 5831 22339 5837
rect 22281 5828 22293 5831
rect 22244 5800 22293 5828
rect 22244 5788 22250 5800
rect 22281 5797 22293 5800
rect 22327 5797 22339 5831
rect 22281 5791 22339 5797
rect 13648 5732 14320 5760
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 15252 5732 15301 5760
rect 15252 5720 15258 5732
rect 15289 5729 15301 5732
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 19429 5763 19487 5769
rect 19429 5760 19441 5763
rect 19392 5732 19441 5760
rect 19392 5720 19398 5732
rect 19429 5729 19441 5732
rect 19475 5729 19487 5763
rect 19429 5723 19487 5729
rect 20901 5763 20959 5769
rect 20901 5729 20913 5763
rect 20947 5760 20959 5763
rect 20990 5760 20996 5772
rect 20947 5732 20996 5760
rect 20947 5729 20959 5732
rect 20901 5723 20959 5729
rect 20990 5720 20996 5732
rect 21048 5720 21054 5772
rect 2590 5652 2596 5704
rect 2648 5692 2654 5704
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2648 5664 3065 5692
rect 2648 5652 2654 5664
rect 3053 5661 3065 5664
rect 3099 5692 3111 5695
rect 3510 5692 3516 5704
rect 3099 5664 3516 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5692 5043 5695
rect 5074 5692 5080 5704
rect 5031 5664 5080 5692
rect 5031 5661 5043 5664
rect 4985 5655 5043 5661
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 6454 5692 6460 5704
rect 6415 5664 6460 5692
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5661 16543 5695
rect 16485 5655 16543 5661
rect 4525 5627 4583 5633
rect 4525 5593 4537 5627
rect 4571 5624 4583 5627
rect 5350 5624 5356 5636
rect 4571 5596 5356 5624
rect 4571 5593 4583 5596
rect 4525 5587 4583 5593
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 6086 5624 6092 5636
rect 6047 5596 6092 5624
rect 6086 5584 6092 5596
rect 6144 5584 6150 5636
rect 2498 5556 2504 5568
rect 2459 5528 2504 5556
rect 2498 5516 2504 5528
rect 2556 5516 2562 5568
rect 3697 5559 3755 5565
rect 3697 5525 3709 5559
rect 3743 5556 3755 5559
rect 4062 5556 4068 5568
rect 3743 5528 4068 5556
rect 3743 5525 3755 5528
rect 3697 5519 3755 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 5905 5559 5963 5565
rect 5905 5525 5917 5559
rect 5951 5556 5963 5559
rect 5994 5556 6000 5568
rect 5951 5528 6000 5556
rect 5951 5525 5963 5528
rect 5905 5519 5963 5525
rect 5994 5516 6000 5528
rect 6052 5556 6058 5568
rect 6656 5556 6684 5655
rect 7653 5627 7711 5633
rect 7653 5593 7665 5627
rect 7699 5624 7711 5627
rect 7834 5624 7840 5636
rect 7699 5596 7840 5624
rect 7699 5593 7711 5596
rect 7653 5587 7711 5593
rect 7834 5584 7840 5596
rect 7892 5584 7898 5636
rect 8570 5624 8576 5636
rect 8531 5596 8576 5624
rect 8570 5584 8576 5596
rect 8628 5584 8634 5636
rect 9490 5624 9496 5636
rect 9451 5596 9496 5624
rect 9490 5584 9496 5596
rect 9548 5584 9554 5636
rect 13722 5624 13728 5636
rect 13683 5596 13728 5624
rect 13722 5584 13728 5596
rect 13780 5584 13786 5636
rect 14090 5584 14096 5636
rect 14148 5624 14154 5636
rect 14737 5627 14795 5633
rect 14737 5624 14749 5627
rect 14148 5596 14749 5624
rect 14148 5584 14154 5596
rect 14737 5593 14749 5596
rect 14783 5624 14795 5627
rect 15562 5624 15568 5636
rect 14783 5596 15568 5624
rect 14783 5593 14795 5596
rect 14737 5587 14795 5593
rect 15562 5584 15568 5596
rect 15620 5624 15626 5636
rect 16390 5624 16396 5636
rect 15620 5596 16396 5624
rect 15620 5584 15626 5596
rect 16390 5584 16396 5596
rect 16448 5624 16454 5636
rect 16500 5624 16528 5655
rect 19242 5652 19248 5704
rect 19300 5692 19306 5704
rect 19705 5695 19763 5701
rect 19705 5692 19717 5695
rect 19300 5664 19717 5692
rect 19300 5652 19306 5664
rect 19705 5661 19717 5664
rect 19751 5692 19763 5695
rect 20622 5692 20628 5704
rect 19751 5664 20628 5692
rect 19751 5661 19763 5664
rect 19705 5655 19763 5661
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 20806 5652 20812 5704
rect 20864 5692 20870 5704
rect 21726 5692 21732 5704
rect 20864 5664 21732 5692
rect 20864 5652 20870 5664
rect 21726 5652 21732 5664
rect 21784 5652 21790 5704
rect 22756 5692 22784 5868
rect 23017 5865 23029 5868
rect 23063 5896 23075 5899
rect 23106 5896 23112 5908
rect 23063 5868 23112 5896
rect 23063 5865 23075 5868
rect 23017 5859 23075 5865
rect 23106 5856 23112 5868
rect 23164 5856 23170 5908
rect 23753 5899 23811 5905
rect 23753 5865 23765 5899
rect 23799 5896 23811 5899
rect 24026 5896 24032 5908
rect 23799 5868 24032 5896
rect 23799 5865 23811 5868
rect 23753 5859 23811 5865
rect 24026 5856 24032 5868
rect 24084 5856 24090 5908
rect 25498 5896 25504 5908
rect 25459 5868 25504 5896
rect 25498 5856 25504 5868
rect 25556 5856 25562 5908
rect 22833 5831 22891 5837
rect 22833 5797 22845 5831
rect 22879 5828 22891 5831
rect 22922 5828 22928 5840
rect 22879 5800 22928 5828
rect 22879 5797 22891 5800
rect 22833 5791 22891 5797
rect 22922 5788 22928 5800
rect 22980 5828 22986 5840
rect 23382 5828 23388 5840
rect 22980 5800 23388 5828
rect 22980 5788 22986 5800
rect 23382 5788 23388 5800
rect 23440 5788 23446 5840
rect 23842 5720 23848 5772
rect 23900 5760 23906 5772
rect 24029 5763 24087 5769
rect 24029 5760 24041 5763
rect 23900 5732 24041 5760
rect 23900 5720 23906 5732
rect 24029 5729 24041 5732
rect 24075 5729 24087 5763
rect 24029 5723 24087 5729
rect 25317 5763 25375 5769
rect 25317 5729 25329 5763
rect 25363 5760 25375 5763
rect 25406 5760 25412 5772
rect 25363 5732 25412 5760
rect 25363 5729 25375 5732
rect 25317 5723 25375 5729
rect 25406 5720 25412 5732
rect 25464 5720 25470 5772
rect 22922 5692 22928 5704
rect 22756 5664 22928 5692
rect 22922 5652 22928 5664
rect 22980 5652 22986 5704
rect 23106 5692 23112 5704
rect 23067 5664 23112 5692
rect 23106 5652 23112 5664
rect 23164 5652 23170 5704
rect 24305 5695 24363 5701
rect 24305 5661 24317 5695
rect 24351 5692 24363 5695
rect 24854 5692 24860 5704
rect 24351 5664 24860 5692
rect 24351 5661 24363 5664
rect 24305 5655 24363 5661
rect 24854 5652 24860 5664
rect 24912 5652 24918 5704
rect 16448 5596 16528 5624
rect 20717 5627 20775 5633
rect 16448 5584 16454 5596
rect 20717 5593 20729 5627
rect 20763 5624 20775 5627
rect 22370 5624 22376 5636
rect 20763 5596 22376 5624
rect 20763 5593 20775 5596
rect 20717 5587 20775 5593
rect 22370 5584 22376 5596
rect 22428 5584 22434 5636
rect 10226 5556 10232 5568
rect 6052 5528 6684 5556
rect 10187 5528 10232 5556
rect 6052 5516 6058 5528
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 13538 5556 13544 5568
rect 13499 5528 13544 5556
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 16209 5559 16267 5565
rect 16209 5556 16221 5559
rect 15344 5528 16221 5556
rect 15344 5516 15350 5528
rect 16209 5525 16221 5528
rect 16255 5525 16267 5559
rect 16209 5519 16267 5525
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 17862 5556 17868 5568
rect 16724 5528 17868 5556
rect 16724 5516 16730 5528
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 18966 5556 18972 5568
rect 18927 5528 18972 5556
rect 18966 5516 18972 5528
rect 19024 5516 19030 5568
rect 19150 5556 19156 5568
rect 19111 5528 19156 5556
rect 19150 5516 19156 5528
rect 19208 5516 19214 5568
rect 22554 5556 22560 5568
rect 22515 5528 22560 5556
rect 22554 5516 22560 5528
rect 22612 5516 22618 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 2682 5352 2688 5364
rect 1995 5324 2688 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 3326 5352 3332 5364
rect 3191 5324 3332 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 4982 5352 4988 5364
rect 4755 5324 4988 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 6546 5352 6552 5364
rect 6507 5324 6552 5352
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 7098 5312 7104 5364
rect 7156 5352 7162 5364
rect 7285 5355 7343 5361
rect 7285 5352 7297 5355
rect 7156 5324 7297 5352
rect 7156 5312 7162 5324
rect 7285 5321 7297 5324
rect 7331 5352 7343 5355
rect 8110 5352 8116 5364
rect 7331 5324 8116 5352
rect 7331 5321 7343 5324
rect 7285 5315 7343 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 8386 5312 8392 5364
rect 8444 5352 8450 5364
rect 8849 5355 8907 5361
rect 8849 5352 8861 5355
rect 8444 5324 8861 5352
rect 8444 5312 8450 5324
rect 8849 5321 8861 5324
rect 8895 5321 8907 5355
rect 9766 5352 9772 5364
rect 9727 5324 9772 5352
rect 8849 5315 8907 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 10321 5355 10379 5361
rect 10321 5321 10333 5355
rect 10367 5352 10379 5355
rect 10870 5352 10876 5364
rect 10367 5324 10876 5352
rect 10367 5321 10379 5324
rect 10321 5315 10379 5321
rect 10870 5312 10876 5324
rect 10928 5312 10934 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11241 5355 11299 5361
rect 11241 5352 11253 5355
rect 11204 5324 11253 5352
rect 11204 5312 11210 5324
rect 11241 5321 11253 5324
rect 11287 5321 11299 5355
rect 11241 5315 11299 5321
rect 12713 5355 12771 5361
rect 12713 5321 12725 5355
rect 12759 5352 12771 5355
rect 14182 5352 14188 5364
rect 12759 5324 14188 5352
rect 12759 5321 12771 5324
rect 12713 5315 12771 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 15378 5352 15384 5364
rect 15339 5324 15384 5352
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 15838 5352 15844 5364
rect 15799 5324 15844 5352
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 16390 5312 16396 5364
rect 16448 5352 16454 5364
rect 16761 5355 16819 5361
rect 16761 5352 16773 5355
rect 16448 5324 16773 5352
rect 16448 5312 16454 5324
rect 16761 5321 16773 5324
rect 16807 5321 16819 5355
rect 17218 5352 17224 5364
rect 17179 5324 17224 5352
rect 16761 5315 16819 5321
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 18874 5312 18880 5364
rect 18932 5352 18938 5364
rect 19061 5355 19119 5361
rect 19061 5352 19073 5355
rect 18932 5324 19073 5352
rect 18932 5312 18938 5324
rect 19061 5321 19073 5324
rect 19107 5321 19119 5355
rect 19061 5315 19119 5321
rect 2133 5287 2191 5293
rect 2133 5253 2145 5287
rect 2179 5284 2191 5287
rect 2222 5284 2228 5296
rect 2179 5256 2228 5284
rect 2179 5253 2191 5256
rect 2133 5247 2191 5253
rect 2222 5244 2228 5256
rect 2280 5244 2286 5296
rect 3694 5284 3700 5296
rect 3655 5256 3700 5284
rect 3694 5244 3700 5256
rect 3752 5244 3758 5296
rect 5261 5287 5319 5293
rect 5261 5253 5273 5287
rect 5307 5253 5319 5287
rect 5261 5247 5319 5253
rect 6273 5287 6331 5293
rect 6273 5253 6285 5287
rect 6319 5284 6331 5287
rect 6454 5284 6460 5296
rect 6319 5256 6460 5284
rect 6319 5253 6331 5256
rect 6273 5247 6331 5253
rect 2682 5216 2688 5228
rect 2643 5188 2688 5216
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 5276 5216 5304 5247
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 9784 5284 9812 5312
rect 14274 5284 14280 5296
rect 9784 5256 10916 5284
rect 14235 5256 14280 5284
rect 7190 5216 7196 5228
rect 5276 5188 7196 5216
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 10778 5216 10784 5228
rect 10739 5188 10784 5216
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 10888 5225 10916 5256
rect 14274 5244 14280 5256
rect 14332 5244 14338 5296
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 13265 5219 13323 5225
rect 13265 5216 13277 5219
rect 11931 5188 13277 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 13265 5185 13277 5188
rect 13311 5216 13323 5219
rect 13633 5219 13691 5225
rect 13633 5216 13645 5219
rect 13311 5188 13645 5216
rect 13311 5185 13323 5188
rect 13265 5179 13323 5185
rect 13633 5185 13645 5188
rect 13679 5216 13691 5219
rect 13998 5216 14004 5228
rect 13679 5188 14004 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 13998 5176 14004 5188
rect 14056 5176 14062 5228
rect 14366 5176 14372 5228
rect 14424 5216 14430 5228
rect 16206 5216 16212 5228
rect 14424 5188 15240 5216
rect 16167 5188 16212 5216
rect 14424 5176 14430 5188
rect 2406 5148 2412 5160
rect 2367 5120 2412 5148
rect 2406 5108 2412 5120
rect 2464 5108 2470 5160
rect 5534 5148 5540 5160
rect 5495 5120 5540 5148
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 7469 5151 7527 5157
rect 7469 5117 7481 5151
rect 7515 5148 7527 5151
rect 7558 5148 7564 5160
rect 7515 5120 7564 5148
rect 7515 5117 7527 5120
rect 7469 5111 7527 5117
rect 7558 5108 7564 5120
rect 7616 5148 7622 5160
rect 8202 5148 8208 5160
rect 7616 5120 8208 5148
rect 7616 5108 7622 5120
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 10226 5108 10232 5160
rect 10284 5148 10290 5160
rect 10686 5148 10692 5160
rect 10284 5120 10692 5148
rect 10284 5108 10290 5120
rect 10686 5108 10692 5120
rect 10744 5148 10750 5160
rect 10744 5120 10824 5148
rect 10744 5108 10750 5120
rect 2498 5040 2504 5092
rect 2556 5080 2562 5092
rect 2593 5083 2651 5089
rect 2593 5080 2605 5083
rect 2556 5052 2605 5080
rect 2556 5040 2562 5052
rect 2593 5049 2605 5052
rect 2639 5049 2651 5083
rect 2593 5043 2651 5049
rect 3513 5083 3571 5089
rect 3513 5049 3525 5083
rect 3559 5080 3571 5083
rect 3970 5080 3976 5092
rect 3559 5052 3976 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 4062 5040 4068 5092
rect 4120 5080 4126 5092
rect 4249 5083 4307 5089
rect 4249 5080 4261 5083
rect 4120 5052 4261 5080
rect 4120 5040 4126 5052
rect 4249 5049 4261 5052
rect 4295 5080 4307 5083
rect 5350 5080 5356 5092
rect 4295 5052 5356 5080
rect 4295 5049 4307 5052
rect 4249 5043 4307 5049
rect 5350 5040 5356 5052
rect 5408 5040 5414 5092
rect 5813 5083 5871 5089
rect 5813 5049 5825 5083
rect 5859 5080 5871 5083
rect 5994 5080 6000 5092
rect 5859 5052 6000 5080
rect 5859 5049 5871 5052
rect 5813 5043 5871 5049
rect 5994 5040 6000 5052
rect 6052 5080 6058 5092
rect 6730 5080 6736 5092
rect 6052 5052 6736 5080
rect 6052 5040 6058 5052
rect 6730 5040 6736 5052
rect 6788 5040 6794 5092
rect 7736 5083 7794 5089
rect 7736 5049 7748 5083
rect 7782 5080 7794 5083
rect 8110 5080 8116 5092
rect 7782 5052 8116 5080
rect 7782 5049 7794 5052
rect 7736 5043 7794 5049
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 10796 5089 10824 5120
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 12161 5151 12219 5157
rect 12161 5148 12173 5151
rect 11388 5120 12173 5148
rect 11388 5108 11394 5120
rect 12161 5117 12173 5120
rect 12207 5148 12219 5151
rect 12250 5148 12256 5160
rect 12207 5120 12256 5148
rect 12207 5117 12219 5120
rect 12161 5111 12219 5117
rect 12250 5108 12256 5120
rect 12308 5148 12314 5160
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12308 5120 13001 5148
rect 12308 5108 12314 5120
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 14093 5151 14151 5157
rect 14093 5117 14105 5151
rect 14139 5148 14151 5151
rect 14458 5148 14464 5160
rect 14139 5120 14464 5148
rect 14139 5117 14151 5120
rect 14093 5111 14151 5117
rect 14458 5108 14464 5120
rect 14516 5148 14522 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14516 5120 14565 5148
rect 14516 5108 14522 5120
rect 14553 5117 14565 5120
rect 14599 5148 14611 5151
rect 15102 5148 15108 5160
rect 14599 5120 15108 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 15102 5108 15108 5120
rect 15160 5108 15166 5160
rect 15212 5148 15240 5188
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 16393 5219 16451 5225
rect 16393 5185 16405 5219
rect 16439 5216 16451 5219
rect 17236 5216 17264 5312
rect 16439 5188 17264 5216
rect 19076 5216 19104 5315
rect 20254 5312 20260 5364
rect 20312 5352 20318 5364
rect 20625 5355 20683 5361
rect 20625 5352 20637 5355
rect 20312 5324 20637 5352
rect 20312 5312 20318 5324
rect 20625 5321 20637 5324
rect 20671 5352 20683 5355
rect 20898 5352 20904 5364
rect 20671 5324 20904 5352
rect 20671 5321 20683 5324
rect 20625 5315 20683 5321
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 23382 5312 23388 5364
rect 23440 5352 23446 5364
rect 23477 5355 23535 5361
rect 23477 5352 23489 5355
rect 23440 5324 23489 5352
rect 23440 5312 23446 5324
rect 23477 5321 23489 5324
rect 23523 5321 23535 5355
rect 23477 5315 23535 5321
rect 23842 5312 23848 5364
rect 23900 5352 23906 5364
rect 24213 5355 24271 5361
rect 24213 5352 24225 5355
rect 23900 5324 24225 5352
rect 23900 5312 23906 5324
rect 24213 5321 24225 5324
rect 24259 5321 24271 5355
rect 24762 5352 24768 5364
rect 24723 5324 24768 5352
rect 24213 5315 24271 5321
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 25406 5352 25412 5364
rect 25367 5324 25412 5352
rect 25406 5312 25412 5324
rect 25464 5312 25470 5364
rect 22097 5287 22155 5293
rect 22097 5253 22109 5287
rect 22143 5284 22155 5287
rect 22186 5284 22192 5296
rect 22143 5256 22192 5284
rect 22143 5253 22155 5256
rect 22097 5247 22155 5253
rect 22186 5244 22192 5256
rect 22244 5244 22250 5296
rect 23106 5284 23112 5296
rect 22664 5256 23112 5284
rect 22664 5225 22692 5256
rect 23106 5244 23112 5256
rect 23164 5284 23170 5296
rect 23937 5287 23995 5293
rect 23937 5284 23949 5287
rect 23164 5256 23949 5284
rect 23164 5244 23170 5256
rect 23937 5253 23949 5256
rect 23983 5284 23995 5287
rect 24118 5284 24124 5296
rect 23983 5256 24124 5284
rect 23983 5253 23995 5256
rect 23937 5247 23995 5253
rect 24118 5244 24124 5256
rect 24176 5244 24182 5296
rect 19245 5219 19303 5225
rect 19245 5216 19257 5219
rect 19076 5188 19257 5216
rect 16439 5185 16451 5188
rect 16393 5179 16451 5185
rect 19245 5185 19257 5188
rect 19291 5185 19303 5219
rect 19245 5179 19303 5185
rect 21545 5219 21603 5225
rect 21545 5185 21557 5219
rect 21591 5216 21603 5219
rect 22649 5219 22707 5225
rect 22649 5216 22661 5219
rect 21591 5188 22661 5216
rect 21591 5185 21603 5188
rect 21545 5179 21603 5185
rect 22649 5185 22661 5188
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 22922 5176 22928 5228
rect 22980 5216 22986 5228
rect 23017 5219 23075 5225
rect 23017 5216 23029 5219
rect 22980 5188 23029 5216
rect 22980 5176 22986 5188
rect 23017 5185 23029 5188
rect 23063 5185 23075 5219
rect 23017 5179 23075 5185
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 24762 5216 24768 5228
rect 23808 5188 24768 5216
rect 23808 5176 23814 5188
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 17497 5151 17555 5157
rect 17497 5148 17509 5151
rect 15212 5120 17509 5148
rect 17497 5117 17509 5120
rect 17543 5117 17555 5151
rect 18046 5148 18052 5160
rect 18007 5120 18052 5148
rect 17497 5111 17555 5117
rect 18046 5108 18052 5120
rect 18104 5148 18110 5160
rect 18601 5151 18659 5157
rect 18601 5148 18613 5151
rect 18104 5120 18613 5148
rect 18104 5108 18110 5120
rect 18601 5117 18613 5120
rect 18647 5117 18659 5151
rect 18601 5111 18659 5117
rect 21913 5151 21971 5157
rect 21913 5117 21925 5151
rect 21959 5148 21971 5151
rect 22373 5151 22431 5157
rect 22373 5148 22385 5151
rect 21959 5120 22385 5148
rect 21959 5117 21971 5120
rect 21913 5111 21971 5117
rect 22373 5117 22385 5120
rect 22419 5148 22431 5151
rect 22738 5148 22744 5160
rect 22419 5120 22744 5148
rect 22419 5117 22431 5120
rect 22373 5111 22431 5117
rect 22738 5108 22744 5120
rect 22796 5108 22802 5160
rect 24578 5148 24584 5160
rect 24539 5120 24584 5148
rect 24578 5108 24584 5120
rect 24636 5108 24642 5160
rect 10781 5083 10839 5089
rect 10781 5049 10793 5083
rect 10827 5049 10839 5083
rect 13170 5080 13176 5092
rect 13131 5052 13176 5080
rect 10781 5043 10839 5049
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 13906 5040 13912 5092
rect 13964 5080 13970 5092
rect 14737 5083 14795 5089
rect 14737 5080 14749 5083
rect 13964 5052 14749 5080
rect 13964 5040 13970 5052
rect 14737 5049 14749 5052
rect 14783 5049 14795 5083
rect 14737 5043 14795 5049
rect 14826 5040 14832 5092
rect 14884 5080 14890 5092
rect 16301 5083 16359 5089
rect 14884 5052 14929 5080
rect 14884 5040 14890 5052
rect 16301 5049 16313 5083
rect 16347 5080 16359 5083
rect 16482 5080 16488 5092
rect 16347 5052 16488 5080
rect 16347 5049 16359 5052
rect 16301 5043 16359 5049
rect 16482 5040 16488 5052
rect 16540 5040 16546 5092
rect 18966 5040 18972 5092
rect 19024 5080 19030 5092
rect 19518 5089 19524 5092
rect 19512 5080 19524 5089
rect 19024 5052 19524 5080
rect 19024 5040 19030 5052
rect 19512 5043 19524 5052
rect 19518 5040 19524 5043
rect 19576 5040 19582 5092
rect 22557 5083 22615 5089
rect 22557 5049 22569 5083
rect 22603 5080 22615 5083
rect 22646 5080 22652 5092
rect 22603 5052 22652 5080
rect 22603 5049 22615 5052
rect 22557 5043 22615 5049
rect 22646 5040 22652 5052
rect 22704 5080 22710 5092
rect 23198 5080 23204 5092
rect 22704 5052 23204 5080
rect 22704 5040 22710 5052
rect 23198 5040 23204 5052
rect 23256 5040 23262 5092
rect 4154 5012 4160 5024
rect 4115 4984 4160 5012
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5718 5012 5724 5024
rect 5123 4984 5724 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 10134 5012 10140 5024
rect 10047 4984 10140 5012
rect 10134 4972 10140 4984
rect 10192 5012 10198 5024
rect 10962 5012 10968 5024
rect 10192 4984 10968 5012
rect 10192 4972 10198 4984
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 1857 4811 1915 4817
rect 1857 4808 1869 4811
rect 1820 4780 1869 4808
rect 1820 4768 1826 4780
rect 1857 4777 1869 4780
rect 1903 4777 1915 4811
rect 1857 4771 1915 4777
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 2590 4808 2596 4820
rect 2363 4780 2596 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 2958 4808 2964 4820
rect 2919 4780 2964 4808
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 4614 4808 4620 4820
rect 4575 4780 4620 4808
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 5534 4808 5540 4820
rect 5495 4780 5540 4808
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 6178 4808 6184 4820
rect 6139 4780 6184 4808
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 7745 4811 7803 4817
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 7926 4808 7932 4820
rect 7791 4780 7932 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8202 4808 8208 4820
rect 8163 4780 8208 4808
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 9398 4808 9404 4820
rect 9359 4780 9404 4808
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 12066 4808 12072 4820
rect 12027 4780 12072 4808
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 12759 4780 12817 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 12805 4777 12817 4780
rect 12851 4808 12863 4811
rect 13170 4808 13176 4820
rect 12851 4780 13176 4808
rect 12851 4777 12863 4780
rect 12805 4771 12863 4777
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 13449 4811 13507 4817
rect 13449 4777 13461 4811
rect 13495 4808 13507 4811
rect 14274 4808 14280 4820
rect 13495 4780 14280 4808
rect 13495 4777 13507 4780
rect 13449 4771 13507 4777
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 17773 4811 17831 4817
rect 17773 4808 17785 4811
rect 14424 4780 17785 4808
rect 14424 4768 14430 4780
rect 17773 4777 17785 4780
rect 17819 4777 17831 4811
rect 17773 4771 17831 4777
rect 18417 4811 18475 4817
rect 18417 4777 18429 4811
rect 18463 4808 18475 4811
rect 19334 4808 19340 4820
rect 18463 4780 19340 4808
rect 18463 4777 18475 4780
rect 18417 4771 18475 4777
rect 19334 4768 19340 4780
rect 19392 4768 19398 4820
rect 21358 4808 21364 4820
rect 19628 4780 21364 4808
rect 19628 4752 19656 4780
rect 21358 4768 21364 4780
rect 21416 4768 21422 4820
rect 22097 4811 22155 4817
rect 22097 4777 22109 4811
rect 22143 4808 22155 4811
rect 22646 4808 22652 4820
rect 22143 4780 22652 4808
rect 22143 4777 22155 4780
rect 22097 4771 22155 4777
rect 22646 4768 22652 4780
rect 22704 4768 22710 4820
rect 25222 4808 25228 4820
rect 25183 4780 25228 4808
rect 25222 4768 25228 4780
rect 25280 4768 25286 4820
rect 25590 4808 25596 4820
rect 25551 4780 25596 4808
rect 25590 4768 25596 4780
rect 25648 4768 25654 4820
rect 2774 4700 2780 4752
rect 2832 4740 2838 4752
rect 3053 4743 3111 4749
rect 2832 4712 2877 4740
rect 2832 4700 2838 4712
rect 3053 4709 3065 4743
rect 3099 4740 3111 4743
rect 4062 4740 4068 4752
rect 3099 4712 4068 4740
rect 3099 4709 3111 4712
rect 3053 4703 3111 4709
rect 2682 4632 2688 4684
rect 2740 4672 2746 4684
rect 3068 4672 3096 4703
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 4430 4740 4436 4752
rect 4391 4712 4436 4740
rect 4430 4700 4436 4712
rect 4488 4740 4494 4752
rect 4798 4740 4804 4752
rect 4488 4712 4804 4740
rect 4488 4700 4494 4712
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 5074 4700 5080 4752
rect 5132 4740 5138 4752
rect 5169 4743 5227 4749
rect 5169 4740 5181 4743
rect 5132 4712 5181 4740
rect 5132 4700 5138 4712
rect 5169 4709 5181 4712
rect 5215 4740 5227 4743
rect 6086 4740 6092 4752
rect 5215 4712 6092 4740
rect 5215 4709 5227 4712
rect 5169 4703 5227 4709
rect 6086 4700 6092 4712
rect 6144 4700 6150 4752
rect 7837 4743 7895 4749
rect 7837 4709 7849 4743
rect 7883 4740 7895 4743
rect 8386 4740 8392 4752
rect 7883 4712 8392 4740
rect 7883 4709 7895 4712
rect 7837 4703 7895 4709
rect 8386 4700 8392 4712
rect 8444 4700 8450 4752
rect 8570 4740 8576 4752
rect 8531 4712 8576 4740
rect 8570 4700 8576 4712
rect 8628 4700 8634 4752
rect 13262 4740 13268 4752
rect 13223 4712 13268 4740
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 13906 4700 13912 4752
rect 13964 4740 13970 4752
rect 14185 4743 14243 4749
rect 14185 4740 14197 4743
rect 13964 4712 14197 4740
rect 13964 4700 13970 4712
rect 14185 4709 14197 4712
rect 14231 4709 14243 4743
rect 14185 4703 14243 4709
rect 18785 4743 18843 4749
rect 18785 4709 18797 4743
rect 18831 4740 18843 4743
rect 19242 4740 19248 4752
rect 18831 4712 19248 4740
rect 18831 4709 18843 4712
rect 18785 4703 18843 4709
rect 19242 4700 19248 4712
rect 19300 4700 19306 4752
rect 19610 4740 19616 4752
rect 19523 4712 19616 4740
rect 19610 4700 19616 4712
rect 19668 4700 19674 4752
rect 19797 4743 19855 4749
rect 19797 4709 19809 4743
rect 19843 4740 19855 4743
rect 20162 4740 20168 4752
rect 19843 4712 20168 4740
rect 19843 4709 19855 4712
rect 19797 4703 19855 4709
rect 20162 4700 20168 4712
rect 20220 4740 20226 4752
rect 20346 4740 20352 4752
rect 20220 4712 20352 4740
rect 20220 4700 20226 4712
rect 20346 4700 20352 4712
rect 20404 4700 20410 4752
rect 21453 4743 21511 4749
rect 21453 4740 21465 4743
rect 20824 4712 21465 4740
rect 2740 4644 3096 4672
rect 3697 4675 3755 4681
rect 2740 4632 2746 4644
rect 3697 4641 3709 4675
rect 3743 4672 3755 4675
rect 4154 4672 4160 4684
rect 3743 4644 4160 4672
rect 3743 4641 3755 4644
rect 3697 4635 3755 4641
rect 4154 4632 4160 4644
rect 4212 4672 4218 4684
rect 5442 4672 5448 4684
rect 4212 4644 5448 4672
rect 4212 4632 4218 4644
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 6638 4672 6644 4684
rect 6319 4644 6644 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6638 4632 6644 4644
rect 6696 4672 6702 4684
rect 7101 4675 7159 4681
rect 7101 4672 7113 4675
rect 6696 4644 7113 4672
rect 6696 4632 6702 4644
rect 7101 4641 7113 4644
rect 7147 4672 7159 4675
rect 8110 4672 8116 4684
rect 7147 4644 8116 4672
rect 7147 4641 7159 4644
rect 7101 4635 7159 4641
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 10025 4675 10083 4681
rect 10025 4672 10037 4675
rect 9732 4644 10037 4672
rect 9732 4632 9738 4644
rect 10025 4641 10037 4644
rect 10071 4641 10083 4675
rect 10025 4635 10083 4641
rect 13722 4632 13728 4684
rect 13780 4672 13786 4684
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 13780 4644 14657 4672
rect 13780 4632 13786 4644
rect 14645 4641 14657 4644
rect 14691 4672 14703 4675
rect 14826 4672 14832 4684
rect 14691 4644 14832 4672
rect 14691 4641 14703 4644
rect 14645 4635 14703 4641
rect 14826 4632 14832 4644
rect 14884 4672 14890 4684
rect 16114 4681 16120 4684
rect 16108 4672 16120 4681
rect 14884 4644 15608 4672
rect 16075 4644 16120 4672
rect 14884 4632 14890 4644
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 1578 4604 1584 4616
rect 1443 4576 1584 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 4982 4604 4988 4616
rect 4755 4576 4988 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4604 6239 4607
rect 6454 4604 6460 4616
rect 6227 4576 6460 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 7742 4604 7748 4616
rect 7703 4576 7748 4604
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 8260 4576 9781 4604
rect 8260 4564 8266 4576
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 13587 4576 14872 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 2501 4539 2559 4545
rect 2501 4505 2513 4539
rect 2547 4536 2559 4539
rect 3050 4536 3056 4548
rect 2547 4508 3056 4536
rect 2547 4505 2559 4508
rect 2501 4499 2559 4505
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 4157 4539 4215 4545
rect 4157 4505 4169 4539
rect 4203 4536 4215 4539
rect 5258 4536 5264 4548
rect 4203 4508 5264 4536
rect 4203 4505 4215 4508
rect 4157 4499 4215 4505
rect 5258 4496 5264 4508
rect 5316 4496 5322 4548
rect 5721 4539 5779 4545
rect 5721 4505 5733 4539
rect 5767 4536 5779 4539
rect 7926 4536 7932 4548
rect 5767 4508 7932 4536
rect 5767 4505 5779 4508
rect 5721 4499 5779 4505
rect 7926 4496 7932 4508
rect 7984 4496 7990 4548
rect 14844 4480 14872 4576
rect 6730 4468 6736 4480
rect 6691 4440 6736 4468
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 7285 4471 7343 4477
rect 7285 4437 7297 4471
rect 7331 4468 7343 4471
rect 7834 4468 7840 4480
rect 7331 4440 7840 4468
rect 7331 4437 7343 4440
rect 7285 4431 7343 4437
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 9125 4471 9183 4477
rect 9125 4468 9137 4471
rect 8352 4440 9137 4468
rect 8352 4428 8358 4440
rect 9125 4437 9137 4440
rect 9171 4468 9183 4471
rect 9582 4468 9588 4480
rect 9171 4440 9588 4468
rect 9171 4437 9183 4440
rect 9125 4431 9183 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 11146 4468 11152 4480
rect 11107 4440 11152 4468
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 11698 4468 11704 4480
rect 11659 4440 11704 4468
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 12342 4428 12348 4480
rect 12400 4468 12406 4480
rect 12805 4471 12863 4477
rect 12805 4468 12817 4471
rect 12400 4440 12817 4468
rect 12400 4428 12406 4440
rect 12805 4437 12817 4440
rect 12851 4437 12863 4471
rect 12986 4468 12992 4480
rect 12947 4440 12992 4468
rect 12805 4431 12863 4437
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 14826 4428 14832 4480
rect 14884 4468 14890 4480
rect 15580 4477 15608 4644
rect 16108 4635 16120 4644
rect 16172 4672 16178 4684
rect 16666 4672 16672 4684
rect 16172 4644 16672 4672
rect 16114 4632 16120 4635
rect 16172 4632 16178 4644
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 18414 4632 18420 4684
rect 18472 4672 18478 4684
rect 18966 4672 18972 4684
rect 18472 4644 18972 4672
rect 18472 4632 18478 4644
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 19153 4675 19211 4681
rect 19153 4641 19165 4675
rect 19199 4672 19211 4675
rect 19518 4672 19524 4684
rect 19199 4644 19524 4672
rect 19199 4641 19211 4644
rect 19153 4635 19211 4641
rect 19518 4632 19524 4644
rect 19576 4672 19582 4684
rect 19889 4675 19947 4681
rect 19889 4672 19901 4675
rect 19576 4644 19901 4672
rect 19576 4632 19582 4644
rect 19889 4641 19901 4644
rect 19935 4672 19947 4675
rect 20254 4672 20260 4684
rect 19935 4644 20260 4672
rect 19935 4641 19947 4644
rect 19889 4635 19947 4641
rect 20254 4632 20260 4644
rect 20312 4632 20318 4684
rect 20824 4616 20852 4712
rect 21453 4709 21465 4712
rect 21499 4709 21511 4743
rect 21453 4703 21511 4709
rect 22824 4743 22882 4749
rect 22824 4709 22836 4743
rect 22870 4740 22882 4743
rect 23106 4740 23112 4752
rect 22870 4712 23112 4740
rect 22870 4709 22882 4712
rect 22824 4703 22882 4709
rect 23106 4700 23112 4712
rect 23164 4700 23170 4752
rect 20898 4632 20904 4684
rect 20956 4672 20962 4684
rect 21545 4675 21603 4681
rect 21545 4672 21557 4675
rect 20956 4644 21557 4672
rect 20956 4632 20962 4644
rect 21545 4641 21557 4644
rect 21591 4641 21603 4675
rect 21545 4635 21603 4641
rect 22094 4632 22100 4684
rect 22152 4672 22158 4684
rect 22557 4675 22615 4681
rect 22557 4672 22569 4675
rect 22152 4644 22569 4672
rect 22152 4632 22158 4644
rect 22557 4641 22569 4644
rect 22603 4672 22615 4675
rect 22646 4672 22652 4684
rect 22603 4644 22652 4672
rect 22603 4641 22615 4644
rect 22557 4635 22615 4641
rect 22646 4632 22652 4644
rect 22704 4632 22710 4684
rect 24946 4632 24952 4684
rect 25004 4672 25010 4684
rect 25041 4675 25099 4681
rect 25041 4672 25053 4675
rect 25004 4644 25053 4672
rect 25004 4632 25010 4644
rect 25041 4641 25053 4644
rect 25087 4641 25099 4675
rect 25041 4635 25099 4641
rect 15654 4564 15660 4616
rect 15712 4604 15718 4616
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15712 4576 15853 4604
rect 15712 4564 15718 4576
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 20806 4604 20812 4616
rect 15841 4567 15899 4573
rect 20272 4576 20812 4604
rect 19337 4539 19395 4545
rect 19337 4505 19349 4539
rect 19383 4536 19395 4539
rect 20272 4536 20300 4576
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 21100 4576 21373 4604
rect 19383 4508 20300 4536
rect 20349 4539 20407 4545
rect 19383 4505 19395 4508
rect 19337 4499 19395 4505
rect 20349 4505 20361 4539
rect 20395 4536 20407 4539
rect 20990 4536 20996 4548
rect 20395 4508 20996 4536
rect 20395 4505 20407 4508
rect 20349 4499 20407 4505
rect 20990 4496 20996 4508
rect 21048 4496 21054 4548
rect 14921 4471 14979 4477
rect 14921 4468 14933 4471
rect 14884 4440 14933 4468
rect 14884 4428 14890 4440
rect 14921 4437 14933 4440
rect 14967 4437 14979 4471
rect 14921 4431 14979 4437
rect 15565 4471 15623 4477
rect 15565 4437 15577 4471
rect 15611 4468 15623 4471
rect 15838 4468 15844 4480
rect 15611 4440 15844 4468
rect 15611 4437 15623 4440
rect 15565 4431 15623 4437
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 17218 4468 17224 4480
rect 17179 4440 17224 4468
rect 17218 4428 17224 4440
rect 17276 4428 17282 4480
rect 19886 4428 19892 4480
rect 19944 4468 19950 4480
rect 20717 4471 20775 4477
rect 20717 4468 20729 4471
rect 19944 4440 20729 4468
rect 19944 4428 19950 4440
rect 20717 4437 20729 4440
rect 20763 4468 20775 4471
rect 21100 4468 21128 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 24578 4604 24584 4616
rect 24539 4576 24584 4604
rect 21361 4567 21419 4573
rect 24578 4564 24584 4576
rect 24636 4564 24642 4616
rect 22370 4468 22376 4480
rect 20763 4440 21128 4468
rect 22331 4440 22376 4468
rect 20763 4437 20775 4440
rect 20717 4431 20775 4437
rect 22370 4428 22376 4440
rect 22428 4428 22434 4480
rect 23474 4428 23480 4480
rect 23532 4468 23538 4480
rect 23937 4471 23995 4477
rect 23937 4468 23949 4471
rect 23532 4440 23949 4468
rect 23532 4428 23538 4440
rect 23937 4437 23949 4440
rect 23983 4437 23995 4471
rect 23937 4431 23995 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2866 4264 2872 4276
rect 2827 4236 2872 4264
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 4982 4264 4988 4276
rect 4943 4236 4988 4264
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 6178 4264 6184 4276
rect 6139 4236 6184 4264
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 6638 4264 6644 4276
rect 6599 4236 6644 4264
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 7561 4267 7619 4273
rect 7561 4233 7573 4267
rect 7607 4264 7619 4267
rect 7742 4264 7748 4276
rect 7607 4236 7748 4264
rect 7607 4233 7619 4236
rect 7561 4227 7619 4233
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 8386 4224 8392 4276
rect 8444 4264 8450 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 8444 4236 8493 4264
rect 8444 4224 8450 4236
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 9122 4264 9128 4276
rect 9083 4236 9128 4264
rect 8481 4227 8539 4233
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 10686 4264 10692 4276
rect 10647 4236 10692 4264
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 13633 4267 13691 4273
rect 13633 4264 13645 4267
rect 13320 4236 13645 4264
rect 13320 4224 13326 4236
rect 13633 4233 13645 4236
rect 13679 4233 13691 4267
rect 13633 4227 13691 4233
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 19610 4264 19616 4276
rect 19383 4236 19616 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 19610 4224 19616 4236
rect 19668 4224 19674 4276
rect 20898 4264 20904 4276
rect 20859 4236 20904 4264
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 22646 4224 22652 4276
rect 22704 4264 22710 4276
rect 22925 4267 22983 4273
rect 22925 4264 22937 4267
rect 22704 4236 22937 4264
rect 22704 4224 22710 4236
rect 22925 4233 22937 4236
rect 22971 4233 22983 4267
rect 22925 4227 22983 4233
rect 23106 4224 23112 4276
rect 23164 4264 23170 4276
rect 23293 4267 23351 4273
rect 23293 4264 23305 4267
rect 23164 4236 23305 4264
rect 23164 4224 23170 4236
rect 23293 4233 23305 4236
rect 23339 4233 23351 4267
rect 23293 4227 23351 4233
rect 24946 4224 24952 4276
rect 25004 4264 25010 4276
rect 25501 4267 25559 4273
rect 25501 4264 25513 4267
rect 25004 4236 25513 4264
rect 25004 4224 25010 4236
rect 25501 4233 25513 4236
rect 25547 4233 25559 4267
rect 25501 4227 25559 4233
rect 2774 4156 2780 4208
rect 2832 4156 2838 4208
rect 6454 4196 6460 4208
rect 5552 4168 6460 4196
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 2314 4128 2320 4140
rect 1903 4100 2320 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 2792 4128 2820 4156
rect 5353 4131 5411 4137
rect 5353 4128 5365 4131
rect 2547 4100 2820 4128
rect 4172 4100 5365 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 1946 4020 1952 4072
rect 2004 4060 2010 4072
rect 2041 4063 2099 4069
rect 2041 4060 2053 4063
rect 2004 4032 2053 4060
rect 2004 4020 2010 4032
rect 2041 4029 2053 4032
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 2961 4063 3019 4069
rect 2961 4029 2973 4063
rect 3007 4029 3019 4063
rect 2961 4023 3019 4029
rect 3228 4063 3286 4069
rect 3228 4029 3240 4063
rect 3274 4060 3286 4063
rect 3510 4060 3516 4072
rect 3274 4032 3516 4060
rect 3274 4029 3286 4032
rect 3228 4023 3286 4029
rect 1854 3952 1860 4004
rect 1912 3992 1918 4004
rect 2590 3992 2596 4004
rect 1912 3964 2596 3992
rect 1912 3952 1918 3964
rect 2590 3952 2596 3964
rect 2648 3952 2654 4004
rect 2976 3992 3004 4023
rect 3510 4020 3516 4032
rect 3568 4020 3574 4072
rect 3602 4020 3608 4072
rect 3660 4060 3666 4072
rect 4172 4060 4200 4100
rect 5353 4097 5365 4100
rect 5399 4128 5411 4131
rect 5552 4128 5580 4168
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 7190 4156 7196 4208
rect 7248 4196 7254 4208
rect 8570 4196 8576 4208
rect 7248 4168 8576 4196
rect 7248 4156 7254 4168
rect 8570 4156 8576 4168
rect 8628 4156 8634 4208
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 19521 4199 19579 4205
rect 9732 4168 11008 4196
rect 9732 4156 9738 4168
rect 7374 4128 7380 4140
rect 5399 4100 5580 4128
rect 7335 4100 7380 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 7374 4088 7380 4100
rect 7432 4128 7438 4140
rect 7929 4131 7987 4137
rect 7929 4128 7941 4131
rect 7432 4100 7941 4128
rect 7432 4088 7438 4100
rect 7929 4097 7941 4100
rect 7975 4097 7987 4131
rect 8110 4128 8116 4140
rect 8071 4100 8116 4128
rect 7929 4091 7987 4097
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 9640 4100 9720 4128
rect 9640 4088 9646 4100
rect 5442 4060 5448 4072
rect 3660 4032 4200 4060
rect 5403 4032 5448 4060
rect 3660 4020 3666 4032
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 9692 4069 9720 4100
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 10100 4100 10425 4128
rect 10100 4088 10106 4100
rect 10413 4097 10425 4100
rect 10459 4097 10471 4131
rect 10980 4128 11008 4168
rect 19521 4165 19533 4199
rect 19567 4165 19579 4199
rect 20254 4196 20260 4208
rect 19521 4159 19579 4165
rect 20088 4168 20260 4196
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 10980 4100 12173 4128
rect 10413 4091 10471 4097
rect 12161 4097 12173 4100
rect 12207 4128 12219 4131
rect 14093 4131 14151 4137
rect 12207 4100 13308 4128
rect 12207 4097 12219 4100
rect 12161 4091 12219 4097
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4029 9735 4063
rect 10428 4060 10456 4091
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10428 4032 10977 4060
rect 9677 4023 9735 4029
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 11606 4060 11612 4072
rect 11287 4032 11612 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 13280 4004 13308 4100
rect 14093 4097 14105 4131
rect 14139 4128 14151 4131
rect 14182 4128 14188 4140
rect 14139 4100 14188 4128
rect 14139 4097 14151 4100
rect 14093 4091 14151 4097
rect 14182 4088 14188 4100
rect 14240 4128 14246 4140
rect 14826 4128 14832 4140
rect 14240 4100 14832 4128
rect 14240 4088 14246 4100
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4128 16727 4131
rect 17954 4128 17960 4140
rect 16715 4100 17960 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18874 4088 18880 4140
rect 18932 4128 18938 4140
rect 19536 4128 19564 4159
rect 19886 4128 19892 4140
rect 18932 4100 18977 4128
rect 19536 4100 19892 4128
rect 18932 4088 18938 4100
rect 19886 4088 19892 4100
rect 19944 4088 19950 4140
rect 20088 4137 20116 4168
rect 20254 4156 20260 4168
rect 20312 4156 20318 4208
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 21453 4131 21511 4137
rect 21453 4097 21465 4131
rect 21499 4128 21511 4131
rect 22465 4131 22523 4137
rect 22465 4128 22477 4131
rect 21499 4100 22477 4128
rect 21499 4097 21511 4100
rect 21453 4091 21511 4097
rect 22465 4097 22477 4100
rect 22511 4128 22523 4131
rect 22554 4128 22560 4140
rect 22511 4100 22560 4128
rect 22511 4097 22523 4100
rect 22465 4091 22523 4097
rect 22554 4088 22560 4100
rect 22612 4088 22618 4140
rect 23014 4088 23020 4140
rect 23072 4128 23078 4140
rect 23845 4131 23903 4137
rect 23845 4128 23857 4131
rect 23072 4100 23857 4128
rect 23072 4088 23078 4100
rect 23845 4097 23857 4100
rect 23891 4097 23903 4131
rect 24854 4128 24860 4140
rect 24815 4100 24860 4128
rect 23845 4091 23903 4097
rect 24854 4088 24860 4100
rect 24912 4128 24918 4140
rect 24912 4100 24992 4128
rect 24912 4088 24918 4100
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 16758 4060 16764 4072
rect 15611 4032 16764 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 16758 4020 16764 4032
rect 16816 4020 16822 4072
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4060 17923 4063
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17911 4032 18061 4060
rect 17911 4029 17923 4032
rect 17865 4023 17923 4029
rect 18049 4029 18061 4032
rect 18095 4060 18107 4063
rect 18138 4060 18144 4072
rect 18095 4032 18144 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 18325 4063 18383 4069
rect 18325 4029 18337 4063
rect 18371 4060 18383 4063
rect 21174 4060 21180 4072
rect 18371 4032 21180 4060
rect 18371 4029 18383 4032
rect 18325 4023 18383 4029
rect 21174 4020 21180 4032
rect 21232 4020 21238 4072
rect 23658 4060 23664 4072
rect 23619 4032 23664 4060
rect 23658 4020 23664 4032
rect 23716 4060 23722 4072
rect 24964 4069 24992 4100
rect 24397 4063 24455 4069
rect 24397 4060 24409 4063
rect 23716 4032 24409 4060
rect 23716 4020 23722 4032
rect 24397 4029 24409 4032
rect 24443 4029 24455 4063
rect 24397 4023 24455 4029
rect 24949 4063 25007 4069
rect 24949 4029 24961 4063
rect 24995 4029 25007 4063
rect 24949 4023 25007 4029
rect 3326 3992 3332 4004
rect 2976 3964 3332 3992
rect 3326 3952 3332 3964
rect 3384 3992 3390 4004
rect 4062 3992 4068 4004
rect 3384 3964 4068 3992
rect 3384 3952 3390 3964
rect 4062 3952 4068 3964
rect 4120 3952 4126 4004
rect 5721 3995 5779 4001
rect 5721 3961 5733 3995
rect 5767 3992 5779 3995
rect 6362 3992 6368 4004
rect 5767 3964 6368 3992
rect 5767 3961 5779 3964
rect 5721 3955 5779 3961
rect 6362 3952 6368 3964
rect 6420 3952 6426 4004
rect 7282 3952 7288 4004
rect 7340 3992 7346 4004
rect 8021 3995 8079 4001
rect 8021 3992 8033 3995
rect 7340 3964 8033 3992
rect 7340 3952 7346 3964
rect 8021 3961 8033 3964
rect 8067 3961 8079 3995
rect 8021 3955 8079 3961
rect 9401 3995 9459 4001
rect 9401 3961 9413 3995
rect 9447 3992 9459 3995
rect 9490 3992 9496 4004
rect 9447 3964 9496 3992
rect 9447 3961 9459 3964
rect 9401 3955 9459 3961
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 10137 3995 10195 4001
rect 9640 3964 9685 3992
rect 9640 3952 9646 3964
rect 10137 3961 10149 3995
rect 10183 3992 10195 3995
rect 11149 3995 11207 4001
rect 11149 3992 11161 3995
rect 10183 3964 11161 3992
rect 10183 3961 10195 3964
rect 10137 3955 10195 3961
rect 11149 3961 11161 3964
rect 11195 3992 11207 3995
rect 11974 3992 11980 4004
rect 11195 3964 11980 3992
rect 11195 3961 11207 3964
rect 11149 3955 11207 3961
rect 11974 3952 11980 3964
rect 12032 3952 12038 4004
rect 12986 3992 12992 4004
rect 12947 3964 12992 3992
rect 12986 3952 12992 3964
rect 13044 3952 13050 4004
rect 13262 3992 13268 4004
rect 13223 3964 13268 3992
rect 13262 3952 13268 3964
rect 13320 3952 13326 4004
rect 14553 3995 14611 4001
rect 14553 3961 14565 3995
rect 14599 3992 14611 3995
rect 15470 3992 15476 4004
rect 14599 3964 15476 3992
rect 14599 3961 14611 3964
rect 14553 3955 14611 3961
rect 15470 3952 15476 3964
rect 15528 3952 15534 4004
rect 16669 3995 16727 4001
rect 16669 3961 16681 3995
rect 16715 3992 16727 3995
rect 18414 3992 18420 4004
rect 16715 3964 18420 3992
rect 16715 3961 16727 3964
rect 16669 3955 16727 3961
rect 18414 3952 18420 3964
rect 18472 3952 18478 4004
rect 19426 3952 19432 4004
rect 19484 3992 19490 4004
rect 22002 4001 22008 4004
rect 19797 3995 19855 4001
rect 19797 3992 19809 3995
rect 19484 3964 19809 3992
rect 19484 3952 19490 3964
rect 19797 3961 19809 3964
rect 19843 3992 19855 3995
rect 21987 3995 22008 4001
rect 19843 3964 20116 3992
rect 19843 3961 19855 3964
rect 19797 3955 19855 3961
rect 1486 3933 1492 3936
rect 1479 3927 1492 3933
rect 1479 3924 1491 3927
rect 1447 3896 1491 3924
rect 1479 3893 1491 3896
rect 1479 3887 1492 3893
rect 1486 3884 1492 3887
rect 1544 3884 1550 3936
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3924 2007 3927
rect 2222 3924 2228 3936
rect 1995 3896 2228 3924
rect 1995 3893 2007 3896
rect 1949 3887 2007 3893
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3924 4399 3927
rect 5166 3924 5172 3936
rect 4387 3896 5172 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 8941 3927 8999 3933
rect 8941 3893 8953 3927
rect 8987 3924 8999 3927
rect 9600 3924 9628 3952
rect 8987 3896 9628 3924
rect 12703 3927 12761 3933
rect 8987 3893 8999 3896
rect 8941 3887 8999 3893
rect 12703 3893 12715 3927
rect 12749 3924 12761 3927
rect 12894 3924 12900 3936
rect 12749 3896 12900 3924
rect 12749 3893 12761 3896
rect 12703 3887 12761 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13173 3927 13231 3933
rect 13173 3893 13185 3927
rect 13219 3924 13231 3927
rect 14267 3927 14325 3933
rect 14267 3924 14279 3927
rect 13219 3896 14279 3924
rect 13219 3893 13231 3896
rect 13173 3887 13231 3893
rect 14267 3893 14279 3896
rect 14313 3924 14325 3927
rect 14366 3924 14372 3936
rect 14313 3896 14372 3924
rect 14313 3893 14325 3896
rect 14267 3887 14325 3893
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 14737 3927 14795 3933
rect 14737 3893 14749 3927
rect 14783 3924 14795 3927
rect 15378 3924 15384 3936
rect 14783 3896 15384 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 15562 3884 15568 3936
rect 15620 3924 15626 3936
rect 15841 3927 15899 3933
rect 15841 3924 15853 3927
rect 15620 3896 15853 3924
rect 15620 3884 15626 3896
rect 15841 3893 15853 3896
rect 15887 3893 15899 3927
rect 15841 3887 15899 3893
rect 16199 3927 16257 3933
rect 16199 3893 16211 3927
rect 16245 3924 16257 3927
rect 16482 3924 16488 3936
rect 16245 3896 16488 3924
rect 16245 3893 16257 3896
rect 16199 3887 16257 3893
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 17126 3924 17132 3936
rect 17087 3896 17132 3924
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 19981 3927 20039 3933
rect 19981 3924 19993 3927
rect 18932 3896 19993 3924
rect 18932 3884 18938 3896
rect 19981 3893 19993 3896
rect 20027 3893 20039 3927
rect 20088 3924 20116 3964
rect 21987 3961 21999 3995
rect 21987 3955 22008 3961
rect 22002 3952 22008 3955
rect 22060 3952 22066 4004
rect 22557 3995 22615 4001
rect 22557 3992 22569 3995
rect 22112 3964 22569 3992
rect 20441 3927 20499 3933
rect 20441 3924 20453 3927
rect 20088 3896 20453 3924
rect 19981 3887 20039 3893
rect 20441 3893 20453 3896
rect 20487 3893 20499 3927
rect 20441 3887 20499 3893
rect 21174 3884 21180 3936
rect 21232 3924 21238 3936
rect 21726 3924 21732 3936
rect 21232 3896 21732 3924
rect 21232 3884 21238 3896
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 21821 3927 21879 3933
rect 21821 3893 21833 3927
rect 21867 3924 21879 3927
rect 22112 3924 22140 3964
rect 22557 3961 22569 3964
rect 22603 3992 22615 3995
rect 22830 3992 22836 4004
rect 22603 3964 22836 3992
rect 22603 3961 22615 3964
rect 22557 3955 22615 3961
rect 22830 3952 22836 3964
rect 22888 3992 22894 4004
rect 23474 3992 23480 4004
rect 22888 3964 23480 3992
rect 22888 3952 22894 3964
rect 23474 3952 23480 3964
rect 23532 3952 23538 4004
rect 25222 3952 25228 4004
rect 25280 3992 25286 4004
rect 25869 3995 25927 4001
rect 25869 3992 25881 3995
rect 25280 3964 25881 3992
rect 25280 3952 25286 3964
rect 25869 3961 25881 3964
rect 25915 3961 25927 3995
rect 25869 3955 25927 3961
rect 21867 3896 22140 3924
rect 21867 3893 21879 3896
rect 21821 3887 21879 3893
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 22465 3927 22523 3933
rect 22465 3924 22477 3927
rect 22244 3896 22477 3924
rect 22244 3884 22250 3896
rect 22465 3893 22477 3896
rect 22511 3893 22523 3927
rect 25130 3924 25136 3936
rect 25091 3896 25136 3924
rect 22465 3887 22523 3893
rect 25130 3884 25136 3896
rect 25188 3884 25194 3936
rect 26234 3924 26240 3936
rect 26195 3896 26240 3924
rect 26234 3884 26240 3896
rect 26292 3884 26298 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1397 3723 1455 3729
rect 1397 3689 1409 3723
rect 1443 3720 1455 3723
rect 1670 3720 1676 3732
rect 1443 3692 1676 3720
rect 1443 3689 1455 3692
rect 1397 3683 1455 3689
rect 1670 3680 1676 3692
rect 1728 3680 1734 3732
rect 2317 3723 2375 3729
rect 2317 3689 2329 3723
rect 2363 3720 2375 3723
rect 2682 3720 2688 3732
rect 2363 3692 2688 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 2961 3723 3019 3729
rect 2961 3689 2973 3723
rect 3007 3720 3019 3723
rect 3050 3720 3056 3732
rect 3007 3692 3056 3720
rect 3007 3689 3019 3692
rect 2961 3683 3019 3689
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 3326 3680 3332 3732
rect 3384 3720 3390 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3384 3692 3433 3720
rect 3384 3680 3390 3692
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 3510 3680 3516 3732
rect 3568 3720 3574 3732
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 3568 3692 3801 3720
rect 3568 3680 3574 3692
rect 3789 3689 3801 3692
rect 3835 3689 3847 3723
rect 3789 3683 3847 3689
rect 4893 3723 4951 3729
rect 4893 3689 4905 3723
rect 4939 3720 4951 3723
rect 5166 3720 5172 3732
rect 4939 3692 5172 3720
rect 4939 3689 4951 3692
rect 4893 3683 4951 3689
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5445 3723 5503 3729
rect 5445 3689 5457 3723
rect 5491 3720 5503 3723
rect 6638 3720 6644 3732
rect 5491 3692 6644 3720
rect 5491 3689 5503 3692
rect 5445 3683 5503 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 7469 3723 7527 3729
rect 7469 3720 7481 3723
rect 7340 3692 7481 3720
rect 7340 3680 7346 3692
rect 7469 3689 7481 3692
rect 7515 3720 7527 3723
rect 7558 3720 7564 3732
rect 7515 3692 7564 3720
rect 7515 3689 7527 3692
rect 7469 3683 7527 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 8536 3692 8585 3720
rect 8536 3680 8542 3692
rect 8573 3689 8585 3692
rect 8619 3689 8631 3723
rect 8573 3683 8631 3689
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9674 3720 9680 3732
rect 9539 3692 9680 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 11517 3723 11575 3729
rect 11517 3720 11529 3723
rect 11112 3692 11529 3720
rect 11112 3680 11118 3692
rect 11517 3689 11529 3692
rect 11563 3689 11575 3723
rect 11517 3683 11575 3689
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 13320 3692 14105 3720
rect 13320 3680 13326 3692
rect 14093 3689 14105 3692
rect 14139 3689 14151 3723
rect 14093 3683 14151 3689
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14608 3692 15025 3720
rect 14608 3680 14614 3692
rect 15013 3689 15025 3692
rect 15059 3720 15071 3723
rect 15838 3720 15844 3732
rect 15059 3692 15844 3720
rect 15059 3689 15071 3692
rect 15013 3683 15071 3689
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 18506 3680 18512 3732
rect 18564 3720 18570 3732
rect 18877 3723 18935 3729
rect 18877 3720 18889 3723
rect 18564 3692 18889 3720
rect 18564 3680 18570 3692
rect 18877 3689 18889 3692
rect 18923 3689 18935 3723
rect 20254 3720 20260 3732
rect 20215 3692 20260 3720
rect 18877 3683 18935 3689
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 20717 3723 20775 3729
rect 20717 3689 20729 3723
rect 20763 3720 20775 3723
rect 20806 3720 20812 3732
rect 20763 3692 20812 3720
rect 20763 3689 20775 3692
rect 20717 3683 20775 3689
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 22278 3720 22284 3732
rect 22239 3692 22284 3720
rect 22278 3680 22284 3692
rect 22336 3680 22342 3732
rect 23474 3680 23480 3732
rect 23532 3720 23538 3732
rect 23937 3723 23995 3729
rect 23937 3720 23949 3723
rect 23532 3692 23949 3720
rect 23532 3680 23538 3692
rect 23937 3689 23949 3692
rect 23983 3689 23995 3723
rect 23937 3683 23995 3689
rect 25225 3723 25283 3729
rect 25225 3689 25237 3723
rect 25271 3720 25283 3723
rect 25314 3720 25320 3732
rect 25271 3692 25320 3720
rect 25271 3689 25283 3692
rect 25225 3683 25283 3689
rect 25314 3680 25320 3692
rect 25372 3680 25378 3732
rect 25406 3680 25412 3732
rect 25464 3720 25470 3732
rect 25593 3723 25651 3729
rect 25593 3720 25605 3723
rect 25464 3692 25605 3720
rect 25464 3680 25470 3692
rect 25593 3689 25605 3692
rect 25639 3689 25651 3723
rect 25593 3683 25651 3689
rect 2777 3655 2835 3661
rect 2777 3621 2789 3655
rect 2823 3652 2835 3655
rect 3694 3652 3700 3664
rect 2823 3624 3700 3652
rect 2823 3621 2835 3624
rect 2777 3615 2835 3621
rect 3694 3612 3700 3624
rect 3752 3612 3758 3664
rect 5804 3655 5862 3661
rect 5804 3621 5816 3655
rect 5850 3652 5862 3655
rect 5994 3652 6000 3664
rect 5850 3624 6000 3652
rect 5850 3621 5862 3624
rect 5804 3615 5862 3621
rect 5994 3612 6000 3624
rect 6052 3652 6058 3664
rect 6730 3652 6736 3664
rect 6052 3624 6736 3652
rect 6052 3612 6058 3624
rect 6730 3612 6736 3624
rect 6788 3612 6794 3664
rect 12253 3655 12311 3661
rect 12253 3621 12265 3655
rect 12299 3652 12311 3655
rect 12980 3655 13038 3661
rect 12980 3652 12992 3655
rect 12299 3624 12992 3652
rect 12299 3621 12311 3624
rect 12253 3615 12311 3621
rect 12980 3621 12992 3624
rect 13026 3652 13038 3655
rect 14182 3652 14188 3664
rect 13026 3624 14188 3652
rect 13026 3621 13038 3624
rect 12980 3615 13038 3621
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 15654 3652 15660 3664
rect 15615 3624 15660 3652
rect 15654 3612 15660 3624
rect 15712 3612 15718 3664
rect 16758 3612 16764 3664
rect 16816 3652 16822 3664
rect 17190 3655 17248 3661
rect 17190 3652 17202 3655
rect 16816 3624 17202 3652
rect 16816 3612 16822 3624
rect 17190 3621 17202 3624
rect 17236 3621 17248 3655
rect 17190 3615 17248 3621
rect 19705 3655 19763 3661
rect 19705 3621 19717 3655
rect 19751 3652 19763 3655
rect 19978 3652 19984 3664
rect 19751 3624 19984 3652
rect 19751 3621 19763 3624
rect 19705 3615 19763 3621
rect 19978 3612 19984 3624
rect 20036 3612 20042 3664
rect 21177 3655 21235 3661
rect 21177 3621 21189 3655
rect 21223 3652 21235 3655
rect 21818 3652 21824 3664
rect 21223 3624 21824 3652
rect 21223 3621 21235 3624
rect 21177 3615 21235 3621
rect 21818 3612 21824 3624
rect 21876 3612 21882 3664
rect 22830 3661 22836 3664
rect 22824 3652 22836 3661
rect 22791 3624 22836 3652
rect 22824 3615 22836 3624
rect 22830 3612 22836 3615
rect 22888 3612 22894 3664
rect 23566 3612 23572 3664
rect 23624 3652 23630 3664
rect 23750 3652 23756 3664
rect 23624 3624 23756 3652
rect 23624 3612 23630 3624
rect 23750 3612 23756 3624
rect 23808 3612 23814 3664
rect 4062 3584 4068 3596
rect 4023 3556 4068 3584
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 6270 3584 6276 3596
rect 4387 3556 6276 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 7929 3587 7987 3593
rect 7929 3553 7941 3587
rect 7975 3584 7987 3587
rect 8665 3587 8723 3593
rect 8665 3584 8677 3587
rect 7975 3556 8677 3584
rect 7975 3553 7987 3556
rect 7929 3547 7987 3553
rect 8665 3553 8677 3556
rect 8711 3553 8723 3587
rect 8665 3547 8723 3553
rect 3050 3516 3056 3528
rect 3011 3488 3056 3516
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 3326 3476 3332 3528
rect 3384 3516 3390 3528
rect 3878 3516 3884 3528
rect 3384 3488 3884 3516
rect 3384 3476 3390 3488
rect 3878 3476 3884 3488
rect 3936 3516 3942 3528
rect 5537 3519 5595 3525
rect 5537 3516 5549 3519
rect 3936 3488 5549 3516
rect 3936 3476 3942 3488
rect 5537 3485 5549 3488
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 2498 3448 2504 3460
rect 2459 3420 2504 3448
rect 2498 3408 2504 3420
rect 2556 3408 2562 3460
rect 1946 3380 1952 3392
rect 1907 3352 1952 3380
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 5552 3380 5580 3479
rect 7944 3460 7972 3547
rect 9122 3544 9128 3596
rect 9180 3544 9186 3596
rect 10404 3587 10462 3593
rect 10404 3553 10416 3587
rect 10450 3584 10462 3587
rect 11146 3584 11152 3596
rect 10450 3556 11152 3584
rect 10450 3553 10462 3556
rect 10404 3547 10462 3553
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3584 12679 3587
rect 13722 3584 13728 3596
rect 12667 3556 13728 3584
rect 12667 3553 12679 3556
rect 12621 3547 12679 3553
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 15562 3544 15568 3596
rect 15620 3584 15626 3596
rect 16942 3584 16948 3596
rect 15620 3556 16948 3584
rect 15620 3544 15626 3556
rect 16942 3544 16948 3556
rect 17000 3544 17006 3596
rect 19426 3584 19432 3596
rect 19387 3556 19432 3584
rect 19426 3544 19432 3556
rect 19484 3544 19490 3596
rect 20901 3587 20959 3593
rect 20901 3553 20913 3587
rect 20947 3584 20959 3587
rect 20990 3584 20996 3596
rect 20947 3556 20996 3584
rect 20947 3553 20959 3556
rect 20901 3547 20959 3553
rect 20990 3544 20996 3556
rect 21048 3584 21054 3596
rect 21634 3584 21640 3596
rect 21048 3556 21640 3584
rect 21048 3544 21054 3556
rect 21634 3544 21640 3556
rect 21692 3544 21698 3596
rect 22005 3587 22063 3593
rect 22005 3553 22017 3587
rect 22051 3584 22063 3587
rect 22186 3584 22192 3596
rect 22051 3556 22192 3584
rect 22051 3553 22063 3556
rect 22005 3547 22063 3553
rect 22186 3544 22192 3556
rect 22244 3544 22250 3596
rect 22557 3587 22615 3593
rect 22557 3553 22569 3587
rect 22603 3584 22615 3587
rect 22646 3584 22652 3596
rect 22603 3556 22652 3584
rect 22603 3553 22615 3556
rect 22557 3547 22615 3553
rect 22646 3544 22652 3556
rect 22704 3544 22710 3596
rect 25038 3584 25044 3596
rect 24999 3556 25044 3584
rect 25038 3544 25044 3556
rect 25096 3544 25102 3596
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 25958 3584 25964 3596
rect 25372 3556 25964 3584
rect 25372 3544 25378 3556
rect 25958 3544 25964 3556
rect 26016 3544 26022 3596
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 9140 3516 9168 3544
rect 8619 3488 9168 3516
rect 9953 3519 10011 3525
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 9999 3488 10149 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 12710 3516 12716 3528
rect 12671 3488 12716 3516
rect 10137 3479 10195 3485
rect 6917 3451 6975 3457
rect 6917 3417 6929 3451
rect 6963 3448 6975 3451
rect 7098 3448 7104 3460
rect 6963 3420 7104 3448
rect 6963 3417 6975 3420
rect 6917 3411 6975 3417
rect 7098 3408 7104 3420
rect 7156 3448 7162 3460
rect 7926 3448 7932 3460
rect 7156 3420 7932 3448
rect 7156 3408 7162 3420
rect 7926 3408 7932 3420
rect 7984 3408 7990 3460
rect 9125 3451 9183 3457
rect 9125 3417 9137 3451
rect 9171 3448 9183 3451
rect 9490 3448 9496 3460
rect 9171 3420 9496 3448
rect 9171 3417 9183 3420
rect 9125 3411 9183 3417
rect 9490 3408 9496 3420
rect 9548 3448 9554 3460
rect 10042 3448 10048 3460
rect 9548 3420 10048 3448
rect 9548 3408 9554 3420
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 6454 3380 6460 3392
rect 5552 3352 6460 3380
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 8110 3380 8116 3392
rect 8071 3352 8116 3380
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 10152 3380 10180 3479
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 15930 3516 15936 3528
rect 15843 3488 15936 3516
rect 15930 3476 15936 3488
rect 15988 3516 15994 3528
rect 19337 3519 19395 3525
rect 15988 3488 16804 3516
rect 15988 3476 15994 3488
rect 15378 3448 15384 3460
rect 15339 3420 15384 3448
rect 15378 3408 15384 3420
rect 15436 3408 15442 3460
rect 14734 3380 14740 3392
rect 9456 3352 10180 3380
rect 14695 3352 14740 3380
rect 9456 3340 9462 3352
rect 14734 3340 14740 3352
rect 14792 3340 14798 3392
rect 15286 3340 15292 3392
rect 15344 3380 15350 3392
rect 16114 3380 16120 3392
rect 15344 3352 16120 3380
rect 15344 3340 15350 3352
rect 16114 3340 16120 3352
rect 16172 3380 16178 3392
rect 16776 3389 16804 3488
rect 19337 3485 19349 3519
rect 19383 3516 19395 3519
rect 20346 3516 20352 3528
rect 19383 3488 20352 3516
rect 19383 3485 19395 3488
rect 19337 3479 19395 3485
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 24854 3448 24860 3460
rect 24815 3420 24860 3448
rect 24854 3408 24860 3420
rect 24912 3408 24918 3460
rect 16301 3383 16359 3389
rect 16301 3380 16313 3383
rect 16172 3352 16313 3380
rect 16172 3340 16178 3352
rect 16301 3349 16313 3352
rect 16347 3349 16359 3383
rect 16301 3343 16359 3349
rect 16761 3383 16819 3389
rect 16761 3349 16773 3383
rect 16807 3380 16819 3383
rect 18325 3383 18383 3389
rect 18325 3380 18337 3383
rect 16807 3352 18337 3380
rect 16807 3349 16819 3352
rect 16761 3343 16819 3349
rect 18325 3349 18337 3352
rect 18371 3349 18383 3383
rect 18325 3343 18383 3349
rect 24026 3340 24032 3392
rect 24084 3380 24090 3392
rect 24489 3383 24547 3389
rect 24489 3380 24501 3383
rect 24084 3352 24501 3380
rect 24084 3340 24090 3352
rect 24489 3349 24501 3352
rect 24535 3349 24547 3383
rect 24489 3343 24547 3349
rect 25774 3340 25780 3392
rect 25832 3380 25838 3392
rect 25961 3383 26019 3389
rect 25961 3380 25973 3383
rect 25832 3352 25973 3380
rect 25832 3340 25838 3352
rect 25961 3349 25973 3352
rect 26007 3349 26019 3383
rect 25961 3343 26019 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 2004 3148 3924 3176
rect 2004 3136 2010 3148
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 1486 2972 1492 2984
rect 1443 2944 1492 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 1486 2932 1492 2944
rect 1544 2932 1550 2984
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 2639 2944 2697 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 2685 2941 2697 2944
rect 2731 2972 2743 2975
rect 3326 2972 3332 2984
rect 2731 2944 3332 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 1670 2904 1676 2916
rect 1631 2876 1676 2904
rect 1670 2864 1676 2876
rect 1728 2864 1734 2916
rect 2952 2907 3010 2913
rect 2952 2873 2964 2907
rect 2998 2904 3010 2907
rect 3142 2904 3148 2916
rect 2998 2876 3148 2904
rect 2998 2873 3010 2876
rect 2952 2867 3010 2873
rect 3142 2864 3148 2876
rect 3200 2864 3206 2916
rect 2225 2839 2283 2845
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 3050 2836 3056 2848
rect 2271 2808 3056 2836
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 3896 2836 3924 3148
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 5258 3176 5264 3188
rect 4120 3148 5264 3176
rect 4120 3136 4126 3148
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 6273 3179 6331 3185
rect 6273 3145 6285 3179
rect 6319 3176 6331 3179
rect 6454 3176 6460 3188
rect 6319 3148 6460 3176
rect 6319 3145 6331 3148
rect 6273 3139 6331 3145
rect 6454 3136 6460 3148
rect 6512 3176 6518 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6512 3148 6561 3176
rect 6512 3136 6518 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 9125 3179 9183 3185
rect 9125 3176 9137 3179
rect 8352 3148 9137 3176
rect 8352 3136 8358 3148
rect 9125 3145 9137 3148
rect 9171 3145 9183 3179
rect 9125 3139 9183 3145
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3040 5779 3043
rect 9140 3040 9168 3139
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 14277 3179 14335 3185
rect 14277 3176 14289 3179
rect 14240 3148 14289 3176
rect 14240 3136 14246 3148
rect 14277 3145 14289 3148
rect 14323 3145 14335 3179
rect 14277 3139 14335 3145
rect 15381 3179 15439 3185
rect 15381 3145 15393 3179
rect 15427 3176 15439 3179
rect 15654 3176 15660 3188
rect 15427 3148 15660 3176
rect 15427 3145 15439 3148
rect 15381 3139 15439 3145
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 16816 3148 16865 3176
rect 16816 3136 16822 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17000 3148 17417 3176
rect 17000 3136 17006 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17770 3176 17776 3188
rect 17731 3148 17776 3176
rect 17405 3139 17463 3145
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18138 3176 18144 3188
rect 18099 3148 18144 3176
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19392 3148 19437 3176
rect 19392 3136 19398 3148
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20438 3176 20444 3188
rect 20036 3148 20444 3176
rect 20036 3136 20042 3148
rect 20438 3136 20444 3148
rect 20496 3176 20502 3188
rect 20717 3179 20775 3185
rect 20717 3176 20729 3179
rect 20496 3148 20729 3176
rect 20496 3136 20502 3148
rect 20717 3145 20729 3148
rect 20763 3145 20775 3179
rect 20990 3176 20996 3188
rect 20951 3148 20996 3176
rect 20717 3139 20775 3145
rect 20990 3136 20996 3148
rect 21048 3136 21054 3188
rect 22370 3176 22376 3188
rect 22331 3148 22376 3176
rect 22370 3136 22376 3148
rect 22428 3136 22434 3188
rect 22830 3136 22836 3188
rect 22888 3176 22894 3188
rect 23385 3179 23443 3185
rect 23385 3176 23397 3179
rect 22888 3148 23397 3176
rect 22888 3136 22894 3148
rect 23385 3145 23397 3148
rect 23431 3145 23443 3179
rect 24946 3176 24952 3188
rect 24907 3148 24952 3176
rect 23385 3139 23443 3145
rect 24946 3136 24952 3148
rect 25004 3136 25010 3188
rect 25038 3136 25044 3188
rect 25096 3176 25102 3188
rect 25777 3179 25835 3185
rect 25777 3176 25789 3179
rect 25096 3148 25789 3176
rect 25096 3136 25102 3148
rect 25777 3145 25789 3148
rect 25823 3145 25835 3179
rect 25777 3139 25835 3145
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 5767 3012 6960 3040
rect 9140 3012 9321 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 6932 2984 6960 3012
rect 9309 3009 9321 3012
rect 9355 3040 9367 3043
rect 17788 3040 17816 3136
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 19061 3111 19119 3117
rect 19061 3108 19073 3111
rect 18012 3080 19073 3108
rect 18012 3068 18018 3080
rect 19061 3077 19073 3080
rect 19107 3077 19119 3111
rect 19702 3108 19708 3120
rect 19663 3080 19708 3108
rect 19061 3071 19119 3077
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 9355 3012 9444 3040
rect 17788 3012 18521 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9416 2984 9444 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 5077 2975 5135 2981
rect 5077 2941 5089 2975
rect 5123 2972 5135 2975
rect 5813 2975 5871 2981
rect 5813 2972 5825 2975
rect 5123 2944 5825 2972
rect 5123 2941 5135 2944
rect 5077 2935 5135 2941
rect 5813 2941 5825 2944
rect 5859 2941 5871 2975
rect 5813 2935 5871 2941
rect 5718 2904 5724 2916
rect 5679 2876 5724 2904
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 5828 2904 5856 2935
rect 6454 2932 6460 2984
rect 6512 2972 6518 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6512 2944 6837 2972
rect 6512 2932 6518 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 6914 2932 6920 2984
rect 6972 2932 6978 2984
rect 7098 2981 7104 2984
rect 7092 2972 7104 2981
rect 7059 2944 7104 2972
rect 7092 2935 7104 2944
rect 7098 2932 7104 2935
rect 7156 2932 7162 2984
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 9456 2944 11253 2972
rect 9456 2932 9462 2944
rect 11241 2941 11253 2944
rect 11287 2972 11299 2975
rect 12161 2975 12219 2981
rect 12161 2972 12173 2975
rect 11287 2944 12173 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 12161 2941 12173 2944
rect 12207 2972 12219 2975
rect 12710 2972 12716 2984
rect 12207 2944 12716 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 12710 2932 12716 2944
rect 12768 2972 12774 2984
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12768 2944 12909 2972
rect 12768 2932 12774 2944
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 12897 2935 12955 2941
rect 13164 2975 13222 2981
rect 13164 2941 13176 2975
rect 13210 2972 13222 2975
rect 13722 2972 13728 2984
rect 13210 2944 13728 2972
rect 13210 2941 13222 2944
rect 13164 2935 13222 2941
rect 9554 2907 9612 2913
rect 9554 2904 9566 2907
rect 5828 2876 7052 2904
rect 4065 2839 4123 2845
rect 4065 2836 4077 2839
rect 3896 2808 4077 2836
rect 4065 2805 4077 2808
rect 4111 2836 4123 2839
rect 4246 2836 4252 2848
rect 4111 2808 4252 2836
rect 4111 2805 4123 2808
rect 4065 2799 4123 2805
rect 4246 2796 4252 2808
rect 4304 2836 4310 2848
rect 4617 2839 4675 2845
rect 4617 2836 4629 2839
rect 4304 2808 4629 2836
rect 4304 2796 4310 2808
rect 4617 2805 4629 2808
rect 4663 2805 4675 2839
rect 7024 2836 7052 2876
rect 8772 2876 9566 2904
rect 8772 2845 8800 2876
rect 9554 2873 9566 2876
rect 9600 2873 9612 2907
rect 9554 2867 9612 2873
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 7024 2808 8217 2836
rect 4617 2799 4675 2805
rect 8205 2805 8217 2808
rect 8251 2836 8263 2839
rect 8757 2839 8815 2845
rect 8757 2836 8769 2839
rect 8251 2808 8769 2836
rect 8251 2805 8263 2808
rect 8205 2799 8263 2805
rect 8757 2805 8769 2808
rect 8803 2805 8815 2839
rect 10686 2836 10692 2848
rect 10647 2808 10692 2836
rect 8757 2799 8815 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 11146 2796 11152 2848
rect 11204 2836 11210 2848
rect 11609 2839 11667 2845
rect 11609 2836 11621 2839
rect 11204 2808 11621 2836
rect 11204 2796 11210 2808
rect 11609 2805 11621 2808
rect 11655 2805 11667 2839
rect 12912 2836 12940 2935
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2972 15255 2975
rect 15473 2975 15531 2981
rect 15473 2972 15485 2975
rect 15243 2944 15485 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 15473 2941 15485 2944
rect 15519 2972 15531 2975
rect 15562 2972 15568 2984
rect 15519 2944 15568 2972
rect 15519 2941 15531 2944
rect 15473 2935 15531 2941
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 19076 2972 19104 3071
rect 19702 3068 19708 3080
rect 19760 3068 19766 3120
rect 22646 3068 22652 3120
rect 22704 3108 22710 3120
rect 23017 3111 23075 3117
rect 23017 3108 23029 3111
rect 22704 3080 23029 3108
rect 22704 3068 22710 3080
rect 23017 3077 23029 3080
rect 23063 3077 23075 3111
rect 24486 3108 24492 3120
rect 24447 3080 24492 3108
rect 23017 3071 23075 3077
rect 24486 3068 24492 3080
rect 24544 3068 24550 3120
rect 19521 3043 19579 3049
rect 19521 3009 19533 3043
rect 19567 3040 19579 3043
rect 20162 3040 20168 3052
rect 19567 3012 20168 3040
rect 19567 3009 19579 3012
rect 19521 3003 19579 3009
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 21450 3040 21456 3052
rect 21411 3012 21456 3040
rect 21450 3000 21456 3012
rect 21508 3000 21514 3052
rect 23934 3040 23940 3052
rect 23895 3012 23940 3040
rect 23934 3000 23940 3012
rect 23992 3000 23998 3052
rect 25317 3043 25375 3049
rect 25317 3009 25329 3043
rect 25363 3040 25375 3043
rect 25682 3040 25688 3052
rect 25363 3012 25688 3040
rect 25363 3009 25375 3012
rect 25317 3003 25375 3009
rect 25682 3000 25688 3012
rect 25740 3000 25746 3052
rect 20257 2975 20315 2981
rect 20257 2972 20269 2975
rect 19076 2944 20269 2972
rect 20257 2941 20269 2944
rect 20303 2972 20315 2975
rect 20530 2972 20536 2984
rect 20303 2944 20536 2972
rect 20303 2941 20315 2944
rect 20257 2935 20315 2941
rect 20530 2932 20536 2944
rect 20588 2932 20594 2984
rect 20714 2932 20720 2984
rect 20772 2972 20778 2984
rect 21177 2975 21235 2981
rect 21177 2972 21189 2975
rect 20772 2944 21189 2972
rect 20772 2932 20778 2944
rect 21177 2941 21189 2944
rect 21223 2972 21235 2975
rect 21913 2975 21971 2981
rect 21913 2972 21925 2975
rect 21223 2944 21925 2972
rect 21223 2941 21235 2944
rect 21177 2935 21235 2941
rect 21913 2941 21925 2944
rect 21959 2941 21971 2975
rect 21913 2935 21971 2941
rect 22370 2932 22376 2984
rect 22428 2972 22434 2984
rect 22465 2975 22523 2981
rect 22465 2972 22477 2975
rect 22428 2944 22477 2972
rect 22428 2932 22434 2944
rect 22465 2941 22477 2944
rect 22511 2941 22523 2975
rect 23750 2972 23756 2984
rect 23711 2944 23756 2972
rect 22465 2935 22523 2941
rect 23750 2932 23756 2944
rect 23808 2932 23814 2984
rect 24946 2932 24952 2984
rect 25004 2972 25010 2984
rect 25041 2975 25099 2981
rect 25041 2972 25053 2975
rect 25004 2944 25053 2972
rect 25004 2932 25010 2944
rect 25041 2941 25053 2944
rect 25087 2941 25099 2975
rect 26234 2972 26240 2984
rect 26195 2944 26240 2972
rect 25041 2935 25099 2941
rect 26234 2932 26240 2944
rect 26292 2932 26298 2984
rect 14734 2864 14740 2916
rect 14792 2904 14798 2916
rect 15718 2907 15776 2913
rect 15718 2904 15730 2907
rect 14792 2876 15730 2904
rect 14792 2864 14798 2876
rect 15718 2873 15730 2876
rect 15764 2904 15776 2907
rect 16666 2904 16672 2916
rect 15764 2876 16672 2904
rect 15764 2873 15776 2876
rect 15718 2867 15776 2873
rect 16666 2864 16672 2876
rect 16724 2864 16730 2916
rect 18690 2904 18696 2916
rect 18651 2876 18696 2904
rect 18690 2864 18696 2876
rect 18748 2864 18754 2916
rect 19702 2904 19708 2916
rect 18984 2876 19708 2904
rect 14921 2839 14979 2845
rect 14921 2836 14933 2839
rect 12912 2808 14933 2836
rect 11609 2799 11667 2805
rect 14921 2805 14933 2808
rect 14967 2836 14979 2839
rect 15197 2839 15255 2845
rect 15197 2836 15209 2839
rect 14967 2808 15209 2836
rect 14967 2805 14979 2808
rect 14921 2799 14979 2805
rect 15197 2805 15209 2808
rect 15243 2805 15255 2839
rect 15197 2799 15255 2805
rect 18601 2839 18659 2845
rect 18601 2805 18613 2839
rect 18647 2836 18659 2839
rect 18984 2836 19012 2876
rect 19702 2864 19708 2876
rect 19760 2864 19766 2916
rect 18647 2808 19012 2836
rect 19337 2839 19395 2845
rect 18647 2805 18659 2808
rect 18601 2799 18659 2805
rect 19337 2805 19349 2839
rect 19383 2836 19395 2839
rect 20162 2836 20168 2848
rect 19383 2808 20168 2836
rect 19383 2805 19395 2808
rect 19337 2799 19395 2805
rect 20162 2796 20168 2808
rect 20220 2796 20226 2848
rect 22646 2836 22652 2848
rect 22607 2808 22652 2836
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1578 2592 1584 2644
rect 1636 2632 1642 2644
rect 1857 2635 1915 2641
rect 1857 2632 1869 2635
rect 1636 2604 1869 2632
rect 1636 2592 1642 2604
rect 1857 2601 1869 2604
rect 1903 2632 1915 2635
rect 3878 2632 3884 2644
rect 1903 2604 2268 2632
rect 3839 2604 3884 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 1397 2567 1455 2573
rect 1397 2533 1409 2567
rect 1443 2564 1455 2567
rect 2130 2564 2136 2576
rect 1443 2536 2136 2564
rect 1443 2533 1455 2536
rect 1397 2527 1455 2533
rect 2130 2524 2136 2536
rect 2188 2524 2194 2576
rect 2240 2428 2268 2604
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 5994 2632 6000 2644
rect 5491 2604 6000 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 7248 2604 7481 2632
rect 7248 2592 7254 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 7926 2632 7932 2644
rect 7469 2595 7527 2601
rect 7576 2604 7932 2632
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 2958 2564 2964 2576
rect 2363 2536 2964 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 2958 2524 2964 2536
rect 3016 2524 3022 2576
rect 3050 2524 3056 2576
rect 3108 2564 3114 2576
rect 3421 2567 3479 2573
rect 3421 2564 3433 2567
rect 3108 2536 3433 2564
rect 3108 2524 3114 2536
rect 3421 2533 3433 2536
rect 3467 2533 3479 2567
rect 3421 2527 3479 2533
rect 3896 2496 3924 2592
rect 4246 2524 4252 2576
rect 4304 2573 4310 2576
rect 7576 2573 7604 2604
rect 7926 2592 7932 2604
rect 7984 2632 7990 2644
rect 8297 2635 8355 2641
rect 8297 2632 8309 2635
rect 7984 2604 8309 2632
rect 7984 2592 7990 2604
rect 8297 2601 8309 2604
rect 8343 2601 8355 2635
rect 9122 2632 9128 2644
rect 9083 2604 9128 2632
rect 8297 2595 8355 2601
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 9398 2592 9404 2644
rect 9456 2632 9462 2644
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 9456 2604 9505 2632
rect 9456 2592 9462 2604
rect 9493 2601 9505 2604
rect 9539 2601 9551 2635
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 9493 2595 9551 2601
rect 4304 2567 4368 2573
rect 4304 2533 4322 2567
rect 4356 2533 4368 2567
rect 4304 2527 4368 2533
rect 7561 2567 7619 2573
rect 7561 2533 7573 2567
rect 7607 2533 7619 2567
rect 7561 2527 7619 2533
rect 4304 2524 4310 2527
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3896 2468 4077 2496
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 6638 2496 6644 2508
rect 6599 2468 6644 2496
rect 4065 2459 4123 2465
rect 6638 2456 6644 2468
rect 6696 2496 6702 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6696 2468 7297 2496
rect 6696 2456 6702 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 7285 2459 7343 2465
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 9508 2496 9536 2595
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 14642 2592 14648 2644
rect 14700 2632 14706 2644
rect 15197 2635 15255 2641
rect 15197 2632 15209 2635
rect 14700 2604 15209 2632
rect 14700 2592 14706 2604
rect 15197 2601 15209 2604
rect 15243 2632 15255 2635
rect 15243 2604 15884 2632
rect 15243 2601 15255 2604
rect 15197 2595 15255 2601
rect 10686 2524 10692 2576
rect 10744 2524 10750 2576
rect 13630 2524 13636 2576
rect 13688 2564 13694 2576
rect 15856 2573 15884 2604
rect 15930 2592 15936 2644
rect 15988 2632 15994 2644
rect 15988 2604 16160 2632
rect 15988 2592 15994 2604
rect 14369 2567 14427 2573
rect 14369 2564 14381 2567
rect 13688 2536 14381 2564
rect 13688 2524 13694 2536
rect 14369 2533 14381 2536
rect 14415 2533 14427 2567
rect 14369 2527 14427 2533
rect 15841 2567 15899 2573
rect 15841 2533 15853 2567
rect 15887 2533 15899 2567
rect 16022 2564 16028 2576
rect 15983 2536 16028 2564
rect 15841 2527 15899 2533
rect 16022 2524 16028 2536
rect 16080 2524 16086 2576
rect 16132 2573 16160 2604
rect 16850 2592 16856 2644
rect 16908 2632 16914 2644
rect 17589 2635 17647 2641
rect 17589 2632 17601 2635
rect 16908 2604 17601 2632
rect 16908 2592 16914 2604
rect 17589 2601 17601 2604
rect 17635 2601 17647 2635
rect 17589 2595 17647 2601
rect 19334 2592 19340 2644
rect 19392 2632 19398 2644
rect 20073 2635 20131 2641
rect 20073 2632 20085 2635
rect 19392 2604 20085 2632
rect 19392 2592 19398 2604
rect 20073 2601 20085 2604
rect 20119 2601 20131 2635
rect 20073 2595 20131 2601
rect 20530 2592 20536 2644
rect 20588 2632 20594 2644
rect 22189 2635 22247 2641
rect 22189 2632 22201 2635
rect 20588 2604 22201 2632
rect 20588 2592 20594 2604
rect 16117 2567 16175 2573
rect 16117 2533 16129 2567
rect 16163 2533 16175 2567
rect 16117 2527 16175 2533
rect 16666 2524 16672 2576
rect 16724 2564 16730 2576
rect 16945 2567 17003 2573
rect 16945 2564 16957 2567
rect 16724 2536 16957 2564
rect 16724 2524 16730 2536
rect 16945 2533 16957 2536
rect 16991 2564 17003 2567
rect 17218 2564 17224 2576
rect 16991 2536 17224 2564
rect 16991 2533 17003 2536
rect 16945 2527 17003 2533
rect 17218 2524 17224 2536
rect 17276 2564 17282 2576
rect 18049 2567 18107 2573
rect 18049 2564 18061 2567
rect 17276 2536 18061 2564
rect 17276 2524 17282 2536
rect 18049 2533 18061 2536
rect 18095 2564 18107 2567
rect 18690 2564 18696 2576
rect 18095 2536 18696 2564
rect 18095 2533 18107 2536
rect 18049 2527 18107 2533
rect 18690 2524 18696 2536
rect 18748 2524 18754 2576
rect 18877 2567 18935 2573
rect 18877 2533 18889 2567
rect 18923 2564 18935 2567
rect 21251 2567 21309 2573
rect 21251 2564 21263 2567
rect 18923 2536 21263 2564
rect 18923 2533 18935 2536
rect 18877 2527 18935 2533
rect 21251 2533 21263 2536
rect 21297 2564 21309 2567
rect 21726 2564 21732 2576
rect 21297 2533 21312 2564
rect 21687 2536 21732 2564
rect 21251 2527 21312 2533
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9508 2468 9781 2496
rect 9769 2465 9781 2468
rect 9815 2465 9827 2499
rect 10025 2499 10083 2505
rect 10025 2496 10037 2499
rect 9769 2459 9827 2465
rect 9876 2468 10037 2496
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2240 2400 2881 2428
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 9122 2388 9128 2440
rect 9180 2428 9186 2440
rect 9876 2428 9904 2468
rect 10025 2465 10037 2468
rect 10071 2496 10083 2499
rect 10704 2496 10732 2524
rect 10071 2468 10732 2496
rect 12621 2499 12679 2505
rect 10071 2465 10083 2468
rect 10025 2459 10083 2465
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 12802 2496 12808 2508
rect 12667 2468 12808 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 12802 2456 12808 2468
rect 12860 2496 12866 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12860 2468 13185 2496
rect 12860 2456 12866 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 14182 2496 14188 2508
rect 14143 2468 14188 2496
rect 13173 2459 13231 2465
rect 14182 2456 14188 2468
rect 14240 2496 14246 2508
rect 14826 2496 14832 2508
rect 14240 2468 14832 2496
rect 14240 2456 14246 2468
rect 14826 2456 14832 2468
rect 14884 2456 14890 2508
rect 16040 2496 16068 2524
rect 16485 2499 16543 2505
rect 16485 2496 16497 2499
rect 16040 2468 16497 2496
rect 16485 2465 16497 2468
rect 16531 2465 16543 2499
rect 16485 2459 16543 2465
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2496 17095 2499
rect 17126 2496 17132 2508
rect 17083 2468 17132 2496
rect 17083 2465 17095 2468
rect 17037 2459 17095 2465
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 18708 2496 18736 2524
rect 18969 2499 19027 2505
rect 18969 2496 18981 2499
rect 18708 2468 18981 2496
rect 18969 2465 18981 2468
rect 19015 2465 19027 2499
rect 18969 2459 19027 2465
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2496 19947 2499
rect 19978 2496 19984 2508
rect 19935 2468 19984 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 20990 2496 20996 2508
rect 20671 2468 20996 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 20990 2456 20996 2468
rect 21048 2456 21054 2508
rect 21284 2496 21312 2527
rect 21726 2524 21732 2536
rect 21784 2524 21790 2576
rect 21836 2573 21864 2604
rect 22189 2601 22201 2604
rect 22235 2601 22247 2635
rect 22189 2595 22247 2601
rect 21821 2567 21879 2573
rect 21821 2533 21833 2567
rect 21867 2533 21879 2567
rect 21821 2527 21879 2533
rect 24210 2524 24216 2576
rect 24268 2564 24274 2576
rect 24305 2567 24363 2573
rect 24305 2564 24317 2567
rect 24268 2536 24317 2564
rect 24268 2524 24274 2536
rect 24305 2533 24317 2536
rect 24351 2533 24363 2567
rect 24305 2527 24363 2533
rect 22557 2499 22615 2505
rect 22557 2496 22569 2499
rect 21284 2468 22569 2496
rect 22557 2465 22569 2468
rect 22603 2465 22615 2499
rect 22557 2459 22615 2465
rect 22741 2499 22799 2505
rect 22741 2465 22753 2499
rect 22787 2496 22799 2499
rect 22922 2496 22928 2508
rect 22787 2468 22928 2496
rect 22787 2465 22799 2468
rect 22741 2459 22799 2465
rect 22922 2456 22928 2468
rect 22980 2496 22986 2508
rect 23293 2499 23351 2505
rect 23293 2496 23305 2499
rect 22980 2468 23305 2496
rect 22980 2456 22986 2468
rect 23293 2465 23305 2468
rect 23339 2465 23351 2499
rect 23293 2459 23351 2465
rect 23474 2456 23480 2508
rect 23532 2496 23538 2508
rect 24029 2499 24087 2505
rect 24029 2496 24041 2499
rect 23532 2468 24041 2496
rect 23532 2456 23538 2468
rect 24029 2465 24041 2468
rect 24075 2496 24087 2499
rect 24765 2499 24823 2505
rect 24765 2496 24777 2499
rect 24075 2468 24777 2496
rect 24075 2465 24087 2468
rect 24029 2459 24087 2465
rect 24765 2465 24777 2468
rect 24811 2465 24823 2499
rect 25130 2496 25136 2508
rect 25091 2468 25136 2496
rect 24765 2459 24823 2465
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 25317 2499 25375 2505
rect 25317 2465 25329 2499
rect 25363 2496 25375 2499
rect 25869 2499 25927 2505
rect 25869 2496 25881 2499
rect 25363 2468 25881 2496
rect 25363 2465 25375 2468
rect 25317 2459 25375 2465
rect 25869 2465 25881 2468
rect 25915 2465 25927 2499
rect 25869 2459 25927 2465
rect 9180 2400 9904 2428
rect 12437 2431 12495 2437
rect 9180 2388 9186 2400
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 12483 2400 14473 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 14461 2397 14473 2400
rect 14507 2428 14519 2431
rect 15286 2428 15292 2440
rect 14507 2400 15292 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 15286 2388 15292 2400
rect 15344 2388 15350 2440
rect 18782 2428 18788 2440
rect 18743 2400 18788 2428
rect 18782 2388 18788 2400
rect 18840 2388 18846 2440
rect 19705 2431 19763 2437
rect 19705 2397 19717 2431
rect 19751 2428 19763 2431
rect 20162 2428 20168 2440
rect 19751 2400 20168 2428
rect 19751 2397 19763 2400
rect 19705 2391 19763 2397
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 21637 2431 21695 2437
rect 21637 2428 21649 2431
rect 20916 2400 21649 2428
rect 7006 2360 7012 2372
rect 6967 2332 7012 2360
rect 7006 2320 7012 2332
rect 7064 2320 7070 2372
rect 12802 2360 12808 2372
rect 12763 2332 12808 2360
rect 12802 2320 12808 2332
rect 12860 2320 12866 2372
rect 13906 2360 13912 2372
rect 13867 2332 13912 2360
rect 13906 2320 13912 2332
rect 13964 2320 13970 2372
rect 15470 2320 15476 2372
rect 15528 2360 15534 2372
rect 15565 2363 15623 2369
rect 15565 2360 15577 2363
rect 15528 2332 15577 2360
rect 15528 2320 15534 2332
rect 15565 2329 15577 2332
rect 15611 2329 15623 2363
rect 18414 2360 18420 2372
rect 18375 2332 18420 2360
rect 15565 2323 15623 2329
rect 18414 2320 18420 2332
rect 18472 2320 18478 2372
rect 20916 2304 20944 2400
rect 21637 2397 21649 2400
rect 21683 2397 21695 2431
rect 23658 2428 23664 2440
rect 23619 2400 23664 2428
rect 21637 2391 21695 2397
rect 23658 2388 23664 2400
rect 23716 2388 23722 2440
rect 25038 2388 25044 2440
rect 25096 2428 25102 2440
rect 25332 2428 25360 2459
rect 25096 2400 25360 2428
rect 25096 2388 25102 2400
rect 20990 2320 20996 2372
rect 21048 2360 21054 2372
rect 21726 2360 21732 2372
rect 21048 2332 21732 2360
rect 21048 2320 21054 2332
rect 21726 2320 21732 2332
rect 21784 2320 21790 2372
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 8662 2292 8668 2304
rect 8623 2264 8668 2292
rect 8662 2252 8668 2264
rect 8720 2252 8726 2304
rect 11698 2292 11704 2304
rect 11659 2264 11704 2292
rect 11698 2252 11704 2264
rect 11756 2252 11762 2304
rect 13630 2292 13636 2304
rect 13591 2264 13636 2292
rect 13630 2252 13636 2264
rect 13688 2252 13694 2304
rect 17218 2292 17224 2304
rect 17179 2264 17224 2292
rect 17218 2252 17224 2264
rect 17276 2252 17282 2304
rect 20898 2292 20904 2304
rect 20859 2264 20904 2292
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 22922 2292 22928 2304
rect 22883 2264 22928 2292
rect 22922 2252 22928 2264
rect 22980 2252 22986 2304
rect 25498 2292 25504 2304
rect 25459 2264 25504 2292
rect 25498 2252 25504 2264
rect 25556 2252 25562 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 11422 2048 11428 2100
rect 11480 2088 11486 2100
rect 16022 2088 16028 2100
rect 11480 2060 16028 2088
rect 11480 2048 11486 2060
rect 16022 2048 16028 2060
rect 16080 2048 16086 2100
rect 13538 1572 13544 1624
rect 13596 1612 13602 1624
rect 15378 1612 15384 1624
rect 13596 1584 15384 1612
rect 13596 1572 13602 1584
rect 15378 1572 15384 1584
rect 15436 1572 15442 1624
rect 22554 1572 22560 1624
rect 22612 1612 22618 1624
rect 23566 1612 23572 1624
rect 22612 1584 23572 1612
rect 22612 1572 22618 1584
rect 23566 1572 23572 1584
rect 23624 1572 23630 1624
rect 5534 1368 5540 1420
rect 5592 1408 5598 1420
rect 6178 1408 6184 1420
rect 5592 1380 6184 1408
rect 5592 1368 5598 1380
rect 6178 1368 6184 1380
rect 6236 1368 6242 1420
rect 4522 660 4528 672
rect 3160 632 4528 660
rect 3160 604 3188 632
rect 4522 620 4528 632
rect 4580 620 4586 672
rect 3142 552 3148 604
rect 3200 552 3206 604
rect 3694 552 3700 604
rect 3752 592 3758 604
rect 3786 592 3792 604
rect 3752 564 3792 592
rect 3752 552 3758 564
rect 3786 552 3792 564
rect 3844 552 3850 604
rect 12158 552 12164 604
rect 12216 592 12222 604
rect 12526 592 12532 604
rect 12216 564 12532 592
rect 12216 552 12222 564
rect 12526 552 12532 564
rect 12584 552 12590 604
rect 18874 552 18880 604
rect 18932 592 18938 604
rect 18966 592 18972 604
rect 18932 564 18972 592
rect 18932 552 18938 564
rect 18966 552 18972 564
rect 19024 552 19030 604
<< via1 >>
rect 22008 26596 22060 26648
rect 23572 26596 23624 26648
rect 14648 26392 14700 26444
rect 23480 26392 23532 26444
rect 3424 26256 3476 26308
rect 11244 26256 11296 26308
rect 22192 26256 22244 26308
rect 23480 26256 23532 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 3056 24828 3108 24880
rect 15936 24828 15988 24880
rect 21180 24828 21232 24880
rect 23480 24828 23532 24880
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 23848 19796 23900 19848
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 23756 19252 23808 19304
rect 26884 19116 26936 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 23480 18819 23532 18828
rect 23480 18785 23489 18819
rect 23489 18785 23523 18819
rect 23523 18785 23532 18819
rect 23480 18776 23532 18785
rect 24584 18819 24636 18828
rect 24584 18785 24593 18819
rect 24593 18785 24627 18819
rect 24627 18785 24636 18819
rect 24584 18776 24636 18785
rect 22836 18708 22888 18760
rect 24124 18572 24176 18624
rect 24216 18572 24268 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 24676 18368 24728 18420
rect 756 18028 808 18080
rect 2044 18071 2096 18080
rect 2044 18037 2053 18071
rect 2053 18037 2087 18071
rect 2087 18037 2096 18071
rect 2044 18028 2096 18037
rect 20168 18071 20220 18080
rect 20168 18037 20177 18071
rect 20177 18037 20211 18071
rect 20211 18037 20220 18071
rect 20168 18028 20220 18037
rect 22376 18028 22428 18080
rect 23296 18028 23348 18080
rect 23480 18028 23532 18080
rect 24032 18028 24084 18080
rect 25412 18028 25464 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 23388 17824 23440 17876
rect 2504 17731 2556 17740
rect 2504 17697 2513 17731
rect 2513 17697 2547 17731
rect 2547 17697 2556 17731
rect 2504 17688 2556 17697
rect 22468 17688 22520 17740
rect 24676 17688 24728 17740
rect 2044 17663 2096 17672
rect 2044 17629 2053 17663
rect 2053 17629 2087 17663
rect 2087 17629 2096 17663
rect 2044 17620 2096 17629
rect 19524 17663 19576 17672
rect 19524 17629 19533 17663
rect 19533 17629 19567 17663
rect 19567 17629 19576 17663
rect 19524 17620 19576 17629
rect 21732 17620 21784 17672
rect 23020 17663 23072 17672
rect 23020 17629 23029 17663
rect 23029 17629 23063 17663
rect 23063 17629 23072 17663
rect 23020 17620 23072 17629
rect 664 17484 716 17536
rect 2596 17484 2648 17536
rect 22560 17484 22612 17536
rect 23572 17484 23624 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2504 17280 2556 17332
rect 22468 17280 22520 17332
rect 2320 17212 2372 17264
rect 23020 17144 23072 17196
rect 1860 16940 1912 16992
rect 25780 17212 25832 17264
rect 24124 17076 24176 17128
rect 22652 17051 22704 17060
rect 2688 16940 2740 16992
rect 3148 16983 3200 16992
rect 3148 16949 3157 16983
rect 3157 16949 3191 16983
rect 3191 16949 3200 16983
rect 3148 16940 3200 16949
rect 20536 16940 20588 16992
rect 20812 16983 20864 16992
rect 20812 16949 20821 16983
rect 20821 16949 20855 16983
rect 20855 16949 20864 16983
rect 20812 16940 20864 16949
rect 21088 16983 21140 16992
rect 21088 16949 21097 16983
rect 21097 16949 21131 16983
rect 21131 16949 21140 16983
rect 21088 16940 21140 16949
rect 21824 16983 21876 16992
rect 21824 16949 21833 16983
rect 21833 16949 21867 16983
rect 21867 16949 21876 16983
rect 22652 17017 22661 17051
rect 22661 17017 22695 17051
rect 22695 17017 22704 17051
rect 22652 17008 22704 17017
rect 23480 17008 23532 17060
rect 22560 16983 22612 16992
rect 21824 16940 21876 16949
rect 22560 16949 22569 16983
rect 22569 16949 22603 16983
rect 22603 16949 22612 16983
rect 22560 16940 22612 16949
rect 23664 16940 23716 16992
rect 24676 16940 24728 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2044 16779 2096 16788
rect 2044 16745 2053 16779
rect 2053 16745 2087 16779
rect 2087 16745 2096 16779
rect 2044 16736 2096 16745
rect 2136 16736 2188 16788
rect 21824 16736 21876 16788
rect 22652 16736 22704 16788
rect 23940 16779 23992 16788
rect 23940 16745 23949 16779
rect 23949 16745 23983 16779
rect 23983 16745 23992 16779
rect 23940 16736 23992 16745
rect 25964 16736 26016 16788
rect 4896 16668 4948 16720
rect 23020 16668 23072 16720
rect 2504 16643 2556 16652
rect 2504 16609 2513 16643
rect 2513 16609 2547 16643
rect 2547 16609 2556 16643
rect 2504 16600 2556 16609
rect 2688 16600 2740 16652
rect 4068 16600 4120 16652
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 10140 16600 10192 16652
rect 15752 16600 15804 16652
rect 17868 16600 17920 16652
rect 18788 16643 18840 16652
rect 18788 16609 18797 16643
rect 18797 16609 18831 16643
rect 18831 16609 18840 16643
rect 18788 16600 18840 16609
rect 21824 16600 21876 16652
rect 23388 16600 23440 16652
rect 25320 16600 25372 16652
rect 5264 16532 5316 16584
rect 22560 16575 22612 16584
rect 22560 16541 22569 16575
rect 22569 16541 22603 16575
rect 22603 16541 22612 16575
rect 22560 16532 22612 16541
rect 21548 16464 21600 16516
rect 1216 16396 1268 16448
rect 2872 16396 2924 16448
rect 2964 16396 3016 16448
rect 10968 16396 11020 16448
rect 14832 16396 14884 16448
rect 21272 16396 21324 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 4068 16192 4120 16244
rect 23020 16192 23072 16244
rect 2228 16124 2280 16176
rect 4804 16124 4856 16176
rect 11796 16124 11848 16176
rect 15660 16124 15712 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 10692 15988 10744 16040
rect 11888 15988 11940 16040
rect 4068 15920 4120 15972
rect 4344 15920 4396 15972
rect 4620 15963 4672 15972
rect 4620 15929 4629 15963
rect 4629 15929 4663 15963
rect 4663 15929 4672 15963
rect 4620 15920 4672 15929
rect 4712 15963 4764 15972
rect 4712 15929 4721 15963
rect 4721 15929 4755 15963
rect 4755 15929 4764 15963
rect 4712 15920 4764 15929
rect 9956 15963 10008 15972
rect 9956 15929 9965 15963
rect 9965 15929 9999 15963
rect 9999 15929 10008 15963
rect 9956 15920 10008 15929
rect 10968 15963 11020 15972
rect 10968 15929 10977 15963
rect 10977 15929 11011 15963
rect 11011 15929 11020 15963
rect 10968 15920 11020 15929
rect 14556 15963 14608 15972
rect 14556 15929 14565 15963
rect 14565 15929 14599 15963
rect 14599 15929 14608 15963
rect 14556 15920 14608 15929
rect 14740 15963 14792 15972
rect 14740 15929 14749 15963
rect 14749 15929 14783 15963
rect 14783 15929 14792 15963
rect 14740 15920 14792 15929
rect 21548 15920 21600 15972
rect 2504 15852 2556 15904
rect 4896 15852 4948 15904
rect 5264 15852 5316 15904
rect 6552 15852 6604 15904
rect 6828 15852 6880 15904
rect 16488 15852 16540 15904
rect 18972 15895 19024 15904
rect 18972 15861 18981 15895
rect 18981 15861 19015 15895
rect 19015 15861 19024 15895
rect 18972 15852 19024 15861
rect 20444 15852 20496 15904
rect 20628 15895 20680 15904
rect 20628 15861 20637 15895
rect 20637 15861 20671 15895
rect 20671 15861 20680 15895
rect 20628 15852 20680 15861
rect 20904 15895 20956 15904
rect 20904 15861 20913 15895
rect 20913 15861 20947 15895
rect 20947 15861 20956 15895
rect 20904 15852 20956 15861
rect 22560 15852 22612 15904
rect 23112 15895 23164 15904
rect 23112 15861 23121 15895
rect 23121 15861 23155 15895
rect 23155 15861 23164 15895
rect 23940 16031 23992 16040
rect 23940 15997 23974 16031
rect 23974 15997 23992 16031
rect 23940 15988 23992 15997
rect 23112 15852 23164 15861
rect 25044 15895 25096 15904
rect 25044 15861 25053 15895
rect 25053 15861 25087 15895
rect 25087 15861 25096 15895
rect 25044 15852 25096 15861
rect 25320 15852 25372 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2964 15691 3016 15700
rect 2964 15657 2973 15691
rect 2973 15657 3007 15691
rect 3007 15657 3016 15691
rect 2964 15648 3016 15657
rect 11888 15691 11940 15700
rect 11888 15657 11897 15691
rect 11897 15657 11931 15691
rect 11931 15657 11940 15691
rect 11888 15648 11940 15657
rect 14556 15648 14608 15700
rect 19984 15648 20036 15700
rect 23020 15648 23072 15700
rect 23940 15648 23992 15700
rect 4896 15623 4948 15632
rect 4896 15589 4905 15623
rect 4905 15589 4939 15623
rect 4939 15589 4948 15623
rect 4896 15580 4948 15589
rect 5448 15580 5500 15632
rect 10600 15580 10652 15632
rect 15660 15623 15712 15632
rect 15660 15589 15669 15623
rect 15669 15589 15703 15623
rect 15703 15589 15712 15623
rect 15660 15580 15712 15589
rect 15844 15623 15896 15632
rect 15844 15589 15853 15623
rect 15853 15589 15887 15623
rect 15887 15589 15896 15623
rect 15844 15580 15896 15589
rect 21824 15580 21876 15632
rect 16580 15512 16632 15564
rect 18144 15555 18196 15564
rect 18144 15521 18153 15555
rect 18153 15521 18187 15555
rect 18187 15521 18196 15555
rect 18144 15512 18196 15521
rect 19340 15512 19392 15564
rect 20996 15512 21048 15564
rect 25044 15512 25096 15564
rect 1860 15444 1912 15496
rect 2504 15444 2556 15496
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 4896 15487 4948 15496
rect 4896 15453 4905 15487
rect 4905 15453 4939 15487
rect 4939 15453 4948 15487
rect 4896 15444 4948 15453
rect 5080 15444 5132 15496
rect 5540 15444 5592 15496
rect 7012 15487 7064 15496
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 8484 15487 8536 15496
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 13084 15444 13136 15496
rect 15476 15444 15528 15496
rect 17592 15444 17644 15496
rect 19432 15444 19484 15496
rect 20904 15487 20956 15496
rect 20904 15453 20913 15487
rect 20913 15453 20947 15487
rect 20947 15453 20956 15487
rect 20904 15444 20956 15453
rect 23940 15487 23992 15496
rect 23940 15453 23949 15487
rect 23949 15453 23983 15487
rect 23983 15453 23992 15487
rect 23940 15444 23992 15453
rect 3424 15376 3476 15428
rect 4068 15376 4120 15428
rect 4620 15376 4672 15428
rect 6276 15376 6328 15428
rect 20720 15376 20772 15428
rect 1860 15351 1912 15360
rect 1860 15317 1869 15351
rect 1869 15317 1903 15351
rect 1903 15317 1912 15351
rect 1860 15308 1912 15317
rect 2596 15308 2648 15360
rect 4344 15308 4396 15360
rect 5356 15351 5408 15360
rect 5356 15317 5365 15351
rect 5365 15317 5399 15351
rect 5399 15317 5408 15351
rect 5356 15308 5408 15317
rect 6000 15308 6052 15360
rect 6460 15351 6512 15360
rect 6460 15317 6469 15351
rect 6469 15317 6503 15351
rect 6503 15317 6512 15351
rect 6460 15308 6512 15317
rect 12992 15308 13044 15360
rect 15384 15351 15436 15360
rect 15384 15317 15393 15351
rect 15393 15317 15427 15351
rect 15427 15317 15436 15351
rect 15384 15308 15436 15317
rect 18328 15351 18380 15360
rect 18328 15317 18337 15351
rect 18337 15317 18371 15351
rect 18371 15317 18380 15351
rect 18328 15308 18380 15317
rect 20352 15351 20404 15360
rect 20352 15317 20361 15351
rect 20361 15317 20395 15351
rect 20395 15317 20404 15351
rect 20352 15308 20404 15317
rect 21548 15308 21600 15360
rect 22560 15308 22612 15360
rect 24952 15308 25004 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2872 15147 2924 15156
rect 2872 15113 2881 15147
rect 2881 15113 2915 15147
rect 2915 15113 2924 15147
rect 2872 15104 2924 15113
rect 4712 15104 4764 15156
rect 5448 15104 5500 15156
rect 9680 15147 9732 15156
rect 9680 15113 9689 15147
rect 9689 15113 9723 15147
rect 9723 15113 9732 15147
rect 9680 15104 9732 15113
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 15476 15104 15528 15156
rect 16396 15104 16448 15156
rect 16580 15104 16632 15156
rect 19248 15104 19300 15156
rect 19432 15104 19484 15156
rect 20996 15147 21048 15156
rect 20996 15113 21005 15147
rect 21005 15113 21039 15147
rect 21039 15113 21048 15147
rect 20996 15104 21048 15113
rect 1768 14968 1820 15020
rect 13912 15036 13964 15088
rect 24676 15036 24728 15088
rect 10600 14968 10652 15020
rect 11152 14968 11204 15020
rect 5264 14900 5316 14952
rect 2044 14875 2096 14884
rect 2044 14841 2053 14875
rect 2053 14841 2087 14875
rect 2087 14841 2096 14875
rect 2044 14832 2096 14841
rect 3148 14832 3200 14884
rect 6736 14832 6788 14884
rect 1584 14807 1636 14816
rect 1584 14773 1593 14807
rect 1593 14773 1627 14807
rect 1627 14773 1636 14807
rect 1584 14764 1636 14773
rect 4988 14807 5040 14816
rect 4988 14773 4997 14807
rect 4997 14773 5031 14807
rect 5031 14773 5040 14807
rect 4988 14764 5040 14773
rect 6644 14807 6696 14816
rect 6644 14773 6653 14807
rect 6653 14773 6687 14807
rect 6687 14773 6696 14807
rect 10140 14900 10192 14952
rect 12808 14900 12860 14952
rect 6920 14832 6972 14884
rect 9680 14832 9732 14884
rect 10508 14832 10560 14884
rect 12348 14832 12400 14884
rect 12992 14875 13044 14884
rect 12992 14841 13001 14875
rect 13001 14841 13035 14875
rect 13035 14841 13044 14875
rect 12992 14832 13044 14841
rect 6644 14764 6696 14773
rect 7840 14764 7892 14816
rect 9128 14764 9180 14816
rect 11888 14764 11940 14816
rect 14556 14968 14608 15020
rect 25044 15011 25096 15020
rect 25044 14977 25053 15011
rect 25053 14977 25087 15011
rect 25087 14977 25096 15011
rect 25044 14968 25096 14977
rect 15108 14943 15160 14952
rect 15108 14909 15117 14943
rect 15117 14909 15151 14943
rect 15151 14909 15160 14943
rect 15108 14900 15160 14909
rect 18236 14900 18288 14952
rect 19432 14900 19484 14952
rect 20904 14900 20956 14952
rect 22100 14943 22152 14952
rect 22100 14909 22109 14943
rect 22109 14909 22143 14943
rect 22143 14909 22152 14943
rect 22100 14900 22152 14909
rect 14832 14832 14884 14884
rect 15660 14832 15712 14884
rect 18144 14832 18196 14884
rect 19248 14832 19300 14884
rect 20352 14832 20404 14884
rect 23296 14832 23348 14884
rect 24308 14875 24360 14884
rect 24308 14841 24317 14875
rect 24317 14841 24351 14875
rect 24351 14841 24360 14875
rect 24308 14832 24360 14841
rect 24860 14832 24912 14884
rect 15108 14764 15160 14816
rect 15568 14764 15620 14816
rect 18696 14807 18748 14816
rect 18696 14773 18705 14807
rect 18705 14773 18739 14807
rect 18739 14773 18748 14807
rect 18696 14764 18748 14773
rect 20628 14764 20680 14816
rect 22652 14764 22704 14816
rect 23112 14764 23164 14816
rect 23940 14764 23992 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2780 14535 2832 14544
rect 2780 14501 2789 14535
rect 2789 14501 2823 14535
rect 2823 14501 2832 14535
rect 3148 14560 3200 14612
rect 5080 14560 5132 14612
rect 7196 14560 7248 14612
rect 10140 14560 10192 14612
rect 10692 14560 10744 14612
rect 11336 14560 11388 14612
rect 15660 14560 15712 14612
rect 19984 14560 20036 14612
rect 20720 14603 20772 14612
rect 20720 14569 20729 14603
rect 20729 14569 20763 14603
rect 20763 14569 20772 14603
rect 20720 14560 20772 14569
rect 22100 14603 22152 14612
rect 22100 14569 22109 14603
rect 22109 14569 22143 14603
rect 22143 14569 22152 14603
rect 22100 14560 22152 14569
rect 25044 14560 25096 14612
rect 2780 14492 2832 14501
rect 4712 14492 4764 14544
rect 7012 14492 7064 14544
rect 7840 14535 7892 14544
rect 7840 14501 7849 14535
rect 7849 14501 7883 14535
rect 7883 14501 7892 14535
rect 7840 14492 7892 14501
rect 11060 14492 11112 14544
rect 3332 14424 3384 14476
rect 10876 14424 10928 14476
rect 11796 14492 11848 14544
rect 12716 14535 12768 14544
rect 12716 14501 12725 14535
rect 12725 14501 12759 14535
rect 12759 14501 12768 14535
rect 12716 14492 12768 14501
rect 16396 14492 16448 14544
rect 16580 14535 16632 14544
rect 16580 14501 16592 14535
rect 16592 14501 16632 14535
rect 16580 14492 16632 14501
rect 20536 14492 20588 14544
rect 21364 14492 21416 14544
rect 2596 14356 2648 14408
rect 2872 14356 2924 14408
rect 4620 14356 4672 14408
rect 11152 14356 11204 14408
rect 15568 14424 15620 14476
rect 16948 14424 17000 14476
rect 20076 14424 20128 14476
rect 24308 14492 24360 14544
rect 25320 14535 25372 14544
rect 25320 14501 25329 14535
rect 25329 14501 25363 14535
rect 25363 14501 25372 14535
rect 25320 14492 25372 14501
rect 12716 14399 12768 14408
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 12992 14356 13044 14408
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 18420 14356 18472 14408
rect 22652 14424 22704 14476
rect 23112 14424 23164 14476
rect 25044 14467 25096 14476
rect 25044 14433 25053 14467
rect 25053 14433 25087 14467
rect 25087 14433 25096 14467
rect 25044 14424 25096 14433
rect 20720 14356 20772 14408
rect 21548 14399 21600 14408
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 1400 14220 1452 14272
rect 2044 14220 2096 14272
rect 3148 14288 3200 14340
rect 7288 14331 7340 14340
rect 7288 14297 7297 14331
rect 7297 14297 7331 14331
rect 7331 14297 7340 14331
rect 7288 14288 7340 14297
rect 10968 14288 11020 14340
rect 14740 14288 14792 14340
rect 15844 14288 15896 14340
rect 22100 14288 22152 14340
rect 2688 14220 2740 14272
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 4252 14220 4304 14229
rect 6092 14263 6144 14272
rect 6092 14229 6101 14263
rect 6101 14229 6135 14263
rect 6135 14229 6144 14263
rect 6092 14220 6144 14229
rect 6920 14220 6972 14272
rect 8392 14220 8444 14272
rect 8576 14263 8628 14272
rect 8576 14229 8585 14263
rect 8585 14229 8619 14263
rect 8619 14229 8628 14263
rect 8576 14220 8628 14229
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 9220 14220 9272 14272
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 11612 14220 11664 14229
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 12256 14263 12308 14272
rect 12256 14229 12265 14263
rect 12265 14229 12299 14263
rect 12299 14229 12308 14263
rect 12256 14220 12308 14229
rect 12440 14220 12492 14272
rect 13176 14263 13228 14272
rect 13176 14229 13185 14263
rect 13185 14229 13219 14263
rect 13219 14229 13228 14263
rect 13176 14220 13228 14229
rect 17684 14263 17736 14272
rect 17684 14229 17693 14263
rect 17693 14229 17727 14263
rect 17727 14229 17736 14263
rect 17684 14220 17736 14229
rect 18236 14220 18288 14272
rect 19892 14263 19944 14272
rect 19892 14229 19901 14263
rect 19901 14229 19935 14263
rect 19935 14229 19944 14263
rect 19892 14220 19944 14229
rect 19984 14220 20036 14272
rect 20904 14220 20956 14272
rect 23664 14220 23716 14272
rect 23940 14263 23992 14272
rect 23940 14229 23949 14263
rect 23949 14229 23983 14263
rect 23983 14229 23992 14263
rect 23940 14220 23992 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2780 14016 2832 14068
rect 4344 14059 4396 14068
rect 4344 14025 4353 14059
rect 4353 14025 4387 14059
rect 4387 14025 4396 14059
rect 4344 14016 4396 14025
rect 4712 14016 4764 14068
rect 6644 14016 6696 14068
rect 7196 14059 7248 14068
rect 7196 14025 7205 14059
rect 7205 14025 7239 14059
rect 7239 14025 7248 14059
rect 7196 14016 7248 14025
rect 10784 14059 10836 14068
rect 10784 14025 10793 14059
rect 10793 14025 10827 14059
rect 10827 14025 10836 14059
rect 10784 14016 10836 14025
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 12716 14016 12768 14068
rect 12808 14016 12860 14068
rect 3148 13991 3200 14000
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 3148 13957 3157 13991
rect 3157 13957 3191 13991
rect 3191 13957 3200 13991
rect 3148 13948 3200 13957
rect 4620 13948 4672 14000
rect 11152 13948 11204 14000
rect 11336 13948 11388 14000
rect 12440 13948 12492 14000
rect 3332 13880 3384 13932
rect 5080 13880 5132 13932
rect 6644 13880 6696 13932
rect 2044 13855 2096 13864
rect 2044 13821 2078 13855
rect 2078 13821 2096 13855
rect 2044 13812 2096 13821
rect 4344 13812 4396 13864
rect 10968 13880 11020 13932
rect 11612 13880 11664 13932
rect 13544 13880 13596 13932
rect 15568 14016 15620 14068
rect 15660 14016 15712 14068
rect 21364 14059 21416 14068
rect 21364 14025 21373 14059
rect 21373 14025 21407 14059
rect 21407 14025 21416 14059
rect 21364 14016 21416 14025
rect 21732 14016 21784 14068
rect 19340 13948 19392 14000
rect 20628 13948 20680 14000
rect 23388 14016 23440 14068
rect 23848 14016 23900 14068
rect 24860 14016 24912 14068
rect 22100 13991 22152 14000
rect 22100 13957 22109 13991
rect 22109 13957 22143 13991
rect 22143 13957 22152 13991
rect 22100 13948 22152 13957
rect 23020 13880 23072 13932
rect 23940 13880 23992 13932
rect 7840 13812 7892 13864
rect 7656 13744 7708 13796
rect 11060 13744 11112 13796
rect 12256 13812 12308 13864
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 13176 13812 13228 13864
rect 11336 13787 11388 13796
rect 11336 13753 11345 13787
rect 11345 13753 11379 13787
rect 11379 13753 11388 13787
rect 11336 13744 11388 13753
rect 14832 13744 14884 13796
rect 18328 13855 18380 13864
rect 18328 13821 18337 13855
rect 18337 13821 18371 13855
rect 18371 13821 18380 13855
rect 18328 13812 18380 13821
rect 19432 13855 19484 13864
rect 19432 13821 19441 13855
rect 19441 13821 19475 13855
rect 19475 13821 19484 13855
rect 24124 13855 24176 13864
rect 19432 13812 19484 13821
rect 19156 13744 19208 13796
rect 1216 13676 1268 13728
rect 1492 13676 1544 13728
rect 4160 13719 4212 13728
rect 4160 13685 4169 13719
rect 4169 13685 4203 13719
rect 4203 13685 4212 13719
rect 4160 13676 4212 13685
rect 4988 13676 5040 13728
rect 6920 13676 6972 13728
rect 7472 13676 7524 13728
rect 7840 13676 7892 13728
rect 10784 13676 10836 13728
rect 14372 13719 14424 13728
rect 14372 13685 14381 13719
rect 14381 13685 14415 13719
rect 14415 13685 14424 13719
rect 14372 13676 14424 13685
rect 16212 13676 16264 13728
rect 16396 13676 16448 13728
rect 16948 13719 17000 13728
rect 16948 13685 16957 13719
rect 16957 13685 16991 13719
rect 16991 13685 17000 13719
rect 16948 13676 17000 13685
rect 17224 13676 17276 13728
rect 24124 13821 24133 13855
rect 24133 13821 24167 13855
rect 24167 13821 24176 13855
rect 24124 13812 24176 13821
rect 22100 13744 22152 13796
rect 22560 13787 22612 13796
rect 22560 13753 22569 13787
rect 22569 13753 22603 13787
rect 22603 13753 22612 13787
rect 22560 13744 22612 13753
rect 24952 13812 25004 13864
rect 19984 13676 20036 13728
rect 22744 13676 22796 13728
rect 24124 13676 24176 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1400 13472 1452 13524
rect 1768 13515 1820 13524
rect 1768 13481 1777 13515
rect 1777 13481 1811 13515
rect 1811 13481 1820 13515
rect 1768 13472 1820 13481
rect 4712 13472 4764 13524
rect 5080 13515 5132 13524
rect 5080 13481 5089 13515
rect 5089 13481 5123 13515
rect 5123 13481 5132 13515
rect 5080 13472 5132 13481
rect 5448 13472 5500 13524
rect 6644 13515 6696 13524
rect 6644 13481 6653 13515
rect 6653 13481 6687 13515
rect 6687 13481 6696 13515
rect 6644 13472 6696 13481
rect 7012 13515 7064 13524
rect 7012 13481 7021 13515
rect 7021 13481 7055 13515
rect 7055 13481 7064 13515
rect 7012 13472 7064 13481
rect 2780 13447 2832 13456
rect 2780 13413 2789 13447
rect 2789 13413 2823 13447
rect 2823 13413 2832 13447
rect 4620 13447 4672 13456
rect 2780 13404 2832 13413
rect 4620 13413 4629 13447
rect 4629 13413 4663 13447
rect 4663 13413 4672 13447
rect 6000 13447 6052 13456
rect 4620 13404 4672 13413
rect 6000 13413 6009 13447
rect 6009 13413 6043 13447
rect 6043 13413 6052 13447
rect 6000 13404 6052 13413
rect 7196 13404 7248 13456
rect 11152 13472 11204 13524
rect 15660 13472 15712 13524
rect 16396 13472 16448 13524
rect 16580 13515 16632 13524
rect 16580 13481 16589 13515
rect 16589 13481 16623 13515
rect 16623 13481 16632 13515
rect 16580 13472 16632 13481
rect 20076 13472 20128 13524
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 21180 13472 21232 13524
rect 24676 13515 24728 13524
rect 24676 13481 24685 13515
rect 24685 13481 24719 13515
rect 24719 13481 24728 13515
rect 24676 13472 24728 13481
rect 7748 13447 7800 13456
rect 7748 13413 7757 13447
rect 7757 13413 7791 13447
rect 7791 13413 7800 13447
rect 7748 13404 7800 13413
rect 1676 13336 1728 13388
rect 3516 13336 3568 13388
rect 5448 13336 5500 13388
rect 7564 13379 7616 13388
rect 7564 13345 7573 13379
rect 7573 13345 7607 13379
rect 7607 13345 7616 13379
rect 7564 13336 7616 13345
rect 7840 13379 7892 13388
rect 7840 13345 7849 13379
rect 7849 13345 7883 13379
rect 7883 13345 7892 13379
rect 7840 13336 7892 13345
rect 9404 13336 9456 13388
rect 12440 13336 12492 13388
rect 13544 13404 13596 13456
rect 16212 13447 16264 13456
rect 16212 13413 16221 13447
rect 16221 13413 16255 13447
rect 16255 13413 16264 13447
rect 16212 13404 16264 13413
rect 17684 13404 17736 13456
rect 12808 13336 12860 13388
rect 17224 13336 17276 13388
rect 20352 13336 20404 13388
rect 22192 13404 22244 13456
rect 23020 13447 23072 13456
rect 23020 13413 23054 13447
rect 23054 13413 23072 13447
rect 23020 13404 23072 13413
rect 25228 13379 25280 13388
rect 25228 13345 25237 13379
rect 25237 13345 25271 13379
rect 25271 13345 25280 13379
rect 25228 13336 25280 13345
rect 2688 13132 2740 13184
rect 4068 13268 4120 13320
rect 5080 13268 5132 13320
rect 6184 13268 6236 13320
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 15844 13268 15896 13320
rect 16304 13268 16356 13320
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 22560 13268 22612 13320
rect 22744 13311 22796 13320
rect 22744 13277 22753 13311
rect 22753 13277 22787 13311
rect 22787 13277 22796 13311
rect 22744 13268 22796 13277
rect 4160 13243 4212 13252
rect 4160 13209 4169 13243
rect 4169 13209 4203 13243
rect 4203 13209 4212 13243
rect 4160 13200 4212 13209
rect 5356 13200 5408 13252
rect 5724 13243 5776 13252
rect 5724 13209 5733 13243
rect 5733 13209 5767 13243
rect 5767 13209 5776 13243
rect 5724 13200 5776 13209
rect 8208 13200 8260 13252
rect 16672 13200 16724 13252
rect 3148 13132 3200 13184
rect 3332 13132 3384 13184
rect 8300 13175 8352 13184
rect 8300 13141 8309 13175
rect 8309 13141 8343 13175
rect 8343 13141 8352 13175
rect 8300 13132 8352 13141
rect 9680 13132 9732 13184
rect 14188 13132 14240 13184
rect 14832 13132 14884 13184
rect 18512 13175 18564 13184
rect 18512 13141 18521 13175
rect 18521 13141 18555 13175
rect 18555 13141 18564 13175
rect 18512 13132 18564 13141
rect 19156 13132 19208 13184
rect 20076 13132 20128 13184
rect 20996 13175 21048 13184
rect 20996 13141 21005 13175
rect 21005 13141 21039 13175
rect 21039 13141 21048 13175
rect 20996 13132 21048 13141
rect 23112 13132 23164 13184
rect 24124 13175 24176 13184
rect 24124 13141 24133 13175
rect 24133 13141 24167 13175
rect 24167 13141 24176 13175
rect 24124 13132 24176 13141
rect 25044 13175 25096 13184
rect 25044 13141 25053 13175
rect 25053 13141 25087 13175
rect 25087 13141 25096 13175
rect 25044 13132 25096 13141
rect 26148 13132 26200 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1676 12971 1728 12980
rect 1676 12937 1685 12971
rect 1685 12937 1719 12971
rect 1719 12937 1728 12971
rect 1676 12928 1728 12937
rect 1860 12928 1912 12980
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 4620 12971 4672 12980
rect 4620 12937 4629 12971
rect 4629 12937 4663 12971
rect 4663 12937 4672 12971
rect 4620 12928 4672 12937
rect 5264 12971 5316 12980
rect 5264 12937 5273 12971
rect 5273 12937 5307 12971
rect 5307 12937 5316 12971
rect 5264 12928 5316 12937
rect 1952 12792 2004 12844
rect 3332 12860 3384 12912
rect 2504 12792 2556 12844
rect 2872 12792 2924 12844
rect 4160 12835 4212 12844
rect 4160 12801 4169 12835
rect 4169 12801 4203 12835
rect 4203 12801 4212 12835
rect 4160 12792 4212 12801
rect 4712 12792 4764 12844
rect 5724 12792 5776 12844
rect 4436 12724 4488 12776
rect 4620 12724 4672 12776
rect 6092 12724 6144 12776
rect 7840 12928 7892 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 10968 12928 11020 12980
rect 13544 12971 13596 12980
rect 13544 12937 13553 12971
rect 13553 12937 13587 12971
rect 13587 12937 13596 12971
rect 13544 12928 13596 12937
rect 14740 12928 14792 12980
rect 15936 12971 15988 12980
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 21180 12928 21232 12980
rect 22192 12971 22244 12980
rect 22192 12937 22201 12971
rect 22201 12937 22235 12971
rect 22235 12937 22244 12971
rect 22192 12928 22244 12937
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 25044 12928 25096 12980
rect 25228 12971 25280 12980
rect 25228 12937 25237 12971
rect 25237 12937 25271 12971
rect 25271 12937 25280 12971
rect 25228 12928 25280 12937
rect 25688 12971 25740 12980
rect 25688 12937 25697 12971
rect 25697 12937 25731 12971
rect 25731 12937 25740 12971
rect 25688 12928 25740 12937
rect 12440 12860 12492 12912
rect 14556 12860 14608 12912
rect 14832 12860 14884 12912
rect 15844 12860 15896 12912
rect 16396 12860 16448 12912
rect 19432 12860 19484 12912
rect 7656 12792 7708 12844
rect 11152 12792 11204 12844
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 16580 12835 16632 12844
rect 16580 12801 16589 12835
rect 16589 12801 16623 12835
rect 16623 12801 16632 12835
rect 16580 12792 16632 12801
rect 17684 12792 17736 12844
rect 18512 12792 18564 12844
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 22560 12792 22612 12844
rect 24492 12792 24544 12844
rect 24952 12792 25004 12844
rect 14648 12724 14700 12776
rect 15660 12724 15712 12776
rect 15844 12724 15896 12776
rect 19984 12724 20036 12776
rect 2504 12699 2556 12708
rect 2504 12665 2513 12699
rect 2513 12665 2547 12699
rect 2547 12665 2556 12699
rect 2504 12656 2556 12665
rect 4160 12699 4212 12708
rect 4160 12665 4169 12699
rect 4169 12665 4203 12699
rect 4203 12665 4212 12699
rect 4160 12656 4212 12665
rect 4804 12656 4856 12708
rect 6000 12656 6052 12708
rect 6184 12656 6236 12708
rect 7932 12656 7984 12708
rect 8300 12699 8352 12708
rect 8300 12665 8312 12699
rect 8312 12665 8352 12699
rect 8300 12656 8352 12665
rect 9772 12656 9824 12708
rect 10968 12656 11020 12708
rect 11060 12656 11112 12708
rect 13636 12656 13688 12708
rect 13820 12656 13872 12708
rect 14372 12656 14424 12708
rect 15936 12656 15988 12708
rect 17776 12699 17828 12708
rect 17776 12665 17785 12699
rect 17785 12665 17819 12699
rect 17819 12665 17828 12699
rect 18880 12699 18932 12708
rect 17776 12656 17828 12665
rect 18880 12665 18889 12699
rect 18889 12665 18923 12699
rect 18923 12665 18932 12699
rect 18880 12656 18932 12665
rect 20720 12724 20772 12776
rect 21548 12724 21600 12776
rect 22652 12724 22704 12776
rect 23388 12724 23440 12776
rect 25504 12767 25556 12776
rect 25504 12733 25513 12767
rect 25513 12733 25547 12767
rect 25547 12733 25556 12767
rect 25504 12724 25556 12733
rect 2688 12588 2740 12640
rect 2780 12588 2832 12640
rect 3332 12588 3384 12640
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 10692 12631 10744 12640
rect 10692 12597 10701 12631
rect 10701 12597 10735 12631
rect 10735 12597 10744 12631
rect 11336 12631 11388 12640
rect 10692 12588 10744 12597
rect 11336 12597 11345 12631
rect 11345 12597 11379 12631
rect 11379 12597 11388 12631
rect 11336 12588 11388 12597
rect 11704 12588 11756 12640
rect 17224 12631 17276 12640
rect 17224 12597 17233 12631
rect 17233 12597 17267 12631
rect 17267 12597 17276 12631
rect 17224 12588 17276 12597
rect 19156 12588 19208 12640
rect 21548 12588 21600 12640
rect 22744 12588 22796 12640
rect 24676 12588 24728 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2044 12384 2096 12436
rect 4068 12384 4120 12436
rect 6092 12384 6144 12436
rect 6460 12384 6512 12436
rect 6644 12384 6696 12436
rect 8300 12427 8352 12436
rect 4804 12316 4856 12368
rect 6184 12359 6236 12368
rect 6184 12325 6193 12359
rect 6193 12325 6227 12359
rect 6227 12325 6236 12359
rect 6184 12316 6236 12325
rect 7104 12316 7156 12368
rect 7288 12316 7340 12368
rect 7656 12316 7708 12368
rect 8300 12393 8309 12427
rect 8309 12393 8343 12427
rect 8343 12393 8352 12427
rect 8300 12384 8352 12393
rect 9312 12427 9364 12436
rect 9312 12393 9321 12427
rect 9321 12393 9355 12427
rect 9355 12393 9364 12427
rect 9312 12384 9364 12393
rect 12808 12384 12860 12436
rect 13544 12384 13596 12436
rect 14096 12384 14148 12436
rect 14372 12384 14424 12436
rect 14740 12427 14792 12436
rect 14740 12393 14749 12427
rect 14749 12393 14783 12427
rect 14783 12393 14792 12427
rect 14740 12384 14792 12393
rect 16304 12384 16356 12436
rect 18788 12427 18840 12436
rect 18788 12393 18797 12427
rect 18797 12393 18831 12427
rect 18831 12393 18840 12427
rect 18788 12384 18840 12393
rect 19156 12427 19208 12436
rect 19156 12393 19165 12427
rect 19165 12393 19199 12427
rect 19199 12393 19208 12427
rect 19156 12384 19208 12393
rect 20260 12384 20312 12436
rect 20536 12384 20588 12436
rect 20628 12384 20680 12436
rect 20996 12384 21048 12436
rect 21640 12384 21692 12436
rect 22652 12384 22704 12436
rect 7932 12316 7984 12368
rect 9864 12316 9916 12368
rect 11060 12316 11112 12368
rect 14280 12316 14332 12368
rect 14464 12316 14516 12368
rect 17684 12316 17736 12368
rect 19340 12316 19392 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 4988 12248 5040 12300
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 10876 12248 10928 12300
rect 11244 12291 11296 12300
rect 11244 12257 11278 12291
rect 11278 12257 11296 12291
rect 11244 12248 11296 12257
rect 13820 12248 13872 12300
rect 17316 12248 17368 12300
rect 18972 12248 19024 12300
rect 21548 12359 21600 12368
rect 21548 12325 21557 12359
rect 21557 12325 21591 12359
rect 21591 12325 21600 12359
rect 21548 12316 21600 12325
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 2504 12180 2556 12232
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 4896 12180 4948 12232
rect 6184 12180 6236 12232
rect 7380 12180 7432 12232
rect 8392 12180 8444 12232
rect 10968 12223 11020 12232
rect 10968 12189 10977 12223
rect 10977 12189 11011 12223
rect 11011 12189 11020 12223
rect 10968 12180 11020 12189
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 15936 12180 15988 12232
rect 19432 12180 19484 12232
rect 3516 12112 3568 12164
rect 5540 12112 5592 12164
rect 1584 12044 1636 12096
rect 3424 12087 3476 12096
rect 3424 12053 3433 12087
rect 3433 12053 3467 12087
rect 3467 12053 3476 12087
rect 3424 12044 3476 12053
rect 6644 12087 6696 12096
rect 6644 12053 6653 12087
rect 6653 12053 6687 12087
rect 6687 12053 6696 12087
rect 6644 12044 6696 12053
rect 7196 12112 7248 12164
rect 8576 12155 8628 12164
rect 8576 12121 8585 12155
rect 8585 12121 8619 12155
rect 8619 12121 8628 12155
rect 8576 12112 8628 12121
rect 10140 12112 10192 12164
rect 13728 12155 13780 12164
rect 13728 12121 13737 12155
rect 13737 12121 13771 12155
rect 13771 12121 13780 12155
rect 13728 12112 13780 12121
rect 20168 12180 20220 12232
rect 20536 12180 20588 12232
rect 22284 12248 22336 12300
rect 22652 12248 22704 12300
rect 22100 12180 22152 12232
rect 23020 12384 23072 12436
rect 24492 12427 24544 12436
rect 24492 12393 24501 12427
rect 24501 12393 24535 12427
rect 24535 12393 24544 12427
rect 24492 12384 24544 12393
rect 23848 12316 23900 12368
rect 25228 12359 25280 12368
rect 25228 12325 25237 12359
rect 25237 12325 25271 12359
rect 25271 12325 25280 12359
rect 25228 12316 25280 12325
rect 23112 12248 23164 12300
rect 20260 12112 20312 12164
rect 23572 12180 23624 12232
rect 25044 12248 25096 12300
rect 25320 12248 25372 12300
rect 24860 12180 24912 12232
rect 23388 12112 23440 12164
rect 7012 12044 7064 12096
rect 8668 12044 8720 12096
rect 9496 12044 9548 12096
rect 12256 12044 12308 12096
rect 15844 12044 15896 12096
rect 18144 12087 18196 12096
rect 18144 12053 18153 12087
rect 18153 12053 18187 12087
rect 18187 12053 18196 12087
rect 18144 12044 18196 12053
rect 20168 12044 20220 12096
rect 20352 12087 20404 12096
rect 20352 12053 20361 12087
rect 20361 12053 20395 12087
rect 20395 12053 20404 12087
rect 20352 12044 20404 12053
rect 20720 12087 20772 12096
rect 20720 12053 20729 12087
rect 20729 12053 20763 12087
rect 20763 12053 20772 12087
rect 20720 12044 20772 12053
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 22376 12044 22428 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1400 11840 1452 11892
rect 1676 11840 1728 11892
rect 2228 11840 2280 11892
rect 3148 11883 3200 11892
rect 3148 11849 3157 11883
rect 3157 11849 3191 11883
rect 3191 11849 3200 11883
rect 3148 11840 3200 11849
rect 4988 11840 5040 11892
rect 7564 11840 7616 11892
rect 8668 11840 8720 11892
rect 10876 11883 10928 11892
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 11244 11840 11296 11892
rect 14280 11840 14332 11892
rect 14832 11840 14884 11892
rect 16212 11840 16264 11892
rect 17684 11840 17736 11892
rect 18972 11883 19024 11892
rect 18972 11849 18981 11883
rect 18981 11849 19015 11883
rect 19015 11849 19024 11883
rect 18972 11840 19024 11849
rect 2412 11772 2464 11824
rect 1860 11636 1912 11688
rect 2320 11611 2372 11620
rect 2320 11577 2329 11611
rect 2329 11577 2363 11611
rect 2363 11577 2372 11611
rect 2320 11568 2372 11577
rect 1860 11500 1912 11552
rect 1952 11500 2004 11552
rect 2688 11500 2740 11552
rect 4988 11704 5040 11756
rect 7380 11704 7432 11756
rect 8024 11772 8076 11824
rect 8116 11772 8168 11824
rect 16580 11772 16632 11824
rect 7932 11747 7984 11756
rect 7932 11713 7941 11747
rect 7941 11713 7975 11747
rect 7975 11713 7984 11747
rect 7932 11704 7984 11713
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 9496 11747 9548 11756
rect 9496 11713 9505 11747
rect 9505 11713 9539 11747
rect 9539 11713 9548 11747
rect 9496 11704 9548 11713
rect 12348 11704 12400 11756
rect 16396 11704 16448 11756
rect 17960 11704 18012 11756
rect 4712 11636 4764 11688
rect 8392 11679 8444 11688
rect 8392 11645 8401 11679
rect 8401 11645 8435 11679
rect 8435 11645 8444 11679
rect 8392 11636 8444 11645
rect 13452 11636 13504 11688
rect 13636 11679 13688 11688
rect 13636 11645 13670 11679
rect 13670 11645 13688 11679
rect 13636 11636 13688 11645
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 18972 11636 19024 11688
rect 19984 11840 20036 11892
rect 20720 11840 20772 11892
rect 21272 11840 21324 11892
rect 22100 11883 22152 11892
rect 22100 11849 22109 11883
rect 22109 11849 22143 11883
rect 22143 11849 22152 11883
rect 24768 11883 24820 11892
rect 22100 11840 22152 11849
rect 24768 11849 24777 11883
rect 24777 11849 24811 11883
rect 24811 11849 24820 11883
rect 24768 11840 24820 11849
rect 25412 11883 25464 11892
rect 25412 11849 25421 11883
rect 25421 11849 25455 11883
rect 25455 11849 25464 11883
rect 25412 11840 25464 11849
rect 23388 11772 23440 11824
rect 23848 11772 23900 11824
rect 25596 11772 25648 11824
rect 24124 11704 24176 11756
rect 22284 11679 22336 11688
rect 22284 11645 22293 11679
rect 22293 11645 22327 11679
rect 22327 11645 22336 11679
rect 22284 11636 22336 11645
rect 23572 11636 23624 11688
rect 25228 11679 25280 11688
rect 25228 11645 25237 11679
rect 25237 11645 25271 11679
rect 25271 11645 25280 11679
rect 25228 11636 25280 11645
rect 3884 11611 3936 11620
rect 3884 11577 3893 11611
rect 3893 11577 3927 11611
rect 3927 11577 3936 11611
rect 3884 11568 3936 11577
rect 4804 11568 4856 11620
rect 5816 11568 5868 11620
rect 7656 11568 7708 11620
rect 7840 11611 7892 11620
rect 7840 11577 7849 11611
rect 7849 11577 7883 11611
rect 7883 11577 7892 11611
rect 7840 11568 7892 11577
rect 13268 11611 13320 11620
rect 4252 11500 4304 11552
rect 5356 11543 5408 11552
rect 5356 11509 5365 11543
rect 5365 11509 5399 11543
rect 5399 11509 5408 11543
rect 5356 11500 5408 11509
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 6644 11500 6696 11552
rect 6828 11500 6880 11552
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 10876 11500 10928 11552
rect 12256 11543 12308 11552
rect 12256 11509 12265 11543
rect 12265 11509 12299 11543
rect 12299 11509 12308 11543
rect 12256 11500 12308 11509
rect 13268 11577 13277 11611
rect 13277 11577 13311 11611
rect 13311 11577 13320 11611
rect 13268 11568 13320 11577
rect 14096 11568 14148 11620
rect 18144 11568 18196 11620
rect 23112 11611 23164 11620
rect 23112 11577 23121 11611
rect 23121 11577 23155 11611
rect 23155 11577 23164 11611
rect 23112 11568 23164 11577
rect 14832 11500 14884 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 17224 11500 17276 11552
rect 17776 11500 17828 11552
rect 18420 11500 18472 11552
rect 19432 11500 19484 11552
rect 22468 11543 22520 11552
rect 22468 11509 22477 11543
rect 22477 11509 22511 11543
rect 22511 11509 22520 11543
rect 22468 11500 22520 11509
rect 24768 11500 24820 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 3424 11296 3476 11348
rect 5356 11296 5408 11348
rect 6828 11296 6880 11348
rect 7932 11296 7984 11348
rect 3976 11228 4028 11280
rect 4252 11271 4304 11280
rect 4252 11237 4261 11271
rect 4261 11237 4295 11271
rect 4295 11237 4304 11271
rect 4252 11228 4304 11237
rect 4712 11271 4764 11280
rect 4712 11237 4721 11271
rect 4721 11237 4755 11271
rect 4755 11237 4764 11271
rect 4712 11228 4764 11237
rect 5448 11228 5500 11280
rect 7380 11271 7432 11280
rect 7380 11237 7389 11271
rect 7389 11237 7423 11271
rect 7423 11237 7432 11271
rect 7380 11228 7432 11237
rect 8300 11296 8352 11348
rect 9404 11296 9456 11348
rect 11428 11339 11480 11348
rect 11428 11305 11437 11339
rect 11437 11305 11471 11339
rect 11471 11305 11480 11339
rect 11428 11296 11480 11305
rect 12256 11296 12308 11348
rect 13636 11296 13688 11348
rect 16672 11296 16724 11348
rect 17316 11296 17368 11348
rect 17960 11339 18012 11348
rect 17960 11305 17969 11339
rect 17969 11305 18003 11339
rect 18003 11305 18012 11339
rect 17960 11296 18012 11305
rect 18144 11296 18196 11348
rect 19340 11339 19392 11348
rect 19340 11305 19349 11339
rect 19349 11305 19383 11339
rect 19383 11305 19392 11339
rect 19340 11296 19392 11305
rect 20260 11339 20312 11348
rect 20260 11305 20269 11339
rect 20269 11305 20303 11339
rect 20303 11305 20312 11339
rect 20260 11296 20312 11305
rect 20720 11339 20772 11348
rect 20720 11305 20729 11339
rect 20729 11305 20763 11339
rect 20763 11305 20772 11339
rect 20720 11296 20772 11305
rect 21640 11339 21692 11348
rect 21640 11305 21649 11339
rect 21649 11305 21683 11339
rect 21683 11305 21692 11339
rect 21640 11296 21692 11305
rect 24124 11296 24176 11348
rect 25044 11339 25096 11348
rect 25044 11305 25053 11339
rect 25053 11305 25087 11339
rect 25087 11305 25096 11339
rect 25044 11296 25096 11305
rect 25412 11339 25464 11348
rect 25412 11305 25421 11339
rect 25421 11305 25455 11339
rect 25455 11305 25464 11339
rect 25412 11296 25464 11305
rect 3424 11160 3476 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 3516 11092 3568 11144
rect 9312 11228 9364 11280
rect 10784 11228 10836 11280
rect 13728 11228 13780 11280
rect 15568 11271 15620 11280
rect 15568 11237 15577 11271
rect 15577 11237 15611 11271
rect 15611 11237 15620 11271
rect 15568 11228 15620 11237
rect 16488 11228 16540 11280
rect 17684 11228 17736 11280
rect 18512 11228 18564 11280
rect 19984 11228 20036 11280
rect 20352 11228 20404 11280
rect 4988 11135 5040 11144
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 2320 11024 2372 11076
rect 7932 11160 7984 11212
rect 9864 11160 9916 11212
rect 11612 11160 11664 11212
rect 14464 11160 14516 11212
rect 14832 11160 14884 11212
rect 15384 11160 15436 11212
rect 19708 11203 19760 11212
rect 8024 11135 8076 11144
rect 8024 11101 8033 11135
rect 8033 11101 8067 11135
rect 8067 11101 8076 11135
rect 8024 11092 8076 11101
rect 9956 11092 10008 11144
rect 10968 11092 11020 11144
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 14280 11092 14332 11144
rect 17224 11092 17276 11144
rect 7748 11024 7800 11076
rect 9772 11067 9824 11076
rect 9772 11033 9781 11067
rect 9781 11033 9815 11067
rect 9815 11033 9824 11067
rect 9772 11024 9824 11033
rect 8576 10999 8628 11008
rect 8576 10965 8585 10999
rect 8585 10965 8619 10999
rect 8619 10965 8628 10999
rect 8576 10956 8628 10965
rect 13544 10956 13596 11008
rect 16948 11024 17000 11076
rect 19708 11169 19717 11203
rect 19717 11169 19751 11203
rect 19751 11169 19760 11203
rect 19708 11160 19760 11169
rect 20168 11160 20220 11212
rect 20720 11160 20772 11212
rect 25596 11160 25648 11212
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 19432 11092 19484 11144
rect 20260 11092 20312 11144
rect 22560 11092 22612 11144
rect 15660 10956 15712 11008
rect 16580 10956 16632 11008
rect 17684 10956 17736 11008
rect 20352 11024 20404 11076
rect 18236 10956 18288 11008
rect 18696 10956 18748 11008
rect 22376 10956 22428 11008
rect 23664 10956 23716 11008
rect 23756 10956 23808 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2964 10752 3016 10804
rect 3976 10795 4028 10804
rect 3976 10761 3985 10795
rect 3985 10761 4019 10795
rect 4019 10761 4028 10795
rect 3976 10752 4028 10761
rect 4988 10795 5040 10804
rect 4988 10761 4997 10795
rect 4997 10761 5031 10795
rect 5031 10761 5040 10795
rect 4988 10752 5040 10761
rect 5264 10752 5316 10804
rect 5540 10752 5592 10804
rect 6828 10752 6880 10804
rect 8024 10752 8076 10804
rect 10876 10795 10928 10804
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 12532 10752 12584 10804
rect 1768 10684 1820 10736
rect 5172 10684 5224 10736
rect 7932 10684 7984 10736
rect 8208 10684 8260 10736
rect 11796 10684 11848 10736
rect 13452 10752 13504 10804
rect 14832 10752 14884 10804
rect 16488 10795 16540 10804
rect 16488 10761 16497 10795
rect 16497 10761 16531 10795
rect 16531 10761 16540 10795
rect 16488 10752 16540 10761
rect 20720 10795 20772 10804
rect 20720 10761 20729 10795
rect 20729 10761 20763 10795
rect 20763 10761 20772 10795
rect 20720 10752 20772 10761
rect 14004 10684 14056 10736
rect 14740 10684 14792 10736
rect 23480 10684 23532 10736
rect 2596 10616 2648 10668
rect 2780 10659 2832 10668
rect 2780 10625 2789 10659
rect 2789 10625 2823 10659
rect 2823 10625 2832 10659
rect 2780 10616 2832 10625
rect 3240 10616 3292 10668
rect 4712 10616 4764 10668
rect 6368 10616 6420 10668
rect 11428 10659 11480 10668
rect 11428 10625 11437 10659
rect 11437 10625 11471 10659
rect 11471 10625 11480 10659
rect 11428 10616 11480 10625
rect 12440 10616 12492 10668
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 15660 10616 15712 10625
rect 20720 10616 20772 10668
rect 3792 10591 3844 10600
rect 3792 10557 3801 10591
rect 3801 10557 3835 10591
rect 3835 10557 3844 10591
rect 4252 10591 4304 10600
rect 3792 10548 3844 10557
rect 4252 10557 4261 10591
rect 4261 10557 4295 10591
rect 4295 10557 4304 10591
rect 4252 10548 4304 10557
rect 5356 10548 5408 10600
rect 8116 10548 8168 10600
rect 8300 10591 8352 10600
rect 8300 10557 8309 10591
rect 8309 10557 8343 10591
rect 8343 10557 8352 10591
rect 8300 10548 8352 10557
rect 8576 10591 8628 10600
rect 8576 10557 8610 10591
rect 8610 10557 8628 10591
rect 8576 10548 8628 10557
rect 13452 10591 13504 10600
rect 13452 10557 13461 10591
rect 13461 10557 13495 10591
rect 13495 10557 13504 10591
rect 13452 10548 13504 10557
rect 14648 10548 14700 10600
rect 2964 10480 3016 10532
rect 7288 10523 7340 10532
rect 7288 10489 7297 10523
rect 7297 10489 7331 10523
rect 7331 10489 7340 10523
rect 7288 10480 7340 10489
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 7380 10412 7432 10464
rect 9680 10455 9732 10464
rect 9680 10421 9689 10455
rect 9689 10421 9723 10455
rect 9723 10421 9732 10455
rect 9680 10412 9732 10421
rect 9864 10412 9916 10464
rect 10692 10455 10744 10464
rect 10692 10421 10701 10455
rect 10701 10421 10735 10455
rect 10735 10421 10744 10455
rect 10692 10412 10744 10421
rect 12532 10480 12584 10532
rect 13360 10480 13412 10532
rect 16028 10523 16080 10532
rect 16028 10489 16037 10523
rect 16037 10489 16071 10523
rect 16071 10489 16080 10523
rect 16028 10480 16080 10489
rect 17132 10480 17184 10532
rect 12256 10455 12308 10464
rect 12256 10421 12265 10455
rect 12265 10421 12299 10455
rect 12299 10421 12308 10455
rect 18144 10548 18196 10600
rect 19708 10548 19760 10600
rect 20076 10591 20128 10600
rect 20076 10557 20085 10591
rect 20085 10557 20119 10591
rect 20119 10557 20128 10591
rect 20076 10548 20128 10557
rect 21548 10548 21600 10600
rect 22376 10616 22428 10668
rect 23664 10591 23716 10600
rect 20904 10480 20956 10532
rect 12256 10412 12308 10421
rect 13728 10412 13780 10464
rect 16396 10412 16448 10464
rect 17224 10412 17276 10464
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 18512 10412 18564 10464
rect 21272 10412 21324 10464
rect 21548 10412 21600 10464
rect 22192 10480 22244 10532
rect 23388 10480 23440 10532
rect 23664 10557 23673 10591
rect 23673 10557 23707 10591
rect 23707 10557 23716 10591
rect 23664 10548 23716 10557
rect 23756 10548 23808 10600
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 25596 10455 25648 10464
rect 25596 10421 25605 10455
rect 25605 10421 25639 10455
rect 25639 10421 25648 10455
rect 25596 10412 25648 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1860 10208 1912 10260
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 3240 10251 3292 10260
rect 2780 10208 2832 10217
rect 3240 10217 3249 10251
rect 3249 10217 3283 10251
rect 3283 10217 3292 10251
rect 3240 10208 3292 10217
rect 4528 10208 4580 10260
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 8116 10208 8168 10260
rect 8300 10251 8352 10260
rect 8300 10217 8309 10251
rect 8309 10217 8343 10251
rect 8343 10217 8352 10251
rect 8300 10208 8352 10217
rect 1400 10140 1452 10192
rect 4804 10183 4856 10192
rect 4804 10149 4813 10183
rect 4813 10149 4847 10183
rect 4847 10149 4856 10183
rect 4804 10140 4856 10149
rect 5540 10140 5592 10192
rect 6460 10140 6512 10192
rect 1768 10072 1820 10124
rect 2780 10072 2832 10124
rect 5172 10072 5224 10124
rect 5448 10072 5500 10124
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 3424 10004 3476 10056
rect 4712 9936 4764 9988
rect 8944 10208 8996 10260
rect 10232 10183 10284 10192
rect 10232 10149 10241 10183
rect 10241 10149 10275 10183
rect 10275 10149 10284 10183
rect 10232 10140 10284 10149
rect 13728 10208 13780 10260
rect 14004 10251 14056 10260
rect 14004 10217 14013 10251
rect 14013 10217 14047 10251
rect 14047 10217 14056 10251
rect 14004 10208 14056 10217
rect 14648 10208 14700 10260
rect 17316 10251 17368 10260
rect 13176 10183 13228 10192
rect 13176 10149 13185 10183
rect 13185 10149 13219 10183
rect 13219 10149 13228 10183
rect 13176 10140 13228 10149
rect 13360 10140 13412 10192
rect 15660 10183 15712 10192
rect 15660 10149 15694 10183
rect 15694 10149 15712 10183
rect 15660 10140 15712 10149
rect 15844 10140 15896 10192
rect 17316 10217 17325 10251
rect 17325 10217 17359 10251
rect 17359 10217 17368 10251
rect 17316 10208 17368 10217
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 18236 10208 18288 10260
rect 18604 10208 18656 10260
rect 20720 10251 20772 10260
rect 20720 10217 20729 10251
rect 20729 10217 20763 10251
rect 20763 10217 20772 10251
rect 20720 10208 20772 10217
rect 22836 10251 22888 10260
rect 22836 10217 22845 10251
rect 22845 10217 22879 10251
rect 22879 10217 22888 10251
rect 22836 10208 22888 10217
rect 23756 10251 23808 10260
rect 23756 10217 23765 10251
rect 23765 10217 23799 10251
rect 23799 10217 23808 10251
rect 23756 10208 23808 10217
rect 17408 10140 17460 10192
rect 18512 10183 18564 10192
rect 18512 10149 18521 10183
rect 18521 10149 18555 10183
rect 18555 10149 18564 10183
rect 18512 10140 18564 10149
rect 21916 10140 21968 10192
rect 9680 10072 9732 10124
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 8668 9979 8720 9988
rect 8668 9945 8677 9979
rect 8677 9945 8711 9979
rect 8711 9945 8720 9979
rect 8668 9936 8720 9945
rect 9496 9936 9548 9988
rect 11980 10072 12032 10124
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 12992 10072 13044 10081
rect 14648 10072 14700 10124
rect 18052 10072 18104 10124
rect 19432 10072 19484 10124
rect 21732 10115 21784 10124
rect 21732 10081 21766 10115
rect 21766 10081 21784 10115
rect 21732 10072 21784 10081
rect 22836 10072 22888 10124
rect 23664 10072 23716 10124
rect 25044 10072 25096 10124
rect 12440 10004 12492 10056
rect 13452 10004 13504 10056
rect 16396 10004 16448 10056
rect 19156 10004 19208 10056
rect 20904 10004 20956 10056
rect 12164 9936 12216 9988
rect 2320 9868 2372 9920
rect 5356 9868 5408 9920
rect 7472 9868 7524 9920
rect 8300 9868 8352 9920
rect 9312 9868 9364 9920
rect 10968 9868 11020 9920
rect 11612 9868 11664 9920
rect 12532 9868 12584 9920
rect 13636 9936 13688 9988
rect 15384 9868 15436 9920
rect 16856 9936 16908 9988
rect 18144 9936 18196 9988
rect 18972 9936 19024 9988
rect 16580 9868 16632 9920
rect 18604 9868 18656 9920
rect 19616 9868 19668 9920
rect 20536 9868 20588 9920
rect 24952 9868 25004 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1860 9664 1912 9716
rect 4528 9664 4580 9716
rect 5448 9664 5500 9716
rect 6460 9707 6512 9716
rect 6460 9673 6469 9707
rect 6469 9673 6503 9707
rect 6503 9673 6512 9707
rect 6460 9664 6512 9673
rect 6828 9664 6880 9716
rect 8576 9664 8628 9716
rect 10324 9707 10376 9716
rect 10324 9673 10333 9707
rect 10333 9673 10367 9707
rect 10367 9673 10376 9707
rect 10324 9664 10376 9673
rect 13268 9664 13320 9716
rect 10876 9639 10928 9648
rect 2964 9528 3016 9580
rect 4160 9571 4212 9580
rect 4160 9537 4169 9571
rect 4169 9537 4203 9571
rect 4203 9537 4212 9571
rect 4160 9528 4212 9537
rect 10876 9605 10885 9639
rect 10885 9605 10919 9639
rect 10919 9605 10928 9639
rect 10876 9596 10928 9605
rect 12440 9596 12492 9648
rect 13360 9596 13412 9648
rect 15660 9664 15712 9716
rect 18236 9664 18288 9716
rect 18788 9664 18840 9716
rect 23388 9664 23440 9716
rect 23664 9664 23716 9716
rect 15108 9596 15160 9648
rect 17960 9596 18012 9648
rect 18512 9596 18564 9648
rect 21180 9596 21232 9648
rect 23572 9596 23624 9648
rect 24124 9639 24176 9648
rect 24124 9605 24133 9639
rect 24133 9605 24167 9639
rect 24167 9605 24176 9639
rect 24124 9596 24176 9605
rect 2412 9460 2464 9512
rect 12348 9528 12400 9580
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 18052 9528 18104 9580
rect 21088 9528 21140 9580
rect 22100 9528 22152 9580
rect 24492 9528 24544 9580
rect 8300 9460 8352 9512
rect 8944 9460 8996 9512
rect 13820 9460 13872 9512
rect 4528 9392 4580 9444
rect 7472 9392 7524 9444
rect 9680 9435 9732 9444
rect 9680 9401 9689 9435
rect 9689 9401 9723 9435
rect 9723 9401 9732 9435
rect 9680 9392 9732 9401
rect 11152 9435 11204 9444
rect 11152 9401 11161 9435
rect 11161 9401 11195 9435
rect 11195 9401 11204 9435
rect 11152 9392 11204 9401
rect 13636 9435 13688 9444
rect 13636 9401 13645 9435
rect 13645 9401 13679 9435
rect 13679 9401 13688 9435
rect 13636 9392 13688 9401
rect 14832 9392 14884 9444
rect 16028 9460 16080 9512
rect 16488 9460 16540 9512
rect 17776 9392 17828 9444
rect 18144 9392 18196 9444
rect 19616 9460 19668 9512
rect 20720 9460 20772 9512
rect 18972 9392 19024 9444
rect 21088 9392 21140 9444
rect 21640 9392 21692 9444
rect 23572 9392 23624 9444
rect 24584 9435 24636 9444
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 3056 9324 3108 9333
rect 4988 9324 5040 9376
rect 9220 9367 9272 9376
rect 9220 9333 9229 9367
rect 9229 9333 9263 9367
rect 9263 9333 9272 9367
rect 9220 9324 9272 9333
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 10968 9324 11020 9376
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 13176 9324 13228 9376
rect 15844 9324 15896 9376
rect 16580 9324 16632 9376
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 20904 9367 20956 9376
rect 20904 9333 20913 9367
rect 20913 9333 20947 9367
rect 20947 9333 20956 9367
rect 20904 9324 20956 9333
rect 21824 9324 21876 9376
rect 24584 9401 24593 9435
rect 24593 9401 24627 9435
rect 24627 9401 24636 9435
rect 24584 9392 24636 9401
rect 24952 9392 25004 9444
rect 25044 9367 25096 9376
rect 25044 9333 25053 9367
rect 25053 9333 25087 9367
rect 25087 9333 25096 9367
rect 25044 9324 25096 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1400 9120 1452 9172
rect 2136 9120 2188 9172
rect 3056 9163 3108 9172
rect 3056 9129 3065 9163
rect 3065 9129 3099 9163
rect 3099 9129 3108 9163
rect 3056 9120 3108 9129
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 4528 9120 4580 9172
rect 4804 9120 4856 9172
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 5632 9120 5684 9172
rect 6368 9163 6420 9172
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 6920 9163 6972 9172
rect 6920 9129 6929 9163
rect 6929 9129 6963 9163
rect 6963 9129 6972 9163
rect 6920 9120 6972 9129
rect 7104 9120 7156 9172
rect 1860 8823 1912 8832
rect 1860 8789 1869 8823
rect 1869 8789 1903 8823
rect 1903 8789 1912 8823
rect 1860 8780 1912 8789
rect 2412 9095 2464 9104
rect 2412 9061 2421 9095
rect 2421 9061 2455 9095
rect 2455 9061 2464 9095
rect 2412 9052 2464 9061
rect 4896 9052 4948 9104
rect 6644 9052 6696 9104
rect 8300 9052 8352 9104
rect 8484 9052 8536 9104
rect 13452 9120 13504 9172
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 14740 9163 14792 9172
rect 14740 9129 14749 9163
rect 14749 9129 14783 9163
rect 14783 9129 14792 9163
rect 14740 9120 14792 9129
rect 18972 9120 19024 9172
rect 20444 9120 20496 9172
rect 23480 9120 23532 9172
rect 24492 9120 24544 9172
rect 24860 9163 24912 9172
rect 24860 9129 24869 9163
rect 24869 9129 24903 9163
rect 24903 9129 24912 9163
rect 24860 9120 24912 9129
rect 26240 9120 26292 9172
rect 9036 9095 9088 9104
rect 4988 8984 5040 9036
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 5080 8916 5132 8968
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 7472 8916 7524 8968
rect 8576 8916 8628 8968
rect 5356 8848 5408 8900
rect 6736 8848 6788 8900
rect 8116 8891 8168 8900
rect 8116 8857 8125 8891
rect 8125 8857 8159 8891
rect 8159 8857 8168 8891
rect 8116 8848 8168 8857
rect 8392 8848 8444 8900
rect 9036 9061 9045 9095
rect 9045 9061 9079 9095
rect 9079 9061 9088 9095
rect 9036 9052 9088 9061
rect 12348 9052 12400 9104
rect 13176 9052 13228 9104
rect 15108 9095 15160 9104
rect 15108 9061 15117 9095
rect 15117 9061 15151 9095
rect 15151 9061 15160 9095
rect 15108 9052 15160 9061
rect 15292 9052 15344 9104
rect 15752 9052 15804 9104
rect 16028 9052 16080 9104
rect 17960 9095 18012 9104
rect 17960 9061 17994 9095
rect 17994 9061 18012 9095
rect 17960 9052 18012 9061
rect 21180 9095 21232 9104
rect 21180 9061 21214 9095
rect 21214 9061 21232 9095
rect 21180 9052 21232 9061
rect 22100 9052 22152 9104
rect 25504 9052 25556 9104
rect 26424 9052 26476 9104
rect 11796 8984 11848 9036
rect 16304 9027 16356 9036
rect 16304 8993 16313 9027
rect 16313 8993 16347 9027
rect 16347 8993 16356 9027
rect 16304 8984 16356 8993
rect 17776 8984 17828 9036
rect 20168 8984 20220 9036
rect 22468 8984 22520 9036
rect 24676 9027 24728 9036
rect 24676 8993 24685 9027
rect 24685 8993 24719 9027
rect 24719 8993 24728 9027
rect 24676 8984 24728 8993
rect 10140 8916 10192 8968
rect 15476 8916 15528 8968
rect 16396 8916 16448 8968
rect 17408 8916 17460 8968
rect 20904 8959 20956 8968
rect 20904 8925 20913 8959
rect 20913 8925 20947 8959
rect 20947 8925 20956 8959
rect 20904 8916 20956 8925
rect 23664 8916 23716 8968
rect 25044 8916 25096 8968
rect 16672 8891 16724 8900
rect 16672 8857 16681 8891
rect 16681 8857 16715 8891
rect 16715 8857 16724 8891
rect 16672 8848 16724 8857
rect 24584 8848 24636 8900
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9404 8780 9456 8789
rect 9680 8780 9732 8832
rect 11612 8823 11664 8832
rect 11612 8789 11621 8823
rect 11621 8789 11655 8823
rect 11655 8789 11664 8823
rect 11612 8780 11664 8789
rect 12440 8823 12492 8832
rect 12440 8789 12449 8823
rect 12449 8789 12483 8823
rect 12483 8789 12492 8823
rect 12440 8780 12492 8789
rect 16488 8780 16540 8832
rect 17040 8823 17092 8832
rect 17040 8789 17049 8823
rect 17049 8789 17083 8823
rect 17083 8789 17092 8823
rect 17040 8780 17092 8789
rect 17592 8823 17644 8832
rect 17592 8789 17601 8823
rect 17601 8789 17635 8823
rect 17635 8789 17644 8823
rect 17592 8780 17644 8789
rect 19432 8780 19484 8832
rect 19708 8823 19760 8832
rect 19708 8789 19717 8823
rect 19717 8789 19751 8823
rect 19751 8789 19760 8823
rect 19708 8780 19760 8789
rect 20168 8780 20220 8832
rect 22376 8780 22428 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1676 8576 1728 8628
rect 1952 8576 2004 8628
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 2964 8576 3016 8628
rect 4988 8619 5040 8628
rect 4988 8585 4997 8619
rect 4997 8585 5031 8619
rect 5031 8585 5040 8619
rect 4988 8576 5040 8585
rect 6460 8576 6512 8628
rect 8208 8619 8260 8628
rect 8208 8585 8217 8619
rect 8217 8585 8251 8619
rect 8251 8585 8260 8619
rect 8208 8576 8260 8585
rect 8944 8576 8996 8628
rect 10140 8576 10192 8628
rect 10784 8576 10836 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 2136 8508 2188 8560
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 4896 8508 4948 8560
rect 9956 8508 10008 8560
rect 5356 8440 5408 8492
rect 5632 8440 5684 8492
rect 5908 8440 5960 8492
rect 6184 8440 6236 8492
rect 6460 8440 6512 8492
rect 6644 8440 6696 8492
rect 8576 8440 8628 8492
rect 11244 8440 11296 8492
rect 11704 8508 11756 8560
rect 12348 8576 12400 8628
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 16120 8619 16172 8628
rect 16120 8585 16129 8619
rect 16129 8585 16163 8619
rect 16163 8585 16172 8619
rect 16120 8576 16172 8585
rect 19984 8576 20036 8628
rect 21364 8576 21416 8628
rect 12624 8551 12676 8560
rect 12624 8517 12633 8551
rect 12633 8517 12667 8551
rect 12667 8517 12676 8551
rect 12624 8508 12676 8517
rect 16396 8551 16448 8560
rect 16396 8517 16405 8551
rect 16405 8517 16439 8551
rect 16439 8517 16448 8551
rect 16396 8508 16448 8517
rect 18144 8551 18196 8560
rect 18144 8517 18153 8551
rect 18153 8517 18187 8551
rect 18187 8517 18196 8551
rect 18144 8508 18196 8517
rect 20720 8508 20772 8560
rect 21640 8551 21692 8560
rect 21640 8517 21649 8551
rect 21649 8517 21683 8551
rect 21683 8517 21692 8551
rect 21640 8508 21692 8517
rect 23664 8576 23716 8628
rect 24676 8576 24728 8628
rect 24860 8619 24912 8628
rect 24860 8585 24869 8619
rect 24869 8585 24903 8619
rect 24903 8585 24912 8619
rect 24860 8576 24912 8585
rect 25136 8619 25188 8628
rect 25136 8585 25145 8619
rect 25145 8585 25179 8619
rect 25179 8585 25188 8619
rect 25136 8576 25188 8585
rect 12716 8440 12768 8492
rect 16304 8440 16356 8492
rect 18972 8440 19024 8492
rect 21180 8440 21232 8492
rect 22376 8440 22428 8492
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 2504 8372 2556 8424
rect 2688 8304 2740 8356
rect 5448 8415 5500 8424
rect 5448 8381 5457 8415
rect 5457 8381 5491 8415
rect 5491 8381 5500 8415
rect 5448 8372 5500 8381
rect 6736 8372 6788 8424
rect 9680 8415 9732 8424
rect 3148 8304 3200 8356
rect 5724 8347 5776 8356
rect 5724 8313 5733 8347
rect 5733 8313 5767 8347
rect 5767 8313 5776 8347
rect 5724 8304 5776 8313
rect 7104 8347 7156 8356
rect 7104 8313 7113 8347
rect 7113 8313 7147 8347
rect 7147 8313 7156 8347
rect 7104 8304 7156 8313
rect 8392 8304 8444 8356
rect 8668 8347 8720 8356
rect 8668 8313 8677 8347
rect 8677 8313 8711 8347
rect 8711 8313 8720 8347
rect 8668 8304 8720 8313
rect 9312 8304 9364 8356
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 9588 8304 9640 8356
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 11888 8304 11940 8356
rect 4712 8236 4764 8288
rect 5264 8236 5316 8288
rect 9680 8236 9732 8288
rect 9864 8236 9916 8288
rect 12164 8236 12216 8288
rect 13176 8236 13228 8288
rect 14096 8415 14148 8424
rect 14096 8381 14130 8415
rect 14130 8381 14148 8415
rect 14096 8372 14148 8381
rect 16120 8372 16172 8424
rect 19984 8372 20036 8424
rect 21916 8415 21968 8424
rect 21916 8381 21925 8415
rect 21925 8381 21959 8415
rect 21959 8381 21968 8415
rect 21916 8372 21968 8381
rect 23480 8372 23532 8424
rect 24952 8415 25004 8424
rect 24952 8381 24961 8415
rect 24961 8381 24995 8415
rect 24995 8381 25004 8415
rect 24952 8372 25004 8381
rect 13820 8236 13872 8288
rect 16304 8236 16356 8288
rect 17592 8304 17644 8356
rect 18604 8347 18656 8356
rect 18604 8313 18613 8347
rect 18613 8313 18647 8347
rect 18647 8313 18656 8347
rect 18604 8304 18656 8313
rect 20444 8304 20496 8356
rect 22376 8304 22428 8356
rect 24216 8304 24268 8356
rect 26792 8304 26844 8356
rect 17408 8236 17460 8288
rect 20904 8236 20956 8288
rect 21548 8236 21600 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1768 8032 1820 8084
rect 2228 8032 2280 8084
rect 2964 8075 3016 8084
rect 2964 8041 2973 8075
rect 2973 8041 3007 8075
rect 3007 8041 3016 8075
rect 2964 8032 3016 8041
rect 4436 8032 4488 8084
rect 5356 8032 5408 8084
rect 4528 7964 4580 8016
rect 6184 7964 6236 8016
rect 6828 8032 6880 8084
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 8208 8032 8260 8084
rect 8576 8032 8628 8084
rect 10968 8032 11020 8084
rect 11796 8032 11848 8084
rect 12716 8075 12768 8084
rect 12716 8041 12725 8075
rect 12725 8041 12759 8075
rect 12759 8041 12768 8075
rect 12716 8032 12768 8041
rect 13728 8032 13780 8084
rect 13820 8032 13872 8084
rect 14832 8032 14884 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 18328 8032 18380 8084
rect 18512 8075 18564 8084
rect 18512 8041 18521 8075
rect 18521 8041 18555 8075
rect 18555 8041 18564 8075
rect 18512 8032 18564 8041
rect 20720 8032 20772 8084
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 23664 8075 23716 8084
rect 23664 8041 23673 8075
rect 23673 8041 23707 8075
rect 23707 8041 23716 8075
rect 23664 8032 23716 8041
rect 7012 7964 7064 8016
rect 13452 8007 13504 8016
rect 13452 7973 13461 8007
rect 13461 7973 13495 8007
rect 13495 7973 13504 8007
rect 13452 7964 13504 7973
rect 15936 8007 15988 8016
rect 15936 7973 15945 8007
rect 15945 7973 15979 8007
rect 15979 7973 15988 8007
rect 15936 7964 15988 7973
rect 17500 7964 17552 8016
rect 19156 7964 19208 8016
rect 19340 7964 19392 8016
rect 21180 8007 21232 8016
rect 5632 7896 5684 7948
rect 6368 7896 6420 7948
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 11336 7896 11388 7948
rect 14096 7896 14148 7948
rect 15660 7939 15712 7948
rect 15660 7905 15669 7939
rect 15669 7905 15703 7939
rect 15703 7905 15712 7939
rect 15660 7896 15712 7905
rect 18236 7896 18288 7948
rect 21180 7973 21189 8007
rect 21189 7973 21223 8007
rect 21223 7973 21232 8007
rect 21180 7964 21232 7973
rect 22376 7964 22428 8016
rect 23848 7964 23900 8016
rect 21548 7896 21600 7948
rect 23572 7896 23624 7948
rect 24124 7896 24176 7948
rect 2964 7871 3016 7880
rect 2964 7837 2973 7871
rect 2973 7837 3007 7871
rect 3007 7837 3016 7871
rect 2964 7828 3016 7837
rect 3148 7828 3200 7880
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 1860 7760 1912 7812
rect 2596 7760 2648 7812
rect 4896 7760 4948 7812
rect 2320 7692 2372 7744
rect 3792 7692 3844 7744
rect 4252 7692 4304 7744
rect 9036 7692 9088 7744
rect 9864 7692 9916 7744
rect 11152 7828 11204 7880
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 17960 7871 18012 7880
rect 17960 7837 17969 7871
rect 17969 7837 18003 7871
rect 18003 7837 18012 7871
rect 17960 7828 18012 7837
rect 13544 7760 13596 7812
rect 15384 7803 15436 7812
rect 15384 7769 15393 7803
rect 15393 7769 15427 7803
rect 15427 7769 15436 7803
rect 15384 7760 15436 7769
rect 17592 7803 17644 7812
rect 17592 7769 17601 7803
rect 17601 7769 17635 7803
rect 17635 7769 17644 7803
rect 17592 7760 17644 7769
rect 10140 7692 10192 7744
rect 11244 7692 11296 7744
rect 12256 7735 12308 7744
rect 12256 7701 12265 7735
rect 12265 7701 12299 7735
rect 12299 7701 12308 7735
rect 12256 7692 12308 7701
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 19156 7735 19208 7744
rect 19156 7701 19165 7735
rect 19165 7701 19199 7735
rect 19199 7701 19208 7735
rect 19156 7692 19208 7701
rect 19524 7692 19576 7744
rect 19892 7692 19944 7744
rect 20904 7760 20956 7812
rect 22744 7828 22796 7880
rect 23112 7828 23164 7880
rect 20444 7735 20496 7744
rect 20444 7701 20453 7735
rect 20453 7701 20487 7735
rect 20487 7701 20496 7735
rect 20444 7692 20496 7701
rect 23112 7735 23164 7744
rect 23112 7701 23121 7735
rect 23121 7701 23155 7735
rect 23155 7701 23164 7735
rect 23112 7692 23164 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2872 7488 2924 7540
rect 3700 7531 3752 7540
rect 3700 7497 3709 7531
rect 3709 7497 3743 7531
rect 3743 7497 3752 7531
rect 3700 7488 3752 7497
rect 4620 7531 4672 7540
rect 4620 7497 4629 7531
rect 4629 7497 4663 7531
rect 4663 7497 4672 7531
rect 4620 7488 4672 7497
rect 5448 7488 5500 7540
rect 6368 7488 6420 7540
rect 4436 7420 4488 7472
rect 4528 7420 4580 7472
rect 2228 7352 2280 7404
rect 3516 7352 3568 7404
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 5448 7352 5500 7404
rect 6276 7352 6328 7404
rect 7564 7352 7616 7404
rect 9496 7488 9548 7540
rect 12900 7488 12952 7540
rect 15844 7488 15896 7540
rect 16120 7531 16172 7540
rect 16120 7497 16129 7531
rect 16129 7497 16163 7531
rect 16163 7497 16172 7531
rect 16120 7488 16172 7497
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 18236 7488 18288 7540
rect 20904 7488 20956 7540
rect 9772 7352 9824 7404
rect 10784 7352 10836 7404
rect 6644 7284 6696 7336
rect 6828 7284 6880 7336
rect 10968 7327 11020 7336
rect 10968 7293 10977 7327
rect 10977 7293 11011 7327
rect 11011 7293 11020 7327
rect 10968 7284 11020 7293
rect 12900 7284 12952 7336
rect 13176 7284 13228 7336
rect 13820 7327 13872 7336
rect 13820 7293 13854 7327
rect 13854 7293 13872 7327
rect 2596 7259 2648 7268
rect 2596 7225 2605 7259
rect 2605 7225 2639 7259
rect 2639 7225 2648 7259
rect 2596 7216 2648 7225
rect 3608 7216 3660 7268
rect 3792 7216 3844 7268
rect 5356 7216 5408 7268
rect 6092 7216 6144 7268
rect 8024 7216 8076 7268
rect 3056 7191 3108 7200
rect 3056 7157 3065 7191
rect 3065 7157 3099 7191
rect 3099 7157 3108 7191
rect 3056 7148 3108 7157
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 6368 7148 6420 7200
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 9220 7191 9272 7200
rect 9220 7157 9229 7191
rect 9229 7157 9263 7191
rect 9263 7157 9272 7191
rect 9220 7148 9272 7157
rect 10140 7148 10192 7200
rect 10876 7191 10928 7200
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 11336 7191 11388 7200
rect 10876 7148 10928 7157
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 13820 7284 13872 7293
rect 14648 7284 14700 7336
rect 18328 7284 18380 7336
rect 18880 7284 18932 7336
rect 19892 7284 19944 7336
rect 22284 7488 22336 7540
rect 23020 7488 23072 7540
rect 24124 7488 24176 7540
rect 25412 7531 25464 7540
rect 25412 7497 25421 7531
rect 25421 7497 25455 7531
rect 25455 7497 25464 7531
rect 25412 7488 25464 7497
rect 22560 7420 22612 7472
rect 23848 7420 23900 7472
rect 22652 7352 22704 7404
rect 23112 7352 23164 7404
rect 22100 7284 22152 7336
rect 22284 7284 22336 7336
rect 16672 7259 16724 7268
rect 16672 7225 16681 7259
rect 16681 7225 16715 7259
rect 16715 7225 16724 7259
rect 16672 7216 16724 7225
rect 19340 7216 19392 7268
rect 19524 7259 19576 7268
rect 19524 7225 19558 7259
rect 19558 7225 19576 7259
rect 19524 7216 19576 7225
rect 23664 7284 23716 7336
rect 23480 7259 23532 7268
rect 13820 7148 13872 7200
rect 14648 7148 14700 7200
rect 16304 7148 16356 7200
rect 16764 7148 16816 7200
rect 18328 7148 18380 7200
rect 20260 7148 20312 7200
rect 20628 7191 20680 7200
rect 20628 7157 20637 7191
rect 20637 7157 20671 7191
rect 20671 7157 20680 7191
rect 20628 7148 20680 7157
rect 22192 7148 22244 7200
rect 23480 7225 23489 7259
rect 23489 7225 23523 7259
rect 23523 7225 23532 7259
rect 23480 7216 23532 7225
rect 23112 7148 23164 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 6276 6987 6328 6996
rect 6276 6953 6285 6987
rect 6285 6953 6319 6987
rect 6319 6953 6328 6987
rect 6276 6944 6328 6953
rect 6644 6987 6696 6996
rect 6644 6953 6653 6987
rect 6653 6953 6687 6987
rect 6687 6953 6696 6987
rect 6644 6944 6696 6953
rect 7932 6987 7984 6996
rect 7932 6953 7941 6987
rect 7941 6953 7975 6987
rect 7975 6953 7984 6987
rect 7932 6944 7984 6953
rect 10968 6944 11020 6996
rect 13452 6944 13504 6996
rect 14096 6944 14148 6996
rect 15660 6944 15712 6996
rect 18512 6944 18564 6996
rect 22652 6944 22704 6996
rect 4712 6876 4764 6928
rect 1768 6851 1820 6860
rect 1768 6817 1802 6851
rect 1802 6817 1820 6851
rect 1768 6808 1820 6817
rect 4160 6808 4212 6860
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 6920 6851 6972 6860
rect 4252 6808 4304 6817
rect 6920 6817 6929 6851
rect 6929 6817 6963 6851
rect 6963 6817 6972 6851
rect 6920 6808 6972 6817
rect 7196 6808 7248 6860
rect 10692 6876 10744 6928
rect 1492 6783 1544 6792
rect 1492 6749 1501 6783
rect 1501 6749 1535 6783
rect 1535 6749 1544 6783
rect 1492 6740 1544 6749
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 5632 6715 5684 6724
rect 5632 6681 5641 6715
rect 5641 6681 5675 6715
rect 5675 6681 5684 6715
rect 5632 6672 5684 6681
rect 6000 6672 6052 6724
rect 7472 6715 7524 6724
rect 7472 6681 7481 6715
rect 7481 6681 7515 6715
rect 7515 6681 7524 6715
rect 7472 6672 7524 6681
rect 2688 6604 2740 6656
rect 3424 6604 3476 6656
rect 8852 6672 8904 6724
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 9312 6604 9364 6656
rect 11060 6808 11112 6860
rect 13544 6808 13596 6860
rect 14004 6808 14056 6860
rect 14648 6851 14700 6860
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 14648 6808 14700 6817
rect 14740 6808 14792 6860
rect 9864 6647 9916 6656
rect 9864 6613 9873 6647
rect 9873 6613 9907 6647
rect 9907 6613 9916 6647
rect 9864 6604 9916 6613
rect 10692 6647 10744 6656
rect 10692 6613 10701 6647
rect 10701 6613 10735 6647
rect 10735 6613 10744 6647
rect 10692 6604 10744 6613
rect 12808 6740 12860 6792
rect 13636 6740 13688 6792
rect 15568 6740 15620 6792
rect 17408 6876 17460 6928
rect 19064 6876 19116 6928
rect 19616 6876 19668 6928
rect 20076 6876 20128 6928
rect 23848 6876 23900 6928
rect 16120 6851 16172 6860
rect 16120 6817 16154 6851
rect 16154 6817 16172 6851
rect 16120 6808 16172 6817
rect 16672 6808 16724 6860
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 19524 6808 19576 6860
rect 20720 6851 20772 6860
rect 19340 6740 19392 6792
rect 20720 6817 20729 6851
rect 20729 6817 20763 6851
rect 20763 6817 20772 6851
rect 20720 6808 20772 6817
rect 21180 6808 21232 6860
rect 22376 6851 22428 6860
rect 22376 6817 22385 6851
rect 22385 6817 22419 6851
rect 22419 6817 22428 6851
rect 22376 6808 22428 6817
rect 13728 6715 13780 6724
rect 13728 6681 13737 6715
rect 13737 6681 13771 6715
rect 13771 6681 13780 6715
rect 13728 6672 13780 6681
rect 13820 6672 13872 6724
rect 20076 6672 20128 6724
rect 22192 6740 22244 6792
rect 23388 6808 23440 6860
rect 25596 6808 25648 6860
rect 22652 6783 22704 6792
rect 22652 6749 22668 6783
rect 22668 6749 22702 6783
rect 22702 6749 22704 6783
rect 22652 6740 22704 6749
rect 25320 6715 25372 6724
rect 25320 6681 25329 6715
rect 25329 6681 25363 6715
rect 25363 6681 25372 6715
rect 25320 6672 25372 6681
rect 11152 6604 11204 6656
rect 11336 6604 11388 6656
rect 14096 6604 14148 6656
rect 17224 6647 17276 6656
rect 17224 6613 17233 6647
rect 17233 6613 17267 6647
rect 17267 6613 17276 6647
rect 17224 6604 17276 6613
rect 19340 6647 19392 6656
rect 19340 6613 19349 6647
rect 19349 6613 19383 6647
rect 19383 6613 19392 6647
rect 19340 6604 19392 6613
rect 20260 6647 20312 6656
rect 20260 6613 20269 6647
rect 20269 6613 20303 6647
rect 20303 6613 20312 6647
rect 20260 6604 20312 6613
rect 20812 6604 20864 6656
rect 21088 6647 21140 6656
rect 21088 6613 21097 6647
rect 21097 6613 21131 6647
rect 21131 6613 21140 6647
rect 21088 6604 21140 6613
rect 22100 6604 22152 6656
rect 22652 6604 22704 6656
rect 24032 6647 24084 6656
rect 24032 6613 24041 6647
rect 24041 6613 24075 6647
rect 24075 6613 24084 6647
rect 24032 6604 24084 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1492 6400 1544 6452
rect 3516 6443 3568 6452
rect 3516 6409 3525 6443
rect 3525 6409 3559 6443
rect 3559 6409 3568 6443
rect 3516 6400 3568 6409
rect 4252 6443 4304 6452
rect 4252 6409 4261 6443
rect 4261 6409 4295 6443
rect 4295 6409 4304 6443
rect 4252 6400 4304 6409
rect 5448 6400 5500 6452
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 8024 6400 8076 6452
rect 10784 6443 10836 6452
rect 10784 6409 10793 6443
rect 10793 6409 10827 6443
rect 10827 6409 10836 6443
rect 10784 6400 10836 6409
rect 13636 6443 13688 6452
rect 13636 6409 13645 6443
rect 13645 6409 13679 6443
rect 13679 6409 13688 6443
rect 13636 6400 13688 6409
rect 17408 6400 17460 6452
rect 18880 6443 18932 6452
rect 18880 6409 18889 6443
rect 18889 6409 18923 6443
rect 18923 6409 18932 6443
rect 18880 6400 18932 6409
rect 19616 6400 19668 6452
rect 20812 6443 20864 6452
rect 20812 6409 20821 6443
rect 20821 6409 20855 6443
rect 20855 6409 20864 6443
rect 20812 6400 20864 6409
rect 22652 6400 22704 6452
rect 5080 6264 5132 6316
rect 7564 6375 7616 6384
rect 7564 6341 7573 6375
rect 7573 6341 7607 6375
rect 7607 6341 7616 6375
rect 12532 6375 12584 6384
rect 7564 6332 7616 6341
rect 12532 6341 12541 6375
rect 12541 6341 12575 6375
rect 12575 6341 12584 6375
rect 12532 6332 12584 6341
rect 23296 6332 23348 6384
rect 2228 6196 2280 6248
rect 2688 6196 2740 6248
rect 8392 6196 8444 6248
rect 9772 6196 9824 6248
rect 11336 6239 11388 6248
rect 11336 6205 11345 6239
rect 11345 6205 11379 6239
rect 11379 6205 11388 6239
rect 11336 6196 11388 6205
rect 3240 6128 3292 6180
rect 5724 6171 5776 6180
rect 5724 6137 5733 6171
rect 5733 6137 5767 6171
rect 5767 6137 5776 6171
rect 5724 6128 5776 6137
rect 9680 6128 9732 6180
rect 10692 6128 10744 6180
rect 13544 6264 13596 6316
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 19248 6264 19300 6316
rect 22376 6264 22428 6316
rect 23388 6264 23440 6316
rect 14096 6239 14148 6248
rect 6000 6060 6052 6112
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 10140 6103 10192 6112
rect 10140 6069 10149 6103
rect 10149 6069 10183 6103
rect 10183 6069 10192 6103
rect 10140 6060 10192 6069
rect 12256 6103 12308 6112
rect 12256 6069 12265 6103
rect 12265 6069 12299 6103
rect 12299 6069 12308 6103
rect 12256 6060 12308 6069
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 16580 6239 16632 6248
rect 16580 6205 16589 6239
rect 16589 6205 16623 6239
rect 16623 6205 16632 6239
rect 16580 6196 16632 6205
rect 18052 6239 18104 6248
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 18880 6196 18932 6248
rect 20260 6196 20312 6248
rect 25596 6239 25648 6248
rect 13084 6171 13136 6180
rect 13084 6137 13093 6171
rect 13093 6137 13127 6171
rect 13127 6137 13136 6171
rect 13084 6128 13136 6137
rect 14004 6128 14056 6180
rect 13176 6060 13228 6112
rect 15384 6060 15436 6112
rect 16120 6128 16172 6180
rect 22560 6171 22612 6180
rect 22560 6137 22569 6171
rect 22569 6137 22603 6171
rect 22603 6137 22612 6171
rect 22560 6128 22612 6137
rect 25596 6205 25605 6239
rect 25605 6205 25639 6239
rect 25639 6205 25648 6239
rect 25596 6196 25648 6205
rect 24032 6128 24084 6180
rect 15568 6060 15620 6112
rect 17316 6103 17368 6112
rect 17316 6069 17325 6103
rect 17325 6069 17359 6103
rect 17359 6069 17368 6103
rect 17316 6060 17368 6069
rect 21180 6060 21232 6112
rect 24124 6060 24176 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1400 5899 1452 5908
rect 1400 5865 1409 5899
rect 1409 5865 1443 5899
rect 1443 5865 1452 5899
rect 1400 5856 1452 5865
rect 2228 5899 2280 5908
rect 2228 5865 2237 5899
rect 2237 5865 2271 5899
rect 2271 5865 2280 5899
rect 2228 5856 2280 5865
rect 4712 5856 4764 5908
rect 4988 5899 5040 5908
rect 4988 5865 4997 5899
rect 4997 5865 5031 5899
rect 5031 5865 5040 5899
rect 4988 5856 5040 5865
rect 5172 5856 5224 5908
rect 6368 5856 6420 5908
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 6920 5856 6972 5908
rect 8944 5899 8996 5908
rect 2872 5788 2924 5840
rect 5080 5831 5132 5840
rect 5080 5797 5089 5831
rect 5089 5797 5123 5831
rect 5123 5797 5132 5831
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 9680 5899 9732 5908
rect 9680 5865 9689 5899
rect 9689 5865 9723 5899
rect 9723 5865 9732 5899
rect 9680 5856 9732 5865
rect 11060 5856 11112 5908
rect 11612 5856 11664 5908
rect 13084 5856 13136 5908
rect 13820 5856 13872 5908
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 19156 5856 19208 5908
rect 20076 5899 20128 5908
rect 20076 5865 20085 5899
rect 20085 5865 20119 5899
rect 20119 5865 20128 5899
rect 20076 5856 20128 5865
rect 22560 5856 22612 5908
rect 5080 5788 5132 5797
rect 8116 5831 8168 5840
rect 8116 5797 8125 5831
rect 8125 5797 8159 5831
rect 8159 5797 8168 5831
rect 8116 5788 8168 5797
rect 3332 5720 3384 5772
rect 4068 5720 4120 5772
rect 4528 5720 4580 5772
rect 8392 5788 8444 5840
rect 10140 5788 10192 5840
rect 11152 5788 11204 5840
rect 10968 5763 11020 5772
rect 10968 5729 11002 5763
rect 11002 5729 11020 5763
rect 10968 5720 11020 5729
rect 13728 5788 13780 5840
rect 14188 5831 14240 5840
rect 14188 5797 14197 5831
rect 14197 5797 14231 5831
rect 14231 5797 14240 5831
rect 14188 5788 14240 5797
rect 15384 5788 15436 5840
rect 17224 5788 17276 5840
rect 21732 5788 21784 5840
rect 22192 5788 22244 5840
rect 15200 5720 15252 5772
rect 19340 5720 19392 5772
rect 20996 5720 21048 5772
rect 2596 5652 2648 5704
rect 3516 5652 3568 5704
rect 5080 5652 5132 5704
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 5356 5584 5408 5636
rect 6092 5627 6144 5636
rect 6092 5593 6101 5627
rect 6101 5593 6135 5627
rect 6135 5593 6144 5627
rect 6092 5584 6144 5593
rect 2504 5559 2556 5568
rect 2504 5525 2513 5559
rect 2513 5525 2547 5559
rect 2547 5525 2556 5559
rect 2504 5516 2556 5525
rect 4068 5516 4120 5568
rect 6000 5516 6052 5568
rect 7840 5584 7892 5636
rect 8576 5627 8628 5636
rect 8576 5593 8585 5627
rect 8585 5593 8619 5627
rect 8619 5593 8628 5627
rect 8576 5584 8628 5593
rect 9496 5627 9548 5636
rect 9496 5593 9505 5627
rect 9505 5593 9539 5627
rect 9539 5593 9548 5627
rect 9496 5584 9548 5593
rect 13728 5627 13780 5636
rect 13728 5593 13737 5627
rect 13737 5593 13771 5627
rect 13771 5593 13780 5627
rect 13728 5584 13780 5593
rect 14096 5584 14148 5636
rect 15568 5584 15620 5636
rect 16396 5584 16448 5636
rect 19248 5652 19300 5704
rect 20628 5652 20680 5704
rect 20812 5652 20864 5704
rect 21732 5652 21784 5704
rect 23112 5856 23164 5908
rect 24032 5856 24084 5908
rect 25504 5899 25556 5908
rect 25504 5865 25513 5899
rect 25513 5865 25547 5899
rect 25547 5865 25556 5899
rect 25504 5856 25556 5865
rect 22928 5788 22980 5840
rect 23388 5788 23440 5840
rect 23848 5720 23900 5772
rect 25412 5720 25464 5772
rect 22928 5652 22980 5704
rect 23112 5695 23164 5704
rect 23112 5661 23121 5695
rect 23121 5661 23155 5695
rect 23155 5661 23164 5695
rect 23112 5652 23164 5661
rect 24860 5652 24912 5704
rect 22376 5584 22428 5636
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 13544 5559 13596 5568
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 15292 5516 15344 5568
rect 16672 5516 16724 5568
rect 17868 5559 17920 5568
rect 17868 5525 17877 5559
rect 17877 5525 17911 5559
rect 17911 5525 17920 5559
rect 17868 5516 17920 5525
rect 18972 5559 19024 5568
rect 18972 5525 18981 5559
rect 18981 5525 19015 5559
rect 19015 5525 19024 5559
rect 18972 5516 19024 5525
rect 19156 5559 19208 5568
rect 19156 5525 19165 5559
rect 19165 5525 19199 5559
rect 19199 5525 19208 5559
rect 19156 5516 19208 5525
rect 22560 5559 22612 5568
rect 22560 5525 22569 5559
rect 22569 5525 22603 5559
rect 22603 5525 22612 5559
rect 22560 5516 22612 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2688 5312 2740 5364
rect 3332 5312 3384 5364
rect 4988 5312 5040 5364
rect 6552 5355 6604 5364
rect 6552 5321 6561 5355
rect 6561 5321 6595 5355
rect 6595 5321 6604 5355
rect 6552 5312 6604 5321
rect 7104 5312 7156 5364
rect 8116 5312 8168 5364
rect 8392 5312 8444 5364
rect 9772 5355 9824 5364
rect 9772 5321 9781 5355
rect 9781 5321 9815 5355
rect 9815 5321 9824 5355
rect 9772 5312 9824 5321
rect 10876 5312 10928 5364
rect 11152 5312 11204 5364
rect 14188 5312 14240 5364
rect 15384 5355 15436 5364
rect 15384 5321 15393 5355
rect 15393 5321 15427 5355
rect 15427 5321 15436 5355
rect 15384 5312 15436 5321
rect 15844 5355 15896 5364
rect 15844 5321 15853 5355
rect 15853 5321 15887 5355
rect 15887 5321 15896 5355
rect 15844 5312 15896 5321
rect 16396 5312 16448 5364
rect 17224 5355 17276 5364
rect 17224 5321 17233 5355
rect 17233 5321 17267 5355
rect 17267 5321 17276 5355
rect 17224 5312 17276 5321
rect 18880 5312 18932 5364
rect 2228 5244 2280 5296
rect 3700 5287 3752 5296
rect 3700 5253 3709 5287
rect 3709 5253 3743 5287
rect 3743 5253 3752 5287
rect 3700 5244 3752 5253
rect 2688 5219 2740 5228
rect 2688 5185 2697 5219
rect 2697 5185 2731 5219
rect 2731 5185 2740 5219
rect 2688 5176 2740 5185
rect 6460 5244 6512 5296
rect 14280 5287 14332 5296
rect 7196 5176 7248 5228
rect 10784 5219 10836 5228
rect 10784 5185 10793 5219
rect 10793 5185 10827 5219
rect 10827 5185 10836 5219
rect 10784 5176 10836 5185
rect 14280 5253 14289 5287
rect 14289 5253 14323 5287
rect 14323 5253 14332 5287
rect 14280 5244 14332 5253
rect 14004 5176 14056 5228
rect 14372 5176 14424 5228
rect 16212 5219 16264 5228
rect 2412 5151 2464 5160
rect 2412 5117 2421 5151
rect 2421 5117 2455 5151
rect 2455 5117 2464 5151
rect 2412 5108 2464 5117
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 7564 5108 7616 5160
rect 8208 5108 8260 5160
rect 10232 5108 10284 5160
rect 10692 5108 10744 5160
rect 2504 5040 2556 5092
rect 3976 5083 4028 5092
rect 3976 5049 3985 5083
rect 3985 5049 4019 5083
rect 4019 5049 4028 5083
rect 3976 5040 4028 5049
rect 4068 5040 4120 5092
rect 5356 5040 5408 5092
rect 6000 5040 6052 5092
rect 6736 5040 6788 5092
rect 8116 5040 8168 5092
rect 11336 5108 11388 5160
rect 12256 5108 12308 5160
rect 14464 5108 14516 5160
rect 15108 5108 15160 5160
rect 16212 5185 16221 5219
rect 16221 5185 16255 5219
rect 16255 5185 16264 5219
rect 16212 5176 16264 5185
rect 20260 5312 20312 5364
rect 20904 5312 20956 5364
rect 23388 5312 23440 5364
rect 23848 5312 23900 5364
rect 24768 5355 24820 5364
rect 24768 5321 24777 5355
rect 24777 5321 24811 5355
rect 24811 5321 24820 5355
rect 24768 5312 24820 5321
rect 25412 5355 25464 5364
rect 25412 5321 25421 5355
rect 25421 5321 25455 5355
rect 25455 5321 25464 5355
rect 25412 5312 25464 5321
rect 22192 5244 22244 5296
rect 23112 5244 23164 5296
rect 24124 5244 24176 5296
rect 22928 5176 22980 5228
rect 23756 5176 23808 5228
rect 24768 5176 24820 5228
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 22744 5108 22796 5160
rect 24584 5151 24636 5160
rect 24584 5117 24593 5151
rect 24593 5117 24627 5151
rect 24627 5117 24636 5151
rect 24584 5108 24636 5117
rect 13176 5083 13228 5092
rect 13176 5049 13185 5083
rect 13185 5049 13219 5083
rect 13219 5049 13228 5083
rect 13176 5040 13228 5049
rect 13912 5040 13964 5092
rect 14832 5083 14884 5092
rect 14832 5049 14841 5083
rect 14841 5049 14875 5083
rect 14875 5049 14884 5083
rect 14832 5040 14884 5049
rect 16488 5040 16540 5092
rect 18972 5040 19024 5092
rect 19524 5083 19576 5092
rect 19524 5049 19558 5083
rect 19558 5049 19576 5083
rect 19524 5040 19576 5049
rect 22652 5040 22704 5092
rect 23204 5040 23256 5092
rect 4160 5015 4212 5024
rect 4160 4981 4169 5015
rect 4169 4981 4203 5015
rect 4203 4981 4212 5015
rect 4160 4972 4212 4981
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 10140 5015 10192 5024
rect 10140 4981 10149 5015
rect 10149 4981 10183 5015
rect 10183 4981 10192 5015
rect 10140 4972 10192 4981
rect 10968 4972 11020 5024
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1768 4768 1820 4820
rect 2596 4768 2648 4820
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 4620 4811 4672 4820
rect 4620 4777 4629 4811
rect 4629 4777 4663 4811
rect 4663 4777 4672 4811
rect 4620 4768 4672 4777
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 6184 4811 6236 4820
rect 6184 4777 6193 4811
rect 6193 4777 6227 4811
rect 6227 4777 6236 4811
rect 6184 4768 6236 4777
rect 7932 4768 7984 4820
rect 8208 4811 8260 4820
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 9404 4811 9456 4820
rect 9404 4777 9413 4811
rect 9413 4777 9447 4811
rect 9447 4777 9456 4811
rect 9404 4768 9456 4777
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 13176 4768 13228 4820
rect 14280 4768 14332 4820
rect 14372 4768 14424 4820
rect 19340 4768 19392 4820
rect 21364 4768 21416 4820
rect 22652 4768 22704 4820
rect 25228 4811 25280 4820
rect 25228 4777 25237 4811
rect 25237 4777 25271 4811
rect 25271 4777 25280 4811
rect 25228 4768 25280 4777
rect 25596 4811 25648 4820
rect 25596 4777 25605 4811
rect 25605 4777 25639 4811
rect 25639 4777 25648 4811
rect 25596 4768 25648 4777
rect 2780 4743 2832 4752
rect 2780 4709 2789 4743
rect 2789 4709 2823 4743
rect 2823 4709 2832 4743
rect 2780 4700 2832 4709
rect 2688 4632 2740 4684
rect 4068 4700 4120 4752
rect 4436 4743 4488 4752
rect 4436 4709 4445 4743
rect 4445 4709 4479 4743
rect 4479 4709 4488 4743
rect 4436 4700 4488 4709
rect 4804 4700 4856 4752
rect 5080 4700 5132 4752
rect 6092 4700 6144 4752
rect 8392 4700 8444 4752
rect 8576 4743 8628 4752
rect 8576 4709 8585 4743
rect 8585 4709 8619 4743
rect 8619 4709 8628 4743
rect 8576 4700 8628 4709
rect 13268 4743 13320 4752
rect 13268 4709 13277 4743
rect 13277 4709 13311 4743
rect 13311 4709 13320 4743
rect 13268 4700 13320 4709
rect 13912 4700 13964 4752
rect 19248 4700 19300 4752
rect 19616 4743 19668 4752
rect 19616 4709 19625 4743
rect 19625 4709 19659 4743
rect 19659 4709 19668 4743
rect 19616 4700 19668 4709
rect 20168 4700 20220 4752
rect 20352 4700 20404 4752
rect 4160 4632 4212 4684
rect 5448 4632 5500 4684
rect 6644 4632 6696 4684
rect 8116 4632 8168 4684
rect 9680 4632 9732 4684
rect 13728 4632 13780 4684
rect 14832 4632 14884 4684
rect 16120 4675 16172 4684
rect 1584 4564 1636 4616
rect 4988 4564 5040 4616
rect 6460 4564 6512 4616
rect 7748 4607 7800 4616
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 8208 4564 8260 4616
rect 3056 4496 3108 4548
rect 5264 4496 5316 4548
rect 7932 4496 7984 4548
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 7840 4428 7892 4480
rect 8300 4428 8352 4480
rect 9588 4428 9640 4480
rect 11152 4471 11204 4480
rect 11152 4437 11161 4471
rect 11161 4437 11195 4471
rect 11195 4437 11204 4471
rect 11152 4428 11204 4437
rect 11704 4471 11756 4480
rect 11704 4437 11713 4471
rect 11713 4437 11747 4471
rect 11747 4437 11756 4471
rect 11704 4428 11756 4437
rect 12348 4428 12400 4480
rect 12992 4471 13044 4480
rect 12992 4437 13001 4471
rect 13001 4437 13035 4471
rect 13035 4437 13044 4471
rect 12992 4428 13044 4437
rect 14832 4428 14884 4480
rect 16120 4641 16154 4675
rect 16154 4641 16172 4675
rect 16120 4632 16172 4641
rect 16672 4632 16724 4684
rect 18420 4632 18472 4684
rect 18972 4632 19024 4684
rect 19524 4632 19576 4684
rect 20260 4632 20312 4684
rect 23112 4700 23164 4752
rect 20904 4632 20956 4684
rect 22100 4632 22152 4684
rect 22652 4632 22704 4684
rect 24952 4632 25004 4684
rect 15660 4564 15712 4616
rect 20812 4564 20864 4616
rect 20996 4539 21048 4548
rect 20996 4505 21005 4539
rect 21005 4505 21039 4539
rect 21039 4505 21048 4539
rect 20996 4496 21048 4505
rect 15844 4428 15896 4480
rect 17224 4471 17276 4480
rect 17224 4437 17233 4471
rect 17233 4437 17267 4471
rect 17267 4437 17276 4471
rect 17224 4428 17276 4437
rect 19892 4428 19944 4480
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 22376 4471 22428 4480
rect 22376 4437 22385 4471
rect 22385 4437 22419 4471
rect 22419 4437 22428 4471
rect 22376 4428 22428 4437
rect 23480 4428 23532 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2872 4267 2924 4276
rect 2872 4233 2881 4267
rect 2881 4233 2915 4267
rect 2915 4233 2924 4267
rect 2872 4224 2924 4233
rect 4988 4267 5040 4276
rect 4988 4233 4997 4267
rect 4997 4233 5031 4267
rect 5031 4233 5040 4267
rect 4988 4224 5040 4233
rect 6184 4267 6236 4276
rect 6184 4233 6193 4267
rect 6193 4233 6227 4267
rect 6227 4233 6236 4267
rect 6184 4224 6236 4233
rect 6644 4267 6696 4276
rect 6644 4233 6653 4267
rect 6653 4233 6687 4267
rect 6687 4233 6696 4267
rect 6644 4224 6696 4233
rect 7748 4224 7800 4276
rect 8392 4224 8444 4276
rect 9128 4267 9180 4276
rect 9128 4233 9137 4267
rect 9137 4233 9171 4267
rect 9171 4233 9180 4267
rect 9128 4224 9180 4233
rect 10692 4267 10744 4276
rect 10692 4233 10701 4267
rect 10701 4233 10735 4267
rect 10735 4233 10744 4267
rect 10692 4224 10744 4233
rect 13268 4224 13320 4276
rect 19616 4224 19668 4276
rect 20904 4267 20956 4276
rect 20904 4233 20913 4267
rect 20913 4233 20947 4267
rect 20947 4233 20956 4267
rect 20904 4224 20956 4233
rect 22652 4224 22704 4276
rect 23112 4224 23164 4276
rect 24952 4224 25004 4276
rect 2780 4156 2832 4208
rect 2320 4088 2372 4140
rect 1952 4020 2004 4072
rect 1860 3952 1912 4004
rect 2596 3952 2648 4004
rect 3516 4020 3568 4072
rect 3608 4020 3660 4072
rect 6460 4156 6512 4208
rect 7196 4156 7248 4208
rect 8576 4156 8628 4208
rect 9680 4156 9732 4208
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 8116 4131 8168 4140
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 9588 4088 9640 4140
rect 5448 4063 5500 4072
rect 5448 4029 5457 4063
rect 5457 4029 5491 4063
rect 5491 4029 5500 4063
rect 5448 4020 5500 4029
rect 10048 4088 10100 4140
rect 11612 4063 11664 4072
rect 11612 4029 11621 4063
rect 11621 4029 11655 4063
rect 11655 4029 11664 4063
rect 11612 4020 11664 4029
rect 14188 4088 14240 4140
rect 14832 4131 14884 4140
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 17960 4088 18012 4140
rect 18880 4131 18932 4140
rect 18880 4097 18889 4131
rect 18889 4097 18923 4131
rect 18923 4097 18932 4131
rect 18880 4088 18932 4097
rect 19892 4088 19944 4140
rect 20260 4156 20312 4208
rect 22560 4088 22612 4140
rect 23020 4088 23072 4140
rect 24860 4131 24912 4140
rect 24860 4097 24869 4131
rect 24869 4097 24903 4131
rect 24903 4097 24912 4131
rect 24860 4088 24912 4097
rect 16764 4063 16816 4072
rect 16764 4029 16773 4063
rect 16773 4029 16807 4063
rect 16807 4029 16816 4063
rect 16764 4020 16816 4029
rect 18144 4020 18196 4072
rect 21180 4020 21232 4072
rect 23664 4063 23716 4072
rect 23664 4029 23673 4063
rect 23673 4029 23707 4063
rect 23707 4029 23716 4063
rect 23664 4020 23716 4029
rect 3332 3952 3384 4004
rect 4068 3952 4120 4004
rect 6368 3952 6420 4004
rect 7288 3952 7340 4004
rect 9496 3952 9548 4004
rect 9588 3995 9640 4004
rect 9588 3961 9597 3995
rect 9597 3961 9631 3995
rect 9631 3961 9640 3995
rect 9588 3952 9640 3961
rect 11980 3952 12032 4004
rect 12992 3995 13044 4004
rect 12992 3961 13001 3995
rect 13001 3961 13035 3995
rect 13035 3961 13044 3995
rect 12992 3952 13044 3961
rect 13268 3995 13320 4004
rect 13268 3961 13277 3995
rect 13277 3961 13311 3995
rect 13311 3961 13320 3995
rect 13268 3952 13320 3961
rect 15476 3952 15528 4004
rect 18420 3952 18472 4004
rect 19432 3952 19484 4004
rect 22008 3995 22060 4004
rect 1492 3927 1544 3936
rect 1492 3893 1525 3927
rect 1525 3893 1544 3927
rect 1492 3884 1544 3893
rect 2228 3884 2280 3936
rect 5172 3884 5224 3936
rect 12900 3884 12952 3936
rect 14372 3884 14424 3936
rect 15384 3884 15436 3936
rect 15568 3884 15620 3936
rect 16488 3884 16540 3936
rect 17132 3927 17184 3936
rect 17132 3893 17141 3927
rect 17141 3893 17175 3927
rect 17175 3893 17184 3927
rect 17132 3884 17184 3893
rect 18880 3884 18932 3936
rect 22008 3961 22033 3995
rect 22033 3961 22060 3995
rect 22008 3952 22060 3961
rect 21180 3884 21232 3936
rect 21732 3884 21784 3936
rect 22836 3952 22888 4004
rect 23480 3952 23532 4004
rect 25228 3952 25280 4004
rect 22192 3884 22244 3936
rect 25136 3927 25188 3936
rect 25136 3893 25145 3927
rect 25145 3893 25179 3927
rect 25179 3893 25188 3927
rect 25136 3884 25188 3893
rect 26240 3927 26292 3936
rect 26240 3893 26249 3927
rect 26249 3893 26283 3927
rect 26283 3893 26292 3927
rect 26240 3884 26292 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1676 3680 1728 3732
rect 2688 3680 2740 3732
rect 3056 3680 3108 3732
rect 3332 3680 3384 3732
rect 3516 3680 3568 3732
rect 5172 3680 5224 3732
rect 6644 3680 6696 3732
rect 7288 3680 7340 3732
rect 7564 3680 7616 3732
rect 8484 3680 8536 3732
rect 9680 3680 9732 3732
rect 11060 3680 11112 3732
rect 13268 3680 13320 3732
rect 14556 3680 14608 3732
rect 15844 3723 15896 3732
rect 15844 3689 15853 3723
rect 15853 3689 15887 3723
rect 15887 3689 15896 3723
rect 15844 3680 15896 3689
rect 18512 3680 18564 3732
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 20812 3680 20864 3732
rect 22284 3723 22336 3732
rect 22284 3689 22293 3723
rect 22293 3689 22327 3723
rect 22327 3689 22336 3723
rect 22284 3680 22336 3689
rect 23480 3680 23532 3732
rect 25320 3680 25372 3732
rect 25412 3680 25464 3732
rect 3700 3612 3752 3664
rect 6000 3612 6052 3664
rect 6736 3612 6788 3664
rect 14188 3612 14240 3664
rect 15660 3655 15712 3664
rect 15660 3621 15669 3655
rect 15669 3621 15703 3655
rect 15703 3621 15712 3655
rect 15660 3612 15712 3621
rect 16764 3612 16816 3664
rect 19984 3612 20036 3664
rect 21824 3612 21876 3664
rect 22836 3655 22888 3664
rect 22836 3621 22870 3655
rect 22870 3621 22888 3655
rect 22836 3612 22888 3621
rect 23572 3612 23624 3664
rect 23756 3612 23808 3664
rect 4068 3587 4120 3596
rect 4068 3553 4077 3587
rect 4077 3553 4111 3587
rect 4111 3553 4120 3587
rect 4068 3544 4120 3553
rect 6276 3544 6328 3596
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3332 3476 3384 3528
rect 3884 3476 3936 3528
rect 2504 3451 2556 3460
rect 2504 3417 2513 3451
rect 2513 3417 2547 3451
rect 2547 3417 2556 3451
rect 2504 3408 2556 3417
rect 1952 3383 2004 3392
rect 1952 3349 1961 3383
rect 1961 3349 1995 3383
rect 1995 3349 2004 3383
rect 1952 3340 2004 3349
rect 9128 3544 9180 3596
rect 11152 3544 11204 3596
rect 13728 3544 13780 3596
rect 15568 3544 15620 3596
rect 16948 3587 17000 3596
rect 16948 3553 16957 3587
rect 16957 3553 16991 3587
rect 16991 3553 17000 3587
rect 16948 3544 17000 3553
rect 19432 3587 19484 3596
rect 19432 3553 19441 3587
rect 19441 3553 19475 3587
rect 19475 3553 19484 3587
rect 19432 3544 19484 3553
rect 20996 3544 21048 3596
rect 21640 3544 21692 3596
rect 22192 3544 22244 3596
rect 22652 3544 22704 3596
rect 25044 3587 25096 3596
rect 25044 3553 25053 3587
rect 25053 3553 25087 3587
rect 25087 3553 25096 3587
rect 25044 3544 25096 3553
rect 25320 3544 25372 3596
rect 25964 3544 26016 3596
rect 12716 3519 12768 3528
rect 7104 3408 7156 3460
rect 7932 3408 7984 3460
rect 9496 3408 9548 3460
rect 10048 3408 10100 3460
rect 6460 3340 6512 3392
rect 8116 3383 8168 3392
rect 8116 3349 8125 3383
rect 8125 3349 8159 3383
rect 8159 3349 8168 3383
rect 8116 3340 8168 3349
rect 9404 3340 9456 3392
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 12716 3476 12768 3485
rect 15936 3519 15988 3528
rect 15936 3485 15945 3519
rect 15945 3485 15979 3519
rect 15979 3485 15988 3519
rect 15936 3476 15988 3485
rect 15384 3451 15436 3460
rect 15384 3417 15393 3451
rect 15393 3417 15427 3451
rect 15427 3417 15436 3451
rect 15384 3408 15436 3417
rect 14740 3383 14792 3392
rect 14740 3349 14749 3383
rect 14749 3349 14783 3383
rect 14783 3349 14792 3383
rect 14740 3340 14792 3349
rect 15292 3340 15344 3392
rect 16120 3340 16172 3392
rect 20352 3476 20404 3528
rect 24860 3451 24912 3460
rect 24860 3417 24869 3451
rect 24869 3417 24903 3451
rect 24903 3417 24912 3451
rect 24860 3408 24912 3417
rect 24032 3340 24084 3392
rect 25780 3340 25832 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1952 3136 2004 3188
rect 1492 2932 1544 2984
rect 3332 2932 3384 2984
rect 1676 2907 1728 2916
rect 1676 2873 1685 2907
rect 1685 2873 1719 2907
rect 1719 2873 1728 2907
rect 1676 2864 1728 2873
rect 3148 2864 3200 2916
rect 3056 2796 3108 2848
rect 4068 3136 4120 3188
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 6460 3136 6512 3188
rect 8300 3136 8352 3188
rect 14188 3136 14240 3188
rect 15660 3136 15712 3188
rect 16764 3136 16816 3188
rect 16948 3136 17000 3188
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 18144 3179 18196 3188
rect 18144 3145 18153 3179
rect 18153 3145 18187 3179
rect 18187 3145 18196 3179
rect 18144 3136 18196 3145
rect 19340 3179 19392 3188
rect 19340 3145 19349 3179
rect 19349 3145 19383 3179
rect 19383 3145 19392 3179
rect 19340 3136 19392 3145
rect 19984 3136 20036 3188
rect 20444 3136 20496 3188
rect 20996 3179 21048 3188
rect 20996 3145 21005 3179
rect 21005 3145 21039 3179
rect 21039 3145 21048 3179
rect 20996 3136 21048 3145
rect 22376 3179 22428 3188
rect 22376 3145 22385 3179
rect 22385 3145 22419 3179
rect 22419 3145 22428 3179
rect 22376 3136 22428 3145
rect 22836 3136 22888 3188
rect 24952 3179 25004 3188
rect 24952 3145 24961 3179
rect 24961 3145 24995 3179
rect 24995 3145 25004 3179
rect 24952 3136 25004 3145
rect 25044 3136 25096 3188
rect 17960 3068 18012 3120
rect 19708 3111 19760 3120
rect 5724 2907 5776 2916
rect 5724 2873 5733 2907
rect 5733 2873 5767 2907
rect 5767 2873 5776 2907
rect 5724 2864 5776 2873
rect 6460 2932 6512 2984
rect 6920 2932 6972 2984
rect 7104 2975 7156 2984
rect 7104 2941 7138 2975
rect 7138 2941 7156 2975
rect 7104 2932 7156 2941
rect 9404 2932 9456 2984
rect 12716 2975 12768 2984
rect 12716 2941 12725 2975
rect 12725 2941 12759 2975
rect 12759 2941 12768 2975
rect 12716 2932 12768 2941
rect 4252 2796 4304 2848
rect 10692 2839 10744 2848
rect 10692 2805 10701 2839
rect 10701 2805 10735 2839
rect 10735 2805 10744 2839
rect 10692 2796 10744 2805
rect 11152 2796 11204 2848
rect 13728 2932 13780 2984
rect 15568 2932 15620 2984
rect 19708 3077 19717 3111
rect 19717 3077 19751 3111
rect 19751 3077 19760 3111
rect 19708 3068 19760 3077
rect 22652 3068 22704 3120
rect 24492 3111 24544 3120
rect 24492 3077 24501 3111
rect 24501 3077 24535 3111
rect 24535 3077 24544 3111
rect 24492 3068 24544 3077
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 21456 3000 21508 3009
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 25688 3000 25740 3052
rect 20536 2932 20588 2984
rect 20720 2932 20772 2984
rect 22376 2932 22428 2984
rect 23756 2975 23808 2984
rect 23756 2941 23765 2975
rect 23765 2941 23799 2975
rect 23799 2941 23808 2975
rect 23756 2932 23808 2941
rect 24952 2932 25004 2984
rect 26240 2975 26292 2984
rect 26240 2941 26249 2975
rect 26249 2941 26283 2975
rect 26283 2941 26292 2975
rect 26240 2932 26292 2941
rect 14740 2864 14792 2916
rect 16672 2864 16724 2916
rect 18696 2907 18748 2916
rect 18696 2873 18705 2907
rect 18705 2873 18739 2907
rect 18739 2873 18748 2907
rect 18696 2864 18748 2873
rect 19708 2864 19760 2916
rect 20168 2839 20220 2848
rect 20168 2805 20177 2839
rect 20177 2805 20211 2839
rect 20211 2805 20220 2839
rect 20168 2796 20220 2805
rect 22652 2839 22704 2848
rect 22652 2805 22661 2839
rect 22661 2805 22695 2839
rect 22695 2805 22704 2839
rect 22652 2796 22704 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1584 2592 1636 2644
rect 3884 2635 3936 2644
rect 2136 2524 2188 2576
rect 3884 2601 3893 2635
rect 3893 2601 3927 2635
rect 3927 2601 3936 2635
rect 3884 2592 3936 2601
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 7196 2592 7248 2644
rect 7932 2635 7984 2644
rect 2964 2567 3016 2576
rect 2964 2533 2973 2567
rect 2973 2533 3007 2567
rect 3007 2533 3016 2567
rect 2964 2524 3016 2533
rect 3056 2567 3108 2576
rect 3056 2533 3065 2567
rect 3065 2533 3099 2567
rect 3099 2533 3108 2567
rect 3056 2524 3108 2533
rect 4252 2524 4304 2576
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 9404 2592 9456 2644
rect 11152 2635 11204 2644
rect 6644 2499 6696 2508
rect 6644 2465 6653 2499
rect 6653 2465 6687 2499
rect 6687 2465 6696 2499
rect 6644 2456 6696 2465
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 14648 2592 14700 2644
rect 10692 2524 10744 2576
rect 13636 2524 13688 2576
rect 15936 2592 15988 2644
rect 16028 2567 16080 2576
rect 16028 2533 16037 2567
rect 16037 2533 16071 2567
rect 16071 2533 16080 2567
rect 16028 2524 16080 2533
rect 16856 2592 16908 2644
rect 19340 2592 19392 2644
rect 20536 2592 20588 2644
rect 16672 2524 16724 2576
rect 17224 2524 17276 2576
rect 18696 2524 18748 2576
rect 21732 2567 21784 2576
rect 9128 2388 9180 2440
rect 12808 2456 12860 2508
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14832 2499 14884 2508
rect 14188 2456 14240 2465
rect 14832 2465 14841 2499
rect 14841 2465 14875 2499
rect 14875 2465 14884 2499
rect 14832 2456 14884 2465
rect 17132 2456 17184 2508
rect 19984 2456 20036 2508
rect 20996 2456 21048 2508
rect 21732 2533 21741 2567
rect 21741 2533 21775 2567
rect 21775 2533 21784 2567
rect 21732 2524 21784 2533
rect 24216 2524 24268 2576
rect 22928 2456 22980 2508
rect 23480 2456 23532 2508
rect 25136 2499 25188 2508
rect 25136 2465 25145 2499
rect 25145 2465 25179 2499
rect 25179 2465 25188 2499
rect 25136 2456 25188 2465
rect 15292 2388 15344 2440
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 20168 2388 20220 2440
rect 7012 2363 7064 2372
rect 7012 2329 7021 2363
rect 7021 2329 7055 2363
rect 7055 2329 7064 2363
rect 7012 2320 7064 2329
rect 12808 2363 12860 2372
rect 12808 2329 12817 2363
rect 12817 2329 12851 2363
rect 12851 2329 12860 2363
rect 12808 2320 12860 2329
rect 13912 2363 13964 2372
rect 13912 2329 13921 2363
rect 13921 2329 13955 2363
rect 13955 2329 13964 2363
rect 13912 2320 13964 2329
rect 15476 2320 15528 2372
rect 18420 2363 18472 2372
rect 18420 2329 18429 2363
rect 18429 2329 18463 2363
rect 18463 2329 18472 2363
rect 18420 2320 18472 2329
rect 23664 2431 23716 2440
rect 23664 2397 23673 2431
rect 23673 2397 23707 2431
rect 23707 2397 23716 2431
rect 23664 2388 23716 2397
rect 25044 2388 25096 2440
rect 20996 2320 21048 2372
rect 21732 2320 21784 2372
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 8668 2295 8720 2304
rect 8668 2261 8677 2295
rect 8677 2261 8711 2295
rect 8711 2261 8720 2295
rect 8668 2252 8720 2261
rect 11704 2295 11756 2304
rect 11704 2261 11713 2295
rect 11713 2261 11747 2295
rect 11747 2261 11756 2295
rect 11704 2252 11756 2261
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 17224 2295 17276 2304
rect 17224 2261 17233 2295
rect 17233 2261 17267 2295
rect 17267 2261 17276 2295
rect 17224 2252 17276 2261
rect 20904 2295 20956 2304
rect 20904 2261 20913 2295
rect 20913 2261 20947 2295
rect 20947 2261 20956 2295
rect 20904 2252 20956 2261
rect 22928 2295 22980 2304
rect 22928 2261 22937 2295
rect 22937 2261 22971 2295
rect 22971 2261 22980 2295
rect 22928 2252 22980 2261
rect 25504 2295 25556 2304
rect 25504 2261 25513 2295
rect 25513 2261 25547 2295
rect 25547 2261 25556 2295
rect 25504 2252 25556 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 11428 2048 11480 2100
rect 16028 2048 16080 2100
rect 13544 1572 13596 1624
rect 15384 1572 15436 1624
rect 22560 1572 22612 1624
rect 23572 1572 23624 1624
rect 5540 1368 5592 1420
rect 6184 1368 6236 1420
rect 4528 620 4580 672
rect 3148 552 3200 604
rect 3700 552 3752 604
rect 3792 552 3844 604
rect 12164 552 12216 604
rect 12532 552 12584 604
rect 18880 552 18932 604
rect 18972 552 19024 604
<< metal2 >>
rect 2778 27704 2834 27713
rect 2778 27639 2834 27648
rect 23478 27704 23534 27713
rect 23478 27639 23534 27648
rect 2226 26344 2282 26353
rect 2226 26279 2282 26288
rect 756 18080 808 18086
rect 2044 18080 2096 18086
rect 756 18022 808 18028
rect 2042 18048 2044 18057
rect 2096 18048 2098 18057
rect 664 17536 716 17542
rect 664 17478 716 17484
rect 676 10713 704 17478
rect 768 12073 796 18022
rect 2042 17983 2098 17992
rect 2044 17672 2096 17678
rect 2042 17640 2044 17649
rect 2096 17640 2098 17649
rect 2042 17575 2098 17584
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1216 16448 1268 16454
rect 1216 16390 1268 16396
rect 1122 14784 1178 14793
rect 1122 14719 1178 14728
rect 754 12064 810 12073
rect 754 11999 810 12008
rect 662 10704 718 10713
rect 662 10639 718 10648
rect 294 10296 350 10305
rect 294 10231 350 10240
rect 308 480 336 10231
rect 1136 4842 1164 14719
rect 1228 13734 1256 16390
rect 1872 15502 1900 16934
rect 2042 16824 2098 16833
rect 2042 16759 2044 16768
rect 2096 16759 2098 16768
rect 2136 16788 2188 16794
rect 2044 16730 2096 16736
rect 2136 16730 2188 16736
rect 2042 16144 2098 16153
rect 2042 16079 2044 16088
rect 2096 16079 2098 16088
rect 2044 16050 2096 16056
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1596 14385 1624 14758
rect 1582 14376 1638 14385
rect 1582 14311 1638 14320
rect 1400 14272 1452 14278
rect 1398 14240 1400 14249
rect 1452 14240 1454 14249
rect 1398 14175 1454 14184
rect 1674 13968 1730 13977
rect 1780 13938 1808 14962
rect 1674 13903 1730 13912
rect 1768 13932 1820 13938
rect 1216 13728 1268 13734
rect 1216 13670 1268 13676
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1400 13524 1452 13530
rect 1400 13466 1452 13472
rect 1412 12306 1440 13466
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1412 11898 1440 12242
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1400 11144 1452 11150
rect 1398 11112 1400 11121
rect 1452 11112 1454 11121
rect 1398 11047 1454 11056
rect 1400 10192 1452 10198
rect 1400 10134 1452 10140
rect 1412 9178 1440 10134
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1504 8129 1532 13670
rect 1688 13394 1716 13903
rect 1768 13874 1820 13880
rect 1780 13530 1808 13874
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1688 12986 1716 13330
rect 1872 12986 1900 15302
rect 2042 14920 2098 14929
rect 2042 14855 2044 14864
rect 2096 14855 2098 14864
rect 2044 14826 2096 14832
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 2056 13870 2084 14214
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1872 12617 1900 12922
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1858 12608 1914 12617
rect 1858 12543 1914 12552
rect 1964 12458 1992 12786
rect 1955 12430 1992 12458
rect 2056 12442 2084 13806
rect 2044 12436 2096 12442
rect 1955 12424 1983 12430
rect 1780 12396 1983 12424
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1490 8120 1546 8129
rect 1490 8055 1546 8064
rect 1398 7984 1454 7993
rect 1398 7919 1454 7928
rect 1412 5914 1440 7919
rect 1492 6792 1544 6798
rect 1596 6769 1624 12038
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1688 8809 1716 11834
rect 1780 10742 1808 12396
rect 2044 12378 2096 12384
rect 1858 12336 1914 12345
rect 2056 12322 2084 12378
rect 1858 12271 1914 12280
rect 1964 12294 2084 12322
rect 1872 11694 1900 12271
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1964 11558 1992 12294
rect 2042 12200 2098 12209
rect 2042 12135 2098 12144
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1768 10736 1820 10742
rect 1768 10678 1820 10684
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 10130 1808 10406
rect 1872 10266 1900 11494
rect 1964 11354 1992 11494
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1950 11248 2006 11257
rect 1950 11183 2006 11192
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 1674 8800 1730 8809
rect 1674 8735 1730 8744
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1492 6734 1544 6740
rect 1582 6760 1638 6769
rect 1504 6458 1532 6734
rect 1582 6695 1638 6704
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 1688 6202 1716 8570
rect 1780 8090 1808 10066
rect 1872 9722 1900 10202
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1872 8673 1900 8774
rect 1858 8664 1914 8673
rect 1964 8634 1992 11183
rect 1858 8599 1914 8608
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1964 8401 1992 8434
rect 1950 8392 2006 8401
rect 1950 8327 2006 8336
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1766 6896 1822 6905
rect 1766 6831 1768 6840
rect 1820 6831 1822 6840
rect 1768 6802 1820 6808
rect 1504 6174 1716 6202
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1504 5794 1532 6174
rect 1674 6080 1730 6089
rect 1674 6015 1730 6024
rect 860 4814 1164 4842
rect 1412 5766 1532 5794
rect 860 480 888 4814
rect 1412 480 1440 5766
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1492 3936 1544 3942
rect 1490 3904 1492 3913
rect 1544 3904 1546 3913
rect 1490 3839 1546 3848
rect 1504 2990 1532 3839
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1596 2650 1624 4558
rect 1688 3738 1716 6015
rect 1780 4826 1808 6802
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1872 4010 1900 7754
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1964 3398 1992 4014
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1964 3194 1992 3334
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1674 2952 1730 2961
rect 1674 2887 1676 2896
rect 1728 2887 1730 2896
rect 1676 2858 1728 2864
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 2056 480 2084 12135
rect 2148 10033 2176 16730
rect 2240 16289 2268 26279
rect 2502 17776 2558 17785
rect 2502 17711 2504 17720
rect 2556 17711 2558 17720
rect 2504 17682 2556 17688
rect 2516 17338 2544 17682
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2320 17264 2372 17270
rect 2320 17206 2372 17212
rect 2226 16280 2282 16289
rect 2226 16215 2282 16224
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2240 11898 2268 16118
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2332 11778 2360 17206
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 2516 15910 2544 16594
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2516 15745 2544 15846
rect 2502 15736 2558 15745
rect 2502 15671 2558 15680
rect 2608 15586 2636 17478
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2700 16658 2728 16934
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 2424 15558 2636 15586
rect 2424 13025 2452 15558
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2410 13016 2466 13025
rect 2410 12951 2466 12960
rect 2516 12850 2544 15438
rect 2792 15416 2820 27639
rect 3422 27024 3478 27033
rect 3422 26959 3478 26968
rect 3436 26314 3464 26959
rect 22008 26648 22060 26654
rect 22008 26590 22060 26596
rect 14648 26444 14700 26450
rect 14648 26386 14700 26392
rect 3424 26308 3476 26314
rect 3424 26250 3476 26256
rect 11244 26308 11296 26314
rect 11244 26250 11296 26256
rect 3054 25664 3110 25673
rect 3054 25599 3110 25608
rect 3068 24886 3096 25599
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 4526 25120 4582 25129
rect 4526 25055 4582 25064
rect 3056 24880 3108 24886
rect 3056 24822 3108 24828
rect 3974 20496 4030 20505
rect 3974 20431 4030 20440
rect 3790 19816 3846 19825
rect 3790 19751 3846 19760
rect 3238 19136 3294 19145
rect 3238 19071 3294 19080
rect 3148 16992 3200 16998
rect 3146 16960 3148 16969
rect 3200 16960 3202 16969
rect 3146 16895 3202 16904
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2884 15586 2912 16390
rect 2976 15706 3004 16390
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2962 15600 3018 15609
rect 2884 15558 2962 15586
rect 2962 15535 3018 15544
rect 2976 15502 3004 15535
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2792 15388 2912 15416
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2778 15328 2834 15337
rect 2608 14521 2636 15302
rect 2778 15263 2834 15272
rect 2792 14550 2820 15263
rect 2884 15162 2912 15388
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2780 14544 2832 14550
rect 2594 14512 2650 14521
rect 2780 14486 2832 14492
rect 2594 14447 2650 14456
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2516 12238 2544 12650
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2502 12064 2558 12073
rect 2502 11999 2558 12008
rect 2240 11750 2360 11778
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 2240 11393 2268 11750
rect 2318 11656 2374 11665
rect 2318 11591 2320 11600
rect 2372 11591 2374 11600
rect 2320 11562 2372 11568
rect 2226 11384 2282 11393
rect 2226 11319 2282 11328
rect 2332 11082 2360 11562
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 2424 10577 2452 11766
rect 2410 10568 2466 10577
rect 2410 10503 2466 10512
rect 2318 10432 2374 10441
rect 2318 10367 2374 10376
rect 2332 10266 2360 10367
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2412 10056 2464 10062
rect 2134 10024 2190 10033
rect 2412 9998 2464 10004
rect 2134 9959 2190 9968
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2136 9172 2188 9178
rect 2188 9132 2268 9160
rect 2136 9114 2188 9120
rect 2136 8560 2188 8566
rect 2136 8502 2188 8508
rect 2148 4321 2176 8502
rect 2240 8090 2268 9132
rect 2332 8974 2360 9862
rect 2424 9518 2452 9998
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2412 9104 2464 9110
rect 2516 9081 2544 11999
rect 2608 10674 2636 14350
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 13190 2728 14214
rect 2792 14074 2820 14486
rect 2884 14414 2912 15098
rect 3148 14884 3200 14890
rect 3148 14826 3200 14832
rect 3054 14648 3110 14657
rect 3160 14618 3188 14826
rect 3054 14583 3110 14592
rect 3148 14612 3200 14618
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2780 13456 2832 13462
rect 2780 13398 2832 13404
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12646 2728 13126
rect 2792 12646 2820 13398
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2412 9046 2464 9052
rect 2502 9072 2558 9081
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2332 8129 2360 8910
rect 2424 8634 2452 9046
rect 2502 9007 2558 9016
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2516 8430 2544 9007
rect 2700 8514 2728 11494
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2792 10266 2820 10610
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2608 8486 2728 8514
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2318 8120 2374 8129
rect 2228 8084 2280 8090
rect 2318 8055 2374 8064
rect 2228 8026 2280 8032
rect 2240 7410 2268 8026
rect 2410 7848 2466 7857
rect 2608 7818 2636 8486
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2410 7783 2466 7792
rect 2596 7812 2648 7818
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2240 7313 2268 7346
rect 2226 7304 2282 7313
rect 2226 7239 2282 7248
rect 2332 6769 2360 7686
rect 2318 6760 2374 6769
rect 2318 6695 2374 6704
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2240 5914 2268 6190
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 2134 4312 2190 4321
rect 2134 4247 2190 4256
rect 2240 3942 2268 5238
rect 2332 4146 2360 6695
rect 2424 5166 2452 7783
rect 2596 7754 2648 7760
rect 2594 7440 2650 7449
rect 2594 7375 2650 7384
rect 2608 7274 2636 7375
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 2700 6662 2728 8298
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6254 2728 6598
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2792 5896 2820 10066
rect 2884 9489 2912 12786
rect 2962 10976 3018 10985
rect 3068 10962 3096 14583
rect 3148 14554 3200 14560
rect 3160 14346 3188 14554
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3160 14006 3188 14282
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 11898 3188 13126
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3018 10934 3096 10962
rect 2962 10911 3018 10920
rect 2976 10810 3004 10911
rect 2964 10804 3016 10810
rect 3252 10792 3280 19071
rect 3804 16561 3832 19751
rect 3882 17912 3938 17921
rect 3882 17847 3938 17856
rect 3790 16552 3846 16561
rect 3790 16487 3846 16496
rect 3698 16416 3754 16425
rect 3698 16351 3754 16360
rect 3712 15745 3740 16351
rect 3790 15872 3846 15881
rect 3790 15807 3846 15816
rect 3330 15736 3386 15745
rect 3330 15671 3386 15680
rect 3698 15736 3754 15745
rect 3698 15671 3754 15680
rect 3344 14906 3372 15671
rect 3424 15428 3476 15434
rect 3424 15370 3476 15376
rect 3436 15337 3464 15370
rect 3422 15328 3478 15337
rect 3422 15263 3478 15272
rect 3804 14929 3832 15807
rect 3790 14920 3846 14929
rect 3344 14878 3464 14906
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3344 13977 3372 14418
rect 3330 13968 3386 13977
rect 3330 13903 3332 13912
rect 3384 13903 3386 13912
rect 3332 13874 3384 13880
rect 3344 13843 3372 13874
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3344 12918 3372 13126
rect 3332 12912 3384 12918
rect 3332 12854 3384 12860
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3344 12345 3372 12582
rect 3330 12336 3386 12345
rect 3330 12271 3386 12280
rect 3436 12186 3464 14878
rect 3790 14855 3846 14864
rect 3896 14657 3924 17847
rect 3988 15745 4016 20431
rect 4434 16688 4490 16697
rect 4068 16652 4120 16658
rect 4434 16623 4436 16632
rect 4068 16594 4120 16600
rect 4488 16623 4490 16632
rect 4436 16594 4488 16600
rect 4080 16250 4108 16594
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4068 15972 4120 15978
rect 4068 15914 4120 15920
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 4080 15881 4108 15914
rect 4066 15872 4122 15881
rect 4066 15807 4122 15816
rect 3974 15736 4030 15745
rect 3974 15671 4030 15680
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 3882 14648 3938 14657
rect 3882 14583 3938 14592
rect 3790 14376 3846 14385
rect 3790 14311 3846 14320
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3528 12986 3556 13330
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3606 12608 3662 12617
rect 3606 12543 3662 12552
rect 2964 10746 3016 10752
rect 3160 10764 3280 10792
rect 3344 12158 3464 12186
rect 3516 12164 3568 12170
rect 2976 10538 3004 10746
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2870 9480 2926 9489
rect 2870 9415 2926 9424
rect 2976 8634 3004 9522
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 9178 3096 9318
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 3068 8344 3096 9114
rect 3160 8480 3188 10764
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3252 10266 3280 10610
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3160 8452 3280 8480
rect 3148 8356 3200 8362
rect 3068 8316 3148 8344
rect 3148 8298 3200 8304
rect 2962 8256 3018 8265
rect 2962 8191 3018 8200
rect 2976 8090 3004 8191
rect 2964 8084 3016 8090
rect 2884 8044 2964 8072
rect 2884 7546 2912 8044
rect 2964 8026 3016 8032
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2976 7188 3004 7822
rect 3056 7200 3108 7206
rect 2976 7160 3056 7188
rect 3056 7142 3108 7148
rect 3068 6089 3096 7142
rect 3054 6080 3110 6089
rect 3054 6015 3110 6024
rect 2700 5868 2820 5896
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2516 5273 2544 5510
rect 2502 5264 2558 5273
rect 2502 5199 2558 5208
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2516 5098 2544 5199
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2608 4826 2636 5646
rect 2700 5370 2728 5868
rect 2792 5828 2820 5868
rect 2872 5840 2924 5846
rect 2792 5800 2872 5828
rect 2872 5782 2924 5788
rect 3160 5409 3188 7822
rect 3252 6186 3280 8452
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3344 5778 3372 12158
rect 3516 12106 3568 12112
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11354 3464 12038
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3436 11218 3464 11290
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3528 11150 3556 12106
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3436 9178 3464 9998
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3620 9024 3648 12543
rect 3698 12336 3754 12345
rect 3698 12271 3754 12280
rect 3712 11393 3740 12271
rect 3698 11384 3754 11393
rect 3698 11319 3754 11328
rect 3528 8996 3648 9024
rect 3528 7585 3556 8996
rect 3712 8537 3740 11319
rect 3804 10690 3832 14311
rect 4080 14249 4108 15370
rect 4356 15366 4384 15914
rect 4434 15872 4490 15881
rect 4434 15807 4490 15816
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4252 14272 4304 14278
rect 4066 14240 4122 14249
rect 4252 14214 4304 14220
rect 4066 14175 4122 14184
rect 3974 13968 4030 13977
rect 3974 13903 4030 13912
rect 3988 12322 4016 13903
rect 4080 13818 4108 14175
rect 4264 13954 4292 14214
rect 4356 14074 4384 15302
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4264 13926 4384 13954
rect 4356 13870 4384 13926
rect 4344 13864 4396 13870
rect 4080 13790 4292 13818
rect 4344 13806 4396 13812
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 4172 13433 4200 13670
rect 4158 13424 4214 13433
rect 4158 13359 4214 13368
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4080 12442 4108 13262
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 4172 12850 4200 13194
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4160 12708 4212 12714
rect 4264 12696 4292 13790
rect 4212 12668 4292 12696
rect 4160 12650 4212 12656
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3988 12294 4200 12322
rect 4066 12200 4122 12209
rect 4066 12135 4122 12144
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3896 11257 3924 11562
rect 3976 11280 4028 11286
rect 3882 11248 3938 11257
rect 4080 11257 4108 12135
rect 4172 12050 4200 12294
rect 4356 12209 4384 13806
rect 4448 12782 4476 15807
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4540 12481 4568 25055
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 7102 24440 7158 24449
rect 10289 24432 10585 24452
rect 7102 24375 7158 24384
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6826 21176 6882 21185
rect 6826 21111 6882 21120
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6840 18601 6868 21111
rect 6826 18592 6882 18601
rect 5622 18524 5918 18544
rect 6826 18527 6882 18536
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6366 16824 6422 16833
rect 6366 16759 6422 16768
rect 4896 16720 4948 16726
rect 4896 16662 4948 16668
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4632 15434 4660 15914
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4724 15162 4752 15914
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4724 14550 4752 15098
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4632 14006 4660 14350
rect 4724 14074 4752 14486
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4724 13530 4752 14010
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4620 13456 4672 13462
rect 4620 13398 4672 13404
rect 4632 12986 4660 13398
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4724 12850 4752 13466
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4526 12472 4582 12481
rect 4526 12407 4582 12416
rect 4342 12200 4398 12209
rect 4342 12135 4398 12144
rect 4172 12022 4384 12050
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4264 11286 4292 11494
rect 4252 11280 4304 11286
rect 3976 11222 4028 11228
rect 4066 11248 4122 11257
rect 3882 11183 3938 11192
rect 3988 10810 4016 11222
rect 4066 11183 4122 11192
rect 4172 11240 4252 11268
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3804 10662 3924 10690
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3804 10305 3832 10542
rect 3790 10296 3846 10305
rect 3790 10231 3846 10240
rect 3698 8528 3754 8537
rect 3698 8463 3754 8472
rect 3698 7848 3754 7857
rect 3698 7783 3754 7792
rect 3514 7576 3570 7585
rect 3712 7546 3740 7783
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3514 7511 3570 7520
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 2778 5400 2834 5409
rect 2688 5364 2740 5370
rect 2778 5335 2834 5344
rect 3146 5400 3202 5409
rect 3344 5370 3372 5714
rect 3146 5335 3202 5344
rect 3332 5364 3384 5370
rect 2688 5306 2740 5312
rect 2792 5250 2820 5335
rect 2700 5234 2820 5250
rect 2688 5228 2820 5234
rect 2740 5222 2820 5228
rect 2688 5170 2740 5176
rect 2962 5128 3018 5137
rect 2962 5063 3018 5072
rect 2778 4856 2834 4865
rect 2596 4820 2648 4826
rect 2976 4826 3004 5063
rect 2964 4820 3016 4826
rect 2778 4791 2834 4800
rect 2596 4762 2648 4768
rect 2792 4758 2820 4791
rect 2884 4780 2964 4808
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2596 4004 2648 4010
rect 2596 3946 2648 3952
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2136 2576 2188 2582
rect 2134 2544 2136 2553
rect 2188 2544 2190 2553
rect 2134 2479 2190 2488
rect 2240 1465 2268 3878
rect 2502 3768 2558 3777
rect 2502 3703 2558 3712
rect 2516 3466 2544 3703
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2504 2304 2556 2310
rect 2502 2272 2504 2281
rect 2556 2272 2558 2281
rect 2502 2207 2558 2216
rect 2226 1456 2282 1465
rect 2226 1391 2282 1400
rect 2608 480 2636 3946
rect 2700 3738 2728 4626
rect 2792 4214 2820 4694
rect 2884 4282 2912 4780
rect 2964 4762 3016 4768
rect 3054 4720 3110 4729
rect 3054 4655 3110 4664
rect 3068 4554 3096 4655
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 3068 3738 3096 4490
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3068 3097 3096 3470
rect 3054 3088 3110 3097
rect 3054 3023 3110 3032
rect 3068 2854 3096 3023
rect 3160 2922 3188 5335
rect 3332 5306 3384 5312
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3344 3738 3372 3946
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3344 3534 3372 3674
rect 3332 3528 3384 3534
rect 3436 3505 3464 6598
rect 3528 6458 3556 7346
rect 3804 7274 3832 7686
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3528 5710 3556 6394
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3528 4078 3556 5646
rect 3620 4078 3648 7210
rect 3790 6488 3846 6497
rect 3790 6423 3846 6432
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3712 5137 3740 5238
rect 3698 5128 3754 5137
rect 3698 5063 3754 5072
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3528 3738 3556 4014
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3712 3670 3740 5063
rect 3804 4185 3832 6423
rect 3896 5001 3924 10662
rect 3974 7168 4030 7177
rect 3974 7103 4030 7112
rect 3988 5545 4016 7103
rect 4080 5778 4108 11183
rect 4172 9586 4200 11240
rect 4252 11222 4304 11228
rect 4250 10704 4306 10713
rect 4250 10639 4306 10648
rect 4264 10606 4292 10639
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4172 7290 4200 9522
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4264 7410 4292 7686
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4172 7262 4292 7290
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 6866 4200 7142
rect 4264 6866 4292 7262
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4172 5953 4200 6802
rect 4264 6458 4292 6802
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4158 5944 4214 5953
rect 4158 5879 4214 5888
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4068 5568 4120 5574
rect 3974 5536 4030 5545
rect 4068 5510 4120 5516
rect 3974 5471 4030 5480
rect 4080 5098 4108 5510
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3882 4992 3938 5001
rect 3882 4927 3938 4936
rect 3790 4176 3846 4185
rect 3790 4111 3846 4120
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3884 3528 3936 3534
rect 3332 3470 3384 3476
rect 3422 3496 3478 3505
rect 3344 2990 3372 3470
rect 3988 3505 4016 5034
rect 4080 4758 4108 5034
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 4172 4690 4200 4966
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4264 4128 4292 6394
rect 4080 4100 4292 4128
rect 4080 4010 4108 4100
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3884 3470 3936 3476
rect 3974 3496 4030 3505
rect 3422 3431 3478 3440
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3148 2916 3200 2922
rect 3148 2858 3200 2864
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 3068 2582 3096 2790
rect 3896 2650 3924 3470
rect 3974 3431 4030 3440
rect 4080 3194 4108 3538
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4066 2680 4122 2689
rect 3884 2644 3936 2650
rect 4066 2615 4122 2624
rect 3884 2586 3936 2592
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 2976 1737 3004 2518
rect 3698 2136 3754 2145
rect 3698 2071 3754 2080
rect 2962 1728 3018 1737
rect 2962 1663 3018 1672
rect 3712 610 3740 2071
rect 4080 2009 4108 2615
rect 4264 2582 4292 2790
rect 4252 2576 4304 2582
rect 4252 2518 4304 2524
rect 4066 2000 4122 2009
rect 4066 1935 4122 1944
rect 3148 604 3200 610
rect 3148 546 3200 552
rect 3700 604 3752 610
rect 3700 546 3752 552
rect 3792 604 3844 610
rect 3792 546 3844 552
rect 3160 480 3188 546
rect 3804 480 3832 546
rect 4356 480 4384 12022
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4448 8090 4476 10406
rect 4540 10266 4568 12407
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4540 9722 4568 10202
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4526 9480 4582 9489
rect 4526 9415 4528 9424
rect 4580 9415 4582 9424
rect 4528 9386 4580 9392
rect 4540 9178 4568 9386
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4448 7478 4476 8026
rect 4540 8022 4568 9114
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4540 7478 4568 7958
rect 4632 7886 4660 12718
rect 4816 12714 4844 16118
rect 4908 15910 4936 16662
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5276 15910 5304 16526
rect 5460 16425 6040 16436
rect 5446 16416 6054 16425
rect 5502 16408 5998 16416
rect 5446 16351 5502 16360
rect 5622 16348 5918 16368
rect 5998 16351 6054 16360
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 4908 15638 4936 15846
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 4896 15496 4948 15502
rect 5080 15496 5132 15502
rect 4948 15456 5028 15484
rect 4896 15438 4948 15444
rect 4894 15328 4950 15337
rect 4894 15263 4950 15272
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4724 11694 4752 12174
rect 4816 11801 4844 12310
rect 4908 12238 4936 15263
rect 5000 14822 5028 15456
rect 5276 15473 5304 15846
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5460 15473 5488 15574
rect 5540 15496 5592 15502
rect 5080 15438 5132 15444
rect 5262 15464 5318 15473
rect 4988 14816 5040 14822
rect 4986 14784 4988 14793
rect 5040 14784 5042 14793
rect 4986 14719 5042 14728
rect 5000 14521 5028 14719
rect 5092 14618 5120 15438
rect 5262 15399 5318 15408
rect 5446 15464 5502 15473
rect 5540 15438 5592 15444
rect 5446 15399 5502 15408
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 4986 14512 5042 14521
rect 4986 14447 5042 14456
rect 5092 13938 5120 14554
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 5000 12889 5028 13670
rect 5092 13530 5120 13874
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5092 13326 5120 13466
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5276 12986 5304 14894
rect 5368 13258 5396 15302
rect 5460 15162 5488 15399
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5446 14784 5502 14793
rect 5446 14719 5502 14728
rect 5460 13530 5488 14719
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5552 13410 5580 15438
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 14385 6040 15302
rect 5998 14376 6054 14385
rect 5998 14311 6054 14320
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5722 13560 5778 13569
rect 5722 13495 5778 13504
rect 5460 13394 5580 13410
rect 5448 13388 5580 13394
rect 5500 13382 5580 13388
rect 5448 13330 5500 13336
rect 5736 13258 5764 13495
rect 6012 13462 6040 14311
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5998 13016 6054 13025
rect 5264 12980 5316 12986
rect 5998 12951 6054 12960
rect 5264 12922 5316 12928
rect 4986 12880 5042 12889
rect 4986 12815 5042 12824
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 5000 11898 5028 12242
rect 5736 12209 5764 12786
rect 6012 12714 6040 12951
rect 6104 12782 6132 14214
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6196 12714 6224 13262
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5722 12200 5778 12209
rect 5540 12164 5592 12170
rect 5722 12135 5778 12144
rect 5540 12106 5592 12112
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4802 11792 4858 11801
rect 5000 11762 5028 11834
rect 4802 11727 4858 11736
rect 4988 11756 5040 11762
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4724 11286 4752 11630
rect 4816 11626 4844 11727
rect 4988 11698 5040 11704
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5368 11354 5396 11494
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 4724 10674 4752 11222
rect 4988 11144 5040 11150
rect 4802 11112 4858 11121
rect 4988 11086 5040 11092
rect 4802 11047 4858 11056
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4816 10198 4844 11047
rect 5000 10810 5028 11086
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4710 10024 4766 10033
rect 4710 9959 4712 9968
rect 4764 9959 4766 9968
rect 4712 9930 4764 9936
rect 4816 9178 4844 10134
rect 5184 10130 5212 10678
rect 5172 10124 5224 10130
rect 5276 10112 5304 10746
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5368 10305 5396 10542
rect 5460 10441 5488 11222
rect 5552 10810 5580 12106
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5828 11393 5856 11562
rect 5908 11552 5960 11558
rect 5906 11520 5908 11529
rect 5960 11520 5962 11529
rect 5906 11455 5962 11464
rect 5814 11384 5870 11393
rect 5814 11319 5870 11328
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5446 10432 5502 10441
rect 5446 10367 5502 10376
rect 5354 10296 5410 10305
rect 5460 10266 5488 10367
rect 5354 10231 5410 10240
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5448 10124 5500 10130
rect 5276 10084 5448 10112
rect 5172 10066 5224 10072
rect 5448 10066 5500 10072
rect 5356 9920 5408 9926
rect 5262 9888 5318 9897
rect 5356 9862 5408 9868
rect 5262 9823 5318 9832
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5170 9344 5226 9353
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4908 8566 4936 9046
rect 5000 9042 5028 9318
rect 5170 9279 5226 9288
rect 5078 9208 5134 9217
rect 5078 9143 5134 9152
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5000 8634 5028 8978
rect 5092 8974 5120 9143
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4632 7546 4660 7822
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4724 6934 4752 8230
rect 4908 7818 4936 8502
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4434 6080 4490 6089
rect 4434 6015 4490 6024
rect 4448 4758 4476 6015
rect 4724 5914 4752 6870
rect 5184 6474 5212 9279
rect 5276 8945 5304 9823
rect 5262 8936 5318 8945
rect 5368 8906 5396 9862
rect 5460 9722 5488 10066
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5262 8871 5318 8880
rect 5356 8900 5408 8906
rect 5276 8294 5304 8871
rect 5356 8842 5408 8848
rect 5460 8786 5488 9658
rect 5552 9178 5580 10134
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5644 8820 5672 9114
rect 5368 8758 5488 8786
rect 5552 8792 5672 8820
rect 5368 8498 5396 8758
rect 5446 8664 5502 8673
rect 5446 8599 5502 8608
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5460 8430 5488 8599
rect 5448 8424 5500 8430
rect 5354 8392 5410 8401
rect 5448 8366 5500 8372
rect 5354 8327 5410 8336
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5368 8090 5396 8327
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5552 7562 5580 8792
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5644 7954 5672 8434
rect 5722 8392 5778 8401
rect 5722 8327 5724 8336
rect 5776 8327 5778 8336
rect 5724 8298 5776 8304
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5920 7834 5948 8434
rect 6012 7993 6040 12242
rect 5998 7984 6054 7993
rect 5998 7919 6054 7928
rect 5920 7806 6040 7834
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5460 7546 5580 7562
rect 5448 7540 5580 7546
rect 5500 7534 5580 7540
rect 5448 7482 5500 7488
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5000 6446 5212 6474
rect 5000 5914 5028 6446
rect 5262 6352 5318 6361
rect 5080 6316 5132 6322
rect 5262 6287 5318 6296
rect 5080 6258 5132 6264
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4540 678 4568 5714
rect 4618 5672 4674 5681
rect 4618 5607 4674 5616
rect 4632 4826 4660 5607
rect 5000 5370 5028 5850
rect 5092 5846 5120 6258
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 4988 5364 5040 5370
rect 4908 5324 4988 5352
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4632 3777 4660 4762
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4618 3768 4674 3777
rect 4618 3703 4674 3712
rect 4816 2281 4844 4694
rect 4802 2272 4858 2281
rect 4802 2207 4858 2216
rect 4528 672 4580 678
rect 4528 614 4580 620
rect 4908 480 4936 5324
rect 4988 5306 5040 5312
rect 4986 4856 5042 4865
rect 4986 4791 5042 4800
rect 5000 4622 5028 4791
rect 5092 4758 5120 5646
rect 5184 5409 5212 5850
rect 5170 5400 5226 5409
rect 5170 5335 5226 5344
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5000 4282 5028 4558
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 5184 3942 5212 5335
rect 5276 4554 5304 6287
rect 5368 5642 5396 7210
rect 5460 6458 5488 7346
rect 5538 7304 5594 7313
rect 5538 7239 5594 7248
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5552 5166 5580 7239
rect 5630 6896 5686 6905
rect 5630 6831 5686 6840
rect 5644 6730 5672 6831
rect 6012 6730 6040 7806
rect 6104 7274 6132 12378
rect 6184 12368 6236 12374
rect 6182 12336 6184 12345
rect 6236 12336 6238 12345
rect 6182 12271 6238 12280
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6196 8498 6224 12174
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6092 7268 6144 7274
rect 6092 7210 6144 7216
rect 6196 7018 6224 7958
rect 6288 7410 6316 15370
rect 6380 10674 6408 16759
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6472 12442 6500 15302
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6564 12322 6592 15846
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6656 14074 6684 14758
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6748 13977 6776 14826
rect 6734 13968 6790 13977
rect 6644 13932 6696 13938
rect 6734 13903 6790 13912
rect 6644 13874 6696 13880
rect 6656 13530 6684 13874
rect 6734 13832 6790 13841
rect 6734 13767 6790 13776
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6656 12442 6684 13466
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6472 12294 6592 12322
rect 6642 12336 6698 12345
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6472 10282 6500 12294
rect 6642 12271 6698 12280
rect 6656 12186 6684 12271
rect 6380 10254 6500 10282
rect 6564 12158 6684 12186
rect 6380 9178 6408 10254
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6472 9722 6500 10134
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6472 8634 6500 8910
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6380 7546 6408 7890
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6274 7032 6330 7041
rect 6196 6990 6274 7018
rect 6274 6967 6276 6976
rect 6328 6967 6330 6976
rect 6276 6938 6328 6944
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5998 6488 6054 6497
rect 6288 6458 6316 6938
rect 5998 6423 6054 6432
rect 6276 6452 6328 6458
rect 5722 6216 5778 6225
rect 5722 6151 5724 6160
rect 5776 6151 5778 6160
rect 5724 6122 5776 6128
rect 6012 6118 6040 6423
rect 6276 6394 6328 6400
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6182 5944 6238 5953
rect 6380 5914 6408 7142
rect 6472 6225 6500 8434
rect 6458 6216 6514 6225
rect 6458 6151 6514 6160
rect 6458 5944 6514 5953
rect 6182 5879 6238 5888
rect 6368 5908 6420 5914
rect 6090 5808 6146 5817
rect 6090 5743 6146 5752
rect 6104 5642 6132 5743
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6090 5536 6146 5545
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5184 3738 5212 3878
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5276 1873 5304 3130
rect 5368 2689 5396 5034
rect 5552 4826 5580 5102
rect 6012 5098 6040 5510
rect 6090 5471 6146 5480
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5448 4684 5500 4690
rect 5500 4644 5580 4672
rect 5448 4626 5500 4632
rect 5446 4176 5502 4185
rect 5446 4111 5502 4120
rect 5460 4078 5488 4111
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5354 2680 5410 2689
rect 5354 2615 5410 2624
rect 5552 2292 5580 4644
rect 5736 4593 5764 4966
rect 6104 4758 6132 5471
rect 6196 4826 6224 5879
rect 6564 5914 6592 12158
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6656 11665 6684 12038
rect 6642 11656 6698 11665
rect 6642 11591 6698 11600
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6656 10033 6684 11494
rect 6642 10024 6698 10033
rect 6642 9959 6698 9968
rect 6656 9110 6684 9959
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6748 8906 6776 13767
rect 6840 11558 6868 15846
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6932 14278 6960 14826
rect 7024 14550 7052 15438
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 12186 6960 13670
rect 7024 13530 7052 14486
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7012 12640 7064 12646
rect 7010 12608 7012 12617
rect 7064 12608 7066 12617
rect 7010 12543 7066 12552
rect 7116 12374 7144 24375
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 7562 18320 7618 18329
rect 7562 18255 7618 18264
rect 7470 16552 7526 16561
rect 7470 16487 7526 16496
rect 7378 16008 7434 16017
rect 7378 15943 7434 15952
rect 7194 14648 7250 14657
rect 7194 14583 7196 14592
rect 7248 14583 7250 14592
rect 7196 14554 7248 14560
rect 7208 14074 7236 14554
rect 7286 14376 7342 14385
rect 7286 14311 7288 14320
rect 7340 14311 7342 14320
rect 7288 14282 7340 14288
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7104 12368 7156 12374
rect 7104 12310 7156 12316
rect 6932 12158 7144 12186
rect 7208 12170 7236 13398
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6840 10810 6868 11290
rect 6918 11112 6974 11121
rect 6918 11047 6974 11056
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6642 8800 6698 8809
rect 6642 8735 6698 8744
rect 6656 8498 6684 8735
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6748 8430 6776 8842
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6840 8090 6868 9658
rect 6932 9217 6960 11047
rect 6918 9208 6974 9217
rect 6918 9143 6920 9152
rect 6972 9143 6974 9152
rect 6920 9114 6972 9120
rect 6932 9083 6960 9114
rect 6918 8528 6974 8537
rect 6918 8463 6974 8472
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6840 7342 6868 8026
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6656 7002 6684 7278
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6458 5879 6514 5888
rect 6552 5908 6604 5914
rect 6368 5850 6420 5856
rect 6472 5710 6500 5879
rect 6840 5896 6868 7142
rect 6932 6866 6960 8463
rect 7024 8022 7052 12038
rect 7116 9178 7144 12158
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7300 10656 7328 12310
rect 7392 12238 7420 15943
rect 7484 13734 7512 16487
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7576 13546 7604 18255
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10322 17776 10378 17785
rect 10322 17711 10378 17720
rect 9862 17640 9918 17649
rect 9862 17575 9918 17584
rect 9678 15736 9734 15745
rect 9678 15671 9734 15680
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7852 14550 7880 14758
rect 7840 14544 7892 14550
rect 7840 14486 7892 14492
rect 7852 13870 7880 14486
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7484 13518 7604 13546
rect 7484 13433 7512 13518
rect 7470 13424 7526 13433
rect 7470 13359 7526 13368
rect 7564 13388 7616 13394
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7392 11286 7420 11698
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7378 10840 7434 10849
rect 7378 10775 7434 10784
rect 7208 10628 7328 10656
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 7116 7177 7144 8298
rect 7102 7168 7158 7177
rect 7102 7103 7158 7112
rect 7208 6866 7236 10628
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7300 10169 7328 10474
rect 7392 10470 7420 10775
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7286 10160 7342 10169
rect 7286 10095 7342 10104
rect 7484 10010 7512 13359
rect 7564 13330 7616 13336
rect 7576 11898 7604 13330
rect 7668 12850 7696 13738
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7852 13410 7880 13670
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7668 11937 7696 12310
rect 7654 11928 7710 11937
rect 7564 11892 7616 11898
rect 7654 11863 7710 11872
rect 7564 11834 7616 11840
rect 7668 11626 7696 11863
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7760 11082 7788 13398
rect 7852 13394 7972 13410
rect 7840 13388 7972 13394
rect 7892 13382 7972 13388
rect 7840 13330 7892 13336
rect 7838 13288 7894 13297
rect 7838 13223 7894 13232
rect 7852 12986 7880 13223
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7944 12714 7972 13382
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7838 11792 7894 11801
rect 7944 11762 7972 12310
rect 8022 12064 8078 12073
rect 8022 11999 8078 12008
rect 8036 11830 8064 11999
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 7838 11727 7894 11736
rect 7932 11756 7984 11762
rect 7852 11626 7880 11727
rect 7932 11698 7984 11704
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 7944 11354 7972 11698
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 8022 11248 8078 11257
rect 7932 11212 7984 11218
rect 8022 11183 8078 11192
rect 7932 11154 7984 11160
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7944 10742 7972 11154
rect 8036 11150 8064 11183
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 8036 10810 8064 11086
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7932 10736 7984 10742
rect 8036 10713 8064 10746
rect 7932 10678 7984 10684
rect 8022 10704 8078 10713
rect 8022 10639 8078 10648
rect 8128 10606 8156 11766
rect 8220 11370 8248 13194
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 13025 8340 13126
rect 8298 13016 8354 13025
rect 8298 12951 8354 12960
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8312 12442 8340 12650
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8404 12322 8432 14214
rect 8312 12294 8432 12322
rect 8312 11506 8340 12294
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11694 8432 12174
rect 8392 11688 8444 11694
rect 8390 11656 8392 11665
rect 8444 11656 8446 11665
rect 8390 11591 8446 11600
rect 8312 11478 8432 11506
rect 8220 11354 8340 11370
rect 8220 11348 8352 11354
rect 8220 11342 8300 11348
rect 8300 11290 8352 11296
rect 8208 10736 8260 10742
rect 8206 10704 8208 10713
rect 8260 10704 8262 10713
rect 8206 10639 8262 10648
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8128 10266 8156 10542
rect 8312 10266 8340 10542
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8404 10010 8432 11478
rect 7392 9982 7512 10010
rect 7944 9982 8432 10010
rect 7286 7440 7342 7449
rect 7286 7375 7342 7384
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 6920 5908 6972 5914
rect 6840 5868 6920 5896
rect 6552 5850 6604 5856
rect 6920 5850 6972 5856
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6472 5302 6500 5646
rect 6564 5370 6592 5850
rect 7208 5522 7236 6802
rect 7116 5494 7236 5522
rect 7010 5400 7066 5409
rect 6552 5364 6604 5370
rect 7116 5370 7144 5494
rect 7010 5335 7066 5344
rect 7104 5364 7156 5370
rect 6552 5306 6604 5312
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 5722 4584 5778 4593
rect 5722 4519 5778 4528
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6196 4282 6224 4762
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6090 4040 6146 4049
rect 6090 3975 6146 3984
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5722 3088 5778 3097
rect 5722 3023 5778 3032
rect 5736 2922 5764 3023
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 6012 2650 6040 3606
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5552 2281 6040 2292
rect 5552 2272 6054 2281
rect 5552 2264 5998 2272
rect 5622 2204 5918 2224
rect 5998 2207 6054 2216
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5998 2136 6054 2145
rect 5998 2071 6054 2080
rect 5262 1864 5318 1873
rect 5262 1799 5318 1808
rect 6012 1601 6040 2071
rect 5998 1592 6054 1601
rect 5998 1527 6054 1536
rect 5540 1420 5592 1426
rect 5540 1362 5592 1368
rect 5552 480 5580 1362
rect 6104 480 6132 3975
rect 6196 1426 6224 4218
rect 6472 4214 6500 4558
rect 6656 4282 6684 4626
rect 6748 4486 6776 5034
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6288 3369 6316 3538
rect 6274 3360 6330 3369
rect 6274 3295 6330 3304
rect 6380 1601 6408 3946
rect 6472 3777 6500 4150
rect 6458 3768 6514 3777
rect 6656 3738 6684 4218
rect 6748 3913 6776 4422
rect 6734 3904 6790 3913
rect 6734 3839 6790 3848
rect 6458 3703 6514 3712
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6748 3670 6776 3839
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 3194 6500 3334
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6472 2990 6500 3130
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6920 2984 6972 2990
rect 7024 2972 7052 5335
rect 7104 5306 7156 5312
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7208 4214 7236 5170
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7116 2990 7144 3402
rect 6972 2944 7052 2972
rect 6920 2926 6972 2932
rect 6642 2544 6698 2553
rect 6642 2479 6644 2488
rect 6696 2479 6698 2488
rect 6644 2450 6696 2456
rect 7024 2378 7052 2944
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7208 2650 7236 4150
rect 7300 4010 7328 7375
rect 7392 4146 7420 9982
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9450 7512 9862
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7484 8974 7512 9386
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7838 8800 7894 8809
rect 7838 8735 7894 8744
rect 7654 8120 7710 8129
rect 7654 8055 7656 8064
rect 7708 8055 7710 8064
rect 7656 8026 7708 8032
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7470 6760 7526 6769
rect 7470 6695 7472 6704
rect 7524 6695 7526 6704
rect 7472 6666 7524 6672
rect 7576 6390 7604 7346
rect 7852 6798 7880 8735
rect 7944 7002 7972 9982
rect 8300 9920 8352 9926
rect 8114 9888 8170 9897
rect 8300 9862 8352 9868
rect 8114 9823 8170 9832
rect 8128 8906 8156 9823
rect 8206 9752 8262 9761
rect 8206 9687 8262 9696
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8220 8634 8248 9687
rect 8312 9518 8340 9862
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8496 9110 8524 15438
rect 9692 15162 9720 15671
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9692 14890 9720 15098
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9770 14784 9826 14793
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8588 13841 8616 14214
rect 8574 13832 8630 13841
rect 8574 13767 8630 13776
rect 8574 13424 8630 13433
rect 8574 13359 8630 13368
rect 8588 13025 8616 13359
rect 8574 13016 8630 13025
rect 8574 12951 8630 12960
rect 8574 12200 8630 12209
rect 8574 12135 8576 12144
rect 8628 12135 8630 12144
rect 8576 12106 8628 12112
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8680 11898 8708 12038
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8588 10606 8616 10950
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8588 9722 8616 10542
rect 8956 10266 8984 14214
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8666 10024 8722 10033
rect 8666 9959 8668 9968
rect 8720 9959 8722 9968
rect 8668 9930 8720 9936
rect 9140 9897 9168 14758
rect 9770 14719 9826 14728
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9126 9888 9182 9897
rect 9126 9823 9182 9832
rect 9232 9761 9260 14214
rect 9784 13841 9812 14719
rect 9770 13832 9826 13841
rect 9770 13767 9826 13776
rect 9310 13560 9366 13569
rect 9310 13495 9366 13504
rect 9324 12442 9352 13495
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9416 12986 9444 13330
rect 9680 13320 9732 13326
rect 9732 13280 9812 13308
rect 9680 13262 9732 13268
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9324 11762 9352 12378
rect 9416 12186 9444 12922
rect 9586 12880 9642 12889
rect 9586 12815 9642 12824
rect 9600 12481 9628 12815
rect 9586 12472 9642 12481
rect 9586 12407 9642 12416
rect 9692 12306 9720 13126
rect 9784 12714 9812 13280
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9876 12374 9904 17575
rect 10336 17105 10364 17711
rect 11058 17232 11114 17241
rect 11058 17167 11114 17176
rect 10046 17096 10102 17105
rect 10046 17031 10102 17040
rect 10322 17096 10378 17105
rect 10322 17031 10378 17040
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9968 15162 9996 15914
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9416 12158 9536 12186
rect 9508 12102 9536 12158
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11762 9536 12038
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 11354 9444 11494
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9324 9926 9352 11222
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9770 11112 9826 11121
rect 9770 11047 9772 11056
rect 9824 11047 9826 11056
rect 9772 11018 9824 11024
rect 9876 10470 9904 11154
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9680 10464 9732 10470
rect 9678 10432 9680 10441
rect 9864 10464 9916 10470
rect 9732 10432 9734 10441
rect 9864 10406 9916 10412
rect 9678 10367 9734 10376
rect 9494 10296 9550 10305
rect 9494 10231 9550 10240
rect 9508 9994 9536 10231
rect 9692 10130 9720 10367
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9218 9752 9274 9761
rect 8576 9716 8628 9722
rect 9218 9687 9274 9696
rect 8576 9658 8628 9664
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8208 8084 8260 8090
rect 8312 8072 8340 9046
rect 8588 8974 8616 9658
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8404 8362 8432 8842
rect 8588 8498 8616 8910
rect 8956 8634 8984 9454
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9036 9104 9088 9110
rect 9034 9072 9036 9081
rect 9088 9072 9090 9081
rect 9034 9007 9090 9016
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8260 8044 8340 8072
rect 8208 8026 8260 8032
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8114 7576 8170 7585
rect 8114 7511 8170 7520
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7576 5166 7604 6326
rect 7852 5642 7880 6734
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7944 4978 7972 6938
rect 8036 6798 8064 7210
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8036 6458 8064 6734
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8128 5930 8156 7511
rect 8220 6361 8248 7890
rect 8404 7721 8432 8298
rect 8588 8090 8616 8434
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8482 7984 8538 7993
rect 8482 7919 8484 7928
rect 8536 7919 8538 7928
rect 8484 7890 8536 7896
rect 8390 7712 8446 7721
rect 8390 7647 8446 7656
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8206 6352 8262 6361
rect 8206 6287 8262 6296
rect 8404 6254 8432 6598
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 7852 4950 7972 4978
rect 8036 5902 8156 5930
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7760 4457 7788 4558
rect 7852 4486 7880 4950
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7944 4554 7972 4762
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7840 4480 7892 4486
rect 7746 4448 7802 4457
rect 7840 4422 7892 4428
rect 7746 4383 7802 4392
rect 7760 4282 7788 4383
rect 7944 4321 7972 4490
rect 7930 4312 7986 4321
rect 7748 4276 7800 4282
rect 7930 4247 7986 4256
rect 7748 4218 7800 4224
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7300 3738 7328 3946
rect 8036 3754 8064 5902
rect 8404 5846 8432 6190
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8482 5808 8538 5817
rect 8128 5370 8156 5782
rect 8404 5370 8432 5782
rect 8482 5743 8538 5752
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8128 4690 8156 5034
rect 8220 4826 8248 5102
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8128 4457 8156 4626
rect 8220 4622 8248 4762
rect 8404 4758 8432 5306
rect 8496 5001 8524 5743
rect 8574 5672 8630 5681
rect 8574 5607 8576 5616
rect 8628 5607 8630 5616
rect 8576 5578 8628 5584
rect 8482 4992 8538 5001
rect 8482 4927 8538 4936
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8114 4448 8170 4457
rect 8114 4383 8170 4392
rect 8128 4146 8156 4383
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7852 3726 8064 3754
rect 7286 3632 7342 3641
rect 7286 3567 7342 3576
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 6642 2272 6698 2281
rect 6642 2207 6698 2216
rect 6366 1592 6422 1601
rect 6366 1527 6422 1536
rect 6184 1420 6236 1426
rect 6184 1362 6236 1368
rect 6656 480 6684 2207
rect 7300 480 7328 3567
rect 7576 921 7604 3674
rect 7562 912 7618 921
rect 7562 847 7618 856
rect 7852 480 7880 3726
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7944 2650 7972 3402
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8128 3097 8156 3334
rect 8220 3210 8248 4558
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 3913 8340 4422
rect 8404 4282 8432 4694
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8298 3904 8354 3913
rect 8298 3839 8354 3848
rect 8496 3738 8524 4927
rect 8576 4752 8628 4758
rect 8574 4720 8576 4729
rect 8628 4720 8630 4729
rect 8574 4655 8630 4664
rect 8574 4312 8630 4321
rect 8574 4247 8630 4256
rect 8588 4214 8616 4247
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8680 3618 8708 8298
rect 9232 8265 9260 9318
rect 9324 8362 9352 9862
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9218 8256 9274 8265
rect 9218 8191 9274 8200
rect 8850 8120 8906 8129
rect 8850 8055 8906 8064
rect 8864 6730 8892 8055
rect 9416 7857 9444 8774
rect 9402 7848 9458 7857
rect 9402 7783 9458 7792
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 6361 8800 6598
rect 8758 6352 8814 6361
rect 8758 6287 8814 6296
rect 8942 6080 8998 6089
rect 8942 6015 8998 6024
rect 8956 5914 8984 6015
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9048 5545 9076 7686
rect 9508 7546 9536 9930
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9692 8945 9720 9386
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9678 8936 9734 8945
rect 9678 8871 9734 8880
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 8430 9720 8774
rect 9784 8537 9812 9318
rect 9770 8528 9826 8537
rect 9770 8463 9826 8472
rect 9680 8424 9732 8430
rect 9678 8392 9680 8401
rect 9732 8392 9734 8401
rect 9588 8356 9640 8362
rect 9678 8327 9734 8336
rect 9588 8298 9640 8304
rect 9600 8242 9628 8298
rect 9876 8294 9904 10406
rect 9968 9489 9996 11086
rect 9954 9480 10010 9489
rect 9954 9415 10010 9424
rect 9954 8936 10010 8945
rect 9954 8871 10010 8880
rect 9968 8673 9996 8871
rect 9954 8664 10010 8673
rect 9954 8599 10010 8608
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9680 8288 9732 8294
rect 9600 8236 9680 8242
rect 9600 8230 9732 8236
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9600 8214 9720 8230
rect 9770 8120 9826 8129
rect 9770 8055 9826 8064
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9784 7410 9812 8055
rect 9864 7744 9916 7750
rect 9862 7712 9864 7721
rect 9916 7712 9918 7721
rect 9862 7647 9918 7656
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9126 7304 9182 7313
rect 9126 7239 9182 7248
rect 9034 5536 9090 5545
rect 9034 5471 9090 5480
rect 8404 3590 8708 3618
rect 8220 3194 8340 3210
rect 8220 3188 8352 3194
rect 8220 3182 8300 3188
rect 8300 3130 8352 3136
rect 8114 3088 8170 3097
rect 8114 3023 8170 3032
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8404 480 8432 3590
rect 8482 3360 8538 3369
rect 8482 3295 8538 3304
rect 8496 2514 8524 3295
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8680 2009 8708 2246
rect 8666 2000 8722 2009
rect 8666 1935 8722 1944
rect 9048 480 9076 5471
rect 9140 4282 9168 7239
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9678 7168 9734 7177
rect 9232 7041 9260 7142
rect 9678 7103 9734 7112
rect 9218 7032 9274 7041
rect 9218 6967 9274 6976
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9140 3602 9168 4218
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9324 2825 9352 6598
rect 9692 6338 9720 7103
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9600 6310 9720 6338
rect 9600 5794 9628 6310
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9692 5914 9720 6122
rect 9784 6118 9812 6190
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9600 5766 9720 5794
rect 9494 5672 9550 5681
rect 9494 5607 9496 5616
rect 9548 5607 9550 5616
rect 9496 5578 9548 5584
rect 9402 5128 9458 5137
rect 9402 5063 9458 5072
rect 9416 4826 9444 5063
rect 9404 4820 9456 4826
rect 9692 4808 9720 5766
rect 9784 5370 9812 6054
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9692 4780 9812 4808
rect 9404 4762 9456 4768
rect 9784 4729 9812 4780
rect 9770 4720 9826 4729
rect 9680 4684 9732 4690
rect 9770 4655 9826 4664
rect 9680 4626 9732 4632
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9600 4146 9628 4422
rect 9692 4214 9720 4626
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9586 4040 9642 4049
rect 9496 4004 9548 4010
rect 9586 3975 9588 3984
rect 9496 3946 9548 3952
rect 9640 3975 9642 3984
rect 9588 3946 9640 3952
rect 9508 3466 9536 3946
rect 9586 3768 9642 3777
rect 9692 3738 9720 4150
rect 9586 3703 9642 3712
rect 9680 3732 9732 3738
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 2990 9444 3334
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9310 2816 9366 2825
rect 9310 2751 9366 2760
rect 9126 2680 9182 2689
rect 9416 2650 9444 2926
rect 9126 2615 9128 2624
rect 9180 2615 9182 2624
rect 9404 2644 9456 2650
rect 9128 2586 9180 2592
rect 9404 2586 9456 2592
rect 9140 2446 9168 2586
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9126 2272 9182 2281
rect 9126 2207 9182 2216
rect 9140 1873 9168 2207
rect 9126 1864 9182 1873
rect 9126 1799 9182 1808
rect 9600 480 9628 3703
rect 9680 3674 9732 3680
rect 9876 2145 9904 6598
rect 9862 2136 9918 2145
rect 9862 2071 9918 2080
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 2042 0 2098 480
rect 2594 0 2650 480
rect 3146 0 3202 480
rect 3790 0 3846 480
rect 4342 0 4398 480
rect 4894 0 4950 480
rect 5538 0 5594 480
rect 6090 0 6146 480
rect 6642 0 6698 480
rect 7286 0 7342 480
rect 7838 0 7894 480
rect 8390 0 8446 480
rect 9034 0 9090 480
rect 9586 0 9642 480
rect 9968 377 9996 8502
rect 10060 4146 10088 17031
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10152 14958 10180 16594
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10600 15632 10652 15638
rect 10600 15574 10652 15580
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10152 14618 10180 14894
rect 10520 14890 10548 15438
rect 10612 15026 10640 15574
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14618 10732 15982
rect 10980 15978 11008 16390
rect 10968 15972 11020 15978
rect 10968 15914 11020 15920
rect 10782 15192 10838 15201
rect 10782 15127 10838 15136
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10796 14074 10824 15127
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10888 14113 10916 14418
rect 10980 14346 11008 15914
rect 11072 14929 11100 17167
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11058 14920 11114 14929
rect 11058 14855 11114 14864
rect 11072 14550 11100 14855
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10874 14104 10930 14113
rect 10784 14068 10836 14074
rect 10874 14039 10930 14048
rect 10784 14010 10836 14016
rect 10784 13728 10836 13734
rect 10888 13716 10916 14039
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10836 13688 10916 13716
rect 10784 13670 10836 13676
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10690 12744 10746 12753
rect 10690 12679 10746 12688
rect 10704 12646 10732 12679
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10152 11393 10180 12106
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10138 11384 10194 11393
rect 10289 11376 10585 11396
rect 10138 11319 10194 11328
rect 10152 11121 10180 11319
rect 10796 11286 10824 13670
rect 10980 12986 11008 13874
rect 11072 13802 11100 14486
rect 11164 14414 11192 14962
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11164 14006 11192 14350
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 11164 13530 11192 13942
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 11164 12850 11192 13466
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 11898 10916 12242
rect 10980 12238 11008 12650
rect 11072 12374 11100 12650
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 11256 12306 11284 26250
rect 14278 23760 14334 23769
rect 14278 23695 14334 23704
rect 14292 21978 14320 23695
rect 14292 21950 14412 21978
rect 13358 18864 13414 18873
rect 14384 18850 14412 21950
rect 13358 18799 13414 18808
rect 14108 18822 14412 18850
rect 12530 18592 12586 18601
rect 12530 18527 12586 18536
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11808 15162 11836 16118
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11900 15706 11928 15982
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11796 15156 11848 15162
rect 11848 15116 11928 15144
rect 11796 15098 11848 15104
rect 11794 15056 11850 15065
rect 11794 14991 11850 15000
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11348 14006 11376 14554
rect 11808 14550 11836 14991
rect 11900 14822 11928 15116
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11336 14000 11388 14006
rect 11336 13942 11388 13948
rect 11348 13802 11376 13942
rect 11624 13938 11652 14214
rect 11808 14074 11836 14486
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11336 12640 11388 12646
rect 11334 12608 11336 12617
rect 11704 12640 11756 12646
rect 11388 12608 11390 12617
rect 11704 12582 11756 12588
rect 11334 12543 11390 12552
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10138 11112 10194 11121
rect 10138 11047 10194 11056
rect 10888 10810 10916 11494
rect 10980 11150 11008 12174
rect 11256 11898 11284 12242
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 11440 10674 11468 11290
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10152 9897 10180 9998
rect 10138 9888 10194 9897
rect 10138 9823 10194 9832
rect 10244 9761 10272 10134
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10230 9752 10286 9761
rect 10336 9722 10364 10066
rect 10230 9687 10286 9696
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10152 8634 10180 8910
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10152 7750 10180 8570
rect 10704 8430 10732 10406
rect 11624 9926 11652 11154
rect 10968 9920 11020 9926
rect 10782 9888 10838 9897
rect 10968 9862 11020 9868
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 10782 9823 10838 9832
rect 10796 8634 10824 9823
rect 10876 9648 10928 9654
rect 10874 9616 10876 9625
rect 10928 9616 10930 9625
rect 10874 9551 10930 9560
rect 10980 9382 11008 9862
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10152 7206 10180 7686
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10690 7168 10746 7177
rect 10152 6118 10180 7142
rect 10289 7100 10585 7120
rect 10690 7103 10746 7112
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10704 6934 10732 7103
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10704 6186 10732 6598
rect 10796 6458 10824 7346
rect 10980 7342 11008 8026
rect 11164 7886 11192 9386
rect 11336 9376 11388 9382
rect 11334 9344 11336 9353
rect 11388 9344 11390 9353
rect 11334 9279 11390 9288
rect 11624 8838 11652 9862
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11256 8344 11284 8434
rect 11256 8316 11468 8344
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11164 7585 11192 7822
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11150 7576 11206 7585
rect 11150 7511 11206 7520
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10152 5846 10180 6054
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10782 5672 10838 5681
rect 10782 5607 10838 5616
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10244 5166 10272 5510
rect 10796 5234 10824 5607
rect 10888 5370 10916 7142
rect 10980 7002 11008 7278
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11072 5914 11100 6802
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11164 5846 11192 6598
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10980 5522 11008 5714
rect 10980 5494 11100 5522
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10152 4865 10180 4966
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10138 4856 10194 4865
rect 10289 4848 10585 4868
rect 10138 4791 10194 4800
rect 10704 4282 10732 5102
rect 10968 5024 11020 5030
rect 11072 4978 11100 5494
rect 11164 5370 11192 5782
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11020 4972 11100 4978
rect 10968 4966 11100 4972
rect 10980 4950 11100 4966
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 11072 3738 11100 4950
rect 11152 4480 11204 4486
rect 11150 4448 11152 4457
rect 11204 4448 11206 4457
rect 11150 4383 11206 4392
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10782 3496 10838 3505
rect 10048 3460 10100 3466
rect 10100 3420 10180 3448
rect 10782 3431 10838 3440
rect 10048 3402 10100 3408
rect 10152 2553 10180 3420
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2582 10732 2790
rect 10692 2576 10744 2582
rect 10138 2544 10194 2553
rect 10692 2518 10744 2524
rect 10138 2479 10194 2488
rect 10152 480 10180 2479
rect 10796 2281 10824 3431
rect 11164 2961 11192 3538
rect 11256 3369 11284 7686
rect 11348 7206 11376 7890
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 6662 11376 7142
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11348 6254 11376 6598
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11242 3360 11298 3369
rect 11242 3295 11298 3304
rect 11150 2952 11206 2961
rect 11150 2887 11206 2896
rect 11164 2854 11192 2887
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11164 2650 11192 2790
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 10782 2272 10838 2281
rect 10782 2207 10838 2216
rect 10796 480 10824 2207
rect 11348 480 11376 5102
rect 11440 2106 11468 8316
rect 11624 8129 11652 8774
rect 11716 8566 11744 12582
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10742 11836 11086
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11992 10130 12020 14214
rect 12268 13870 12296 14214
rect 12256 13864 12308 13870
rect 12360 13852 12388 14826
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12452 14006 12480 14214
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12440 13864 12492 13870
rect 12360 13824 12440 13852
rect 12256 13806 12308 13812
rect 12440 13806 12492 13812
rect 12452 13394 12480 13806
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12268 11642 12296 12038
rect 12348 11756 12400 11762
rect 12452 11744 12480 12854
rect 12400 11716 12480 11744
rect 12348 11698 12400 11704
rect 12268 11614 12388 11642
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12070 11384 12126 11393
rect 12268 11354 12296 11494
rect 12070 11319 12126 11328
rect 12256 11348 12308 11354
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11808 8634 11836 8978
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11610 8120 11666 8129
rect 11808 8090 11836 8570
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11610 8055 11666 8064
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11624 4078 11652 5850
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11716 4185 11744 4422
rect 11702 4176 11758 4185
rect 11702 4111 11758 4120
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11428 2100 11480 2106
rect 11428 2042 11480 2048
rect 11716 1465 11744 2246
rect 11702 1456 11758 1465
rect 11702 1391 11758 1400
rect 11900 480 11928 8298
rect 12084 5352 12112 11319
rect 12256 11290 12308 11296
rect 12254 10976 12310 10985
rect 12254 10911 12310 10920
rect 12162 10704 12218 10713
rect 12162 10639 12218 10648
rect 12176 9994 12204 10639
rect 12268 10470 12296 10911
rect 12360 10690 12388 11614
rect 12544 10810 12572 18527
rect 13084 15496 13136 15502
rect 12898 15464 12954 15473
rect 13084 15438 13136 15444
rect 12898 15399 12954 15408
rect 12808 14952 12860 14958
rect 12714 14920 12770 14929
rect 12808 14894 12860 14900
rect 12714 14855 12770 14864
rect 12728 14550 12756 14855
rect 12716 14544 12768 14550
rect 12716 14486 12768 14492
rect 12716 14408 12768 14414
rect 12714 14376 12716 14385
rect 12768 14376 12770 14385
rect 12714 14311 12770 14320
rect 12728 14074 12756 14311
rect 12820 14074 12848 14894
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12714 13832 12770 13841
rect 12714 13767 12770 13776
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12360 10674 12480 10690
rect 12360 10668 12492 10674
rect 12360 10662 12440 10668
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12360 9586 12388 10662
rect 12440 10610 12492 10616
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12452 9654 12480 9998
rect 12544 9926 12572 10474
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12360 9110 12388 9522
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12360 8634 12388 9046
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12452 8430 12480 8774
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 11992 5324 12112 5352
rect 11992 4010 12020 5324
rect 12070 5264 12126 5273
rect 12070 5199 12126 5208
rect 12084 4826 12112 5199
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 12176 610 12204 8230
rect 12452 7993 12480 8366
rect 12544 8265 12572 9862
rect 12728 8616 12756 13767
rect 12820 13394 12848 14010
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12820 12442 12848 13330
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12728 8588 12848 8616
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12636 8401 12664 8502
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12622 8392 12678 8401
rect 12622 8327 12678 8336
rect 12530 8256 12586 8265
rect 12530 8191 12586 8200
rect 12728 8090 12756 8434
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12438 7984 12494 7993
rect 12438 7919 12494 7928
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 7313 12296 7686
rect 12254 7304 12310 7313
rect 12254 7239 12310 7248
rect 12820 6798 12848 8588
rect 12912 7546 12940 15399
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 15201 13032 15302
rect 12990 15192 13046 15201
rect 12990 15127 13046 15136
rect 13004 14890 13032 15127
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 12850 13032 14350
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13004 9897 13032 10066
rect 12990 9888 13046 9897
rect 12990 9823 13046 9832
rect 12990 9752 13046 9761
rect 12990 9687 13046 9696
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12912 7342 12940 7482
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 13004 6644 13032 9687
rect 13096 7018 13124 15438
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13188 13870 13216 14214
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13280 11257 13308 11562
rect 13266 11248 13322 11257
rect 13266 11183 13322 11192
rect 13266 10840 13322 10849
rect 13266 10775 13322 10784
rect 13176 10192 13228 10198
rect 13280 10180 13308 10775
rect 13372 10538 13400 18799
rect 13912 15088 13964 15094
rect 13912 15030 13964 15036
rect 14002 15056 14058 15065
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13556 13462 13584 13874
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13556 12986 13584 13398
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13556 12442 13584 12922
rect 13740 12714 13860 12730
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13740 12708 13872 12714
rect 13740 12702 13820 12708
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13452 11688 13504 11694
rect 13556 11676 13584 12378
rect 13648 11694 13676 12650
rect 13740 12170 13768 12702
rect 13820 12650 13872 12656
rect 13924 12594 13952 15030
rect 14002 14991 14058 15000
rect 13832 12566 13952 12594
rect 13832 12306 13860 12566
rect 14016 12458 14044 14991
rect 13924 12430 14044 12458
rect 14108 12442 14136 18822
rect 14278 18728 14334 18737
rect 14278 18663 14334 18672
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14096 12436 14148 12442
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13504 11648 13584 11676
rect 13636 11688 13688 11694
rect 13452 11630 13504 11636
rect 13636 11630 13688 11636
rect 13464 10810 13492 11630
rect 13648 11354 13676 11630
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13464 10305 13492 10542
rect 13450 10296 13506 10305
rect 13450 10231 13506 10240
rect 13360 10192 13412 10198
rect 13280 10152 13360 10180
rect 13176 10134 13228 10140
rect 13360 10134 13412 10140
rect 13188 9738 13216 10134
rect 13372 9761 13400 10134
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13358 9752 13414 9761
rect 13188 9722 13308 9738
rect 13188 9716 13320 9722
rect 13188 9710 13268 9716
rect 13188 9625 13216 9710
rect 13358 9687 13414 9696
rect 13268 9658 13320 9664
rect 13360 9648 13412 9654
rect 13174 9616 13230 9625
rect 13360 9590 13412 9596
rect 13174 9551 13230 9560
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13188 9110 13216 9318
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13188 8294 13216 9046
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13188 7342 13216 8230
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13096 6990 13308 7018
rect 12820 6616 13032 6644
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12268 5166 12296 6054
rect 12544 5681 12572 6326
rect 12530 5672 12586 5681
rect 12530 5607 12586 5616
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12360 3641 12388 4422
rect 12346 3632 12402 3641
rect 12346 3567 12402 3576
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12728 2990 12756 3470
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12820 2514 12848 6616
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12990 5944 13046 5953
rect 13096 5914 13124 6122
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12990 5879 13046 5888
rect 13084 5908 13136 5914
rect 13004 5794 13032 5879
rect 13084 5850 13136 5856
rect 13004 5766 13124 5794
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13004 4010 13032 4422
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 3097 12940 3878
rect 12898 3088 12954 3097
rect 12898 3023 12954 3032
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12806 2408 12862 2417
rect 12806 2343 12808 2352
rect 12860 2343 12862 2352
rect 12808 2314 12860 2320
rect 13004 1329 13032 3946
rect 12990 1320 13046 1329
rect 12990 1255 13046 1264
rect 12164 604 12216 610
rect 12164 546 12216 552
rect 12532 604 12584 610
rect 12532 546 12584 552
rect 12544 480 12572 546
rect 13096 480 13124 5766
rect 13188 5098 13216 6054
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13188 4826 13216 5034
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13280 4758 13308 6990
rect 13372 6361 13400 9590
rect 13464 9178 13492 9998
rect 13556 9586 13584 10950
rect 13740 10470 13768 11222
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13450 8528 13506 8537
rect 13450 8463 13506 8472
rect 13464 8022 13492 8463
rect 13452 8016 13504 8022
rect 13452 7958 13504 7964
rect 13464 7002 13492 7958
rect 13556 7818 13584 9522
rect 13648 9450 13676 9930
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13740 8090 13768 10202
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13832 8294 13860 9454
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 8090 13860 8230
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13832 7342 13860 8026
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13726 6896 13782 6905
rect 13544 6860 13596 6866
rect 13726 6831 13782 6840
rect 13544 6802 13596 6808
rect 13358 6352 13414 6361
rect 13556 6322 13584 6802
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6458 13676 6734
rect 13740 6730 13768 6831
rect 13832 6730 13860 7142
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13358 6287 13414 6296
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 5574 13584 6258
rect 13740 5846 13768 6666
rect 13818 6624 13874 6633
rect 13818 6559 13874 6568
rect 13832 5914 13860 6559
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13726 5672 13782 5681
rect 13726 5607 13728 5616
rect 13780 5607 13782 5616
rect 13728 5578 13780 5584
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13280 4282 13308 4694
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13280 3738 13308 3946
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13556 1630 13584 5510
rect 13924 5098 13952 12430
rect 14096 12378 14148 12384
rect 14094 12336 14150 12345
rect 14094 12271 14150 12280
rect 14108 12238 14136 12271
rect 14096 12232 14148 12238
rect 14200 12220 14228 13126
rect 14292 12374 14320 18663
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14568 15706 14596 15914
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14568 15026 14596 15642
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14660 14600 14688 26386
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15936 24880 15988 24886
rect 15936 24822 15988 24828
rect 21180 24880 21232 24886
rect 21180 24822 21232 24828
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14738 22536 14794 22545
rect 14738 22471 14794 22480
rect 14752 15978 14780 22471
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14844 16114 14872 16390
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14844 14890 14872 16050
rect 15672 15638 15700 16118
rect 15660 15632 15712 15638
rect 15566 15600 15622 15609
rect 15660 15574 15712 15580
rect 15566 15535 15622 15544
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14568 14572 14688 14600
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14384 12714 14412 13670
rect 14462 13152 14518 13161
rect 14462 13087 14518 13096
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14476 12594 14504 13087
rect 14568 12918 14596 14572
rect 14844 14498 14872 14826
rect 15120 14822 15148 14894
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 14660 14470 14872 14498
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14660 12782 14688 14470
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14752 12986 14780 14282
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14832 13796 14884 13802
rect 14832 13738 14884 13744
rect 14844 13190 14872 13738
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14832 12912 14884 12918
rect 14738 12880 14794 12889
rect 14832 12854 14884 12860
rect 14738 12815 14740 12824
rect 14792 12815 14794 12824
rect 14740 12786 14792 12792
rect 14648 12776 14700 12782
rect 14700 12724 14780 12730
rect 14648 12718 14780 12724
rect 14660 12702 14780 12718
rect 14476 12566 14688 12594
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14280 12232 14332 12238
rect 14200 12192 14280 12220
rect 14096 12174 14148 12180
rect 14280 12174 14332 12180
rect 14108 11626 14136 12174
rect 14292 11898 14320 12174
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14384 11098 14412 12378
rect 14464 12368 14516 12374
rect 14464 12310 14516 12316
rect 14476 11218 14504 12310
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 14016 10266 14044 10678
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14002 9208 14058 9217
rect 14002 9143 14058 9152
rect 14096 9172 14148 9178
rect 14016 8537 14044 9143
rect 14096 9114 14148 9120
rect 14002 8528 14058 8537
rect 14002 8463 14058 8472
rect 14108 8430 14136 9114
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14186 8392 14242 8401
rect 14108 7954 14136 8366
rect 14186 8327 14242 8336
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14108 7002 14136 7890
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14016 6186 14044 6802
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6254 14136 6598
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 14016 5234 14044 6122
rect 14108 5642 14136 6190
rect 14200 5846 14228 8327
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14200 5370 14228 5782
rect 14292 5545 14320 11086
rect 14384 11070 14504 11098
rect 14278 5536 14334 5545
rect 14278 5471 14334 5480
rect 14370 5400 14426 5409
rect 14188 5364 14240 5370
rect 14370 5335 14426 5344
rect 14188 5306 14240 5312
rect 14280 5296 14332 5302
rect 14278 5264 14280 5273
rect 14332 5264 14334 5273
rect 14004 5228 14056 5234
rect 14384 5234 14412 5335
rect 14278 5199 14334 5208
rect 14372 5228 14424 5234
rect 14004 5170 14056 5176
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13924 4758 13952 5034
rect 14292 4826 14320 5199
rect 14372 5170 14424 5176
rect 14476 5166 14504 11070
rect 14660 10606 14688 12566
rect 14752 12442 14780 12702
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14844 11898 14872 12854
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14844 11558 14872 11834
rect 15198 11792 15254 11801
rect 15198 11727 15254 11736
rect 14832 11552 14884 11558
rect 15212 11529 15240 11727
rect 14832 11494 14884 11500
rect 15198 11520 15254 11529
rect 15198 11455 15254 11464
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14844 10810 14872 11154
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14660 10266 14688 10542
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14554 9344 14610 9353
rect 14554 9279 14610 9288
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13740 3602 13768 4626
rect 14384 4321 14412 4762
rect 14370 4312 14426 4321
rect 14370 4247 14426 4256
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14200 3670 14228 4082
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14188 3664 14240 3670
rect 14384 3641 14412 3878
rect 14568 3738 14596 9279
rect 14660 7342 14688 10066
rect 14752 9178 14780 10678
rect 14830 10160 14886 10169
rect 14830 10095 14886 10104
rect 14844 9625 14872 10095
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15108 9648 15160 9654
rect 14830 9616 14886 9625
rect 15108 9590 15160 9596
rect 14830 9551 14886 9560
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14738 8120 14794 8129
rect 14844 8090 14872 9386
rect 15120 9110 15148 9590
rect 15304 9110 15332 14350
rect 15396 11218 15424 15302
rect 15488 15162 15516 15438
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15580 15042 15608 15535
rect 15488 15014 15608 15042
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15396 8344 15424 9862
rect 15488 8974 15516 15014
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 14482 15608 14758
rect 15672 14618 15700 14826
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15580 14074 15608 14418
rect 15672 14074 15700 14554
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15672 12782 15700 13466
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15566 11656 15622 11665
rect 15566 11591 15622 11600
rect 15580 11286 15608 11591
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15672 10849 15700 10950
rect 15658 10840 15714 10849
rect 15658 10775 15714 10784
rect 15672 10674 15700 10775
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15672 10198 15700 10610
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15672 9722 15700 10134
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15764 9194 15792 16594
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15856 14346 15884 15574
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15856 12918 15884 13262
rect 15948 12986 15976 24822
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20258 24304 20314 24313
rect 20258 24239 20314 24248
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 20074 23352 20130 23361
rect 19996 23310 20074 23338
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 16118 20360 16174 20369
rect 16118 20295 16174 20304
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15856 12102 15884 12718
rect 15948 12714 15976 12922
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15856 11393 15884 12038
rect 15842 11384 15898 11393
rect 15842 11319 15898 11328
rect 15844 10192 15896 10198
rect 15844 10134 15896 10140
rect 15856 9382 15884 10134
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15672 9166 15792 9194
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15304 8316 15424 8344
rect 14738 8055 14794 8064
rect 14832 8084 14884 8090
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14660 6866 14688 7142
rect 14752 6866 14780 8055
rect 14832 8026 14884 8032
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 5794 15332 8316
rect 15382 8256 15438 8265
rect 15382 8191 15438 8200
rect 15396 7818 15424 8191
rect 15672 8106 15700 9166
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15764 8634 15792 9046
rect 15948 8673 15976 12174
rect 16026 10568 16082 10577
rect 16026 10503 16028 10512
rect 16080 10503 16082 10512
rect 16028 10474 16080 10480
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16040 9110 16068 9454
rect 16132 9432 16160 20295
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 16486 19816 16542 19825
rect 16486 19751 16542 19760
rect 16500 16153 16528 19751
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 16854 17232 16910 17241
rect 16854 17167 16910 17176
rect 16210 16144 16266 16153
rect 16210 16079 16266 16088
rect 16486 16144 16542 16153
rect 16486 16079 16542 16088
rect 16224 13734 16252 16079
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16302 15056 16358 15065
rect 16302 14991 16358 15000
rect 16316 14385 16344 14991
rect 16408 14550 16436 15098
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16302 14376 16358 14385
rect 16302 14311 16358 14320
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16224 11898 16252 13398
rect 16316 13326 16344 14311
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16408 13530 16436 13670
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16500 13002 16528 15846
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16592 15162 16620 15506
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16592 13530 16620 14486
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16316 12974 16528 13002
rect 16316 12442 16344 12974
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16408 11762 16436 12854
rect 16500 12832 16528 12974
rect 16580 12844 16632 12850
rect 16500 12804 16580 12832
rect 16580 12786 16632 12792
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16500 10810 16528 11222
rect 16592 11014 16620 11766
rect 16684 11354 16712 13194
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10062 16436 10406
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16868 9994 16896 17167
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 17314 16552 17370 16561
rect 17314 16487 17370 16496
rect 17328 15473 17356 16487
rect 17592 15496 17644 15502
rect 17314 15464 17370 15473
rect 17592 15438 17644 15444
rect 17314 15399 17370 15408
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16960 13734 16988 14418
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 13394 17264 13670
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17236 12646 17264 13330
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 12288 17264 12582
rect 17316 12300 17368 12306
rect 17236 12260 17316 12288
rect 17236 11558 17264 12260
rect 17316 12242 17368 12248
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 16960 11082 16988 11494
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16488 9512 16540 9518
rect 16592 9500 16620 9862
rect 16540 9472 16620 9500
rect 16854 9480 16910 9489
rect 16488 9454 16540 9460
rect 16132 9404 16252 9432
rect 16854 9415 16910 9424
rect 16118 9208 16174 9217
rect 16118 9143 16174 9152
rect 16028 9104 16080 9110
rect 16028 9046 16080 9052
rect 15934 8664 15990 8673
rect 15752 8628 15804 8634
rect 16132 8634 16160 9143
rect 15934 8599 15990 8608
rect 16120 8628 16172 8634
rect 15752 8570 15804 8576
rect 16120 8570 16172 8576
rect 16132 8430 16160 8570
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 15842 8256 15898 8265
rect 15842 8191 15898 8200
rect 15672 8078 15792 8106
rect 15856 8090 15884 8191
rect 15934 8120 15990 8129
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15672 7002 15700 7890
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15474 6488 15530 6497
rect 15474 6423 15530 6432
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15396 5846 15424 6054
rect 15488 5914 15516 6423
rect 15580 6118 15608 6734
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15212 5778 15332 5794
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15200 5772 15332 5778
rect 15252 5766 15332 5772
rect 15200 5714 15252 5720
rect 15212 5658 15240 5714
rect 15212 5630 15424 5658
rect 15580 5642 15608 6054
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15108 5160 15160 5166
rect 15108 5102 15160 5108
rect 14832 5092 14884 5098
rect 14832 5034 14884 5040
rect 14844 4690 14872 5034
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 15120 4593 15148 5102
rect 15304 4865 15332 5510
rect 15396 5370 15424 5630
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15290 4856 15346 4865
rect 15290 4791 15346 4800
rect 15474 4856 15530 4865
rect 15474 4791 15530 4800
rect 14646 4584 14702 4593
rect 14646 4519 14702 4528
rect 15106 4584 15162 4593
rect 15106 4519 15162 4528
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14188 3606 14240 3612
rect 14370 3632 14426 3641
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13740 2990 13768 3538
rect 14200 3194 14228 3606
rect 14370 3567 14426 3576
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 14660 2650 14688 4519
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14844 4146 14872 4422
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 15488 4010 15516 4791
rect 15580 4570 15608 5578
rect 15660 4616 15712 4622
rect 15580 4564 15660 4570
rect 15580 4558 15712 4564
rect 15580 4542 15700 4558
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15396 3466 15424 3878
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 14752 2922 14780 3334
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 14648 2644 14700 2650
rect 14292 2604 14648 2632
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13648 2310 13676 2518
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 13910 2408 13966 2417
rect 13910 2343 13912 2352
rect 13964 2343 13966 2352
rect 13912 2314 13964 2320
rect 13636 2304 13688 2310
rect 13634 2272 13636 2281
rect 13688 2272 13690 2281
rect 13634 2207 13690 2216
rect 14200 1737 14228 2450
rect 14186 1728 14242 1737
rect 14186 1663 14242 1672
rect 13544 1624 13596 1630
rect 13544 1566 13596 1572
rect 13634 912 13690 921
rect 13634 847 13690 856
rect 13648 480 13676 847
rect 14292 480 14320 2604
rect 14648 2586 14700 2592
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 14844 480 14872 2450
rect 15304 2446 15332 3334
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15396 1737 15424 3402
rect 15488 2378 15516 3946
rect 15580 3942 15608 4542
rect 15658 4040 15714 4049
rect 15658 3975 15714 3984
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15580 3602 15608 3878
rect 15672 3670 15700 3975
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15580 2990 15608 3538
rect 15672 3194 15700 3606
rect 15764 3233 15792 8078
rect 15844 8084 15896 8090
rect 15934 8055 15990 8064
rect 15844 8026 15896 8032
rect 15856 7546 15884 8026
rect 15948 8022 15976 8055
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 16224 7732 16252 9404
rect 16868 9382 16896 9415
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16302 9072 16358 9081
rect 16302 9007 16304 9016
rect 16356 9007 16358 9016
rect 16304 8978 16356 8984
rect 16316 8498 16344 8978
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16408 8566 16436 8910
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 7886 16344 8230
rect 16304 7880 16356 7886
rect 16302 7848 16304 7857
rect 16356 7848 16358 7857
rect 16302 7783 16358 7792
rect 16224 7704 16344 7732
rect 16118 7576 16174 7585
rect 15844 7540 15896 7546
rect 16174 7520 16252 7528
rect 16118 7511 16120 7520
rect 15844 7482 15896 7488
rect 16172 7500 16252 7520
rect 16120 7482 16172 7488
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 15842 6216 15898 6225
rect 16132 6186 16160 6802
rect 15842 6151 15898 6160
rect 16120 6180 16172 6186
rect 15856 5370 15884 6151
rect 16120 6122 16172 6128
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 16224 5234 16252 7500
rect 16316 7206 16344 7704
rect 16500 7313 16528 8774
rect 16486 7304 16542 7313
rect 16486 7239 16542 7248
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16592 6440 16620 9318
rect 16670 8936 16726 8945
rect 16670 8871 16672 8880
rect 16724 8871 16726 8880
rect 16854 8936 16910 8945
rect 16854 8871 16910 8880
rect 16672 8842 16724 8848
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16684 7274 16712 7686
rect 16762 7440 16818 7449
rect 16762 7375 16818 7384
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16684 6866 16712 7210
rect 16776 7206 16804 7375
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16500 6412 16620 6440
rect 16500 5681 16528 6412
rect 16578 6352 16634 6361
rect 16868 6322 16896 8871
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 17052 8401 17080 8774
rect 17038 8392 17094 8401
rect 17038 8327 17094 8336
rect 16578 6287 16634 6296
rect 16856 6316 16908 6322
rect 16592 6254 16620 6287
rect 16856 6258 16908 6264
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 17144 5681 17172 10474
rect 17236 10470 17264 11086
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17236 10146 17264 10406
rect 17328 10266 17356 11290
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17408 10192 17460 10198
rect 17236 10118 17356 10146
rect 17408 10134 17460 10140
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 5846 17264 6598
rect 17328 6225 17356 10118
rect 17420 10033 17448 10134
rect 17406 10024 17462 10033
rect 17406 9959 17462 9968
rect 17604 9704 17632 15438
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17696 13462 17724 14214
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17696 12374 17724 12786
rect 17774 12744 17830 12753
rect 17774 12679 17776 12688
rect 17828 12679 17830 12688
rect 17776 12650 17828 12656
rect 17684 12368 17736 12374
rect 17684 12310 17736 12316
rect 17696 11898 17724 12310
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17696 11286 17724 11834
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17696 10266 17724 10950
rect 17788 10470 17816 11494
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17604 9676 17724 9704
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17420 8294 17448 8910
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17604 8362 17632 8774
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 6934 17448 8230
rect 17512 8022 17540 8053
rect 17500 8016 17552 8022
rect 17498 7984 17500 7993
rect 17552 7984 17554 7993
rect 17498 7919 17554 7928
rect 17512 7546 17540 7919
rect 17604 7818 17632 8298
rect 17592 7812 17644 7818
rect 17592 7754 17644 7760
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17696 7041 17724 9676
rect 17788 9450 17816 10406
rect 17776 9444 17828 9450
rect 17776 9386 17828 9392
rect 17788 9042 17816 9386
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17880 7970 17908 16594
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18156 14890 18184 15506
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 18248 14278 18276 14894
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17972 11354 18000 11698
rect 18052 11688 18104 11694
rect 18050 11656 18052 11665
rect 18104 11656 18106 11665
rect 18156 11626 18184 12038
rect 18050 11591 18106 11600
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 18050 11520 18106 11529
rect 18050 11455 18106 11464
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 18064 11257 18092 11455
rect 18156 11354 18184 11562
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18050 11248 18106 11257
rect 18050 11183 18106 11192
rect 18064 10130 18092 11183
rect 18156 10606 18184 11290
rect 18248 11014 18276 14214
rect 18340 13977 18368 15302
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18326 13968 18382 13977
rect 18326 13903 18382 13912
rect 18328 13864 18380 13870
rect 18326 13832 18328 13841
rect 18380 13832 18382 13841
rect 18326 13767 18382 13776
rect 18432 12617 18460 14350
rect 18602 13696 18658 13705
rect 18602 13631 18658 13640
rect 18616 13297 18644 13631
rect 18602 13288 18658 13297
rect 18602 13223 18658 13232
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12850 18552 13126
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18418 12608 18474 12617
rect 18474 12566 18552 12594
rect 18418 12543 18474 12552
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17972 9110 18000 9590
rect 18064 9586 18092 10066
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18156 9450 18184 9930
rect 18248 9722 18276 10202
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 17880 7942 18000 7970
rect 17682 7032 17738 7041
rect 17682 6967 17738 6976
rect 17408 6928 17460 6934
rect 17408 6870 17460 6876
rect 17420 6458 17448 6870
rect 17880 6866 17908 7942
rect 17972 7886 18000 7942
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 18050 6352 18106 6361
rect 18050 6287 18106 6296
rect 18064 6254 18092 6287
rect 18052 6248 18104 6254
rect 17314 6216 17370 6225
rect 18052 6190 18104 6196
rect 17314 6151 17370 6160
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 16486 5672 16542 5681
rect 16396 5636 16448 5642
rect 16486 5607 16542 5616
rect 17130 5672 17186 5681
rect 17130 5607 17186 5616
rect 16396 5578 16448 5584
rect 16408 5370 16436 5578
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16500 5098 16528 5607
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16684 4690 16712 5510
rect 17236 5370 17264 5782
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 15844 4480 15896 4486
rect 15896 4440 15976 4468
rect 15844 4422 15896 4428
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15750 3224 15806 3233
rect 15660 3188 15712 3194
rect 15750 3159 15806 3168
rect 15660 3130 15712 3136
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15382 1728 15438 1737
rect 15382 1663 15438 1672
rect 15384 1624 15436 1630
rect 15384 1566 15436 1572
rect 15396 480 15424 1566
rect 15856 1465 15884 3674
rect 15948 3534 15976 4440
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15948 2650 15976 3470
rect 16132 3398 16160 4626
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16500 3777 16528 3878
rect 16486 3768 16542 3777
rect 16486 3703 16542 3712
rect 16776 3670 16804 4014
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 16776 3194 16804 3606
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16960 3194 16988 3538
rect 16764 3188 16816 3194
rect 16948 3188 17000 3194
rect 16816 3148 16896 3176
rect 16764 3130 16816 3136
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 16578 2816 16634 2825
rect 16578 2751 16634 2760
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16028 2576 16080 2582
rect 16026 2544 16028 2553
rect 16080 2544 16082 2553
rect 16026 2479 16082 2488
rect 16028 2100 16080 2106
rect 16028 2042 16080 2048
rect 15842 1456 15898 1465
rect 15842 1391 15898 1400
rect 16040 480 16068 2042
rect 16592 480 16620 2751
rect 16684 2582 16712 2858
rect 16868 2650 16896 3148
rect 16948 3130 17000 3136
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 17144 2514 17172 3878
rect 17236 2582 17264 4422
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 16946 2136 17002 2145
rect 16946 2071 17002 2080
rect 16960 1465 16988 2071
rect 17144 1601 17172 2450
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17130 1592 17186 1601
rect 17130 1527 17186 1536
rect 16946 1456 17002 1465
rect 16946 1391 17002 1400
rect 17130 1456 17186 1465
rect 17130 1391 17186 1400
rect 17144 480 17172 1391
rect 17236 1193 17264 2246
rect 17328 2009 17356 6054
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17880 3890 17908 5510
rect 18052 5160 18104 5166
rect 18050 5128 18052 5137
rect 18104 5128 18106 5137
rect 18050 5063 18106 5072
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17972 4026 18000 4082
rect 18156 4078 18184 8502
rect 18248 8265 18276 9658
rect 18234 8256 18290 8265
rect 18234 8191 18290 8200
rect 18340 8090 18368 11086
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18248 7857 18276 7890
rect 18234 7848 18290 7857
rect 18234 7783 18290 7792
rect 18248 7546 18276 7783
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18340 7342 18368 8026
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18144 4072 18196 4078
rect 17972 3998 18092 4026
rect 18144 4014 18196 4020
rect 17880 3862 18000 3890
rect 17774 3224 17830 3233
rect 17774 3159 17776 3168
rect 17828 3159 17830 3168
rect 17776 3130 17828 3136
rect 17972 3126 18000 3862
rect 18064 3346 18092 3998
rect 18142 3360 18198 3369
rect 18064 3318 18142 3346
rect 18142 3295 18198 3304
rect 18156 3194 18184 3295
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 17774 2952 17830 2961
rect 17774 2887 17830 2896
rect 17314 2000 17370 2009
rect 17314 1935 17370 1944
rect 17222 1184 17278 1193
rect 17222 1119 17278 1128
rect 17788 480 17816 2887
rect 18248 2689 18276 4966
rect 18340 4049 18368 7142
rect 18432 4690 18460 11494
rect 18524 11286 18552 12566
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 10198 18552 10406
rect 18616 10266 18644 13223
rect 18708 11098 18736 14758
rect 18800 12850 18828 16594
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18800 12442 18828 12786
rect 18878 12744 18934 12753
rect 18878 12679 18880 12688
rect 18932 12679 18934 12688
rect 18880 12650 18932 12656
rect 18788 12436 18840 12442
rect 18984 12424 19012 15846
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19352 15450 19380 15506
rect 19260 15422 19380 15450
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19260 15162 19288 15422
rect 19444 15162 19472 15438
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19444 15065 19472 15098
rect 19430 15056 19486 15065
rect 19430 14991 19486 15000
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19156 13796 19208 13802
rect 19156 13738 19208 13744
rect 19168 13190 19196 13738
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19168 12646 19196 13126
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 12442 19196 12582
rect 18788 12378 18840 12384
rect 18892 12396 19012 12424
rect 19156 12436 19208 12442
rect 18708 11070 18828 11098
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18512 10192 18564 10198
rect 18512 10134 18564 10140
rect 18524 9654 18552 10134
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 18524 8090 18552 9590
rect 18616 8362 18644 9862
rect 18708 9489 18736 10950
rect 18800 9722 18828 11070
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18786 9616 18842 9625
rect 18786 9551 18842 9560
rect 18694 9480 18750 9489
rect 18694 9415 18750 9424
rect 18604 8356 18656 8362
rect 18800 8344 18828 9551
rect 18892 8537 18920 12396
rect 19156 12378 19208 12384
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18984 11898 19012 12242
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18984 9994 19012 11630
rect 19260 11234 19288 14826
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19352 12889 19380 13942
rect 19444 13870 19472 14894
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19432 12912 19484 12918
rect 19338 12880 19394 12889
rect 19432 12854 19484 12860
rect 19338 12815 19394 12824
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19352 11354 19380 12310
rect 19444 12238 19472 12854
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19260 11206 19380 11234
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 18972 9988 19024 9994
rect 18972 9930 19024 9936
rect 19168 9602 19196 9998
rect 19352 9738 19380 11206
rect 19444 11150 19472 11494
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19137 9574 19196 9602
rect 19260 9710 19380 9738
rect 18972 9444 19024 9450
rect 18972 9386 19024 9392
rect 18984 9178 19012 9386
rect 19137 9194 19165 9574
rect 18972 9172 19024 9178
rect 19137 9166 19196 9194
rect 18972 9114 19024 9120
rect 18878 8528 18934 8537
rect 18984 8498 19012 9114
rect 18878 8463 18934 8472
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18800 8316 19012 8344
rect 18604 8298 18656 8304
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18524 7002 18552 8026
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18892 6458 18920 7278
rect 18984 6780 19012 8316
rect 19168 8022 19196 9166
rect 19156 8016 19208 8022
rect 19156 7958 19208 7964
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 19062 7168 19118 7177
rect 19062 7103 19118 7112
rect 19076 6934 19104 7103
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 18984 6752 19104 6780
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18892 6254 18920 6394
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18786 5536 18842 5545
rect 18786 5471 18842 5480
rect 18510 4992 18566 5001
rect 18510 4927 18566 4936
rect 18420 4684 18472 4690
rect 18420 4626 18472 4632
rect 18326 4040 18382 4049
rect 18326 3975 18382 3984
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 18432 3233 18460 3946
rect 18524 3738 18552 4927
rect 18800 4434 18828 5471
rect 18892 5370 18920 6190
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 18984 5098 19012 5510
rect 18972 5092 19024 5098
rect 18972 5034 19024 5040
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18878 4448 18934 4457
rect 18800 4406 18878 4434
rect 18878 4383 18934 4392
rect 18892 4146 18920 4383
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18892 3942 18920 4082
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18418 3224 18474 3233
rect 18418 3159 18474 3168
rect 18234 2680 18290 2689
rect 18234 2615 18290 2624
rect 18432 2378 18460 3159
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 18708 2582 18736 2858
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 18788 2440 18840 2446
rect 18786 2408 18788 2417
rect 18840 2408 18842 2417
rect 18420 2372 18472 2378
rect 18786 2343 18842 2352
rect 18420 2314 18472 2320
rect 18326 1592 18382 1601
rect 18326 1527 18382 1536
rect 18340 480 18368 1527
rect 18984 610 19012 4626
rect 19076 921 19104 6752
rect 19168 5914 19196 7686
rect 19260 6322 19288 9710
rect 19444 8838 19472 10066
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19352 7274 19380 7958
rect 19536 7834 19564 17614
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19996 15706 20024 23310
rect 20074 23287 20130 23296
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14618 20024 15642
rect 20074 15192 20130 15201
rect 20074 15127 20130 15136
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 20088 14482 20116 15127
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19892 14272 19944 14278
rect 19892 14214 19944 14220
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19904 14113 19932 14214
rect 19890 14104 19946 14113
rect 19890 14039 19946 14048
rect 19996 13734 20024 14214
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19996 12782 20024 13670
rect 20088 13530 20116 14418
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19996 11898 20024 12718
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19720 10606 19748 11154
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19628 9518 19656 9862
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19708 8832 19760 8838
rect 19706 8800 19708 8809
rect 19760 8800 19762 8809
rect 19706 8735 19762 8744
rect 19996 8634 20024 11222
rect 20088 10690 20116 13126
rect 20180 12238 20208 18022
rect 20272 12442 20300 24239
rect 20350 21584 20406 21593
rect 20350 21519 20406 21528
rect 20364 16017 20392 21519
rect 21192 17105 21220 24822
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21178 17096 21234 17105
rect 21178 17031 21234 17040
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 20350 16008 20406 16017
rect 20350 15943 20406 15952
rect 20364 15586 20392 15943
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20456 15745 20484 15846
rect 20442 15736 20498 15745
rect 20442 15671 20498 15680
rect 20364 15558 20484 15586
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20364 14890 20392 15302
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 11218 20208 12038
rect 20272 11354 20300 12106
rect 20364 12102 20392 13330
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20364 11286 20392 12038
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20088 10662 20208 10690
rect 20076 10600 20128 10606
rect 20074 10568 20076 10577
rect 20128 10568 20130 10577
rect 20074 10503 20130 10512
rect 20074 9616 20130 9625
rect 20074 9551 20130 9560
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19996 8430 20024 8570
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 20088 8242 20116 9551
rect 20180 9042 20208 10662
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 19996 8214 20116 8242
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19444 7806 19564 7834
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19338 7032 19394 7041
rect 19338 6967 19394 6976
rect 19352 6798 19380 6967
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 19352 5778 19380 6598
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19248 5704 19300 5710
rect 19248 5646 19300 5652
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19168 4185 19196 5510
rect 19260 4758 19288 5646
rect 19352 4826 19380 5714
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 19338 4720 19394 4729
rect 19338 4655 19394 4664
rect 19154 4176 19210 4185
rect 19154 4111 19210 4120
rect 19352 3194 19380 4655
rect 19444 4010 19472 7806
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19536 7274 19564 7686
rect 19904 7342 19932 7686
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 19536 6866 19564 7210
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19616 6928 19668 6934
rect 19616 6870 19668 6876
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19628 6458 19656 6870
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5092 19576 5098
rect 19524 5034 19576 5040
rect 19536 4690 19564 5034
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19616 4752 19668 4758
rect 19616 4694 19668 4700
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19628 4282 19656 4694
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19904 4146 19932 4422
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19522 4040 19578 4049
rect 19432 4004 19484 4010
rect 19522 3975 19578 3984
rect 19432 3946 19484 3952
rect 19430 3768 19486 3777
rect 19430 3703 19486 3712
rect 19444 3602 19472 3703
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19338 2816 19394 2825
rect 19338 2751 19394 2760
rect 19352 2650 19380 2751
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19444 2553 19472 3538
rect 19430 2544 19486 2553
rect 19430 2479 19486 2488
rect 19062 912 19118 921
rect 19062 847 19118 856
rect 18880 604 18932 610
rect 18880 546 18932 552
rect 18972 604 19024 610
rect 18972 546 19024 552
rect 18892 480 18920 546
rect 19536 480 19564 3975
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19996 3670 20024 8214
rect 20074 7712 20130 7721
rect 20074 7647 20130 7656
rect 20088 6934 20116 7647
rect 20180 7177 20208 8774
rect 20272 7206 20300 11086
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20260 7200 20312 7206
rect 20166 7168 20222 7177
rect 20260 7142 20312 7148
rect 20166 7103 20222 7112
rect 20364 7041 20392 11018
rect 20456 9178 20484 15558
rect 20548 14550 20576 16934
rect 20628 15904 20680 15910
rect 20626 15872 20628 15881
rect 20680 15872 20682 15881
rect 20626 15807 20682 15816
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20640 14006 20668 14758
rect 20732 14618 20760 15370
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20640 12442 20668 13942
rect 20732 13530 20760 14350
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20548 12322 20576 12378
rect 20548 12294 20668 12322
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20548 10010 20576 12174
rect 20640 10305 20668 12294
rect 20732 12102 20760 12718
rect 20824 12481 20852 16934
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20916 15502 20944 15846
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20916 14958 20944 15438
rect 21008 15162 21036 15506
rect 21100 15473 21128 16934
rect 21086 15464 21142 15473
rect 21086 15399 21142 15408
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20904 14952 20956 14958
rect 20904 14894 20956 14900
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20810 12472 20866 12481
rect 20810 12407 20866 12416
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11898 20760 12038
rect 20916 11937 20944 14214
rect 21192 13530 21220 17031
rect 21548 16516 21600 16522
rect 21548 16458 21600 16464
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 21008 12442 21036 13126
rect 21192 12986 21220 13466
rect 21284 13002 21312 16390
rect 21560 15978 21588 16458
rect 21548 15972 21600 15978
rect 21548 15914 21600 15920
rect 21454 15872 21510 15881
rect 21454 15807 21510 15816
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21376 14074 21404 14486
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21180 12980 21232 12986
rect 21284 12974 21404 13002
rect 21180 12922 21232 12928
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 21270 12336 21326 12345
rect 21270 12271 21272 12280
rect 21324 12271 21326 12280
rect 21272 12242 21324 12248
rect 20902 11928 20958 11937
rect 20720 11892 20772 11898
rect 21284 11898 21312 12242
rect 20902 11863 20958 11872
rect 21272 11892 21324 11898
rect 20720 11834 20772 11840
rect 21272 11834 21324 11840
rect 20718 11656 20774 11665
rect 20718 11591 20774 11600
rect 20732 11354 20760 11591
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20810 11248 20866 11257
rect 20720 11212 20772 11218
rect 20810 11183 20866 11192
rect 20720 11154 20772 11160
rect 20732 10810 20760 11154
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20626 10296 20682 10305
rect 20732 10266 20760 10610
rect 20626 10231 20682 10240
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20548 9982 20668 10010
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20456 8362 20484 9114
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20456 7585 20484 7686
rect 20442 7576 20498 7585
rect 20442 7511 20498 7520
rect 20350 7032 20406 7041
rect 20350 6967 20406 6976
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 20088 5914 20116 6666
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 6254 20300 6598
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 20272 5370 20300 6190
rect 20442 5672 20498 5681
rect 20442 5607 20498 5616
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20166 4856 20222 4865
rect 20166 4791 20222 4800
rect 20180 4758 20208 4791
rect 20168 4752 20220 4758
rect 20074 4720 20130 4729
rect 20168 4694 20220 4700
rect 20352 4752 20404 4758
rect 20352 4694 20404 4700
rect 20074 4655 20130 4664
rect 20260 4684 20312 4690
rect 19984 3664 20036 3670
rect 19984 3606 20036 3612
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19708 3120 19760 3126
rect 19706 3088 19708 3097
rect 19760 3088 19762 3097
rect 19706 3023 19762 3032
rect 19720 2922 19748 3023
rect 19708 2916 19760 2922
rect 19708 2858 19760 2864
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19996 2514 20024 3130
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20088 480 20116 4655
rect 20260 4626 20312 4632
rect 20166 4312 20222 4321
rect 20166 4247 20222 4256
rect 20180 3058 20208 4247
rect 20272 4214 20300 4626
rect 20260 4208 20312 4214
rect 20260 4150 20312 4156
rect 20272 3913 20300 4150
rect 20258 3904 20314 3913
rect 20258 3839 20314 3848
rect 20272 3738 20300 3839
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20364 3534 20392 4694
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20456 3194 20484 5607
rect 20548 4842 20576 9862
rect 20640 9500 20668 9982
rect 20824 9761 20852 11183
rect 21086 10704 21142 10713
rect 21086 10639 21142 10648
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 20916 10062 20944 10474
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20810 9752 20866 9761
rect 20810 9687 20866 9696
rect 20810 9616 20866 9625
rect 20810 9551 20866 9560
rect 20720 9512 20772 9518
rect 20640 9472 20720 9500
rect 20720 9454 20772 9460
rect 20824 8945 20852 9551
rect 20916 9382 20944 9998
rect 20994 9888 21050 9897
rect 20994 9823 21050 9832
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20916 8974 20944 9318
rect 20904 8968 20956 8974
rect 20810 8936 20866 8945
rect 20904 8910 20956 8916
rect 20810 8871 20866 8880
rect 20810 8664 20866 8673
rect 20810 8599 20866 8608
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20732 8090 20760 8502
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20640 5710 20668 7142
rect 20718 6896 20774 6905
rect 20718 6831 20720 6840
rect 20772 6831 20774 6840
rect 20720 6802 20772 6808
rect 20824 6746 20852 8599
rect 20916 8294 20944 8910
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20916 7818 20944 8230
rect 20904 7812 20956 7818
rect 20904 7754 20956 7760
rect 20916 7546 20944 7754
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 20902 7304 20958 7313
rect 20902 7239 20958 7248
rect 20732 6718 20852 6746
rect 20628 5704 20680 5710
rect 20732 5692 20760 6718
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20824 6458 20852 6598
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20812 5704 20864 5710
rect 20732 5664 20812 5692
rect 20628 5646 20680 5652
rect 20812 5646 20864 5652
rect 20916 5522 20944 7239
rect 21008 5953 21036 9823
rect 21100 9586 21128 10639
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21100 9450 21128 9522
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 21192 9110 21220 9590
rect 21180 9104 21232 9110
rect 21180 9046 21232 9052
rect 21192 8498 21220 9046
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 21192 8022 21220 8434
rect 21180 8016 21232 8022
rect 21180 7958 21232 7964
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 20994 5944 21050 5953
rect 20994 5879 21050 5888
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 20732 5494 20944 5522
rect 20548 4814 20668 4842
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 20180 2446 20208 2790
rect 20548 2650 20576 2926
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 20640 480 20668 4814
rect 20732 2990 20760 5494
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20916 4690 20944 5306
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20824 3738 20852 4558
rect 20916 4282 20944 4626
rect 21008 4554 21036 5714
rect 21100 4729 21128 6598
rect 21192 6118 21220 6802
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21086 4720 21142 4729
rect 21086 4655 21142 4664
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 21192 4078 21220 6054
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 21008 3194 21036 3538
rect 20996 3188 21048 3194
rect 20996 3130 21048 3136
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20996 2508 21048 2514
rect 20996 2450 21048 2456
rect 21008 2378 21036 2450
rect 20996 2372 21048 2378
rect 20996 2314 21048 2320
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 20916 1873 20944 2246
rect 21008 2145 21036 2314
rect 21192 2281 21220 3878
rect 21178 2272 21234 2281
rect 21178 2207 21234 2216
rect 20994 2136 21050 2145
rect 20994 2071 21050 2080
rect 20902 1864 20958 1873
rect 20902 1799 20958 1808
rect 21284 480 21312 10406
rect 21376 9217 21404 12974
rect 21362 9208 21418 9217
rect 21362 9143 21418 9152
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21376 8401 21404 8570
rect 21362 8392 21418 8401
rect 21362 8327 21418 8336
rect 21376 4826 21404 8327
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 21468 3058 21496 15807
rect 21560 15366 21588 15914
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21560 14414 21588 15302
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21744 14074 21772 17614
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21836 16794 21864 16934
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 21824 16652 21876 16658
rect 21824 16594 21876 16600
rect 21836 15638 21864 16594
rect 21824 15632 21876 15638
rect 21824 15574 21876 15580
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21560 12782 21588 13262
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21560 12374 21588 12582
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21548 12368 21600 12374
rect 21548 12310 21600 12316
rect 21652 11354 21680 12378
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21560 10470 21588 10542
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21560 8401 21588 10406
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 21744 10033 21772 10066
rect 21730 10024 21786 10033
rect 21730 9959 21786 9968
rect 21730 9888 21786 9897
rect 21730 9823 21786 9832
rect 21640 9444 21692 9450
rect 21640 9386 21692 9392
rect 21652 9081 21680 9386
rect 21638 9072 21694 9081
rect 21638 9007 21694 9016
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21546 8392 21602 8401
rect 21546 8327 21602 8336
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21560 8090 21588 8230
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 21560 5545 21588 7890
rect 21546 5536 21602 5545
rect 21546 5471 21602 5480
rect 21652 3602 21680 8502
rect 21744 5846 21772 9823
rect 21836 9625 21864 15574
rect 21914 13424 21970 13433
rect 21914 13359 21970 13368
rect 21928 10198 21956 13359
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21822 9616 21878 9625
rect 21822 9551 21878 9560
rect 21824 9376 21876 9382
rect 21876 9336 21956 9364
rect 21824 9318 21876 9324
rect 21822 8800 21878 8809
rect 21822 8735 21878 8744
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21744 3942 21772 5646
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 21836 3670 21864 8735
rect 21928 8430 21956 9336
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 22020 4128 22048 26590
rect 23492 26450 23520 27639
rect 23570 27024 23626 27033
rect 23570 26959 23626 26968
rect 23584 26654 23612 26959
rect 23572 26648 23624 26654
rect 23572 26590 23624 26596
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 23478 26344 23534 26353
rect 22192 26308 22244 26314
rect 23478 26279 23480 26288
rect 22192 26250 22244 26256
rect 23532 26279 23534 26288
rect 23480 26250 23532 26256
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22112 14618 22140 14894
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 22112 14346 22140 14554
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 22100 14000 22152 14006
rect 22098 13968 22100 13977
rect 22152 13968 22154 13977
rect 22098 13903 22154 13912
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 22112 12345 22140 13738
rect 22204 13462 22232 26250
rect 23478 25664 23534 25673
rect 23478 25599 23534 25608
rect 23492 24886 23520 25599
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 23480 24880 23532 24886
rect 23480 24822 23532 24828
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 23202 23080 23258 23089
rect 23202 23015 23258 23024
rect 22926 22128 22982 22137
rect 22926 22063 22982 22072
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22282 16688 22338 16697
rect 22282 16623 22338 16632
rect 22192 13456 22244 13462
rect 22192 13398 22244 13404
rect 22204 12986 22232 13398
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22098 12336 22154 12345
rect 22296 12306 22324 16623
rect 22098 12271 22154 12280
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22100 12232 22152 12238
rect 22388 12186 22416 18022
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22480 17338 22508 17682
rect 22742 17640 22798 17649
rect 22742 17575 22798 17584
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22100 12174 22152 12180
rect 22112 11898 22140 12174
rect 22204 12158 22416 12186
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22098 11792 22154 11801
rect 22098 11727 22154 11736
rect 22112 10418 22140 11727
rect 22204 10538 22232 12158
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22296 11694 22324 12038
rect 22388 11801 22416 12038
rect 22374 11792 22430 11801
rect 22374 11727 22430 11736
rect 22284 11688 22336 11694
rect 22480 11642 22508 17274
rect 22572 16998 22600 17478
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22664 16794 22692 17002
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22756 16697 22784 17575
rect 22742 16688 22798 16697
rect 22742 16623 22798 16632
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22572 15910 22600 16526
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22572 13802 22600 15302
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22664 14482 22692 14758
rect 22652 14476 22704 14482
rect 22704 14436 22784 14464
rect 22652 14418 22704 14424
rect 22560 13796 22612 13802
rect 22560 13738 22612 13744
rect 22756 13734 22784 14436
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22756 13326 22784 13670
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22572 12850 22600 13262
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22284 11630 22336 11636
rect 22192 10532 22244 10538
rect 22192 10474 22244 10480
rect 22112 10390 22232 10418
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22112 9110 22140 9522
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 22204 7449 22232 10390
rect 22296 9897 22324 11630
rect 22388 11614 22508 11642
rect 22388 11393 22416 11614
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22374 11384 22430 11393
rect 22374 11319 22430 11328
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22388 10674 22416 10950
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22282 9888 22338 9897
rect 22282 9823 22338 9832
rect 22480 9353 22508 11494
rect 22572 11150 22600 12786
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22664 12442 22692 12718
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22652 12436 22704 12442
rect 22652 12378 22704 12384
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22466 9344 22522 9353
rect 22466 9279 22522 9288
rect 22468 9036 22520 9042
rect 22468 8978 22520 8984
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22388 8498 22416 8774
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22388 8362 22416 8434
rect 22376 8356 22428 8362
rect 22376 8298 22428 8304
rect 22388 8022 22416 8298
rect 22376 8016 22428 8022
rect 22376 7958 22428 7964
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22190 7440 22246 7449
rect 22190 7375 22246 7384
rect 22296 7342 22324 7482
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22112 6662 22140 7278
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22204 6798 22232 7142
rect 22388 6866 22416 7958
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22112 4690 22140 6598
rect 22204 5846 22232 6734
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22282 5944 22338 5953
rect 22282 5879 22338 5888
rect 22192 5840 22244 5846
rect 22192 5782 22244 5788
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 21928 4100 22048 4128
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 21640 3596 21692 3602
rect 21640 3538 21692 3544
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21732 2576 21784 2582
rect 21928 2564 21956 4100
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 22020 3505 22048 3946
rect 22204 3942 22232 5238
rect 22192 3936 22244 3942
rect 22296 3924 22324 5879
rect 22388 5642 22416 6258
rect 22376 5636 22428 5642
rect 22376 5578 22428 5584
rect 22376 4480 22428 4486
rect 22374 4448 22376 4457
rect 22428 4448 22430 4457
rect 22374 4383 22430 4392
rect 22296 3896 22416 3924
rect 22192 3878 22244 3884
rect 22204 3602 22232 3878
rect 22282 3768 22338 3777
rect 22282 3703 22284 3712
rect 22336 3703 22338 3712
rect 22284 3674 22336 3680
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22006 3496 22062 3505
rect 22006 3431 22062 3440
rect 22388 3194 22416 3896
rect 22376 3188 22428 3194
rect 22376 3130 22428 3136
rect 22388 2990 22416 3130
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 22374 2816 22430 2825
rect 22480 2802 22508 8978
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22572 6186 22600 7414
rect 22664 7410 22692 12242
rect 22756 8129 22784 12582
rect 22848 10962 22876 18702
rect 22940 11393 22968 22063
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23032 17202 23060 17614
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23032 16726 23060 17138
rect 23020 16720 23072 16726
rect 23020 16662 23072 16668
rect 23032 16250 23060 16662
rect 23216 16425 23244 23015
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 23662 22264 23718 22273
rect 23662 22199 23718 22208
rect 23478 21040 23534 21049
rect 23478 20975 23534 20984
rect 23492 19394 23520 20975
rect 23400 19366 23520 19394
rect 23296 18080 23348 18086
rect 23296 18022 23348 18028
rect 23202 16416 23258 16425
rect 23202 16351 23258 16360
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23032 15706 23060 16186
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23124 14822 23152 15846
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 23032 13462 23060 13874
rect 23020 13456 23072 13462
rect 23020 13398 23072 13404
rect 23032 12442 23060 13398
rect 23124 13190 23152 14418
rect 23216 14249 23244 16351
rect 23308 15042 23336 18022
rect 23400 17882 23428 19366
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23492 18086 23520 18770
rect 23676 18442 23704 22199
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 23938 20360 23994 20369
rect 23938 20295 23994 20304
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23584 18414 23704 18442
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23388 17876 23440 17882
rect 23388 17818 23440 17824
rect 23400 16658 23428 17818
rect 23584 17649 23612 18414
rect 23570 17640 23626 17649
rect 23570 17575 23626 17584
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23480 17060 23532 17066
rect 23480 17002 23532 17008
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23492 15201 23520 17002
rect 23478 15192 23534 15201
rect 23478 15127 23534 15136
rect 23308 15014 23520 15042
rect 23296 14884 23348 14890
rect 23296 14826 23348 14832
rect 23202 14240 23258 14249
rect 23202 14175 23258 14184
rect 23202 14104 23258 14113
rect 23202 14039 23258 14048
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 23124 12306 23152 13126
rect 23216 12322 23244 14039
rect 23308 13841 23336 14826
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23294 13832 23350 13841
rect 23294 13767 23350 13776
rect 23400 12986 23428 14010
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23400 12782 23428 12922
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23492 12617 23520 15014
rect 23478 12608 23534 12617
rect 23478 12543 23534 12552
rect 23386 12336 23442 12345
rect 23112 12300 23164 12306
rect 23216 12294 23336 12322
rect 23112 12242 23164 12248
rect 23202 12200 23258 12209
rect 23202 12135 23258 12144
rect 23018 12064 23074 12073
rect 23018 11999 23074 12008
rect 22926 11384 22982 11393
rect 22926 11319 22982 11328
rect 22848 10934 22968 10962
rect 22834 10840 22890 10849
rect 22834 10775 22890 10784
rect 22848 10266 22876 10775
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 22742 8120 22798 8129
rect 22742 8055 22798 8064
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22664 7002 22692 7346
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22664 6662 22692 6734
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 22664 6458 22692 6598
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22560 6180 22612 6186
rect 22560 6122 22612 6128
rect 22572 5914 22600 6122
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22560 5568 22612 5574
rect 22560 5510 22612 5516
rect 22572 4146 22600 5510
rect 22756 5166 22784 7822
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22652 5092 22704 5098
rect 22652 5034 22704 5040
rect 22664 4826 22692 5034
rect 22652 4820 22704 4826
rect 22652 4762 22704 4768
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22664 4282 22692 4626
rect 22652 4276 22704 4282
rect 22652 4218 22704 4224
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22664 3602 22692 4218
rect 22848 4128 22876 10066
rect 22940 5846 22968 10934
rect 23032 7546 23060 11999
rect 23112 11620 23164 11626
rect 23112 11562 23164 11568
rect 23124 11121 23152 11562
rect 23110 11112 23166 11121
rect 23110 11047 23166 11056
rect 23124 7886 23152 11047
rect 23112 7880 23164 7886
rect 23112 7822 23164 7828
rect 23112 7744 23164 7750
rect 23112 7686 23164 7692
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23018 7440 23074 7449
rect 23124 7410 23152 7686
rect 23018 7375 23074 7384
rect 23112 7404 23164 7410
rect 22928 5840 22980 5846
rect 22928 5782 22980 5788
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 22940 5234 22968 5646
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 22940 4321 22968 5170
rect 22926 4312 22982 4321
rect 22926 4247 22982 4256
rect 23032 4146 23060 7375
rect 23112 7346 23164 7352
rect 23124 7206 23152 7346
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 23110 6352 23166 6361
rect 23110 6287 23166 6296
rect 23124 5914 23152 6287
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 23124 5302 23152 5646
rect 23112 5296 23164 5302
rect 23112 5238 23164 5244
rect 23124 4758 23152 5238
rect 23216 5098 23244 12135
rect 23308 8401 23336 12294
rect 23584 12322 23612 17478
rect 23664 16992 23716 16998
rect 23664 16934 23716 16940
rect 23676 14278 23704 16934
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23768 13716 23796 19246
rect 23860 14074 23888 19790
rect 23952 17105 23980 20295
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 26884 19168 26936 19174
rect 26884 19110 26936 19116
rect 24582 18864 24638 18873
rect 24582 18799 24584 18808
rect 24636 18799 24638 18808
rect 24584 18770 24636 18776
rect 24596 18714 24624 18770
rect 24596 18686 24716 18714
rect 24124 18624 24176 18630
rect 24124 18566 24176 18572
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 23938 17096 23994 17105
rect 23938 17031 23994 17040
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 23952 16046 23980 16730
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23952 15706 23980 15982
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 23952 14822 23980 15438
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23952 13938 23980 14214
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 23768 13688 23888 13716
rect 23860 12730 23888 13688
rect 23768 12702 23888 12730
rect 23584 12294 23704 12322
rect 23386 12271 23442 12280
rect 23400 12170 23428 12271
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 23388 12164 23440 12170
rect 23388 12106 23440 12112
rect 23584 12073 23612 12174
rect 23570 12064 23626 12073
rect 23570 11999 23626 12008
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 23400 10538 23428 11766
rect 23584 11694 23612 11999
rect 23572 11688 23624 11694
rect 23572 11630 23624 11636
rect 23676 11506 23704 12294
rect 23768 11676 23796 12702
rect 23938 12472 23994 12481
rect 23938 12407 23994 12416
rect 23848 12368 23900 12374
rect 23848 12310 23900 12316
rect 23860 11830 23888 12310
rect 23848 11824 23900 11830
rect 23848 11766 23900 11772
rect 23768 11648 23888 11676
rect 23584 11478 23704 11506
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 23388 10532 23440 10538
rect 23388 10474 23440 10480
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23294 8392 23350 8401
rect 23294 8327 23350 8336
rect 23400 8242 23428 9658
rect 23492 9178 23520 10678
rect 23584 10305 23612 11478
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23756 11008 23808 11014
rect 23756 10950 23808 10956
rect 23676 10606 23704 10950
rect 23768 10606 23796 10950
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23570 10296 23626 10305
rect 23570 10231 23626 10240
rect 23676 10130 23704 10542
rect 23768 10266 23796 10542
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 23570 10024 23626 10033
rect 23570 9959 23626 9968
rect 23584 9654 23612 9959
rect 23676 9722 23704 10066
rect 23754 10024 23810 10033
rect 23754 9959 23810 9968
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23584 9450 23612 9590
rect 23572 9444 23624 9450
rect 23572 9386 23624 9392
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23492 8430 23520 9114
rect 23768 9058 23796 9959
rect 23584 9030 23796 9058
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23400 8214 23520 8242
rect 23492 7426 23520 8214
rect 23584 7954 23612 9030
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23676 8634 23704 8910
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23662 8528 23718 8537
rect 23662 8463 23718 8472
rect 23676 8090 23704 8463
rect 23754 8392 23810 8401
rect 23754 8327 23810 8336
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23400 7398 23520 7426
rect 23400 7154 23428 7398
rect 23676 7342 23704 8026
rect 23664 7336 23716 7342
rect 23478 7304 23534 7313
rect 23664 7278 23716 7284
rect 23478 7239 23480 7248
rect 23532 7239 23534 7248
rect 23480 7210 23532 7216
rect 23400 7126 23704 7154
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23296 6384 23348 6390
rect 23296 6326 23348 6332
rect 23204 5092 23256 5098
rect 23204 5034 23256 5040
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 23124 4282 23152 4694
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 23020 4140 23072 4146
rect 22848 4100 22968 4128
rect 22836 4004 22888 4010
rect 22836 3946 22888 3952
rect 22848 3670 22876 3946
rect 22836 3664 22888 3670
rect 22836 3606 22888 3612
rect 22652 3596 22704 3602
rect 22652 3538 22704 3544
rect 22664 3126 22692 3538
rect 22848 3194 22876 3606
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 22652 3120 22704 3126
rect 22652 3062 22704 3068
rect 22650 2952 22706 2961
rect 22650 2887 22706 2896
rect 22664 2854 22692 2887
rect 22652 2848 22704 2854
rect 22480 2774 22600 2802
rect 22652 2790 22704 2796
rect 22374 2751 22430 2760
rect 21784 2536 21956 2564
rect 21732 2518 21784 2524
rect 21744 2378 21772 2518
rect 21732 2372 21784 2378
rect 21732 2314 21784 2320
rect 21822 606 21878 615
rect 21822 541 21878 550
rect 21836 480 21864 541
rect 22388 480 22416 2751
rect 22572 1630 22600 2774
rect 22940 2514 22968 4100
rect 23020 4082 23072 4088
rect 23018 4040 23074 4049
rect 23018 3975 23074 3984
rect 23308 3992 23336 6326
rect 23400 6322 23428 6802
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 23400 5370 23428 5782
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 23676 5114 23704 7126
rect 23768 5234 23796 8327
rect 23860 8022 23888 11648
rect 23952 8498 23980 12407
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23848 8016 23900 8022
rect 23848 7958 23900 7964
rect 24044 7698 24072 18022
rect 24136 17785 24164 18566
rect 24122 17776 24178 17785
rect 24122 17711 24178 17720
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24136 15065 24164 17070
rect 24122 15056 24178 15065
rect 24122 14991 24178 15000
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 24136 13734 24164 13806
rect 24124 13728 24176 13734
rect 24124 13670 24176 13676
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 24136 11762 24164 13126
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 24136 11354 24164 11698
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 24136 7954 24164 9590
rect 24228 8362 24256 18566
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18426 24716 18686
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24766 18320 24822 18329
rect 24766 18255 24822 18264
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 16998 24716 17682
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24676 15088 24728 15094
rect 24676 15030 24728 15036
rect 24308 14884 24360 14890
rect 24308 14826 24360 14832
rect 24320 14550 24348 14826
rect 24308 14544 24360 14550
rect 24308 14486 24360 14492
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 13530 24716 15030
rect 24780 14906 24808 18255
rect 25412 18080 25464 18086
rect 25412 18022 25464 18028
rect 24858 17640 24914 17649
rect 24858 17575 24914 17584
rect 24872 15065 24900 17575
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 25332 15910 25360 16594
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25056 15570 25084 15846
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 24952 15360 25004 15366
rect 24952 15302 25004 15308
rect 24858 15056 24914 15065
rect 24858 14991 24914 15000
rect 24780 14890 24900 14906
rect 24780 14884 24912 14890
rect 24780 14878 24860 14884
rect 24860 14826 24912 14832
rect 24766 14376 24822 14385
rect 24766 14311 24822 14320
rect 24676 13524 24728 13530
rect 24676 13466 24728 13472
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 24504 12442 24532 12786
rect 24688 12646 24716 13466
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24780 11898 24808 14311
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24872 12238 24900 14010
rect 24964 13870 24992 15302
rect 25056 15026 25084 15506
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25056 14618 25084 14962
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 25332 14550 25360 15846
rect 25320 14544 25372 14550
rect 25320 14486 25372 14492
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 24964 12850 24992 13806
rect 25056 13190 25084 14418
rect 25318 13968 25374 13977
rect 25318 13903 25374 13912
rect 25226 13832 25282 13841
rect 25226 13767 25282 13776
rect 25240 13394 25268 13767
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 25056 12986 25084 13126
rect 25240 12986 25268 13330
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25134 12880 25190 12889
rect 24952 12844 25004 12850
rect 25134 12815 25190 12824
rect 24952 12786 25004 12792
rect 25148 12424 25176 12815
rect 25226 12608 25282 12617
rect 25226 12543 25282 12552
rect 24964 12396 25176 12424
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24780 11558 24808 11834
rect 24964 11778 24992 12396
rect 25240 12374 25268 12543
rect 25228 12368 25280 12374
rect 25228 12310 25280 12316
rect 25332 12306 25360 13903
rect 25424 12628 25452 18022
rect 26054 17776 26110 17785
rect 26054 17711 26110 17720
rect 25780 17264 25832 17270
rect 25780 17206 25832 17212
rect 25594 15600 25650 15609
rect 25594 15535 25650 15544
rect 25504 12776 25556 12782
rect 25502 12744 25504 12753
rect 25556 12744 25558 12753
rect 25502 12679 25558 12688
rect 25424 12600 25544 12628
rect 25410 12336 25466 12345
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 25320 12300 25372 12306
rect 25410 12271 25466 12280
rect 25320 12242 25372 12248
rect 24872 11750 24992 11778
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24872 11370 24900 11750
rect 24780 11342 24900 11370
rect 25056 11354 25084 12242
rect 25424 11898 25452 12271
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 25410 11656 25466 11665
rect 25044 11348 25096 11354
rect 24674 10976 24730 10985
rect 24289 10908 24585 10928
rect 24674 10911 24730 10920
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10169 24716 10911
rect 24674 10160 24730 10169
rect 24674 10095 24730 10104
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24492 9580 24544 9586
rect 24492 9522 24544 9528
rect 24504 9178 24532 9522
rect 24584 9444 24636 9450
rect 24584 9386 24636 9392
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24596 8906 24624 9386
rect 24676 9036 24728 9042
rect 24676 8978 24728 8984
rect 24584 8900 24636 8906
rect 24584 8842 24636 8848
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24688 8634 24716 8978
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24674 8528 24730 8537
rect 24674 8463 24730 8472
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 24214 8256 24270 8265
rect 24214 8191 24270 8200
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 23952 7670 24072 7698
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23860 6934 23888 7414
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23846 6760 23902 6769
rect 23846 6695 23902 6704
rect 23860 5778 23888 6695
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 23860 5370 23888 5714
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23676 5086 23796 5114
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23492 4010 23520 4422
rect 23662 4176 23718 4185
rect 23662 4111 23718 4120
rect 23676 4078 23704 4111
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23480 4004 23532 4010
rect 22928 2508 22980 2514
rect 22928 2450 22980 2456
rect 22928 2304 22980 2310
rect 22928 2246 22980 2252
rect 22560 1624 22612 1630
rect 22560 1566 22612 1572
rect 22940 1465 22968 2246
rect 22926 1456 22982 1465
rect 22926 1391 22982 1400
rect 23032 480 23060 3975
rect 23308 3964 23428 3992
rect 23294 3768 23350 3777
rect 23294 3703 23350 3712
rect 23308 3505 23336 3703
rect 23294 3496 23350 3505
rect 23294 3431 23350 3440
rect 23400 2496 23428 3964
rect 23480 3946 23532 3952
rect 23478 3904 23534 3913
rect 23478 3839 23534 3848
rect 23492 3738 23520 3839
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23768 3670 23796 5086
rect 23572 3664 23624 3670
rect 23572 3606 23624 3612
rect 23756 3664 23808 3670
rect 23756 3606 23808 3612
rect 23480 2508 23532 2514
rect 23400 2468 23480 2496
rect 23480 2450 23532 2456
rect 23584 1737 23612 3606
rect 23952 3058 23980 7670
rect 24136 7546 24164 7890
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24032 6656 24084 6662
rect 24032 6598 24084 6604
rect 24044 6186 24072 6598
rect 24032 6180 24084 6186
rect 24032 6122 24084 6128
rect 24044 5914 24072 6122
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 24032 5908 24084 5914
rect 24032 5850 24084 5856
rect 24030 5808 24086 5817
rect 24030 5743 24086 5752
rect 24044 5114 24072 5743
rect 24136 5302 24164 6054
rect 24124 5296 24176 5302
rect 24124 5238 24176 5244
rect 24044 5086 24164 5114
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 24044 3233 24072 3334
rect 24030 3224 24086 3233
rect 24030 3159 24086 3168
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 23756 2984 23808 2990
rect 23754 2952 23756 2961
rect 23808 2952 23810 2961
rect 23754 2887 23810 2896
rect 23664 2440 23716 2446
rect 23662 2408 23664 2417
rect 23716 2408 23718 2417
rect 23662 2343 23718 2352
rect 23570 1728 23626 1737
rect 23570 1663 23626 1672
rect 23572 1624 23624 1630
rect 23572 1566 23624 1572
rect 23584 480 23612 1566
rect 24136 480 24164 5086
rect 24228 2582 24256 8191
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24584 5160 24636 5166
rect 24584 5102 24636 5108
rect 24596 4622 24624 5102
rect 24688 5001 24716 8463
rect 24780 8344 24808 11342
rect 25044 11290 25096 11296
rect 25240 11257 25268 11630
rect 25410 11591 25466 11600
rect 25424 11354 25452 11591
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 25226 11248 25282 11257
rect 25226 11183 25282 11192
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 25056 10130 25084 10406
rect 25134 10296 25190 10305
rect 25134 10231 25190 10240
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24964 9450 24992 9862
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 25056 9382 25084 10066
rect 25044 9376 25096 9382
rect 24950 9344 25006 9353
rect 25044 9318 25096 9324
rect 24950 9279 25006 9288
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24872 8634 24900 9114
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24964 8430 24992 9279
rect 25056 8974 25084 9318
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25148 8634 25176 10231
rect 25410 9616 25466 9625
rect 25410 9551 25466 9560
rect 25318 9072 25374 9081
rect 25318 9007 25374 9016
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24780 8316 24900 8344
rect 24766 8256 24822 8265
rect 24766 8191 24822 8200
rect 24780 5370 24808 8191
rect 24872 8072 24900 8316
rect 24872 8044 25084 8072
rect 24950 7984 25006 7993
rect 24950 7919 25006 7928
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24674 4992 24730 5001
rect 24674 4927 24730 4936
rect 24584 4616 24636 4622
rect 24582 4584 24584 4593
rect 24636 4584 24638 4593
rect 24582 4519 24638 4528
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24492 3120 24544 3126
rect 24490 3088 24492 3097
rect 24544 3088 24546 3097
rect 24490 3023 24546 3032
rect 24216 2576 24268 2582
rect 24216 2518 24268 2524
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24780 480 24808 5170
rect 24872 4146 24900 5646
rect 24964 4690 24992 7919
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 24964 4282 24992 4626
rect 24952 4276 25004 4282
rect 24952 4218 25004 4224
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24950 3768 25006 3777
rect 24950 3703 25006 3712
rect 24858 3496 24914 3505
rect 24858 3431 24860 3440
rect 24912 3431 24914 3440
rect 24860 3402 24912 3408
rect 24964 3194 24992 3703
rect 25056 3602 25084 8044
rect 25226 7576 25282 7585
rect 25226 7511 25282 7520
rect 25134 5672 25190 5681
rect 25134 5607 25190 5616
rect 25148 3942 25176 5607
rect 25240 4826 25268 7511
rect 25332 7154 25360 9007
rect 25424 7546 25452 9551
rect 25516 9110 25544 12600
rect 25608 11830 25636 15535
rect 25686 13016 25742 13025
rect 25686 12951 25688 12960
rect 25740 12951 25742 12960
rect 25688 12922 25740 12928
rect 25596 11824 25648 11830
rect 25596 11766 25648 11772
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25608 10470 25636 11154
rect 25686 10568 25742 10577
rect 25686 10503 25742 10512
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25608 10033 25636 10406
rect 25594 10024 25650 10033
rect 25594 9959 25650 9968
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 25502 8936 25558 8945
rect 25502 8871 25558 8880
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25332 7126 25452 7154
rect 25318 7032 25374 7041
rect 25318 6967 25374 6976
rect 25332 6730 25360 6967
rect 25320 6724 25372 6730
rect 25320 6666 25372 6672
rect 25318 6352 25374 6361
rect 25318 6287 25374 6296
rect 25228 4820 25280 4826
rect 25228 4762 25280 4768
rect 25228 4004 25280 4010
rect 25228 3946 25280 3952
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 25044 3596 25096 3602
rect 25044 3538 25096 3544
rect 25056 3194 25084 3538
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 24964 2990 24992 3130
rect 24952 2984 25004 2990
rect 24952 2926 25004 2932
rect 25134 2544 25190 2553
rect 25134 2479 25136 2488
rect 25188 2479 25190 2488
rect 25136 2450 25188 2456
rect 25044 2440 25096 2446
rect 25042 2408 25044 2417
rect 25096 2408 25098 2417
rect 25042 2343 25098 2352
rect 25240 1873 25268 3946
rect 25332 3738 25360 6287
rect 25424 5778 25452 7126
rect 25516 5914 25544 8871
rect 25596 6860 25648 6866
rect 25596 6802 25648 6808
rect 25608 6254 25636 6802
rect 25596 6248 25648 6254
rect 25594 6216 25596 6225
rect 25648 6216 25650 6225
rect 25594 6151 25650 6160
rect 25504 5908 25556 5914
rect 25504 5850 25556 5856
rect 25412 5772 25464 5778
rect 25412 5714 25464 5720
rect 25424 5370 25452 5714
rect 25412 5364 25464 5370
rect 25412 5306 25464 5312
rect 25594 5264 25650 5273
rect 25594 5199 25650 5208
rect 25410 5128 25466 5137
rect 25410 5063 25466 5072
rect 25424 3738 25452 5063
rect 25608 4826 25636 5199
rect 25596 4820 25648 4826
rect 25596 4762 25648 4768
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25412 3732 25464 3738
rect 25412 3674 25464 3680
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25226 1864 25282 1873
rect 25226 1799 25282 1808
rect 25332 480 25360 3538
rect 25700 3058 25728 10503
rect 25792 8537 25820 17206
rect 25964 16788 26016 16794
rect 25964 16730 26016 16736
rect 25870 15736 25926 15745
rect 25870 15671 25926 15680
rect 25778 8528 25834 8537
rect 25778 8463 25834 8472
rect 25884 5409 25912 15671
rect 25870 5400 25926 5409
rect 25870 5335 25926 5344
rect 25976 3602 26004 16730
rect 25964 3596 26016 3602
rect 25964 3538 26016 3544
rect 25780 3392 25832 3398
rect 25780 3334 25832 3340
rect 25688 3052 25740 3058
rect 25688 2994 25740 3000
rect 25504 2304 25556 2310
rect 25504 2246 25556 2252
rect 25516 1601 25544 2246
rect 25502 1592 25558 1601
rect 25502 1527 25558 1536
rect 25792 1329 25820 3334
rect 26068 2122 26096 17711
rect 26330 15464 26386 15473
rect 26330 15399 26386 15408
rect 26238 13696 26294 13705
rect 26238 13631 26294 13640
rect 26148 13184 26200 13190
rect 26148 13126 26200 13132
rect 26160 5817 26188 13126
rect 26252 9178 26280 13631
rect 26344 9330 26372 15399
rect 26344 9302 26556 9330
rect 26330 9208 26386 9217
rect 26240 9172 26292 9178
rect 26330 9143 26386 9152
rect 26240 9114 26292 9120
rect 26146 5808 26202 5817
rect 26146 5743 26202 5752
rect 26240 3936 26292 3942
rect 26240 3878 26292 3884
rect 26252 3641 26280 3878
rect 26238 3632 26294 3641
rect 26238 3567 26294 3576
rect 26240 2984 26292 2990
rect 26238 2952 26240 2961
rect 26292 2952 26294 2961
rect 26238 2887 26294 2896
rect 25884 2094 26096 2122
rect 25778 1320 25834 1329
rect 25778 1255 25834 1264
rect 25884 480 25912 2094
rect 9954 368 10010 377
rect 9954 303 10010 312
rect 10138 0 10194 480
rect 10782 0 10838 480
rect 11334 0 11390 480
rect 11886 0 11942 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14278 0 14334 480
rect 14830 0 14886 480
rect 15382 0 15438 480
rect 16026 0 16082 480
rect 16578 0 16634 480
rect 17130 0 17186 480
rect 17774 0 17830 480
rect 18326 0 18382 480
rect 18878 0 18934 480
rect 19522 0 19578 480
rect 20074 0 20130 480
rect 20626 0 20682 480
rect 21270 0 21326 480
rect 21822 0 21878 480
rect 22374 0 22430 480
rect 23018 0 23074 480
rect 23570 0 23626 480
rect 24122 0 24178 480
rect 24766 0 24822 480
rect 25318 0 25374 480
rect 25870 0 25926 480
rect 26344 377 26372 9143
rect 26424 9104 26476 9110
rect 26424 9046 26476 9052
rect 26436 2961 26464 9046
rect 26422 2952 26478 2961
rect 26422 2887 26478 2896
rect 26528 480 26556 9302
rect 26792 8356 26844 8362
rect 26792 8298 26844 8304
rect 26804 2281 26832 8298
rect 26896 4842 26924 19110
rect 27618 5400 27674 5409
rect 27618 5335 27674 5344
rect 26896 4814 27108 4842
rect 26790 2272 26846 2281
rect 26790 2207 26846 2216
rect 27080 480 27108 4814
rect 27632 480 27660 5335
rect 26330 368 26386 377
rect 26330 303 26386 312
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 2778 27648 2834 27704
rect 23478 27648 23534 27704
rect 2226 26288 2282 26344
rect 2042 18028 2044 18048
rect 2044 18028 2096 18048
rect 2096 18028 2098 18048
rect 2042 17992 2098 18028
rect 2042 17620 2044 17640
rect 2044 17620 2096 17640
rect 2096 17620 2098 17640
rect 2042 17584 2098 17620
rect 1122 14728 1178 14784
rect 754 12008 810 12064
rect 662 10648 718 10704
rect 294 10240 350 10296
rect 2042 16788 2098 16824
rect 2042 16768 2044 16788
rect 2044 16768 2096 16788
rect 2096 16768 2098 16788
rect 2042 16108 2098 16144
rect 2042 16088 2044 16108
rect 2044 16088 2096 16108
rect 2096 16088 2098 16108
rect 1582 14320 1638 14376
rect 1398 14220 1400 14240
rect 1400 14220 1452 14240
rect 1452 14220 1454 14240
rect 1398 14184 1454 14220
rect 1674 13912 1730 13968
rect 1398 11092 1400 11112
rect 1400 11092 1452 11112
rect 1452 11092 1454 11112
rect 1398 11056 1454 11092
rect 2042 14884 2098 14920
rect 2042 14864 2044 14884
rect 2044 14864 2096 14884
rect 2096 14864 2098 14884
rect 1858 12552 1914 12608
rect 1490 8064 1546 8120
rect 1398 7928 1454 7984
rect 1858 12280 1914 12336
rect 2042 12144 2098 12200
rect 1950 11192 2006 11248
rect 1674 8744 1730 8800
rect 1582 6704 1638 6760
rect 1858 8608 1914 8664
rect 1950 8336 2006 8392
rect 1766 6860 1822 6896
rect 1766 6840 1768 6860
rect 1768 6840 1820 6860
rect 1820 6840 1822 6860
rect 1674 6024 1730 6080
rect 1490 3884 1492 3904
rect 1492 3884 1544 3904
rect 1544 3884 1546 3904
rect 1490 3848 1546 3884
rect 1674 2916 1730 2952
rect 1674 2896 1676 2916
rect 1676 2896 1728 2916
rect 1728 2896 1730 2916
rect 2502 17740 2558 17776
rect 2502 17720 2504 17740
rect 2504 17720 2556 17740
rect 2556 17720 2558 17740
rect 2226 16224 2282 16280
rect 2502 15680 2558 15736
rect 2410 12960 2466 13016
rect 3422 26968 3478 27024
rect 3054 25608 3110 25664
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 4526 25064 4582 25120
rect 3974 20440 4030 20496
rect 3790 19760 3846 19816
rect 3238 19080 3294 19136
rect 3146 16940 3148 16960
rect 3148 16940 3200 16960
rect 3200 16940 3202 16960
rect 3146 16904 3202 16940
rect 2962 15544 3018 15600
rect 2778 15272 2834 15328
rect 2594 14456 2650 14512
rect 2502 12008 2558 12064
rect 2318 11620 2374 11656
rect 2318 11600 2320 11620
rect 2320 11600 2372 11620
rect 2372 11600 2374 11620
rect 2226 11328 2282 11384
rect 2410 10512 2466 10568
rect 2318 10376 2374 10432
rect 2134 9968 2190 10024
rect 3054 14592 3110 14648
rect 2502 9016 2558 9072
rect 2318 8064 2374 8120
rect 2410 7792 2466 7848
rect 2226 7248 2282 7304
rect 2318 6704 2374 6760
rect 2134 4256 2190 4312
rect 2594 7384 2650 7440
rect 2962 10920 3018 10976
rect 3882 17856 3938 17912
rect 3790 16496 3846 16552
rect 3698 16360 3754 16416
rect 3790 15816 3846 15872
rect 3330 15680 3386 15736
rect 3698 15680 3754 15736
rect 3422 15272 3478 15328
rect 3330 13932 3386 13968
rect 3330 13912 3332 13932
rect 3332 13912 3384 13932
rect 3384 13912 3386 13932
rect 3330 12280 3386 12336
rect 3790 14864 3846 14920
rect 4434 16652 4490 16688
rect 4434 16632 4436 16652
rect 4436 16632 4488 16652
rect 4488 16632 4490 16652
rect 4066 15816 4122 15872
rect 3974 15680 4030 15736
rect 3882 14592 3938 14648
rect 3790 14320 3846 14376
rect 3606 12552 3662 12608
rect 2870 9424 2926 9480
rect 2962 8200 3018 8256
rect 3054 6024 3110 6080
rect 2502 5208 2558 5264
rect 3698 12280 3754 12336
rect 3698 11328 3754 11384
rect 4434 15816 4490 15872
rect 4066 14184 4122 14240
rect 3974 13912 4030 13968
rect 4158 13368 4214 13424
rect 4066 12144 4122 12200
rect 3882 11192 3938 11248
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 7102 24384 7158 24440
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6826 21120 6882 21176
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 6826 18536 6882 18592
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6366 16768 6422 16824
rect 4526 12416 4582 12472
rect 4342 12144 4398 12200
rect 4066 11192 4122 11248
rect 3790 10240 3846 10296
rect 3698 8472 3754 8528
rect 3698 7792 3754 7848
rect 3514 7520 3570 7576
rect 2778 5344 2834 5400
rect 3146 5344 3202 5400
rect 2962 5072 3018 5128
rect 2778 4800 2834 4856
rect 2134 2524 2136 2544
rect 2136 2524 2188 2544
rect 2188 2524 2190 2544
rect 2134 2488 2190 2524
rect 2502 3712 2558 3768
rect 2502 2252 2504 2272
rect 2504 2252 2556 2272
rect 2556 2252 2558 2272
rect 2502 2216 2558 2252
rect 2226 1400 2282 1456
rect 3054 4664 3110 4720
rect 3054 3032 3110 3088
rect 3790 6432 3846 6488
rect 3698 5072 3754 5128
rect 3974 7112 4030 7168
rect 4250 10648 4306 10704
rect 4158 5888 4214 5944
rect 3974 5480 4030 5536
rect 3882 4936 3938 4992
rect 3790 4120 3846 4176
rect 3422 3440 3478 3496
rect 3974 3440 4030 3496
rect 4066 2624 4122 2680
rect 3698 2080 3754 2136
rect 2962 1672 3018 1728
rect 4066 1944 4122 2000
rect 4526 9444 4582 9480
rect 4526 9424 4528 9444
rect 4528 9424 4580 9444
rect 4580 9424 4582 9444
rect 5446 16360 5502 16416
rect 5998 16360 6054 16416
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 4894 15272 4950 15328
rect 4986 14764 4988 14784
rect 4988 14764 5040 14784
rect 5040 14764 5042 14784
rect 4986 14728 5042 14764
rect 5262 15408 5318 15464
rect 5446 15408 5502 15464
rect 4986 14456 5042 14512
rect 5446 14728 5502 14784
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5998 14320 6054 14376
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5722 13504 5778 13560
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5998 12960 6054 13016
rect 4986 12824 5042 12880
rect 5722 12144 5778 12200
rect 4802 11736 4858 11792
rect 4802 11056 4858 11112
rect 4710 9988 4766 10024
rect 4710 9968 4712 9988
rect 4712 9968 4764 9988
rect 4764 9968 4766 9988
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5906 11500 5908 11520
rect 5908 11500 5960 11520
rect 5960 11500 5962 11520
rect 5906 11464 5962 11500
rect 5814 11328 5870 11384
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5446 10376 5502 10432
rect 5354 10240 5410 10296
rect 5262 9832 5318 9888
rect 5170 9288 5226 9344
rect 5078 9152 5134 9208
rect 4434 6024 4490 6080
rect 5262 8880 5318 8936
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5446 8608 5502 8664
rect 5354 8336 5410 8392
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5722 8356 5778 8392
rect 5722 8336 5724 8356
rect 5724 8336 5776 8356
rect 5776 8336 5778 8356
rect 5998 7928 6054 7984
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5262 6296 5318 6352
rect 4618 5616 4674 5672
rect 4618 3712 4674 3768
rect 4802 2216 4858 2272
rect 4986 4800 5042 4856
rect 5170 5344 5226 5400
rect 5538 7248 5594 7304
rect 5630 6840 5686 6896
rect 6182 12316 6184 12336
rect 6184 12316 6236 12336
rect 6236 12316 6238 12336
rect 6182 12280 6238 12316
rect 6734 13912 6790 13968
rect 6734 13776 6790 13832
rect 6642 12280 6698 12336
rect 6274 6996 6330 7032
rect 6274 6976 6276 6996
rect 6276 6976 6328 6996
rect 6328 6976 6330 6996
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5998 6432 6054 6488
rect 5722 6180 5778 6216
rect 5722 6160 5724 6180
rect 5724 6160 5776 6180
rect 5776 6160 5778 6180
rect 6182 5888 6238 5944
rect 6458 6160 6514 6216
rect 6090 5752 6146 5808
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 6090 5480 6146 5536
rect 5446 4120 5502 4176
rect 5354 2624 5410 2680
rect 6458 5888 6514 5944
rect 6642 11600 6698 11656
rect 6642 9968 6698 10024
rect 7010 12588 7012 12608
rect 7012 12588 7064 12608
rect 7064 12588 7066 12608
rect 7010 12552 7066 12588
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 7562 18264 7618 18320
rect 7470 16496 7526 16552
rect 7378 15952 7434 16008
rect 7194 14612 7250 14648
rect 7194 14592 7196 14612
rect 7196 14592 7248 14612
rect 7248 14592 7250 14612
rect 7286 14340 7342 14376
rect 7286 14320 7288 14340
rect 7288 14320 7340 14340
rect 7340 14320 7342 14340
rect 6918 11056 6974 11112
rect 6642 8744 6698 8800
rect 6918 9172 6974 9208
rect 6918 9152 6920 9172
rect 6920 9152 6972 9172
rect 6972 9152 6974 9172
rect 6918 8472 6974 8528
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10322 17720 10378 17776
rect 9862 17584 9918 17640
rect 9678 15680 9734 15736
rect 7470 13368 7526 13424
rect 7378 10784 7434 10840
rect 7102 7112 7158 7168
rect 7286 10104 7342 10160
rect 7654 11872 7710 11928
rect 7838 13232 7894 13288
rect 7838 11736 7894 11792
rect 8022 12008 8078 12064
rect 8022 11192 8078 11248
rect 8022 10648 8078 10704
rect 8298 12960 8354 13016
rect 8390 11636 8392 11656
rect 8392 11636 8444 11656
rect 8444 11636 8446 11656
rect 8390 11600 8446 11636
rect 8206 10684 8208 10704
rect 8208 10684 8260 10704
rect 8260 10684 8262 10704
rect 8206 10648 8262 10684
rect 7286 7384 7342 7440
rect 7010 5344 7066 5400
rect 5722 4528 5778 4584
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6090 3984 6146 4040
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5722 3032 5778 3088
rect 5998 2216 6054 2272
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5998 2080 6054 2136
rect 5262 1808 5318 1864
rect 5998 1536 6054 1592
rect 6274 3304 6330 3360
rect 6458 3712 6514 3768
rect 6734 3848 6790 3904
rect 6642 2508 6698 2544
rect 6642 2488 6644 2508
rect 6644 2488 6696 2508
rect 6696 2488 6698 2508
rect 7838 8744 7894 8800
rect 7654 8084 7710 8120
rect 7654 8064 7656 8084
rect 7656 8064 7708 8084
rect 7708 8064 7710 8084
rect 7470 6724 7526 6760
rect 7470 6704 7472 6724
rect 7472 6704 7524 6724
rect 7524 6704 7526 6724
rect 8114 9832 8170 9888
rect 8206 9696 8262 9752
rect 8574 13776 8630 13832
rect 8574 13368 8630 13424
rect 8574 12960 8630 13016
rect 8574 12164 8630 12200
rect 8574 12144 8576 12164
rect 8576 12144 8628 12164
rect 8628 12144 8630 12164
rect 8666 9988 8722 10024
rect 8666 9968 8668 9988
rect 8668 9968 8720 9988
rect 8720 9968 8722 9988
rect 9770 14728 9826 14784
rect 9126 9832 9182 9888
rect 9770 13776 9826 13832
rect 9310 13504 9366 13560
rect 9586 12824 9642 12880
rect 9586 12416 9642 12472
rect 11058 17176 11114 17232
rect 10046 17040 10102 17096
rect 10322 17040 10378 17096
rect 9770 11076 9826 11112
rect 9770 11056 9772 11076
rect 9772 11056 9824 11076
rect 9824 11056 9826 11076
rect 9678 10412 9680 10432
rect 9680 10412 9732 10432
rect 9732 10412 9734 10432
rect 9678 10376 9734 10412
rect 9494 10240 9550 10296
rect 9218 9696 9274 9752
rect 9034 9052 9036 9072
rect 9036 9052 9088 9072
rect 9088 9052 9090 9072
rect 9034 9016 9090 9052
rect 8114 7520 8170 7576
rect 8482 7948 8538 7984
rect 8482 7928 8484 7948
rect 8484 7928 8536 7948
rect 8536 7928 8538 7948
rect 8390 7656 8446 7712
rect 8206 6296 8262 6352
rect 7746 4392 7802 4448
rect 7930 4256 7986 4312
rect 8482 5752 8538 5808
rect 8574 5636 8630 5672
rect 8574 5616 8576 5636
rect 8576 5616 8628 5636
rect 8628 5616 8630 5636
rect 8482 4936 8538 4992
rect 8114 4392 8170 4448
rect 7286 3576 7342 3632
rect 6642 2216 6698 2272
rect 6366 1536 6422 1592
rect 7562 856 7618 912
rect 8298 3848 8354 3904
rect 8574 4700 8576 4720
rect 8576 4700 8628 4720
rect 8628 4700 8630 4720
rect 8574 4664 8630 4700
rect 8574 4256 8630 4312
rect 9218 8200 9274 8256
rect 8850 8064 8906 8120
rect 9402 7792 9458 7848
rect 8758 6296 8814 6352
rect 8942 6024 8998 6080
rect 9678 8880 9734 8936
rect 9770 8472 9826 8528
rect 9678 8372 9680 8392
rect 9680 8372 9732 8392
rect 9732 8372 9734 8392
rect 9678 8336 9734 8372
rect 9954 9424 10010 9480
rect 9954 8880 10010 8936
rect 9954 8608 10010 8664
rect 9770 8064 9826 8120
rect 9862 7692 9864 7712
rect 9864 7692 9916 7712
rect 9916 7692 9918 7712
rect 9862 7656 9918 7692
rect 9126 7248 9182 7304
rect 9034 5480 9090 5536
rect 8114 3032 8170 3088
rect 8482 3304 8538 3360
rect 8666 1944 8722 2000
rect 9678 7112 9734 7168
rect 9218 6976 9274 7032
rect 9494 5636 9550 5672
rect 9494 5616 9496 5636
rect 9496 5616 9548 5636
rect 9548 5616 9550 5636
rect 9402 5072 9458 5128
rect 9770 4664 9826 4720
rect 9586 4004 9642 4040
rect 9586 3984 9588 4004
rect 9588 3984 9640 4004
rect 9640 3984 9642 4004
rect 9586 3712 9642 3768
rect 9310 2760 9366 2816
rect 9126 2644 9182 2680
rect 9126 2624 9128 2644
rect 9128 2624 9180 2644
rect 9180 2624 9182 2644
rect 9126 2216 9182 2272
rect 9126 1808 9182 1864
rect 9862 2080 9918 2136
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10782 15136 10838 15192
rect 11058 14864 11114 14920
rect 10874 14048 10930 14104
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10690 12688 10746 12744
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10138 11328 10194 11384
rect 14278 23704 14334 23760
rect 13358 18808 13414 18864
rect 12530 18536 12586 18592
rect 11794 15000 11850 15056
rect 11334 12588 11336 12608
rect 11336 12588 11388 12608
rect 11388 12588 11390 12608
rect 11334 12552 11390 12588
rect 10138 11056 10194 11112
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10138 9832 10194 9888
rect 10230 9696 10286 9752
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10782 9832 10838 9888
rect 10874 9596 10876 9616
rect 10876 9596 10928 9616
rect 10928 9596 10930 9616
rect 10874 9560 10930 9596
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10690 7112 10746 7168
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 11334 9324 11336 9344
rect 11336 9324 11388 9344
rect 11388 9324 11390 9344
rect 11334 9288 11390 9324
rect 11150 7520 11206 7576
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10782 5616 10838 5672
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10138 4800 10194 4856
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 11150 4428 11152 4448
rect 11152 4428 11204 4448
rect 11204 4428 11206 4448
rect 11150 4392 11206 4428
rect 10782 3440 10838 3496
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10138 2488 10194 2544
rect 11242 3304 11298 3360
rect 11150 2896 11206 2952
rect 10782 2216 10838 2272
rect 12070 11328 12126 11384
rect 11610 8064 11666 8120
rect 11702 4120 11758 4176
rect 11702 1400 11758 1456
rect 12254 10920 12310 10976
rect 12162 10648 12218 10704
rect 12898 15408 12954 15464
rect 12714 14864 12770 14920
rect 12714 14356 12716 14376
rect 12716 14356 12768 14376
rect 12768 14356 12770 14376
rect 12714 14320 12770 14356
rect 12714 13776 12770 13832
rect 12070 5208 12126 5264
rect 12622 8336 12678 8392
rect 12530 8200 12586 8256
rect 12438 7928 12494 7984
rect 12254 7248 12310 7304
rect 12990 15136 13046 15192
rect 12990 9832 13046 9888
rect 12990 9696 13046 9752
rect 13266 11192 13322 11248
rect 13266 10784 13322 10840
rect 14002 15000 14058 15056
rect 14278 18672 14334 18728
rect 13450 10240 13506 10296
rect 13358 9696 13414 9752
rect 13174 9560 13230 9616
rect 12530 5616 12586 5672
rect 12346 3576 12402 3632
rect 12990 5888 13046 5944
rect 12898 3032 12954 3088
rect 12806 2372 12862 2408
rect 12806 2352 12808 2372
rect 12808 2352 12860 2372
rect 12860 2352 12862 2372
rect 12990 1264 13046 1320
rect 13450 8472 13506 8528
rect 13726 6840 13782 6896
rect 13358 6296 13414 6352
rect 13818 6568 13874 6624
rect 13726 5636 13782 5672
rect 13726 5616 13728 5636
rect 13728 5616 13780 5636
rect 13780 5616 13782 5636
rect 14094 12280 14150 12336
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14738 22480 14794 22536
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15566 15544 15622 15600
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14462 13096 14518 13152
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14738 12844 14794 12880
rect 14738 12824 14740 12844
rect 14740 12824 14792 12844
rect 14792 12824 14794 12844
rect 14002 9152 14058 9208
rect 14002 8472 14058 8528
rect 14186 8336 14242 8392
rect 14278 5480 14334 5536
rect 14370 5344 14426 5400
rect 14278 5244 14280 5264
rect 14280 5244 14332 5264
rect 14332 5244 14334 5264
rect 14278 5208 14334 5244
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15198 11736 15254 11792
rect 15198 11464 15254 11520
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14554 9288 14610 9344
rect 14370 4256 14426 4312
rect 14830 10104 14886 10160
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14830 9560 14886 9616
rect 14738 8064 14794 8120
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15566 11600 15622 11656
rect 15658 10784 15714 10840
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20258 24248 20314 24304
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 16118 20304 16174 20360
rect 15842 11328 15898 11384
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15382 8200 15438 8256
rect 16026 10532 16082 10568
rect 16026 10512 16028 10532
rect 16028 10512 16080 10532
rect 16080 10512 16082 10532
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 16486 19760 16542 19816
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 16854 17176 16910 17232
rect 16210 16088 16266 16144
rect 16486 16088 16542 16144
rect 16302 15000 16358 15056
rect 16302 14320 16358 14376
rect 17314 16496 17370 16552
rect 17314 15408 17370 15464
rect 16854 9424 16910 9480
rect 16118 9152 16174 9208
rect 15934 8608 15990 8664
rect 15842 8200 15898 8256
rect 15474 6432 15530 6488
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15290 4800 15346 4856
rect 15474 4800 15530 4856
rect 14646 4528 14702 4584
rect 15106 4528 15162 4584
rect 14370 3576 14426 3632
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 13910 2372 13966 2408
rect 13910 2352 13912 2372
rect 13912 2352 13964 2372
rect 13964 2352 13966 2372
rect 13634 2252 13636 2272
rect 13636 2252 13688 2272
rect 13688 2252 13690 2272
rect 13634 2216 13690 2252
rect 14186 1672 14242 1728
rect 13634 856 13690 912
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15658 3984 15714 4040
rect 15934 8064 15990 8120
rect 16302 9036 16358 9072
rect 16302 9016 16304 9036
rect 16304 9016 16356 9036
rect 16356 9016 16358 9036
rect 16302 7828 16304 7848
rect 16304 7828 16356 7848
rect 16356 7828 16358 7848
rect 16302 7792 16358 7828
rect 16118 7540 16174 7576
rect 16118 7520 16120 7540
rect 16120 7520 16172 7540
rect 16172 7520 16174 7540
rect 15842 6160 15898 6216
rect 16486 7248 16542 7304
rect 16670 8900 16726 8936
rect 16670 8880 16672 8900
rect 16672 8880 16724 8900
rect 16724 8880 16726 8900
rect 16854 8880 16910 8936
rect 16762 7384 16818 7440
rect 16578 6296 16634 6352
rect 17038 8336 17094 8392
rect 17406 9968 17462 10024
rect 17774 12708 17830 12744
rect 17774 12688 17776 12708
rect 17776 12688 17828 12708
rect 17828 12688 17830 12708
rect 17498 7964 17500 7984
rect 17500 7964 17552 7984
rect 17552 7964 17554 7984
rect 17498 7928 17554 7964
rect 18050 11636 18052 11656
rect 18052 11636 18104 11656
rect 18104 11636 18106 11656
rect 18050 11600 18106 11636
rect 18050 11464 18106 11520
rect 18050 11192 18106 11248
rect 18326 13912 18382 13968
rect 18326 13812 18328 13832
rect 18328 13812 18380 13832
rect 18380 13812 18382 13832
rect 18326 13776 18382 13812
rect 18602 13640 18658 13696
rect 18602 13232 18658 13288
rect 18418 12552 18474 12608
rect 17682 6976 17738 7032
rect 18050 6296 18106 6352
rect 17314 6160 17370 6216
rect 16486 5616 16542 5672
rect 17130 5616 17186 5672
rect 15750 3168 15806 3224
rect 15382 1672 15438 1728
rect 16486 3712 16542 3768
rect 16578 2760 16634 2816
rect 16026 2524 16028 2544
rect 16028 2524 16080 2544
rect 16080 2524 16082 2544
rect 16026 2488 16082 2524
rect 15842 1400 15898 1456
rect 16946 2080 17002 2136
rect 17130 1536 17186 1592
rect 16946 1400 17002 1456
rect 17130 1400 17186 1456
rect 18050 5108 18052 5128
rect 18052 5108 18104 5128
rect 18104 5108 18106 5128
rect 18050 5072 18106 5108
rect 18234 8200 18290 8256
rect 18234 7792 18290 7848
rect 17774 3188 17830 3224
rect 17774 3168 17776 3188
rect 17776 3168 17828 3188
rect 17828 3168 17830 3188
rect 18142 3304 18198 3360
rect 17774 2896 17830 2952
rect 17314 1944 17370 2000
rect 17222 1128 17278 1184
rect 18878 12708 18934 12744
rect 18878 12688 18880 12708
rect 18880 12688 18932 12708
rect 18932 12688 18934 12708
rect 19430 15000 19486 15056
rect 18786 9560 18842 9616
rect 18694 9424 18750 9480
rect 19338 12824 19394 12880
rect 18878 8472 18934 8528
rect 19062 7112 19118 7168
rect 18786 5480 18842 5536
rect 18510 4936 18566 4992
rect 18326 3984 18382 4040
rect 18878 4392 18934 4448
rect 18418 3168 18474 3224
rect 18234 2624 18290 2680
rect 18786 2388 18788 2408
rect 18788 2388 18840 2408
rect 18840 2388 18842 2408
rect 18786 2352 18842 2388
rect 18326 1536 18382 1592
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 20074 23296 20130 23352
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 20074 15136 20130 15192
rect 19890 14048 19946 14104
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19706 8780 19708 8800
rect 19708 8780 19760 8800
rect 19760 8780 19762 8800
rect 19706 8744 19762 8780
rect 20350 21528 20406 21584
rect 21178 17040 21234 17096
rect 20350 15952 20406 16008
rect 20442 15680 20498 15736
rect 20074 10548 20076 10568
rect 20076 10548 20128 10568
rect 20128 10548 20130 10568
rect 20074 10512 20130 10548
rect 20074 9560 20130 9616
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19338 6976 19394 7032
rect 19338 4664 19394 4720
rect 19154 4120 19210 4176
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19522 3984 19578 4040
rect 19430 3712 19486 3768
rect 19338 2760 19394 2816
rect 19430 2488 19486 2544
rect 19062 856 19118 912
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20074 7656 20130 7712
rect 20166 7112 20222 7168
rect 20626 15852 20628 15872
rect 20628 15852 20680 15872
rect 20680 15852 20682 15872
rect 20626 15816 20682 15852
rect 21086 15408 21142 15464
rect 20810 12416 20866 12472
rect 21454 15816 21510 15872
rect 21270 12300 21326 12336
rect 21270 12280 21272 12300
rect 21272 12280 21324 12300
rect 21324 12280 21326 12300
rect 20902 11872 20958 11928
rect 20718 11600 20774 11656
rect 20810 11192 20866 11248
rect 20626 10240 20682 10296
rect 20442 7520 20498 7576
rect 20350 6976 20406 7032
rect 20442 5616 20498 5672
rect 20166 4800 20222 4856
rect 20074 4664 20130 4720
rect 19706 3068 19708 3088
rect 19708 3068 19760 3088
rect 19760 3068 19762 3088
rect 19706 3032 19762 3068
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20166 4256 20222 4312
rect 20258 3848 20314 3904
rect 21086 10648 21142 10704
rect 20810 9696 20866 9752
rect 20810 9560 20866 9616
rect 20994 9832 21050 9888
rect 20810 8880 20866 8936
rect 20810 8608 20866 8664
rect 20718 6860 20774 6896
rect 20718 6840 20720 6860
rect 20720 6840 20772 6860
rect 20772 6840 20774 6860
rect 20902 7248 20958 7304
rect 20994 5888 21050 5944
rect 21086 4664 21142 4720
rect 21178 2216 21234 2272
rect 20994 2080 21050 2136
rect 20902 1808 20958 1864
rect 21362 9152 21418 9208
rect 21362 8336 21418 8392
rect 21730 9968 21786 10024
rect 21730 9832 21786 9888
rect 21638 9016 21694 9072
rect 21546 8336 21602 8392
rect 21546 5480 21602 5536
rect 21914 13368 21970 13424
rect 21822 9560 21878 9616
rect 21822 8744 21878 8800
rect 23570 26968 23626 27024
rect 23478 26308 23534 26344
rect 23478 26288 23480 26308
rect 23480 26288 23532 26308
rect 23532 26288 23534 26308
rect 22098 13948 22100 13968
rect 22100 13948 22152 13968
rect 22152 13948 22154 13968
rect 22098 13912 22154 13948
rect 23478 25608 23534 25664
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 23202 23024 23258 23080
rect 22926 22072 22982 22128
rect 22282 16632 22338 16688
rect 22098 12280 22154 12336
rect 22742 17584 22798 17640
rect 22098 11736 22154 11792
rect 22374 11736 22430 11792
rect 22742 16632 22798 16688
rect 22374 11328 22430 11384
rect 22282 9832 22338 9888
rect 22466 9288 22522 9344
rect 22190 7384 22246 7440
rect 22282 5888 22338 5944
rect 22374 4428 22376 4448
rect 22376 4428 22428 4448
rect 22428 4428 22430 4448
rect 22374 4392 22430 4428
rect 22282 3732 22338 3768
rect 22282 3712 22284 3732
rect 22284 3712 22336 3732
rect 22336 3712 22338 3732
rect 22006 3440 22062 3496
rect 22374 2760 22430 2816
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 23662 22208 23718 22264
rect 23478 20984 23534 21040
rect 23202 16360 23258 16416
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 23938 20304 23994 20360
rect 23570 17584 23626 17640
rect 23478 15136 23534 15192
rect 23202 14184 23258 14240
rect 23202 14048 23258 14104
rect 23294 13776 23350 13832
rect 23478 12552 23534 12608
rect 23202 12144 23258 12200
rect 23018 12008 23074 12064
rect 22926 11328 22982 11384
rect 22834 10784 22890 10840
rect 22742 8064 22798 8120
rect 23110 11056 23166 11112
rect 23018 7384 23074 7440
rect 22926 4256 22982 4312
rect 23110 6296 23166 6352
rect 23386 12280 23442 12336
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24582 18828 24638 18864
rect 24582 18808 24584 18828
rect 24584 18808 24636 18828
rect 24636 18808 24638 18828
rect 23938 17040 23994 17096
rect 23570 12008 23626 12064
rect 23938 12416 23994 12472
rect 23294 8336 23350 8392
rect 23570 10240 23626 10296
rect 23570 9968 23626 10024
rect 23754 9968 23810 10024
rect 23662 8472 23718 8528
rect 23754 8336 23810 8392
rect 23478 7268 23534 7304
rect 23478 7248 23480 7268
rect 23480 7248 23532 7268
rect 23532 7248 23534 7268
rect 22650 2896 22706 2952
rect 21822 550 21878 606
rect 23018 3984 23074 4040
rect 24122 17720 24178 17776
rect 24122 15000 24178 15056
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24766 18264 24822 18320
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24858 17584 24914 17640
rect 24858 15000 24914 15056
rect 24766 14320 24822 14376
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 25318 13912 25374 13968
rect 25226 13776 25282 13832
rect 25134 12824 25190 12880
rect 25226 12552 25282 12608
rect 26054 17720 26110 17776
rect 25594 15544 25650 15600
rect 25502 12724 25504 12744
rect 25504 12724 25556 12744
rect 25556 12724 25558 12744
rect 25502 12688 25558 12724
rect 25410 12280 25466 12336
rect 24674 10920 24730 10976
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24674 10104 24730 10160
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24674 8472 24730 8528
rect 24214 8200 24270 8256
rect 23846 6704 23902 6760
rect 23662 4120 23718 4176
rect 22926 1400 22982 1456
rect 23294 3712 23350 3768
rect 23294 3440 23350 3496
rect 23478 3848 23534 3904
rect 24030 5752 24086 5808
rect 24030 3168 24086 3224
rect 23754 2932 23756 2952
rect 23756 2932 23808 2952
rect 23808 2932 23810 2952
rect 23754 2896 23810 2932
rect 23662 2388 23664 2408
rect 23664 2388 23716 2408
rect 23716 2388 23718 2408
rect 23662 2352 23718 2388
rect 23570 1672 23626 1728
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 25410 11600 25466 11656
rect 25226 11192 25282 11248
rect 25134 10240 25190 10296
rect 24950 9288 25006 9344
rect 25410 9560 25466 9616
rect 25318 9016 25374 9072
rect 24766 8200 24822 8256
rect 24950 7928 25006 7984
rect 24674 4936 24730 4992
rect 24582 4564 24584 4584
rect 24584 4564 24636 4584
rect 24636 4564 24638 4584
rect 24582 4528 24638 4564
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24490 3068 24492 3088
rect 24492 3068 24544 3088
rect 24544 3068 24546 3088
rect 24490 3032 24546 3068
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24950 3712 25006 3768
rect 24858 3460 24914 3496
rect 24858 3440 24860 3460
rect 24860 3440 24912 3460
rect 24912 3440 24914 3460
rect 25226 7520 25282 7576
rect 25134 5616 25190 5672
rect 25686 12980 25742 13016
rect 25686 12960 25688 12980
rect 25688 12960 25740 12980
rect 25740 12960 25742 12980
rect 25686 10512 25742 10568
rect 25594 9968 25650 10024
rect 25502 8880 25558 8936
rect 25318 6976 25374 7032
rect 25318 6296 25374 6352
rect 25134 2508 25190 2544
rect 25134 2488 25136 2508
rect 25136 2488 25188 2508
rect 25188 2488 25190 2508
rect 25042 2388 25044 2408
rect 25044 2388 25096 2408
rect 25096 2388 25098 2408
rect 25042 2352 25098 2388
rect 25594 6196 25596 6216
rect 25596 6196 25648 6216
rect 25648 6196 25650 6216
rect 25594 6160 25650 6196
rect 25594 5208 25650 5264
rect 25410 5072 25466 5128
rect 25226 1808 25282 1864
rect 25870 15680 25926 15736
rect 25778 8472 25834 8528
rect 25870 5344 25926 5400
rect 25502 1536 25558 1592
rect 26330 15408 26386 15464
rect 26238 13640 26294 13696
rect 26330 9152 26386 9208
rect 26146 5752 26202 5808
rect 26238 3576 26294 3632
rect 26238 2932 26240 2952
rect 26240 2932 26292 2952
rect 26292 2932 26294 2952
rect 26238 2896 26294 2932
rect 25778 1264 25834 1320
rect 9954 312 10010 368
rect 26422 2896 26478 2952
rect 27618 5344 27674 5400
rect 26790 2216 26846 2272
rect 26330 312 26386 368
<< metal3 >>
rect 0 27706 480 27736
rect 2773 27706 2839 27709
rect 0 27704 2839 27706
rect 0 27648 2778 27704
rect 2834 27648 2839 27704
rect 0 27646 2839 27648
rect 0 27616 480 27646
rect 2773 27643 2839 27646
rect 23473 27706 23539 27709
rect 27520 27706 28000 27736
rect 23473 27704 28000 27706
rect 23473 27648 23478 27704
rect 23534 27648 28000 27704
rect 23473 27646 28000 27648
rect 23473 27643 23539 27646
rect 27520 27616 28000 27646
rect 0 27026 480 27056
rect 3417 27026 3483 27029
rect 0 27024 3483 27026
rect 0 26968 3422 27024
rect 3478 26968 3483 27024
rect 0 26966 3483 26968
rect 0 26936 480 26966
rect 3417 26963 3483 26966
rect 23565 27026 23631 27029
rect 27520 27026 28000 27056
rect 23565 27024 28000 27026
rect 23565 26968 23570 27024
rect 23626 26968 28000 27024
rect 23565 26966 28000 26968
rect 23565 26963 23631 26966
rect 27520 26936 28000 26966
rect 0 26346 480 26376
rect 2221 26346 2287 26349
rect 0 26344 2287 26346
rect 0 26288 2226 26344
rect 2282 26288 2287 26344
rect 0 26286 2287 26288
rect 0 26256 480 26286
rect 2221 26283 2287 26286
rect 23473 26346 23539 26349
rect 27520 26346 28000 26376
rect 23473 26344 28000 26346
rect 23473 26288 23478 26344
rect 23534 26288 28000 26344
rect 23473 26286 28000 26288
rect 23473 26283 23539 26286
rect 27520 26256 28000 26286
rect 0 25666 480 25696
rect 3049 25666 3115 25669
rect 0 25664 3115 25666
rect 0 25608 3054 25664
rect 3110 25608 3115 25664
rect 0 25606 3115 25608
rect 0 25576 480 25606
rect 3049 25603 3115 25606
rect 23473 25666 23539 25669
rect 27520 25666 28000 25696
rect 23473 25664 28000 25666
rect 23473 25608 23478 25664
rect 23534 25608 28000 25664
rect 23473 25606 28000 25608
rect 23473 25603 23539 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 27520 25576 28000 25606
rect 19610 25535 19930 25536
rect 19374 25196 19380 25260
rect 19444 25258 19450 25260
rect 19444 25198 24778 25258
rect 19444 25196 19450 25198
rect 0 25122 480 25152
rect 4521 25122 4587 25125
rect 0 25120 4587 25122
rect 0 25064 4526 25120
rect 4582 25064 4587 25120
rect 0 25062 4587 25064
rect 24718 25122 24778 25198
rect 24718 25062 26802 25122
rect 0 25032 480 25062
rect 4521 25059 4587 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 26742 24986 26802 25062
rect 27520 24986 28000 25016
rect 26742 24926 28000 24986
rect 27520 24896 28000 24926
rect 10277 24512 10597 24513
rect 0 24442 480 24472
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 7097 24442 7163 24445
rect 0 24440 7163 24442
rect 0 24384 7102 24440
rect 7158 24384 7163 24440
rect 0 24382 7163 24384
rect 0 24352 480 24382
rect 7097 24379 7163 24382
rect 20253 24306 20319 24309
rect 27520 24306 28000 24336
rect 20253 24304 28000 24306
rect 20253 24248 20258 24304
rect 20314 24248 28000 24304
rect 20253 24246 28000 24248
rect 20253 24243 20319 24246
rect 27520 24216 28000 24246
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 0 23762 480 23792
rect 14273 23762 14339 23765
rect 0 23760 14339 23762
rect 0 23704 14278 23760
rect 14334 23704 14339 23760
rect 0 23702 14339 23704
rect 0 23672 480 23702
rect 14273 23699 14339 23702
rect 27520 23626 28000 23656
rect 23476 23566 28000 23626
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 20069 23354 20135 23357
rect 23476 23354 23536 23566
rect 27520 23536 28000 23566
rect 20069 23352 23536 23354
rect 20069 23296 20074 23352
rect 20130 23296 23536 23352
rect 20069 23294 23536 23296
rect 20069 23291 20135 23294
rect 0 23082 480 23112
rect 23197 23082 23263 23085
rect 0 23022 3066 23082
rect 0 22992 480 23022
rect 3006 22538 3066 23022
rect 23197 23080 26802 23082
rect 23197 23024 23202 23080
rect 23258 23024 26802 23080
rect 23197 23022 26802 23024
rect 23197 23019 23263 23022
rect 26742 22946 26802 23022
rect 27520 22946 28000 22976
rect 26742 22886 28000 22946
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 27520 22856 28000 22886
rect 24277 22815 24597 22816
rect 14733 22538 14799 22541
rect 3006 22536 14799 22538
rect 3006 22480 14738 22536
rect 14794 22480 14799 22536
rect 3006 22478 14799 22480
rect 14733 22475 14799 22478
rect 0 22402 480 22432
rect 0 22342 3066 22402
rect 0 22312 480 22342
rect 3006 22130 3066 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 23657 22266 23723 22269
rect 27520 22266 28000 22296
rect 23657 22264 28000 22266
rect 23657 22208 23662 22264
rect 23718 22208 28000 22264
rect 23657 22206 28000 22208
rect 23657 22203 23723 22206
rect 27520 22176 28000 22206
rect 22921 22130 22987 22133
rect 3006 22128 22987 22130
rect 3006 22072 22926 22128
rect 22982 22072 22987 22128
rect 3006 22070 22987 22072
rect 22921 22067 22987 22070
rect 0 21858 480 21888
rect 0 21798 2698 21858
rect 0 21768 480 21798
rect 2638 21722 2698 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 2638 21662 2882 21722
rect 2822 21450 2882 21662
rect 20345 21586 20411 21589
rect 27520 21586 28000 21616
rect 20345 21584 28000 21586
rect 20345 21528 20350 21584
rect 20406 21528 28000 21584
rect 20345 21526 28000 21528
rect 20345 21523 20411 21526
rect 27520 21496 28000 21526
rect 9622 21450 9628 21452
rect 2822 21390 9628 21450
rect 9622 21388 9628 21390
rect 9692 21388 9698 21452
rect 10277 21248 10597 21249
rect 0 21178 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 6821 21178 6887 21181
rect 0 21176 6887 21178
rect 0 21120 6826 21176
rect 6882 21120 6887 21176
rect 0 21118 6887 21120
rect 0 21088 480 21118
rect 6821 21115 6887 21118
rect 23473 21042 23539 21045
rect 27520 21042 28000 21072
rect 23473 21040 28000 21042
rect 23473 20984 23478 21040
rect 23534 20984 28000 21040
rect 23473 20982 28000 20984
rect 23473 20979 23539 20982
rect 27520 20952 28000 20982
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 0 20498 480 20528
rect 3969 20498 4035 20501
rect 0 20496 4035 20498
rect 0 20440 3974 20496
rect 4030 20440 4035 20496
rect 0 20438 4035 20440
rect 0 20408 480 20438
rect 3969 20435 4035 20438
rect 9622 20300 9628 20364
rect 9692 20362 9698 20364
rect 16113 20362 16179 20365
rect 9692 20360 16179 20362
rect 9692 20304 16118 20360
rect 16174 20304 16179 20360
rect 9692 20302 16179 20304
rect 9692 20300 9698 20302
rect 16113 20299 16179 20302
rect 23933 20362 23999 20365
rect 27520 20362 28000 20392
rect 23933 20360 28000 20362
rect 23933 20304 23938 20360
rect 23994 20304 28000 20360
rect 23933 20302 28000 20304
rect 23933 20299 23999 20302
rect 27520 20272 28000 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 19818 480 19848
rect 3785 19818 3851 19821
rect 0 19816 3851 19818
rect 0 19760 3790 19816
rect 3846 19760 3851 19816
rect 0 19758 3851 19760
rect 0 19728 480 19758
rect 3785 19755 3851 19758
rect 16481 19818 16547 19821
rect 16481 19816 24962 19818
rect 16481 19760 16486 19816
rect 16542 19760 24962 19816
rect 16481 19758 24962 19760
rect 16481 19755 16547 19758
rect 24902 19682 24962 19758
rect 27520 19682 28000 19712
rect 24902 19622 28000 19682
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 27520 19592 28000 19622
rect 24277 19551 24597 19552
rect 0 19138 480 19168
rect 3233 19138 3299 19141
rect 0 19136 3299 19138
rect 0 19080 3238 19136
rect 3294 19080 3299 19136
rect 0 19078 3299 19080
rect 0 19048 480 19078
rect 3233 19075 3299 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 27520 19002 28000 19032
rect 24902 18942 28000 19002
rect 13353 18866 13419 18869
rect 24577 18866 24643 18869
rect 13353 18864 24643 18866
rect 13353 18808 13358 18864
rect 13414 18808 24582 18864
rect 24638 18808 24643 18864
rect 13353 18806 24643 18808
rect 13353 18803 13419 18806
rect 24577 18803 24643 18806
rect 14273 18730 14339 18733
rect 24902 18730 24962 18942
rect 27520 18912 28000 18942
rect 14273 18728 24962 18730
rect 14273 18672 14278 18728
rect 14334 18672 24962 18728
rect 14273 18670 24962 18672
rect 14273 18667 14339 18670
rect 0 18594 480 18624
rect 6821 18594 6887 18597
rect 12525 18594 12591 18597
rect 0 18534 1410 18594
rect 0 18504 480 18534
rect 1350 18322 1410 18534
rect 6821 18592 12591 18594
rect 6821 18536 6826 18592
rect 6882 18536 12530 18592
rect 12586 18536 12591 18592
rect 6821 18534 12591 18536
rect 6821 18531 6887 18534
rect 12525 18531 12591 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 7557 18322 7623 18325
rect 1350 18320 7623 18322
rect 1350 18264 7562 18320
rect 7618 18264 7623 18320
rect 1350 18262 7623 18264
rect 7557 18259 7623 18262
rect 24761 18322 24827 18325
rect 27520 18322 28000 18352
rect 24761 18320 28000 18322
rect 24761 18264 24766 18320
rect 24822 18264 28000 18320
rect 24761 18262 28000 18264
rect 24761 18259 24827 18262
rect 27520 18232 28000 18262
rect 2037 18052 2103 18053
rect 2037 18050 2084 18052
rect 1992 18048 2084 18050
rect 1992 17992 2042 18048
rect 1992 17990 2084 17992
rect 2037 17988 2084 17990
rect 2148 17988 2154 18052
rect 2037 17987 2103 17988
rect 10277 17984 10597 17985
rect 0 17914 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 3877 17914 3943 17917
rect 0 17912 3943 17914
rect 0 17856 3882 17912
rect 3938 17856 3943 17912
rect 0 17854 3943 17856
rect 0 17824 480 17854
rect 3877 17851 3943 17854
rect 2497 17778 2563 17781
rect 10317 17778 10383 17781
rect 2497 17776 10383 17778
rect 2497 17720 2502 17776
rect 2558 17720 10322 17776
rect 10378 17720 10383 17776
rect 2497 17718 10383 17720
rect 2497 17715 2563 17718
rect 10317 17715 10383 17718
rect 24117 17778 24183 17781
rect 26049 17778 26115 17781
rect 24117 17776 26115 17778
rect 24117 17720 24122 17776
rect 24178 17720 26054 17776
rect 26110 17720 26115 17776
rect 24117 17718 26115 17720
rect 24117 17715 24183 17718
rect 26049 17715 26115 17718
rect 2037 17642 2103 17645
rect 9857 17642 9923 17645
rect 2037 17640 9923 17642
rect 2037 17584 2042 17640
rect 2098 17584 9862 17640
rect 9918 17584 9923 17640
rect 2037 17582 9923 17584
rect 2037 17579 2103 17582
rect 9857 17579 9923 17582
rect 22737 17642 22803 17645
rect 23565 17642 23631 17645
rect 22737 17640 23631 17642
rect 22737 17584 22742 17640
rect 22798 17584 23570 17640
rect 23626 17584 23631 17640
rect 22737 17582 23631 17584
rect 22737 17579 22803 17582
rect 23565 17579 23631 17582
rect 24853 17642 24919 17645
rect 27520 17642 28000 17672
rect 24853 17640 28000 17642
rect 24853 17584 24858 17640
rect 24914 17584 28000 17640
rect 24853 17582 28000 17584
rect 24853 17579 24919 17582
rect 27520 17552 28000 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 0 17234 480 17264
rect 11053 17234 11119 17237
rect 0 17232 11119 17234
rect 0 17176 11058 17232
rect 11114 17176 11119 17232
rect 0 17174 11119 17176
rect 0 17144 480 17174
rect 11053 17171 11119 17174
rect 16849 17234 16915 17237
rect 16849 17232 24962 17234
rect 16849 17176 16854 17232
rect 16910 17176 24962 17232
rect 16849 17174 24962 17176
rect 16849 17171 16915 17174
rect 10041 17098 10107 17101
rect 10317 17098 10383 17101
rect 21173 17098 21239 17101
rect 10041 17096 21239 17098
rect 10041 17040 10046 17096
rect 10102 17040 10322 17096
rect 10378 17040 21178 17096
rect 21234 17040 21239 17096
rect 10041 17038 21239 17040
rect 10041 17035 10107 17038
rect 10317 17035 10383 17038
rect 21173 17035 21239 17038
rect 23933 17100 23999 17101
rect 23933 17096 23980 17100
rect 24044 17098 24050 17100
rect 23933 17040 23938 17096
rect 23933 17036 23980 17040
rect 24044 17038 24090 17098
rect 24044 17036 24050 17038
rect 23933 17035 23999 17036
rect 3141 16962 3207 16965
rect 6310 16962 6316 16964
rect 3141 16960 6316 16962
rect 3141 16904 3146 16960
rect 3202 16904 6316 16960
rect 3141 16902 6316 16904
rect 3141 16899 3207 16902
rect 6310 16900 6316 16902
rect 6380 16900 6386 16964
rect 24902 16962 24962 17174
rect 27520 16962 28000 16992
rect 24902 16902 28000 16962
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 27520 16872 28000 16902
rect 19610 16831 19930 16832
rect 2037 16826 2103 16829
rect 6361 16826 6427 16829
rect 2037 16824 6427 16826
rect 2037 16768 2042 16824
rect 2098 16768 6366 16824
rect 6422 16768 6427 16824
rect 2037 16766 6427 16768
rect 2037 16763 2103 16766
rect 6361 16763 6427 16766
rect 4429 16690 4495 16693
rect 22277 16690 22343 16693
rect 22737 16690 22803 16693
rect 4429 16688 22803 16690
rect 4429 16632 4434 16688
rect 4490 16632 22282 16688
rect 22338 16632 22742 16688
rect 22798 16632 22803 16688
rect 4429 16630 22803 16632
rect 4429 16627 4495 16630
rect 22277 16627 22343 16630
rect 22737 16627 22803 16630
rect 0 16554 480 16584
rect 3785 16554 3851 16557
rect 7465 16554 7531 16557
rect 17309 16554 17375 16557
rect 0 16494 1410 16554
rect 0 16464 480 16494
rect 1350 16010 1410 16494
rect 3785 16552 7531 16554
rect 3785 16496 3790 16552
rect 3846 16496 7470 16552
rect 7526 16496 7531 16552
rect 3785 16494 7531 16496
rect 3785 16491 3851 16494
rect 7465 16491 7531 16494
rect 7606 16494 17234 16554
rect 3693 16418 3759 16421
rect 5441 16418 5507 16421
rect 3693 16416 5507 16418
rect 3693 16360 3698 16416
rect 3754 16360 5446 16416
rect 5502 16360 5507 16416
rect 3693 16358 5507 16360
rect 3693 16355 3759 16358
rect 5441 16355 5507 16358
rect 5993 16418 6059 16421
rect 7606 16418 7666 16494
rect 5993 16416 7666 16418
rect 5993 16360 5998 16416
rect 6054 16360 7666 16416
rect 5993 16358 7666 16360
rect 17174 16418 17234 16494
rect 17309 16552 24962 16554
rect 17309 16496 17314 16552
rect 17370 16496 24962 16552
rect 17309 16494 24962 16496
rect 17309 16491 17375 16494
rect 23197 16418 23263 16421
rect 17174 16416 23263 16418
rect 17174 16360 23202 16416
rect 23258 16360 23263 16416
rect 17174 16358 23263 16360
rect 5993 16355 6059 16358
rect 23197 16355 23263 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 2221 16282 2287 16285
rect 2446 16282 2452 16284
rect 2221 16280 2452 16282
rect 2221 16224 2226 16280
rect 2282 16224 2452 16280
rect 2221 16222 2452 16224
rect 2221 16219 2287 16222
rect 2446 16220 2452 16222
rect 2516 16220 2522 16284
rect 24902 16282 24962 16494
rect 27520 16282 28000 16312
rect 24902 16222 28000 16282
rect 27520 16192 28000 16222
rect 2037 16146 2103 16149
rect 16205 16146 16271 16149
rect 16481 16146 16547 16149
rect 2037 16144 16547 16146
rect 2037 16088 2042 16144
rect 2098 16088 16210 16144
rect 16266 16088 16486 16144
rect 16542 16088 16547 16144
rect 2037 16086 16547 16088
rect 2037 16083 2103 16086
rect 16205 16083 16271 16086
rect 16481 16083 16547 16086
rect 7373 16010 7439 16013
rect 20345 16010 20411 16013
rect 1350 16008 7439 16010
rect 1350 15952 7378 16008
rect 7434 15952 7439 16008
rect 1350 15950 7439 15952
rect 7373 15947 7439 15950
rect 7606 16008 20411 16010
rect 7606 15952 20350 16008
rect 20406 15952 20411 16008
rect 7606 15950 20411 15952
rect 0 15874 480 15904
rect 3785 15874 3851 15877
rect 0 15872 3851 15874
rect 0 15816 3790 15872
rect 3846 15816 3851 15872
rect 0 15814 3851 15816
rect 0 15784 480 15814
rect 3785 15811 3851 15814
rect 4061 15874 4127 15877
rect 4429 15874 4495 15877
rect 7606 15874 7666 15950
rect 20345 15947 20411 15950
rect 4061 15872 7666 15874
rect 4061 15816 4066 15872
rect 4122 15816 4434 15872
rect 4490 15816 7666 15872
rect 4061 15814 7666 15816
rect 20621 15874 20687 15877
rect 21449 15874 21515 15877
rect 20621 15872 21515 15874
rect 20621 15816 20626 15872
rect 20682 15816 21454 15872
rect 21510 15816 21515 15872
rect 20621 15814 21515 15816
rect 4061 15811 4127 15814
rect 4429 15811 4495 15814
rect 20621 15811 20687 15814
rect 21449 15811 21515 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 2497 15738 2563 15741
rect 3325 15738 3391 15741
rect 3693 15738 3759 15741
rect 2497 15736 3759 15738
rect 2497 15680 2502 15736
rect 2558 15680 3330 15736
rect 3386 15680 3698 15736
rect 3754 15680 3759 15736
rect 2497 15678 3759 15680
rect 2497 15675 2563 15678
rect 3325 15675 3391 15678
rect 3693 15675 3759 15678
rect 3969 15738 4035 15741
rect 9673 15738 9739 15741
rect 3969 15736 9739 15738
rect 3969 15680 3974 15736
rect 4030 15680 9678 15736
rect 9734 15680 9739 15736
rect 3969 15678 9739 15680
rect 3969 15675 4035 15678
rect 9673 15675 9739 15678
rect 20437 15738 20503 15741
rect 25865 15738 25931 15741
rect 20437 15736 25931 15738
rect 20437 15680 20442 15736
rect 20498 15680 25870 15736
rect 25926 15680 25931 15736
rect 20437 15678 25931 15680
rect 20437 15675 20503 15678
rect 25865 15675 25931 15678
rect 2957 15602 3023 15605
rect 15561 15602 15627 15605
rect 2957 15600 15627 15602
rect 2957 15544 2962 15600
rect 3018 15544 15566 15600
rect 15622 15544 15627 15600
rect 2957 15542 15627 15544
rect 2957 15539 3023 15542
rect 15561 15539 15627 15542
rect 25589 15602 25655 15605
rect 27520 15602 28000 15632
rect 25589 15600 28000 15602
rect 25589 15544 25594 15600
rect 25650 15544 28000 15600
rect 25589 15542 28000 15544
rect 25589 15539 25655 15542
rect 27520 15512 28000 15542
rect 5257 15468 5323 15469
rect 5206 15404 5212 15468
rect 5276 15466 5323 15468
rect 5441 15466 5507 15469
rect 12893 15466 12959 15469
rect 17309 15466 17375 15469
rect 5276 15464 5368 15466
rect 5318 15408 5368 15464
rect 5276 15406 5368 15408
rect 5441 15464 17375 15466
rect 5441 15408 5446 15464
rect 5502 15408 12898 15464
rect 12954 15408 17314 15464
rect 17370 15408 17375 15464
rect 5441 15406 17375 15408
rect 5276 15404 5323 15406
rect 5257 15403 5323 15404
rect 5441 15403 5507 15406
rect 12893 15403 12959 15406
rect 17309 15403 17375 15406
rect 21081 15466 21147 15469
rect 26325 15466 26391 15469
rect 21081 15464 26391 15466
rect 21081 15408 21086 15464
rect 21142 15408 26330 15464
rect 26386 15408 26391 15464
rect 21081 15406 26391 15408
rect 21081 15403 21147 15406
rect 26325 15403 26391 15406
rect 0 15330 480 15360
rect 2773 15330 2839 15333
rect 0 15328 2839 15330
rect 0 15272 2778 15328
rect 2834 15272 2839 15328
rect 0 15270 2839 15272
rect 0 15240 480 15270
rect 2773 15267 2839 15270
rect 3417 15330 3483 15333
rect 4889 15330 4955 15333
rect 3417 15328 4955 15330
rect 3417 15272 3422 15328
rect 3478 15272 4894 15328
rect 4950 15272 4955 15328
rect 3417 15270 4955 15272
rect 3417 15267 3483 15270
rect 4889 15267 4955 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 10777 15194 10843 15197
rect 12985 15194 13051 15197
rect 20069 15194 20135 15197
rect 23473 15194 23539 15197
rect 10777 15192 13051 15194
rect 10777 15136 10782 15192
rect 10838 15136 12990 15192
rect 13046 15136 13051 15192
rect 10777 15134 13051 15136
rect 10777 15131 10843 15134
rect 12985 15131 13051 15134
rect 15334 15134 19626 15194
rect 6678 15058 6684 15060
rect 3558 14998 6684 15058
rect 2037 14922 2103 14925
rect 3558 14922 3618 14998
rect 6678 14996 6684 14998
rect 6748 15058 6754 15060
rect 11789 15058 11855 15061
rect 13997 15058 14063 15061
rect 15334 15058 15394 15134
rect 6748 15056 11855 15058
rect 6748 15000 11794 15056
rect 11850 15000 11855 15056
rect 6748 14998 11855 15000
rect 6748 14996 6754 14998
rect 11789 14995 11855 14998
rect 12022 15056 15394 15058
rect 12022 15000 14002 15056
rect 14058 15000 15394 15056
rect 12022 14998 15394 15000
rect 16297 15058 16363 15061
rect 19425 15058 19491 15061
rect 16297 15056 19491 15058
rect 16297 15000 16302 15056
rect 16358 15000 19430 15056
rect 19486 15000 19491 15056
rect 16297 14998 19491 15000
rect 19566 15058 19626 15134
rect 20069 15192 23539 15194
rect 20069 15136 20074 15192
rect 20130 15136 23478 15192
rect 23534 15136 23539 15192
rect 20069 15134 23539 15136
rect 20069 15131 20135 15134
rect 23473 15131 23539 15134
rect 24117 15058 24183 15061
rect 24853 15058 24919 15061
rect 19566 15056 24183 15058
rect 19566 15000 24122 15056
rect 24178 15000 24183 15056
rect 19566 14998 24183 15000
rect 2037 14920 3618 14922
rect 2037 14864 2042 14920
rect 2098 14864 3618 14920
rect 2037 14862 3618 14864
rect 3785 14922 3851 14925
rect 11053 14922 11119 14925
rect 12022 14922 12082 14998
rect 13997 14995 14063 14998
rect 16297 14995 16363 14998
rect 19425 14995 19491 14998
rect 24117 14995 24183 14998
rect 24304 15056 24919 15058
rect 24304 15000 24858 15056
rect 24914 15000 24919 15056
rect 24304 14998 24919 15000
rect 3785 14920 5274 14922
rect 3785 14864 3790 14920
rect 3846 14864 5274 14920
rect 3785 14862 5274 14864
rect 2037 14859 2103 14862
rect 3785 14859 3851 14862
rect 1117 14786 1183 14789
rect 4981 14786 5047 14789
rect 1117 14784 5047 14786
rect 1117 14728 1122 14784
rect 1178 14728 4986 14784
rect 5042 14728 5047 14784
rect 1117 14726 5047 14728
rect 5214 14786 5274 14862
rect 11053 14920 12082 14922
rect 11053 14864 11058 14920
rect 11114 14864 12082 14920
rect 11053 14862 12082 14864
rect 12709 14922 12775 14925
rect 24304 14922 24364 14998
rect 24853 14995 24919 14998
rect 27520 14922 28000 14952
rect 12709 14920 24364 14922
rect 12709 14864 12714 14920
rect 12770 14864 24364 14920
rect 12709 14862 24364 14864
rect 24718 14862 28000 14922
rect 11053 14859 11119 14862
rect 12709 14859 12775 14862
rect 5441 14786 5507 14789
rect 9765 14786 9831 14789
rect 5214 14784 9831 14786
rect 5214 14728 5446 14784
rect 5502 14728 9770 14784
rect 9826 14728 9831 14784
rect 5214 14726 9831 14728
rect 1117 14723 1183 14726
rect 4981 14723 5047 14726
rect 5441 14723 5507 14726
rect 9765 14723 9831 14726
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 3049 14650 3115 14653
rect 0 14648 3115 14650
rect 0 14592 3054 14648
rect 3110 14592 3115 14648
rect 0 14590 3115 14592
rect 0 14560 480 14590
rect 3049 14587 3115 14590
rect 3877 14650 3943 14653
rect 7189 14650 7255 14653
rect 3877 14648 7255 14650
rect 3877 14592 3882 14648
rect 3938 14592 7194 14648
rect 7250 14592 7255 14648
rect 3877 14590 7255 14592
rect 3877 14587 3943 14590
rect 7189 14587 7255 14590
rect 21582 14588 21588 14652
rect 21652 14650 21658 14652
rect 24718 14650 24778 14862
rect 27520 14832 28000 14862
rect 21652 14590 24778 14650
rect 21652 14588 21658 14590
rect 2589 14516 2655 14517
rect 2589 14512 2636 14516
rect 2700 14514 2706 14516
rect 4981 14514 5047 14517
rect 2589 14456 2594 14512
rect 2589 14452 2636 14456
rect 2700 14454 2746 14514
rect 4981 14512 12634 14514
rect 4981 14456 4986 14512
rect 5042 14456 12634 14512
rect 4981 14454 12634 14456
rect 2700 14452 2706 14454
rect 2589 14451 2655 14452
rect 4981 14451 5047 14454
rect 1577 14378 1643 14381
rect 3785 14378 3851 14381
rect 1577 14376 3851 14378
rect 1577 14320 1582 14376
rect 1638 14320 3790 14376
rect 3846 14320 3851 14376
rect 1577 14318 3851 14320
rect 1577 14315 1643 14318
rect 3785 14315 3851 14318
rect 5993 14378 6059 14381
rect 7281 14378 7347 14381
rect 5993 14376 7347 14378
rect 5993 14320 5998 14376
rect 6054 14320 7286 14376
rect 7342 14320 7347 14376
rect 5993 14318 7347 14320
rect 12574 14378 12634 14454
rect 12709 14378 12775 14381
rect 16297 14378 16363 14381
rect 12574 14376 16363 14378
rect 12574 14320 12714 14376
rect 12770 14320 16302 14376
rect 16358 14320 16363 14376
rect 12574 14318 16363 14320
rect 5993 14315 6059 14318
rect 7281 14315 7347 14318
rect 12709 14315 12775 14318
rect 16297 14315 16363 14318
rect 24761 14378 24827 14381
rect 27520 14378 28000 14408
rect 24761 14376 28000 14378
rect 24761 14320 24766 14376
rect 24822 14320 28000 14376
rect 24761 14318 28000 14320
rect 24761 14315 24827 14318
rect 27520 14288 28000 14318
rect 1393 14242 1459 14245
rect 4061 14242 4127 14245
rect 1393 14240 4127 14242
rect 1393 14184 1398 14240
rect 1454 14184 4066 14240
rect 4122 14184 4127 14240
rect 1393 14182 4127 14184
rect 1393 14179 1459 14182
rect 4061 14179 4127 14182
rect 23197 14244 23263 14245
rect 23197 14240 23244 14244
rect 23308 14242 23314 14244
rect 23197 14184 23202 14240
rect 23197 14180 23244 14184
rect 23308 14182 23354 14242
rect 23308 14180 23314 14182
rect 23197 14179 23263 14180
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 10869 14106 10935 14109
rect 6134 14104 10935 14106
rect 6134 14048 10874 14104
rect 10930 14048 10935 14104
rect 6134 14046 10935 14048
rect 0 13970 480 14000
rect 1669 13970 1735 13973
rect 0 13968 1735 13970
rect 0 13912 1674 13968
rect 1730 13912 1735 13968
rect 0 13910 1735 13912
rect 0 13880 480 13910
rect 1669 13907 1735 13910
rect 3325 13970 3391 13973
rect 3969 13970 4035 13973
rect 6134 13970 6194 14046
rect 10869 14043 10935 14046
rect 19885 14106 19951 14109
rect 23197 14106 23263 14109
rect 19885 14104 23263 14106
rect 19885 14048 19890 14104
rect 19946 14048 23202 14104
rect 23258 14048 23263 14104
rect 19885 14046 23263 14048
rect 19885 14043 19951 14046
rect 23197 14043 23263 14046
rect 3325 13968 6194 13970
rect 3325 13912 3330 13968
rect 3386 13912 3974 13968
rect 4030 13912 6194 13968
rect 3325 13910 6194 13912
rect 6729 13970 6795 13973
rect 18321 13970 18387 13973
rect 18638 13970 18644 13972
rect 6729 13968 9690 13970
rect 6729 13912 6734 13968
rect 6790 13912 9690 13968
rect 6729 13910 9690 13912
rect 3325 13907 3391 13910
rect 3969 13907 4035 13910
rect 6729 13907 6795 13910
rect 6729 13834 6795 13837
rect 8569 13834 8635 13837
rect 6729 13832 8635 13834
rect 6729 13776 6734 13832
rect 6790 13776 8574 13832
rect 8630 13776 8635 13832
rect 6729 13774 8635 13776
rect 6729 13771 6795 13774
rect 8569 13771 8635 13774
rect 5717 13562 5783 13565
rect 9305 13562 9371 13565
rect 5717 13560 9371 13562
rect 5717 13504 5722 13560
rect 5778 13504 9310 13560
rect 9366 13504 9371 13560
rect 5717 13502 9371 13504
rect 5717 13499 5783 13502
rect 9305 13499 9371 13502
rect 2262 13364 2268 13428
rect 2332 13426 2338 13428
rect 4153 13426 4219 13429
rect 2332 13424 4219 13426
rect 2332 13368 4158 13424
rect 4214 13368 4219 13424
rect 2332 13366 4219 13368
rect 2332 13364 2338 13366
rect 4153 13363 4219 13366
rect 7465 13426 7531 13429
rect 8569 13426 8635 13429
rect 7465 13424 8635 13426
rect 7465 13368 7470 13424
rect 7526 13368 8574 13424
rect 8630 13368 8635 13424
rect 7465 13366 8635 13368
rect 9630 13426 9690 13910
rect 18321 13968 18644 13970
rect 18321 13912 18326 13968
rect 18382 13912 18644 13968
rect 18321 13910 18644 13912
rect 18321 13907 18387 13910
rect 18638 13908 18644 13910
rect 18708 13908 18714 13972
rect 22093 13970 22159 13973
rect 25313 13970 25379 13973
rect 22093 13968 25379 13970
rect 22093 13912 22098 13968
rect 22154 13912 25318 13968
rect 25374 13912 25379 13968
rect 22093 13910 25379 13912
rect 22093 13907 22159 13910
rect 25313 13907 25379 13910
rect 9765 13834 9831 13837
rect 12709 13834 12775 13837
rect 18321 13834 18387 13837
rect 23289 13834 23355 13837
rect 25221 13834 25287 13837
rect 9765 13832 18387 13834
rect 9765 13776 9770 13832
rect 9826 13776 12714 13832
rect 12770 13776 18326 13832
rect 18382 13776 18387 13832
rect 9765 13774 18387 13776
rect 9765 13771 9831 13774
rect 12709 13771 12775 13774
rect 18321 13771 18387 13774
rect 19382 13774 20178 13834
rect 18597 13698 18663 13701
rect 19382 13698 19442 13774
rect 18597 13696 19442 13698
rect 18597 13640 18602 13696
rect 18658 13640 19442 13696
rect 18597 13638 19442 13640
rect 18597 13635 18663 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 20118 13562 20178 13774
rect 23289 13832 25287 13834
rect 23289 13776 23294 13832
rect 23350 13776 25226 13832
rect 25282 13776 25287 13832
rect 23289 13774 25287 13776
rect 23289 13771 23355 13774
rect 25221 13771 25287 13774
rect 26233 13698 26299 13701
rect 27520 13698 28000 13728
rect 26233 13696 28000 13698
rect 26233 13640 26238 13696
rect 26294 13640 28000 13696
rect 26233 13638 28000 13640
rect 26233 13635 26299 13638
rect 27520 13608 28000 13638
rect 23974 13562 23980 13564
rect 20118 13502 23980 13562
rect 23974 13500 23980 13502
rect 24044 13500 24050 13564
rect 21909 13426 21975 13429
rect 9630 13424 21975 13426
rect 9630 13368 21914 13424
rect 21970 13368 21975 13424
rect 9630 13366 21975 13368
rect 7465 13363 7531 13366
rect 8569 13363 8635 13366
rect 21909 13363 21975 13366
rect 0 13290 480 13320
rect 7833 13290 7899 13293
rect 18597 13290 18663 13293
rect 0 13230 6194 13290
rect 0 13200 480 13230
rect 6134 13154 6194 13230
rect 7833 13288 18663 13290
rect 7833 13232 7838 13288
rect 7894 13232 18602 13288
rect 18658 13232 18663 13288
rect 7833 13230 18663 13232
rect 7833 13227 7899 13230
rect 18597 13227 18663 13230
rect 14457 13154 14523 13157
rect 6134 13152 14523 13154
rect 6134 13096 14462 13152
rect 14518 13096 14523 13152
rect 6134 13094 14523 13096
rect 14457 13091 14523 13094
rect 15334 13094 23674 13154
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 2405 13018 2471 13021
rect 1350 13016 2471 13018
rect 1350 12960 2410 13016
rect 2466 12960 2471 13016
rect 1350 12958 2471 12960
rect 0 12746 480 12776
rect 1350 12746 1410 12958
rect 2405 12955 2471 12958
rect 5993 13018 6059 13021
rect 8293 13018 8359 13021
rect 5993 13016 8359 13018
rect 5993 12960 5998 13016
rect 6054 12960 8298 13016
rect 8354 12960 8359 13016
rect 5993 12958 8359 12960
rect 5993 12955 6059 12958
rect 8293 12955 8359 12958
rect 8569 13018 8635 13021
rect 8569 13016 11162 13018
rect 8569 12960 8574 13016
rect 8630 12960 11162 13016
rect 8569 12958 11162 12960
rect 8569 12955 8635 12958
rect 4981 12882 5047 12885
rect 9581 12882 9647 12885
rect 11102 12882 11162 12958
rect 14733 12882 14799 12885
rect 15334 12882 15394 13094
rect 4981 12880 5780 12882
rect 4981 12824 4986 12880
rect 5042 12824 5780 12880
rect 4981 12822 5780 12824
rect 4981 12819 5047 12822
rect 0 12686 1410 12746
rect 5720 12746 5780 12822
rect 9581 12880 10978 12882
rect 9581 12824 9586 12880
rect 9642 12824 10978 12880
rect 9581 12822 10978 12824
rect 11102 12880 15394 12882
rect 11102 12824 14738 12880
rect 14794 12824 15394 12880
rect 11102 12822 15394 12824
rect 19333 12882 19399 12885
rect 23422 12882 23428 12884
rect 19333 12880 23428 12882
rect 19333 12824 19338 12880
rect 19394 12824 23428 12880
rect 19333 12822 23428 12824
rect 9581 12819 9647 12822
rect 10685 12746 10751 12749
rect 5720 12744 10751 12746
rect 5720 12688 10690 12744
rect 10746 12688 10751 12744
rect 5720 12686 10751 12688
rect 10918 12746 10978 12822
rect 14733 12819 14799 12822
rect 19333 12819 19399 12822
rect 23422 12820 23428 12822
rect 23492 12820 23498 12884
rect 23614 12882 23674 13094
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 25681 13018 25747 13021
rect 27520 13018 28000 13048
rect 25681 13016 28000 13018
rect 25681 12960 25686 13016
rect 25742 12960 28000 13016
rect 25681 12958 28000 12960
rect 25681 12955 25747 12958
rect 27520 12928 28000 12958
rect 25129 12882 25195 12885
rect 23614 12880 25195 12882
rect 23614 12824 25134 12880
rect 25190 12824 25195 12880
rect 23614 12822 25195 12824
rect 25129 12819 25195 12822
rect 17769 12746 17835 12749
rect 10918 12744 17835 12746
rect 10918 12688 17774 12744
rect 17830 12688 17835 12744
rect 10918 12686 17835 12688
rect 0 12656 480 12686
rect 10685 12683 10751 12686
rect 17769 12683 17835 12686
rect 18873 12746 18939 12749
rect 25497 12746 25563 12749
rect 18873 12744 25563 12746
rect 18873 12688 18878 12744
rect 18934 12688 25502 12744
rect 25558 12688 25563 12744
rect 18873 12686 25563 12688
rect 18873 12683 18939 12686
rect 25497 12683 25563 12686
rect 1853 12610 1919 12613
rect 3601 12610 3667 12613
rect 7005 12610 7071 12613
rect 1853 12608 1962 12610
rect 1853 12552 1858 12608
rect 1914 12552 1962 12608
rect 1853 12547 1962 12552
rect 3601 12608 7071 12610
rect 3601 12552 3606 12608
rect 3662 12552 7010 12608
rect 7066 12552 7071 12608
rect 3601 12550 7071 12552
rect 3601 12547 3667 12550
rect 7005 12547 7071 12550
rect 11329 12610 11395 12613
rect 18413 12610 18479 12613
rect 11329 12608 18479 12610
rect 11329 12552 11334 12608
rect 11390 12552 18418 12608
rect 18474 12552 18479 12608
rect 11329 12550 18479 12552
rect 11329 12547 11395 12550
rect 18413 12547 18479 12550
rect 23473 12610 23539 12613
rect 25221 12610 25287 12613
rect 23473 12608 25287 12610
rect 23473 12552 23478 12608
rect 23534 12552 25226 12608
rect 25282 12552 25287 12608
rect 23473 12550 25287 12552
rect 23473 12547 23539 12550
rect 25221 12547 25287 12550
rect 1902 12341 1962 12547
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 4521 12474 4587 12477
rect 9581 12474 9647 12477
rect 4521 12472 9647 12474
rect 4521 12416 4526 12472
rect 4582 12416 9586 12472
rect 9642 12416 9647 12472
rect 4521 12414 9647 12416
rect 4521 12411 4587 12414
rect 9581 12411 9647 12414
rect 20805 12474 20871 12477
rect 23933 12474 23999 12477
rect 20805 12472 23999 12474
rect 20805 12416 20810 12472
rect 20866 12416 23938 12472
rect 23994 12416 23999 12472
rect 20805 12414 23999 12416
rect 20805 12411 20871 12414
rect 23933 12411 23999 12414
rect 1853 12336 1962 12341
rect 1853 12280 1858 12336
rect 1914 12280 1962 12336
rect 1853 12278 1962 12280
rect 3325 12338 3391 12341
rect 3693 12338 3759 12341
rect 6177 12340 6243 12341
rect 3325 12336 3759 12338
rect 3325 12280 3330 12336
rect 3386 12280 3698 12336
rect 3754 12280 3759 12336
rect 3325 12278 3759 12280
rect 1853 12275 1919 12278
rect 3325 12275 3391 12278
rect 3693 12275 3759 12278
rect 6126 12276 6132 12340
rect 6196 12338 6243 12340
rect 6637 12340 6703 12341
rect 6637 12338 6684 12340
rect 6196 12336 6288 12338
rect 6238 12280 6288 12336
rect 6196 12278 6288 12280
rect 6592 12336 6684 12338
rect 6592 12280 6642 12336
rect 6592 12278 6684 12280
rect 6196 12276 6243 12278
rect 6177 12275 6243 12276
rect 6637 12276 6684 12278
rect 6748 12276 6754 12340
rect 14089 12338 14155 12341
rect 21265 12338 21331 12341
rect 14089 12336 21331 12338
rect 14089 12280 14094 12336
rect 14150 12280 21270 12336
rect 21326 12280 21331 12336
rect 14089 12278 21331 12280
rect 6637 12275 6703 12276
rect 14089 12275 14155 12278
rect 21265 12275 21331 12278
rect 22093 12338 22159 12341
rect 23381 12338 23447 12341
rect 22093 12336 23447 12338
rect 22093 12280 22098 12336
rect 22154 12280 23386 12336
rect 23442 12280 23447 12336
rect 22093 12278 23447 12280
rect 22093 12275 22159 12278
rect 23381 12275 23447 12278
rect 25405 12338 25471 12341
rect 27520 12338 28000 12368
rect 25405 12336 28000 12338
rect 25405 12280 25410 12336
rect 25466 12280 28000 12336
rect 25405 12278 28000 12280
rect 25405 12275 25471 12278
rect 27520 12248 28000 12278
rect 2037 12202 2103 12205
rect 2262 12202 2268 12204
rect 2037 12200 2268 12202
rect 2037 12144 2042 12200
rect 2098 12144 2268 12200
rect 2037 12142 2268 12144
rect 2037 12139 2103 12142
rect 2262 12140 2268 12142
rect 2332 12140 2338 12204
rect 4061 12202 4127 12205
rect 4337 12202 4403 12205
rect 4061 12200 4403 12202
rect 4061 12144 4066 12200
rect 4122 12144 4342 12200
rect 4398 12144 4403 12200
rect 4061 12142 4403 12144
rect 4061 12139 4127 12142
rect 4337 12139 4403 12142
rect 5717 12202 5783 12205
rect 8569 12202 8635 12205
rect 23197 12204 23263 12205
rect 23197 12202 23244 12204
rect 5717 12200 8635 12202
rect 5717 12144 5722 12200
rect 5778 12144 8574 12200
rect 8630 12144 8635 12200
rect 5717 12142 8635 12144
rect 5717 12139 5783 12142
rect 8569 12139 8635 12142
rect 14414 12142 15394 12202
rect 23152 12200 23244 12202
rect 23152 12144 23202 12200
rect 23152 12142 23244 12144
rect 0 12066 480 12096
rect 749 12066 815 12069
rect 0 12064 815 12066
rect 0 12008 754 12064
rect 810 12008 815 12064
rect 0 12006 815 12008
rect 0 11976 480 12006
rect 749 12003 815 12006
rect 2497 12066 2563 12069
rect 2630 12066 2636 12068
rect 2497 12064 2636 12066
rect 2497 12008 2502 12064
rect 2558 12008 2636 12064
rect 2497 12006 2636 12008
rect 2497 12003 2563 12006
rect 2630 12004 2636 12006
rect 2700 12004 2706 12068
rect 8017 12066 8083 12069
rect 14414 12066 14474 12142
rect 8017 12064 14474 12066
rect 8017 12008 8022 12064
rect 8078 12008 14474 12064
rect 8017 12006 14474 12008
rect 15334 12066 15394 12142
rect 23197 12140 23244 12142
rect 23308 12140 23314 12204
rect 23197 12139 23263 12140
rect 23013 12066 23079 12069
rect 23565 12066 23631 12069
rect 15334 12064 23631 12066
rect 15334 12008 23018 12064
rect 23074 12008 23570 12064
rect 23626 12008 23631 12064
rect 15334 12006 23631 12008
rect 8017 12003 8083 12006
rect 23013 12003 23079 12006
rect 23565 12003 23631 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 7649 11930 7715 11933
rect 11094 11930 11100 11932
rect 7649 11928 11100 11930
rect 7649 11872 7654 11928
rect 7710 11872 11100 11928
rect 7649 11870 11100 11872
rect 7649 11867 7715 11870
rect 11094 11868 11100 11870
rect 11164 11868 11170 11932
rect 19190 11930 19196 11932
rect 15334 11870 19196 11930
rect 4797 11794 4863 11797
rect 7833 11794 7899 11797
rect 15193 11794 15259 11797
rect 4797 11792 15259 11794
rect 4797 11736 4802 11792
rect 4858 11736 7838 11792
rect 7894 11736 15198 11792
rect 15254 11736 15259 11792
rect 4797 11734 15259 11736
rect 4797 11731 4863 11734
rect 7833 11731 7899 11734
rect 15193 11731 15259 11734
rect 2313 11658 2379 11661
rect 6637 11658 6703 11661
rect 2313 11656 6703 11658
rect 2313 11600 2318 11656
rect 2374 11600 6642 11656
rect 6698 11600 6703 11656
rect 2313 11598 6703 11600
rect 2313 11595 2379 11598
rect 6637 11595 6703 11598
rect 8385 11658 8451 11661
rect 15334 11658 15394 11870
rect 19190 11868 19196 11870
rect 19260 11930 19266 11932
rect 20897 11930 20963 11933
rect 19260 11928 20963 11930
rect 19260 11872 20902 11928
rect 20958 11872 20963 11928
rect 19260 11870 20963 11872
rect 19260 11868 19266 11870
rect 20897 11867 20963 11870
rect 22093 11794 22159 11797
rect 22369 11794 22435 11797
rect 22093 11792 22435 11794
rect 22093 11736 22098 11792
rect 22154 11736 22374 11792
rect 22430 11736 22435 11792
rect 22093 11734 22435 11736
rect 22093 11731 22159 11734
rect 22369 11731 22435 11734
rect 8385 11656 15394 11658
rect 8385 11600 8390 11656
rect 8446 11600 15394 11656
rect 8385 11598 15394 11600
rect 15561 11658 15627 11661
rect 18045 11658 18111 11661
rect 20713 11658 20779 11661
rect 15561 11656 20779 11658
rect 15561 11600 15566 11656
rect 15622 11600 18050 11656
rect 18106 11600 20718 11656
rect 20774 11600 20779 11656
rect 15561 11598 20779 11600
rect 8385 11595 8451 11598
rect 15561 11595 15627 11598
rect 18045 11595 18111 11598
rect 20713 11595 20779 11598
rect 25405 11658 25471 11661
rect 27520 11658 28000 11688
rect 25405 11656 28000 11658
rect 25405 11600 25410 11656
rect 25466 11600 28000 11656
rect 25405 11598 28000 11600
rect 25405 11595 25471 11598
rect 27520 11568 28000 11598
rect 5901 11522 5967 11525
rect 6126 11522 6132 11524
rect 5901 11520 6132 11522
rect 5901 11464 5906 11520
rect 5962 11464 6132 11520
rect 5901 11462 6132 11464
rect 5901 11459 5967 11462
rect 6126 11460 6132 11462
rect 6196 11460 6202 11524
rect 15193 11522 15259 11525
rect 18045 11522 18111 11525
rect 15193 11520 18111 11522
rect 15193 11464 15198 11520
rect 15254 11464 18050 11520
rect 18106 11464 18111 11520
rect 15193 11462 18111 11464
rect 15193 11459 15259 11462
rect 18045 11459 18111 11462
rect 10277 11456 10597 11457
rect 0 11386 480 11416
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 2221 11386 2287 11389
rect 0 11384 2287 11386
rect 0 11328 2226 11384
rect 2282 11328 2287 11384
rect 0 11326 2287 11328
rect 0 11296 480 11326
rect 2221 11323 2287 11326
rect 3693 11386 3759 11389
rect 5809 11386 5875 11389
rect 10133 11386 10199 11389
rect 3693 11384 5875 11386
rect 3693 11328 3698 11384
rect 3754 11328 5814 11384
rect 5870 11328 5875 11384
rect 3693 11326 5875 11328
rect 3693 11323 3759 11326
rect 5809 11323 5875 11326
rect 7790 11384 10199 11386
rect 7790 11328 10138 11384
rect 10194 11328 10199 11384
rect 7790 11326 10199 11328
rect 1945 11250 2011 11253
rect 3877 11250 3943 11253
rect 1945 11248 3943 11250
rect 1945 11192 1950 11248
rect 2006 11192 3882 11248
rect 3938 11192 3943 11248
rect 1945 11190 3943 11192
rect 1945 11187 2011 11190
rect 3877 11187 3943 11190
rect 4061 11250 4127 11253
rect 7790 11250 7850 11326
rect 10133 11323 10199 11326
rect 12065 11386 12131 11389
rect 15837 11386 15903 11389
rect 22369 11386 22435 11389
rect 12065 11384 15903 11386
rect 12065 11328 12070 11384
rect 12126 11328 15842 11384
rect 15898 11328 15903 11384
rect 12065 11326 15903 11328
rect 12065 11323 12131 11326
rect 15837 11323 15903 11326
rect 20670 11384 22435 11386
rect 20670 11328 22374 11384
rect 22430 11328 22435 11384
rect 20670 11326 22435 11328
rect 4061 11248 7850 11250
rect 4061 11192 4066 11248
rect 4122 11192 7850 11248
rect 4061 11190 7850 11192
rect 8017 11250 8083 11253
rect 13261 11250 13327 11253
rect 8017 11248 13327 11250
rect 8017 11192 8022 11248
rect 8078 11192 13266 11248
rect 13322 11192 13327 11248
rect 8017 11190 13327 11192
rect 4061 11187 4127 11190
rect 8017 11187 8083 11190
rect 13261 11187 13327 11190
rect 18045 11250 18111 11253
rect 20670 11250 20730 11326
rect 22369 11323 22435 11326
rect 22921 11386 22987 11389
rect 23054 11386 23060 11388
rect 22921 11384 23060 11386
rect 22921 11328 22926 11384
rect 22982 11328 23060 11384
rect 22921 11326 23060 11328
rect 22921 11323 22987 11326
rect 23054 11324 23060 11326
rect 23124 11324 23130 11388
rect 18045 11248 20730 11250
rect 18045 11192 18050 11248
rect 18106 11192 20730 11248
rect 18045 11190 20730 11192
rect 20805 11250 20871 11253
rect 25221 11250 25287 11253
rect 20805 11248 25287 11250
rect 20805 11192 20810 11248
rect 20866 11192 25226 11248
rect 25282 11192 25287 11248
rect 20805 11190 25287 11192
rect 18045 11187 18111 11190
rect 20805 11187 20871 11190
rect 25221 11187 25287 11190
rect 1393 11114 1459 11117
rect 4797 11114 4863 11117
rect 6913 11114 6979 11117
rect 9765 11114 9831 11117
rect 1393 11112 4863 11114
rect 1393 11056 1398 11112
rect 1454 11056 4802 11112
rect 4858 11056 4863 11112
rect 1393 11054 4863 11056
rect 1393 11051 1459 11054
rect 4797 11051 4863 11054
rect 5398 11054 6194 11114
rect 2957 10978 3023 10981
rect 5398 10978 5458 11054
rect 2957 10976 5458 10978
rect 2957 10920 2962 10976
rect 3018 10920 5458 10976
rect 2957 10918 5458 10920
rect 6134 10978 6194 11054
rect 6913 11112 9831 11114
rect 6913 11056 6918 11112
rect 6974 11056 9770 11112
rect 9826 11056 9831 11112
rect 6913 11054 9831 11056
rect 6913 11051 6979 11054
rect 9765 11051 9831 11054
rect 10133 11114 10199 11117
rect 23105 11114 23171 11117
rect 10133 11112 23171 11114
rect 10133 11056 10138 11112
rect 10194 11056 23110 11112
rect 23166 11056 23171 11112
rect 10133 11054 23171 11056
rect 10133 11051 10199 11054
rect 23105 11051 23171 11054
rect 12249 10978 12315 10981
rect 6134 10976 12315 10978
rect 6134 10920 12254 10976
rect 12310 10920 12315 10976
rect 6134 10918 12315 10920
rect 2957 10915 3023 10918
rect 12249 10915 12315 10918
rect 24669 10978 24735 10981
rect 27520 10978 28000 11008
rect 24669 10976 28000 10978
rect 24669 10920 24674 10976
rect 24730 10920 28000 10976
rect 24669 10918 28000 10920
rect 24669 10915 24735 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 27520 10888 28000 10918
rect 24277 10847 24597 10848
rect 7373 10842 7439 10845
rect 13261 10842 13327 10845
rect 7373 10840 13327 10842
rect 7373 10784 7378 10840
rect 7434 10784 13266 10840
rect 13322 10784 13327 10840
rect 7373 10782 13327 10784
rect 7373 10779 7439 10782
rect 13261 10779 13327 10782
rect 15653 10842 15719 10845
rect 22829 10842 22895 10845
rect 15653 10840 22895 10842
rect 15653 10784 15658 10840
rect 15714 10784 22834 10840
rect 22890 10784 22895 10840
rect 15653 10782 22895 10784
rect 15653 10779 15719 10782
rect 22829 10779 22895 10782
rect 0 10706 480 10736
rect 657 10706 723 10709
rect 0 10704 723 10706
rect 0 10648 662 10704
rect 718 10648 723 10704
rect 0 10646 723 10648
rect 0 10616 480 10646
rect 657 10643 723 10646
rect 4245 10706 4311 10709
rect 8017 10706 8083 10709
rect 4245 10704 8083 10706
rect 4245 10648 4250 10704
rect 4306 10648 8022 10704
rect 8078 10648 8083 10704
rect 4245 10646 8083 10648
rect 4245 10643 4311 10646
rect 8017 10643 8083 10646
rect 8201 10706 8267 10709
rect 12157 10706 12223 10709
rect 21081 10706 21147 10709
rect 8201 10704 12223 10706
rect 8201 10648 8206 10704
rect 8262 10648 12162 10704
rect 12218 10648 12223 10704
rect 8201 10646 12223 10648
rect 8201 10643 8267 10646
rect 12157 10643 12223 10646
rect 19428 10704 21147 10706
rect 19428 10648 21086 10704
rect 21142 10648 21147 10704
rect 19428 10646 21147 10648
rect 2405 10570 2471 10573
rect 16021 10570 16087 10573
rect 2405 10568 16087 10570
rect 2405 10512 2410 10568
rect 2466 10512 16026 10568
rect 16082 10512 16087 10568
rect 2405 10510 16087 10512
rect 2405 10507 2471 10510
rect 16021 10507 16087 10510
rect 2313 10434 2379 10437
rect 2446 10434 2452 10436
rect 2313 10432 2452 10434
rect 2313 10376 2318 10432
rect 2374 10376 2452 10432
rect 2313 10374 2452 10376
rect 2313 10371 2379 10374
rect 2446 10372 2452 10374
rect 2516 10372 2522 10436
rect 5441 10434 5507 10437
rect 9673 10434 9739 10437
rect 5441 10432 9739 10434
rect 5441 10376 5446 10432
rect 5502 10376 9678 10432
rect 9734 10376 9739 10432
rect 5441 10374 9739 10376
rect 5441 10371 5507 10374
rect 9673 10371 9739 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 289 10298 355 10301
rect 3785 10298 3851 10301
rect 289 10296 3851 10298
rect 289 10240 294 10296
rect 350 10240 3790 10296
rect 3846 10240 3851 10296
rect 289 10238 3851 10240
rect 289 10235 355 10238
rect 3785 10235 3851 10238
rect 5349 10298 5415 10301
rect 9489 10298 9555 10301
rect 5349 10296 9555 10298
rect 5349 10240 5354 10296
rect 5410 10240 9494 10296
rect 9550 10240 9555 10296
rect 5349 10238 9555 10240
rect 5349 10235 5415 10238
rect 9489 10235 9555 10238
rect 13445 10298 13511 10301
rect 19428 10298 19488 10646
rect 21081 10643 21147 10646
rect 20069 10570 20135 10573
rect 25681 10570 25747 10573
rect 20069 10568 25747 10570
rect 20069 10512 20074 10568
rect 20130 10512 25686 10568
rect 25742 10512 25747 10568
rect 20069 10510 25747 10512
rect 20069 10507 20135 10510
rect 25681 10507 25747 10510
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 13445 10296 19488 10298
rect 13445 10240 13450 10296
rect 13506 10240 19488 10296
rect 13445 10238 19488 10240
rect 13445 10235 13511 10238
rect 20294 10236 20300 10300
rect 20364 10298 20370 10300
rect 20621 10298 20687 10301
rect 23565 10300 23631 10301
rect 23565 10298 23612 10300
rect 20364 10296 20687 10298
rect 20364 10240 20626 10296
rect 20682 10240 20687 10296
rect 20364 10238 20687 10240
rect 23520 10296 23612 10298
rect 23520 10240 23570 10296
rect 23520 10238 23612 10240
rect 20364 10236 20370 10238
rect 20621 10235 20687 10238
rect 23565 10236 23612 10238
rect 23676 10236 23682 10300
rect 25129 10298 25195 10301
rect 27520 10298 28000 10328
rect 25129 10296 28000 10298
rect 25129 10240 25134 10296
rect 25190 10240 28000 10296
rect 25129 10238 28000 10240
rect 23565 10235 23631 10236
rect 25129 10235 25195 10238
rect 27520 10208 28000 10238
rect 7281 10162 7347 10165
rect 14825 10162 14891 10165
rect 24669 10162 24735 10165
rect 7281 10160 14891 10162
rect 7281 10104 7286 10160
rect 7342 10104 14830 10160
rect 14886 10104 14891 10160
rect 7281 10102 14891 10104
rect 7281 10099 7347 10102
rect 14825 10099 14891 10102
rect 17174 10160 24735 10162
rect 17174 10104 24674 10160
rect 24730 10104 24735 10160
rect 17174 10102 24735 10104
rect 0 10026 480 10056
rect 2129 10026 2195 10029
rect 0 10024 2195 10026
rect 0 9968 2134 10024
rect 2190 9968 2195 10024
rect 0 9966 2195 9968
rect 0 9936 480 9966
rect 2129 9963 2195 9966
rect 4705 10026 4771 10029
rect 6637 10026 6703 10029
rect 4705 10024 6703 10026
rect 4705 9968 4710 10024
rect 4766 9968 6642 10024
rect 6698 9968 6703 10024
rect 4705 9966 6703 9968
rect 4705 9963 4771 9966
rect 6637 9963 6703 9966
rect 8661 10026 8727 10029
rect 17174 10026 17234 10102
rect 24669 10099 24735 10102
rect 8661 10024 17234 10026
rect 8661 9968 8666 10024
rect 8722 9968 17234 10024
rect 8661 9966 17234 9968
rect 17401 10026 17467 10029
rect 21582 10026 21588 10028
rect 17401 10024 21588 10026
rect 17401 9968 17406 10024
rect 17462 9968 21588 10024
rect 17401 9966 21588 9968
rect 8661 9963 8727 9966
rect 17401 9963 17467 9966
rect 21582 9964 21588 9966
rect 21652 9964 21658 10028
rect 21725 10026 21791 10029
rect 23565 10026 23631 10029
rect 21725 10024 23631 10026
rect 21725 9968 21730 10024
rect 21786 9968 23570 10024
rect 23626 9968 23631 10024
rect 21725 9966 23631 9968
rect 21725 9963 21791 9966
rect 23565 9963 23631 9966
rect 23749 10026 23815 10029
rect 25589 10026 25655 10029
rect 23749 10024 25655 10026
rect 23749 9968 23754 10024
rect 23810 9968 25594 10024
rect 25650 9968 25655 10024
rect 23749 9966 25655 9968
rect 23749 9963 23815 9966
rect 25589 9963 25655 9966
rect 5257 9892 5323 9893
rect 5206 9890 5212 9892
rect 5166 9830 5212 9890
rect 5276 9888 5323 9892
rect 5318 9832 5323 9888
rect 5206 9828 5212 9830
rect 5276 9828 5323 9832
rect 5257 9827 5323 9828
rect 8109 9890 8175 9893
rect 9121 9890 9187 9893
rect 10133 9890 10199 9893
rect 8109 9888 10199 9890
rect 8109 9832 8114 9888
rect 8170 9832 9126 9888
rect 9182 9832 10138 9888
rect 10194 9832 10199 9888
rect 8109 9830 10199 9832
rect 8109 9827 8175 9830
rect 9121 9827 9187 9830
rect 10133 9827 10199 9830
rect 10777 9890 10843 9893
rect 12985 9890 13051 9893
rect 20989 9890 21055 9893
rect 10777 9888 13051 9890
rect 10777 9832 10782 9888
rect 10838 9832 12990 9888
rect 13046 9832 13051 9888
rect 10777 9830 13051 9832
rect 10777 9827 10843 9830
rect 12985 9827 13051 9830
rect 15334 9888 21055 9890
rect 15334 9832 20994 9888
rect 21050 9832 21055 9888
rect 15334 9830 21055 9832
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 8201 9754 8267 9757
rect 9213 9754 9279 9757
rect 10225 9754 10291 9757
rect 8201 9752 10291 9754
rect 8201 9696 8206 9752
rect 8262 9696 9218 9752
rect 9274 9696 10230 9752
rect 10286 9696 10291 9752
rect 8201 9694 10291 9696
rect 8201 9691 8267 9694
rect 9213 9691 9279 9694
rect 10225 9691 10291 9694
rect 12985 9754 13051 9757
rect 13353 9754 13419 9757
rect 12985 9752 13419 9754
rect 12985 9696 12990 9752
rect 13046 9696 13358 9752
rect 13414 9696 13419 9752
rect 12985 9694 13419 9696
rect 12985 9691 13051 9694
rect 13353 9691 13419 9694
rect 10869 9618 10935 9621
rect 13169 9618 13235 9621
rect 10869 9616 13235 9618
rect 10869 9560 10874 9616
rect 10930 9560 13174 9616
rect 13230 9560 13235 9616
rect 10869 9558 13235 9560
rect 10869 9555 10935 9558
rect 13169 9555 13235 9558
rect 14825 9618 14891 9621
rect 15334 9618 15394 9830
rect 20989 9827 21055 9830
rect 21725 9890 21791 9893
rect 22277 9890 22343 9893
rect 21725 9888 22343 9890
rect 21725 9832 21730 9888
rect 21786 9832 22282 9888
rect 22338 9832 22343 9888
rect 21725 9830 22343 9832
rect 21725 9827 21791 9830
rect 22277 9827 22343 9830
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 20110 9692 20116 9756
rect 20180 9754 20186 9756
rect 20805 9754 20871 9757
rect 20180 9752 20871 9754
rect 20180 9696 20810 9752
rect 20866 9696 20871 9752
rect 20180 9694 20871 9696
rect 20180 9692 20186 9694
rect 20805 9691 20871 9694
rect 14825 9616 15394 9618
rect 14825 9560 14830 9616
rect 14886 9560 15394 9616
rect 14825 9558 15394 9560
rect 14825 9555 14891 9558
rect 18638 9556 18644 9620
rect 18708 9618 18714 9620
rect 18781 9618 18847 9621
rect 18708 9616 18847 9618
rect 18708 9560 18786 9616
rect 18842 9560 18847 9616
rect 18708 9558 18847 9560
rect 18708 9556 18714 9558
rect 18781 9555 18847 9558
rect 19006 9556 19012 9620
rect 19076 9618 19082 9620
rect 20069 9618 20135 9621
rect 19076 9616 20135 9618
rect 19076 9560 20074 9616
rect 20130 9560 20135 9616
rect 19076 9558 20135 9560
rect 19076 9556 19082 9558
rect 20069 9555 20135 9558
rect 20805 9618 20871 9621
rect 21817 9618 21883 9621
rect 20805 9616 21883 9618
rect 20805 9560 20810 9616
rect 20866 9560 21822 9616
rect 21878 9560 21883 9616
rect 20805 9558 21883 9560
rect 20805 9555 20871 9558
rect 21817 9555 21883 9558
rect 25405 9618 25471 9621
rect 27520 9618 28000 9648
rect 25405 9616 28000 9618
rect 25405 9560 25410 9616
rect 25466 9560 28000 9616
rect 25405 9558 28000 9560
rect 25405 9555 25471 9558
rect 27520 9528 28000 9558
rect 0 9482 480 9512
rect 2865 9482 2931 9485
rect 0 9480 2931 9482
rect 0 9424 2870 9480
rect 2926 9424 2931 9480
rect 0 9422 2931 9424
rect 0 9392 480 9422
rect 2865 9419 2931 9422
rect 4521 9482 4587 9485
rect 9949 9482 10015 9485
rect 16849 9482 16915 9485
rect 4521 9480 16915 9482
rect 4521 9424 4526 9480
rect 4582 9424 9954 9480
rect 10010 9424 16854 9480
rect 16910 9424 16915 9480
rect 4521 9422 16915 9424
rect 4521 9419 4587 9422
rect 9949 9419 10015 9422
rect 16849 9419 16915 9422
rect 18689 9480 18755 9485
rect 18689 9424 18694 9480
rect 18750 9424 18755 9480
rect 18689 9419 18755 9424
rect 5165 9346 5231 9349
rect 11329 9346 11395 9349
rect 14549 9346 14615 9349
rect 5165 9344 9322 9346
rect 5165 9288 5170 9344
rect 5226 9288 9322 9344
rect 5165 9286 9322 9288
rect 5165 9283 5231 9286
rect 5073 9210 5139 9213
rect 6913 9210 6979 9213
rect 5073 9208 6979 9210
rect 5073 9152 5078 9208
rect 5134 9152 6918 9208
rect 6974 9152 6979 9208
rect 5073 9150 6979 9152
rect 5073 9147 5139 9150
rect 6913 9147 6979 9150
rect 2497 9074 2563 9077
rect 9029 9074 9095 9077
rect 2497 9072 9095 9074
rect 2497 9016 2502 9072
rect 2558 9016 9034 9072
rect 9090 9016 9095 9072
rect 2497 9014 9095 9016
rect 9262 9074 9322 9286
rect 11329 9344 14615 9346
rect 11329 9288 11334 9344
rect 11390 9288 14554 9344
rect 14610 9288 14615 9344
rect 11329 9286 14615 9288
rect 18692 9346 18752 9419
rect 22461 9348 22527 9349
rect 18822 9346 18828 9348
rect 18692 9286 18828 9346
rect 11329 9283 11395 9286
rect 14549 9283 14615 9286
rect 18822 9284 18828 9286
rect 18892 9284 18898 9348
rect 22461 9344 22508 9348
rect 22572 9346 22578 9348
rect 22461 9288 22466 9344
rect 22461 9284 22508 9288
rect 22572 9286 22618 9346
rect 22572 9284 22578 9286
rect 23054 9284 23060 9348
rect 23124 9346 23130 9348
rect 24945 9346 25011 9349
rect 23124 9344 25011 9346
rect 23124 9288 24950 9344
rect 25006 9288 25011 9344
rect 23124 9286 25011 9288
rect 23124 9284 23130 9286
rect 22461 9283 22527 9284
rect 24945 9283 25011 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 11094 9148 11100 9212
rect 11164 9210 11170 9212
rect 13997 9210 14063 9213
rect 16113 9210 16179 9213
rect 11164 9208 14063 9210
rect 11164 9152 14002 9208
rect 14058 9152 14063 9208
rect 11164 9150 14063 9152
rect 11164 9148 11170 9150
rect 13997 9147 14063 9150
rect 14230 9208 16179 9210
rect 14230 9152 16118 9208
rect 16174 9152 16179 9208
rect 14230 9150 16179 9152
rect 14230 9074 14290 9150
rect 16113 9147 16179 9150
rect 21357 9210 21423 9213
rect 26325 9210 26391 9213
rect 21357 9208 26391 9210
rect 21357 9152 21362 9208
rect 21418 9152 26330 9208
rect 26386 9152 26391 9208
rect 21357 9150 26391 9152
rect 21357 9147 21423 9150
rect 26325 9147 26391 9150
rect 16297 9074 16363 9077
rect 9262 9014 14290 9074
rect 14414 9072 16363 9074
rect 14414 9016 16302 9072
rect 16358 9016 16363 9072
rect 14414 9014 16363 9016
rect 2497 9011 2563 9014
rect 9029 9011 9095 9014
rect 5257 8938 5323 8941
rect 5257 8936 6056 8938
rect 5257 8880 5262 8936
rect 5318 8880 6056 8936
rect 5257 8878 6056 8880
rect 5257 8875 5323 8878
rect 0 8802 480 8832
rect 1669 8802 1735 8805
rect 0 8800 1735 8802
rect 0 8744 1674 8800
rect 1730 8744 1735 8800
rect 0 8742 1735 8744
rect 0 8712 480 8742
rect 1669 8739 1735 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 1853 8666 1919 8669
rect 5441 8666 5507 8669
rect 1853 8664 5507 8666
rect 1853 8608 1858 8664
rect 1914 8608 5446 8664
rect 5502 8608 5507 8664
rect 1853 8606 5507 8608
rect 5996 8666 6056 8878
rect 6494 8876 6500 8940
rect 6564 8938 6570 8940
rect 9673 8938 9739 8941
rect 6564 8936 9739 8938
rect 6564 8880 9678 8936
rect 9734 8880 9739 8936
rect 6564 8878 9739 8880
rect 6564 8876 6570 8878
rect 9673 8875 9739 8878
rect 9949 8938 10015 8941
rect 14414 8938 14474 9014
rect 16297 9011 16363 9014
rect 21633 9074 21699 9077
rect 25313 9074 25379 9077
rect 21633 9072 25379 9074
rect 21633 9016 21638 9072
rect 21694 9016 25318 9072
rect 25374 9016 25379 9072
rect 21633 9014 25379 9016
rect 21633 9011 21699 9014
rect 25313 9011 25379 9014
rect 16665 8938 16731 8941
rect 9949 8936 14474 8938
rect 9949 8880 9954 8936
rect 10010 8880 14474 8936
rect 9949 8878 14474 8880
rect 14598 8936 16731 8938
rect 14598 8880 16670 8936
rect 16726 8880 16731 8936
rect 14598 8878 16731 8880
rect 9949 8875 10015 8878
rect 6126 8740 6132 8804
rect 6196 8802 6202 8804
rect 6637 8802 6703 8805
rect 6196 8800 6703 8802
rect 6196 8744 6642 8800
rect 6698 8744 6703 8800
rect 6196 8742 6703 8744
rect 6196 8740 6202 8742
rect 6637 8739 6703 8742
rect 7833 8802 7899 8805
rect 14598 8802 14658 8878
rect 16665 8875 16731 8878
rect 16849 8938 16915 8941
rect 20805 8938 20871 8941
rect 16849 8936 20871 8938
rect 16849 8880 16854 8936
rect 16910 8880 20810 8936
rect 20866 8880 20871 8936
rect 16849 8878 20871 8880
rect 16849 8875 16915 8878
rect 20805 8875 20871 8878
rect 25497 8938 25563 8941
rect 27520 8938 28000 8968
rect 25497 8936 28000 8938
rect 25497 8880 25502 8936
rect 25558 8880 28000 8936
rect 25497 8878 28000 8880
rect 25497 8875 25563 8878
rect 27520 8848 28000 8878
rect 7833 8800 14658 8802
rect 7833 8744 7838 8800
rect 7894 8744 14658 8800
rect 7833 8742 14658 8744
rect 19701 8802 19767 8805
rect 21817 8802 21883 8805
rect 19701 8800 21883 8802
rect 19701 8744 19706 8800
rect 19762 8744 21822 8800
rect 21878 8744 21883 8800
rect 19701 8742 21883 8744
rect 7833 8739 7899 8742
rect 19701 8739 19767 8742
rect 21817 8739 21883 8742
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 9949 8666 10015 8669
rect 5996 8664 10015 8666
rect 5996 8608 9954 8664
rect 10010 8608 10015 8664
rect 5996 8606 10015 8608
rect 1853 8603 1919 8606
rect 5398 8603 5507 8606
rect 9949 8603 10015 8606
rect 15929 8666 15995 8669
rect 20805 8666 20871 8669
rect 15929 8664 20871 8666
rect 15929 8608 15934 8664
rect 15990 8608 20810 8664
rect 20866 8608 20871 8664
rect 15929 8606 20871 8608
rect 15929 8603 15995 8606
rect 20805 8603 20871 8606
rect 3693 8532 3759 8533
rect 3693 8528 3740 8532
rect 3804 8530 3810 8532
rect 5398 8530 5458 8603
rect 6913 8530 6979 8533
rect 3693 8472 3698 8528
rect 3693 8468 3740 8472
rect 3804 8470 3850 8530
rect 5398 8528 6979 8530
rect 5398 8472 6918 8528
rect 6974 8472 6979 8528
rect 5398 8470 6979 8472
rect 3804 8468 3810 8470
rect 3693 8467 3759 8468
rect 6913 8467 6979 8470
rect 9765 8530 9831 8533
rect 13445 8530 13511 8533
rect 9765 8528 13511 8530
rect 9765 8472 9770 8528
rect 9826 8472 13450 8528
rect 13506 8472 13511 8528
rect 9765 8470 13511 8472
rect 9765 8467 9831 8470
rect 13445 8467 13511 8470
rect 13997 8530 14063 8533
rect 18873 8530 18939 8533
rect 23657 8530 23723 8533
rect 13997 8528 18706 8530
rect 13997 8472 14002 8528
rect 14058 8472 18706 8528
rect 13997 8470 18706 8472
rect 13997 8467 14063 8470
rect 1945 8394 2011 8397
rect 5349 8394 5415 8397
rect 1945 8392 5415 8394
rect 1945 8336 1950 8392
rect 2006 8336 5354 8392
rect 5410 8336 5415 8392
rect 1945 8334 5415 8336
rect 1945 8331 2011 8334
rect 5349 8331 5415 8334
rect 5717 8394 5783 8397
rect 9673 8394 9739 8397
rect 5717 8392 9739 8394
rect 5717 8336 5722 8392
rect 5778 8336 9678 8392
rect 9734 8336 9739 8392
rect 5717 8334 9739 8336
rect 5717 8331 5783 8334
rect 9673 8331 9739 8334
rect 10910 8332 10916 8396
rect 10980 8394 10986 8396
rect 12617 8394 12683 8397
rect 10980 8392 12683 8394
rect 10980 8336 12622 8392
rect 12678 8336 12683 8392
rect 10980 8334 12683 8336
rect 10980 8332 10986 8334
rect 12617 8331 12683 8334
rect 14181 8394 14247 8397
rect 17033 8394 17099 8397
rect 14181 8392 17099 8394
rect 14181 8336 14186 8392
rect 14242 8336 17038 8392
rect 17094 8336 17099 8392
rect 14181 8334 17099 8336
rect 18646 8394 18706 8470
rect 18873 8528 23723 8530
rect 18873 8472 18878 8528
rect 18934 8472 23662 8528
rect 23718 8472 23723 8528
rect 18873 8470 23723 8472
rect 18873 8467 18939 8470
rect 23657 8467 23723 8470
rect 24669 8530 24735 8533
rect 25773 8530 25839 8533
rect 24669 8528 25839 8530
rect 24669 8472 24674 8528
rect 24730 8472 25778 8528
rect 25834 8472 25839 8528
rect 24669 8470 25839 8472
rect 24669 8467 24735 8470
rect 25773 8467 25839 8470
rect 21357 8394 21423 8397
rect 18646 8392 21423 8394
rect 18646 8336 21362 8392
rect 21418 8336 21423 8392
rect 18646 8334 21423 8336
rect 14181 8331 14247 8334
rect 17033 8331 17099 8334
rect 21357 8331 21423 8334
rect 21541 8392 21607 8397
rect 21541 8336 21546 8392
rect 21602 8336 21607 8392
rect 21541 8331 21607 8336
rect 23289 8394 23355 8397
rect 23749 8394 23815 8397
rect 23289 8392 23815 8394
rect 23289 8336 23294 8392
rect 23350 8336 23754 8392
rect 23810 8336 23815 8392
rect 23289 8334 23815 8336
rect 23289 8331 23355 8334
rect 23749 8331 23815 8334
rect 2957 8258 3023 8261
rect 9213 8258 9279 8261
rect 2957 8256 9279 8258
rect 2957 8200 2962 8256
rect 3018 8200 9218 8256
rect 9274 8200 9279 8256
rect 2957 8198 9279 8200
rect 2957 8195 3023 8198
rect 9213 8195 9279 8198
rect 12525 8258 12591 8261
rect 15377 8258 15443 8261
rect 12525 8256 15443 8258
rect 12525 8200 12530 8256
rect 12586 8200 15382 8256
rect 15438 8200 15443 8256
rect 12525 8198 15443 8200
rect 12525 8195 12591 8198
rect 15377 8195 15443 8198
rect 15837 8258 15903 8261
rect 18229 8258 18295 8261
rect 15837 8256 18295 8258
rect 15837 8200 15842 8256
rect 15898 8200 18234 8256
rect 18290 8200 18295 8256
rect 15837 8198 18295 8200
rect 21544 8258 21604 8331
rect 24209 8258 24275 8261
rect 21544 8256 24275 8258
rect 21544 8200 24214 8256
rect 24270 8200 24275 8256
rect 21544 8198 24275 8200
rect 15837 8195 15903 8198
rect 18229 8195 18295 8198
rect 24209 8195 24275 8198
rect 24761 8258 24827 8261
rect 27520 8258 28000 8288
rect 24761 8256 28000 8258
rect 24761 8200 24766 8256
rect 24822 8200 28000 8256
rect 24761 8198 28000 8200
rect 24761 8195 24827 8198
rect 10277 8192 10597 8193
rect 0 8122 480 8152
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8198
rect 19610 8127 19930 8128
rect 1485 8122 1551 8125
rect 0 8120 1551 8122
rect 0 8064 1490 8120
rect 1546 8064 1551 8120
rect 0 8062 1551 8064
rect 0 8032 480 8062
rect 1485 8059 1551 8062
rect 2313 8122 2379 8125
rect 7649 8122 7715 8125
rect 2313 8120 7715 8122
rect 2313 8064 2318 8120
rect 2374 8064 7654 8120
rect 7710 8064 7715 8120
rect 2313 8062 7715 8064
rect 2313 8059 2379 8062
rect 7649 8059 7715 8062
rect 8845 8122 8911 8125
rect 9765 8122 9831 8125
rect 8845 8120 9831 8122
rect 8845 8064 8850 8120
rect 8906 8064 9770 8120
rect 9826 8064 9831 8120
rect 8845 8062 9831 8064
rect 8845 8059 8911 8062
rect 9765 8059 9831 8062
rect 11605 8122 11671 8125
rect 14733 8122 14799 8125
rect 15929 8122 15995 8125
rect 11605 8120 15995 8122
rect 11605 8064 11610 8120
rect 11666 8064 14738 8120
rect 14794 8064 15934 8120
rect 15990 8064 15995 8120
rect 11605 8062 15995 8064
rect 11605 8059 11671 8062
rect 14733 8059 14799 8062
rect 15929 8059 15995 8062
rect 22737 8122 22803 8125
rect 22870 8122 22876 8124
rect 22737 8120 22876 8122
rect 22737 8064 22742 8120
rect 22798 8064 22876 8120
rect 22737 8062 22876 8064
rect 22737 8059 22803 8062
rect 22870 8060 22876 8062
rect 22940 8060 22946 8124
rect 1393 7986 1459 7989
rect 5993 7986 6059 7989
rect 1393 7984 6059 7986
rect 1393 7928 1398 7984
rect 1454 7928 5998 7984
rect 6054 7928 6059 7984
rect 1393 7926 6059 7928
rect 1393 7923 1459 7926
rect 5993 7923 6059 7926
rect 8477 7986 8543 7989
rect 12433 7986 12499 7989
rect 17493 7986 17559 7989
rect 24945 7986 25011 7989
rect 8477 7984 12499 7986
rect 8477 7928 8482 7984
rect 8538 7928 12438 7984
rect 12494 7928 12499 7984
rect 8477 7926 12499 7928
rect 8477 7923 8543 7926
rect 12433 7923 12499 7926
rect 14598 7984 25011 7986
rect 14598 7928 17498 7984
rect 17554 7928 24950 7984
rect 25006 7928 25011 7984
rect 14598 7926 25011 7928
rect 2405 7850 2471 7853
rect 3693 7850 3759 7853
rect 9397 7850 9463 7853
rect 14598 7850 14658 7926
rect 17493 7923 17559 7926
rect 24945 7923 25011 7926
rect 16297 7850 16363 7853
rect 2405 7848 9463 7850
rect 2405 7792 2410 7848
rect 2466 7792 3698 7848
rect 3754 7792 9402 7848
rect 9458 7792 9463 7848
rect 2405 7790 9463 7792
rect 2405 7787 2471 7790
rect 3693 7787 3759 7790
rect 9397 7787 9463 7790
rect 9584 7790 14658 7850
rect 14782 7848 16363 7850
rect 14782 7792 16302 7848
rect 16358 7792 16363 7848
rect 14782 7790 16363 7792
rect 8385 7714 8451 7717
rect 9584 7714 9644 7790
rect 8385 7712 9644 7714
rect 8385 7656 8390 7712
rect 8446 7656 9644 7712
rect 8385 7654 9644 7656
rect 9857 7714 9923 7717
rect 14782 7714 14842 7790
rect 16297 7787 16363 7790
rect 18086 7788 18092 7852
rect 18156 7850 18162 7852
rect 18229 7850 18295 7853
rect 19374 7850 19380 7852
rect 18156 7848 19380 7850
rect 18156 7792 18234 7848
rect 18290 7792 19380 7848
rect 18156 7790 19380 7792
rect 18156 7788 18162 7790
rect 18229 7787 18295 7790
rect 19374 7788 19380 7790
rect 19444 7788 19450 7852
rect 20069 7716 20135 7717
rect 20069 7714 20116 7716
rect 9857 7712 14842 7714
rect 9857 7656 9862 7712
rect 9918 7656 14842 7712
rect 9857 7654 14842 7656
rect 20024 7712 20116 7714
rect 20024 7656 20074 7712
rect 20024 7654 20116 7656
rect 8385 7651 8451 7654
rect 9857 7651 9923 7654
rect 20069 7652 20116 7654
rect 20180 7652 20186 7716
rect 20069 7651 20135 7652
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 3509 7578 3575 7581
rect 1350 7576 3575 7578
rect 1350 7520 3514 7576
rect 3570 7520 3575 7576
rect 1350 7518 3575 7520
rect 0 7442 480 7472
rect 1350 7442 1410 7518
rect 3509 7515 3575 7518
rect 8109 7578 8175 7581
rect 11145 7578 11211 7581
rect 8109 7576 11211 7578
rect 8109 7520 8114 7576
rect 8170 7520 11150 7576
rect 11206 7520 11211 7576
rect 8109 7518 11211 7520
rect 8109 7515 8175 7518
rect 11145 7515 11211 7518
rect 16113 7578 16179 7581
rect 20437 7578 20503 7581
rect 16113 7576 20503 7578
rect 16113 7520 16118 7576
rect 16174 7520 20442 7576
rect 20498 7520 20503 7576
rect 16113 7518 20503 7520
rect 16113 7515 16179 7518
rect 20437 7515 20503 7518
rect 25221 7578 25287 7581
rect 27520 7578 28000 7608
rect 25221 7576 28000 7578
rect 25221 7520 25226 7576
rect 25282 7520 28000 7576
rect 25221 7518 28000 7520
rect 25221 7515 25287 7518
rect 27520 7488 28000 7518
rect 0 7382 1410 7442
rect 2589 7442 2655 7445
rect 7281 7442 7347 7445
rect 10910 7442 10916 7444
rect 2589 7440 7347 7442
rect 2589 7384 2594 7440
rect 2650 7384 7286 7440
rect 7342 7384 7347 7440
rect 2589 7382 7347 7384
rect 0 7352 480 7382
rect 2589 7379 2655 7382
rect 7281 7379 7347 7382
rect 7422 7382 10916 7442
rect 2221 7306 2287 7309
rect 5533 7306 5599 7309
rect 7422 7306 7482 7382
rect 10910 7380 10916 7382
rect 10980 7380 10986 7444
rect 16757 7442 16823 7445
rect 22185 7442 22251 7445
rect 23013 7442 23079 7445
rect 16757 7440 21098 7442
rect 16757 7384 16762 7440
rect 16818 7384 21098 7440
rect 16757 7382 21098 7384
rect 16757 7379 16823 7382
rect 2221 7304 5599 7306
rect 2221 7248 2226 7304
rect 2282 7248 5538 7304
rect 5594 7248 5599 7304
rect 2221 7246 5599 7248
rect 2221 7243 2287 7246
rect 5533 7243 5599 7246
rect 5720 7246 7482 7306
rect 9121 7306 9187 7309
rect 12249 7306 12315 7309
rect 9121 7304 12315 7306
rect 9121 7248 9126 7304
rect 9182 7248 12254 7304
rect 12310 7248 12315 7304
rect 9121 7246 12315 7248
rect 3969 7170 4035 7173
rect 5720 7170 5780 7246
rect 9121 7243 9187 7246
rect 12249 7243 12315 7246
rect 16481 7306 16547 7309
rect 20897 7306 20963 7309
rect 16481 7304 20963 7306
rect 16481 7248 16486 7304
rect 16542 7248 20902 7304
rect 20958 7248 20963 7304
rect 16481 7246 20963 7248
rect 21038 7306 21098 7382
rect 22185 7440 23079 7442
rect 22185 7384 22190 7440
rect 22246 7384 23018 7440
rect 23074 7384 23079 7440
rect 22185 7382 23079 7384
rect 22185 7379 22251 7382
rect 23013 7379 23079 7382
rect 23473 7306 23539 7309
rect 21038 7304 23539 7306
rect 21038 7248 23478 7304
rect 23534 7248 23539 7304
rect 21038 7246 23539 7248
rect 16481 7243 16547 7246
rect 20897 7243 20963 7246
rect 23473 7243 23539 7246
rect 3969 7168 5780 7170
rect 3969 7112 3974 7168
rect 4030 7112 5780 7168
rect 3969 7110 5780 7112
rect 7097 7170 7163 7173
rect 9673 7170 9739 7173
rect 7097 7168 9739 7170
rect 7097 7112 7102 7168
rect 7158 7112 9678 7168
rect 9734 7112 9739 7168
rect 7097 7110 9739 7112
rect 3969 7107 4035 7110
rect 7097 7107 7163 7110
rect 9673 7107 9739 7110
rect 10685 7170 10751 7173
rect 19057 7170 19123 7173
rect 20161 7172 20227 7173
rect 20110 7170 20116 7172
rect 10685 7168 19123 7170
rect 10685 7112 10690 7168
rect 10746 7112 19062 7168
rect 19118 7112 19123 7168
rect 10685 7110 19123 7112
rect 20070 7110 20116 7170
rect 20180 7168 20227 7172
rect 20222 7112 20227 7168
rect 10685 7107 10751 7110
rect 19057 7107 19123 7110
rect 20110 7108 20116 7110
rect 20180 7108 20227 7112
rect 20161 7107 20227 7108
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 6269 7034 6335 7037
rect 9213 7034 9279 7037
rect 6269 7032 9279 7034
rect 6269 6976 6274 7032
rect 6330 6976 9218 7032
rect 9274 6976 9279 7032
rect 6269 6974 9279 6976
rect 6269 6971 6335 6974
rect 9213 6971 9279 6974
rect 17677 7034 17743 7037
rect 19333 7034 19399 7037
rect 17677 7032 19399 7034
rect 17677 6976 17682 7032
rect 17738 6976 19338 7032
rect 19394 6976 19399 7032
rect 17677 6974 19399 6976
rect 17677 6971 17743 6974
rect 19333 6971 19399 6974
rect 20345 7034 20411 7037
rect 21766 7034 21772 7036
rect 20345 7032 21772 7034
rect 20345 6976 20350 7032
rect 20406 6976 21772 7032
rect 20345 6974 21772 6976
rect 20345 6971 20411 6974
rect 21766 6972 21772 6974
rect 21836 6972 21842 7036
rect 25313 7034 25379 7037
rect 27520 7034 28000 7064
rect 25313 7032 28000 7034
rect 25313 6976 25318 7032
rect 25374 6976 28000 7032
rect 25313 6974 28000 6976
rect 25313 6971 25379 6974
rect 27520 6944 28000 6974
rect 1761 6898 1827 6901
rect 5625 6898 5691 6901
rect 1761 6896 5691 6898
rect 1761 6840 1766 6896
rect 1822 6840 5630 6896
rect 5686 6840 5691 6896
rect 1761 6838 5691 6840
rect 1761 6835 1827 6838
rect 5625 6835 5691 6838
rect 13721 6898 13787 6901
rect 20713 6898 20779 6901
rect 13721 6896 20779 6898
rect 13721 6840 13726 6896
rect 13782 6840 20718 6896
rect 20774 6840 20779 6896
rect 13721 6838 20779 6840
rect 13721 6835 13787 6838
rect 20713 6835 20779 6838
rect 0 6762 480 6792
rect 1577 6762 1643 6765
rect 0 6760 1643 6762
rect 0 6704 1582 6760
rect 1638 6704 1643 6760
rect 0 6702 1643 6704
rect 0 6672 480 6702
rect 1577 6699 1643 6702
rect 2313 6762 2379 6765
rect 7465 6762 7531 6765
rect 23841 6762 23907 6765
rect 2313 6760 7298 6762
rect 2313 6704 2318 6760
rect 2374 6704 7298 6760
rect 2313 6702 7298 6704
rect 2313 6699 2379 6702
rect 7238 6626 7298 6702
rect 7465 6760 23907 6762
rect 7465 6704 7470 6760
rect 7526 6704 23846 6760
rect 23902 6704 23907 6760
rect 7465 6702 23907 6704
rect 7465 6699 7531 6702
rect 23841 6699 23907 6702
rect 13813 6626 13879 6629
rect 7238 6624 13879 6626
rect 7238 6568 13818 6624
rect 13874 6568 13879 6624
rect 7238 6566 13879 6568
rect 13813 6563 13879 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 3785 6490 3851 6493
rect 5390 6490 5396 6492
rect 3785 6488 5396 6490
rect 3785 6432 3790 6488
rect 3846 6432 5396 6488
rect 3785 6430 5396 6432
rect 3785 6427 3851 6430
rect 5390 6428 5396 6430
rect 5460 6428 5466 6492
rect 5993 6490 6059 6493
rect 15469 6492 15535 6493
rect 5993 6488 13232 6490
rect 5993 6432 5998 6488
rect 6054 6432 13232 6488
rect 5993 6430 13232 6432
rect 5993 6427 6059 6430
rect 5257 6354 5323 6357
rect 8201 6354 8267 6357
rect 8753 6354 8819 6357
rect 5257 6352 8819 6354
rect 5257 6296 5262 6352
rect 5318 6296 8206 6352
rect 8262 6296 8758 6352
rect 8814 6296 8819 6352
rect 5257 6294 8819 6296
rect 5257 6291 5323 6294
rect 8201 6291 8267 6294
rect 8753 6291 8819 6294
rect 0 6218 480 6248
rect 3366 6218 3372 6220
rect 0 6158 3372 6218
rect 0 6128 480 6158
rect 3366 6156 3372 6158
rect 3436 6156 3442 6220
rect 5717 6218 5783 6221
rect 6453 6218 6519 6221
rect 13172 6218 13232 6430
rect 15469 6488 15516 6492
rect 15580 6490 15586 6492
rect 15469 6432 15474 6488
rect 15469 6428 15516 6432
rect 15580 6430 15626 6490
rect 15580 6428 15586 6430
rect 15469 6427 15535 6428
rect 13353 6354 13419 6357
rect 16573 6354 16639 6357
rect 18045 6354 18111 6357
rect 23105 6356 23171 6357
rect 20110 6354 20116 6356
rect 13353 6352 16639 6354
rect 13353 6296 13358 6352
rect 13414 6296 16578 6352
rect 16634 6296 16639 6352
rect 13353 6294 16639 6296
rect 13353 6291 13419 6294
rect 16573 6291 16639 6294
rect 16806 6352 20116 6354
rect 16806 6296 18050 6352
rect 18106 6296 20116 6352
rect 16806 6294 20116 6296
rect 15837 6218 15903 6221
rect 16806 6218 16866 6294
rect 18045 6291 18111 6294
rect 20110 6292 20116 6294
rect 20180 6292 20186 6356
rect 23054 6292 23060 6356
rect 23124 6354 23171 6356
rect 25313 6354 25379 6357
rect 27520 6354 28000 6384
rect 23124 6352 23216 6354
rect 23166 6296 23216 6352
rect 23124 6294 23216 6296
rect 25313 6352 28000 6354
rect 25313 6296 25318 6352
rect 25374 6296 28000 6352
rect 25313 6294 28000 6296
rect 23124 6292 23171 6294
rect 23105 6291 23171 6292
rect 25313 6291 25379 6294
rect 27520 6264 28000 6294
rect 17309 6218 17375 6221
rect 25589 6218 25655 6221
rect 5717 6216 10748 6218
rect 5717 6160 5722 6216
rect 5778 6160 6458 6216
rect 6514 6160 10748 6216
rect 5717 6158 10748 6160
rect 13172 6158 15762 6218
rect 5717 6155 5783 6158
rect 6453 6155 6519 6158
rect 1669 6082 1735 6085
rect 3049 6082 3115 6085
rect 1669 6080 3115 6082
rect 1669 6024 1674 6080
rect 1730 6024 3054 6080
rect 3110 6024 3115 6080
rect 1669 6022 3115 6024
rect 1669 6019 1735 6022
rect 3049 6019 3115 6022
rect 4429 6082 4495 6085
rect 8937 6082 9003 6085
rect 4429 6080 9003 6082
rect 4429 6024 4434 6080
rect 4490 6024 8942 6080
rect 8998 6024 9003 6080
rect 4429 6022 9003 6024
rect 4429 6019 4495 6022
rect 8937 6019 9003 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 4153 5946 4219 5949
rect 6177 5946 6243 5949
rect 4153 5944 6243 5946
rect 4153 5888 4158 5944
rect 4214 5888 6182 5944
rect 6238 5888 6243 5944
rect 4153 5886 6243 5888
rect 4153 5883 4219 5886
rect 6177 5883 6243 5886
rect 6310 5884 6316 5948
rect 6380 5946 6386 5948
rect 6453 5946 6519 5949
rect 6862 5946 6868 5948
rect 6380 5944 6868 5946
rect 6380 5888 6458 5944
rect 6514 5888 6868 5944
rect 6380 5886 6868 5888
rect 6380 5884 6386 5886
rect 6453 5883 6519 5886
rect 6862 5884 6868 5886
rect 6932 5884 6938 5948
rect 10688 5946 10748 6158
rect 15702 6082 15762 6158
rect 15837 6216 16866 6218
rect 15837 6160 15842 6216
rect 15898 6160 16866 6216
rect 15837 6158 16866 6160
rect 16944 6216 25655 6218
rect 16944 6160 17314 6216
rect 17370 6160 25594 6216
rect 25650 6160 25655 6216
rect 16944 6158 25655 6160
rect 15837 6155 15903 6158
rect 16944 6082 17004 6158
rect 17309 6155 17375 6158
rect 25589 6155 25655 6158
rect 15702 6022 17004 6082
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 12985 5946 13051 5949
rect 10688 5944 13051 5946
rect 10688 5888 12990 5944
rect 13046 5888 13051 5944
rect 10688 5886 13051 5888
rect 12985 5883 13051 5886
rect 20989 5946 21055 5949
rect 22277 5946 22343 5949
rect 20989 5944 22343 5946
rect 20989 5888 20994 5944
rect 21050 5888 22282 5944
rect 22338 5888 22343 5944
rect 20989 5886 22343 5888
rect 20989 5883 21055 5886
rect 22277 5883 22343 5886
rect 6085 5810 6151 5813
rect 8477 5810 8543 5813
rect 6085 5808 8543 5810
rect 6085 5752 6090 5808
rect 6146 5752 8482 5808
rect 8538 5752 8543 5808
rect 6085 5750 8543 5752
rect 6085 5747 6151 5750
rect 8477 5747 8543 5750
rect 24025 5810 24091 5813
rect 26141 5810 26207 5813
rect 24025 5808 26207 5810
rect 24025 5752 24030 5808
rect 24086 5752 26146 5808
rect 26202 5752 26207 5808
rect 24025 5750 26207 5752
rect 24025 5747 24091 5750
rect 26141 5747 26207 5750
rect 4613 5674 4679 5677
rect 8569 5674 8635 5677
rect 4613 5672 8635 5674
rect 4613 5616 4618 5672
rect 4674 5616 8574 5672
rect 8630 5616 8635 5672
rect 4613 5614 8635 5616
rect 4613 5611 4679 5614
rect 8569 5611 8635 5614
rect 9489 5674 9555 5677
rect 10777 5674 10843 5677
rect 12525 5674 12591 5677
rect 9489 5672 12591 5674
rect 9489 5616 9494 5672
rect 9550 5616 10782 5672
rect 10838 5616 12530 5672
rect 12586 5616 12591 5672
rect 9489 5614 12591 5616
rect 9489 5611 9555 5614
rect 10777 5611 10843 5614
rect 12525 5611 12591 5614
rect 13721 5674 13787 5677
rect 16481 5674 16547 5677
rect 13721 5672 16547 5674
rect 13721 5616 13726 5672
rect 13782 5616 16486 5672
rect 16542 5616 16547 5672
rect 13721 5614 16547 5616
rect 13721 5611 13787 5614
rect 16481 5611 16547 5614
rect 17125 5674 17191 5677
rect 20437 5674 20503 5677
rect 17125 5672 20503 5674
rect 17125 5616 17130 5672
rect 17186 5616 20442 5672
rect 20498 5616 20503 5672
rect 17125 5614 20503 5616
rect 17125 5611 17191 5614
rect 20437 5611 20503 5614
rect 25129 5674 25195 5677
rect 27520 5674 28000 5704
rect 25129 5672 28000 5674
rect 25129 5616 25134 5672
rect 25190 5616 28000 5672
rect 25129 5614 28000 5616
rect 25129 5611 25195 5614
rect 27520 5584 28000 5614
rect 0 5538 480 5568
rect 3969 5538 4035 5541
rect 0 5536 4035 5538
rect 0 5480 3974 5536
rect 4030 5480 4035 5536
rect 0 5478 4035 5480
rect 0 5448 480 5478
rect 3969 5475 4035 5478
rect 6085 5538 6151 5541
rect 9029 5538 9095 5541
rect 14273 5540 14339 5541
rect 6085 5536 9095 5538
rect 6085 5480 6090 5536
rect 6146 5480 9034 5536
rect 9090 5480 9095 5536
rect 6085 5478 9095 5480
rect 6085 5475 6151 5478
rect 9029 5475 9095 5478
rect 14222 5476 14228 5540
rect 14292 5538 14339 5540
rect 18781 5538 18847 5541
rect 21541 5538 21607 5541
rect 14292 5536 14384 5538
rect 14334 5480 14384 5536
rect 14292 5478 14384 5480
rect 18781 5536 21607 5538
rect 18781 5480 18786 5536
rect 18842 5480 21546 5536
rect 21602 5480 21607 5536
rect 18781 5478 21607 5480
rect 14292 5476 14339 5478
rect 14273 5475 14339 5476
rect 18781 5475 18847 5478
rect 21541 5475 21607 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 2773 5402 2839 5405
rect 3141 5402 3207 5405
rect 5165 5402 5231 5405
rect 2773 5400 5231 5402
rect 2773 5344 2778 5400
rect 2834 5344 3146 5400
rect 3202 5344 5170 5400
rect 5226 5344 5231 5400
rect 2773 5342 5231 5344
rect 2773 5339 2839 5342
rect 3141 5339 3207 5342
rect 5165 5339 5231 5342
rect 7005 5402 7071 5405
rect 14365 5402 14431 5405
rect 7005 5400 14431 5402
rect 7005 5344 7010 5400
rect 7066 5344 14370 5400
rect 14426 5344 14431 5400
rect 7005 5342 14431 5344
rect 7005 5339 7071 5342
rect 14365 5339 14431 5342
rect 25865 5402 25931 5405
rect 27613 5402 27679 5405
rect 25865 5400 27679 5402
rect 25865 5344 25870 5400
rect 25926 5344 27618 5400
rect 27674 5344 27679 5400
rect 25865 5342 27679 5344
rect 25865 5339 25931 5342
rect 27613 5339 27679 5342
rect 2497 5266 2563 5269
rect 12065 5266 12131 5269
rect 2497 5264 12131 5266
rect 2497 5208 2502 5264
rect 2558 5208 12070 5264
rect 12126 5208 12131 5264
rect 2497 5206 12131 5208
rect 2497 5203 2563 5206
rect 12065 5203 12131 5206
rect 14273 5266 14339 5269
rect 25589 5266 25655 5269
rect 14273 5264 25655 5266
rect 14273 5208 14278 5264
rect 14334 5208 25594 5264
rect 25650 5208 25655 5264
rect 14273 5206 25655 5208
rect 14273 5203 14339 5206
rect 25589 5203 25655 5206
rect 2957 5132 3023 5133
rect 2957 5130 3004 5132
rect 2912 5128 3004 5130
rect 2912 5072 2962 5128
rect 2912 5070 3004 5072
rect 2957 5068 3004 5070
rect 3068 5068 3074 5132
rect 3693 5130 3759 5133
rect 9397 5130 9463 5133
rect 3693 5128 9463 5130
rect 3693 5072 3698 5128
rect 3754 5072 9402 5128
rect 9458 5072 9463 5128
rect 3693 5070 9463 5072
rect 2957 5067 3023 5068
rect 3693 5067 3759 5070
rect 9397 5067 9463 5070
rect 10136 5070 10748 5130
rect 3877 4994 3943 4997
rect 1350 4992 3943 4994
rect 1350 4936 3882 4992
rect 3938 4936 3943 4992
rect 1350 4934 3943 4936
rect 0 4858 480 4888
rect 1350 4858 1410 4934
rect 3877 4931 3943 4934
rect 8477 4994 8543 4997
rect 10136 4994 10196 5070
rect 8477 4992 10196 4994
rect 8477 4936 8482 4992
rect 8538 4936 10196 4992
rect 8477 4934 10196 4936
rect 10688 4994 10748 5070
rect 17902 5068 17908 5132
rect 17972 5130 17978 5132
rect 18045 5130 18111 5133
rect 25405 5130 25471 5133
rect 17972 5128 18111 5130
rect 17972 5072 18050 5128
rect 18106 5072 18111 5128
rect 17972 5070 18111 5072
rect 17972 5068 17978 5070
rect 18045 5067 18111 5070
rect 18646 5128 25471 5130
rect 18646 5072 25410 5128
rect 25466 5072 25471 5128
rect 18646 5070 25471 5072
rect 18505 4994 18571 4997
rect 10688 4992 18571 4994
rect 10688 4936 18510 4992
rect 18566 4936 18571 4992
rect 10688 4934 18571 4936
rect 8477 4931 8543 4934
rect 18505 4931 18571 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 0 4798 1410 4858
rect 0 4768 480 4798
rect 2078 4796 2084 4860
rect 2148 4858 2154 4860
rect 2773 4858 2839 4861
rect 2148 4856 2839 4858
rect 2148 4800 2778 4856
rect 2834 4800 2839 4856
rect 2148 4798 2839 4800
rect 2148 4796 2154 4798
rect 2773 4795 2839 4798
rect 4981 4858 5047 4861
rect 10133 4858 10199 4861
rect 4981 4856 10199 4858
rect 4981 4800 4986 4856
rect 5042 4800 10138 4856
rect 10194 4800 10199 4856
rect 4981 4798 10199 4800
rect 4981 4795 5047 4798
rect 10133 4795 10199 4798
rect 14222 4796 14228 4860
rect 14292 4858 14298 4860
rect 15285 4858 15351 4861
rect 14292 4856 15351 4858
rect 14292 4800 15290 4856
rect 15346 4800 15351 4856
rect 14292 4798 15351 4800
rect 14292 4796 14298 4798
rect 15285 4795 15351 4798
rect 15469 4858 15535 4861
rect 18646 4858 18706 5070
rect 25405 5067 25471 5070
rect 24669 4994 24735 4997
rect 27520 4994 28000 5024
rect 24669 4992 28000 4994
rect 24669 4936 24674 4992
rect 24730 4936 28000 4992
rect 24669 4934 28000 4936
rect 24669 4931 24735 4934
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 27520 4904 28000 4934
rect 19610 4863 19930 4864
rect 15469 4856 18706 4858
rect 15469 4800 15474 4856
rect 15530 4800 18706 4856
rect 15469 4798 18706 4800
rect 20161 4858 20227 4861
rect 20294 4858 20300 4860
rect 20161 4856 20300 4858
rect 20161 4800 20166 4856
rect 20222 4800 20300 4856
rect 20161 4798 20300 4800
rect 15469 4795 15535 4798
rect 20161 4795 20227 4798
rect 20294 4796 20300 4798
rect 20364 4796 20370 4860
rect 3049 4722 3115 4725
rect 8569 4722 8635 4725
rect 3049 4720 8635 4722
rect 3049 4664 3054 4720
rect 3110 4664 8574 4720
rect 8630 4664 8635 4720
rect 3049 4662 8635 4664
rect 3049 4659 3115 4662
rect 8569 4659 8635 4662
rect 9765 4722 9831 4725
rect 9765 4720 17234 4722
rect 9765 4664 9770 4720
rect 9826 4664 17234 4720
rect 9765 4662 17234 4664
rect 9765 4659 9831 4662
rect 5717 4586 5783 4589
rect 14641 4586 14707 4589
rect 5717 4584 14707 4586
rect 5717 4528 5722 4584
rect 5778 4528 14646 4584
rect 14702 4528 14707 4584
rect 5717 4526 14707 4528
rect 5717 4523 5783 4526
rect 14641 4523 14707 4526
rect 15101 4586 15167 4589
rect 17174 4586 17234 4662
rect 19190 4660 19196 4724
rect 19260 4722 19266 4724
rect 19333 4722 19399 4725
rect 19260 4720 19399 4722
rect 19260 4664 19338 4720
rect 19394 4664 19399 4720
rect 19260 4662 19399 4664
rect 19260 4660 19266 4662
rect 19333 4659 19399 4662
rect 20069 4722 20135 4725
rect 21081 4722 21147 4725
rect 20069 4720 21147 4722
rect 20069 4664 20074 4720
rect 20130 4664 21086 4720
rect 21142 4664 21147 4720
rect 20069 4662 21147 4664
rect 20069 4659 20135 4662
rect 21081 4659 21147 4662
rect 23606 4660 23612 4724
rect 23676 4722 23682 4724
rect 23676 4662 24778 4722
rect 23676 4660 23682 4662
rect 24577 4586 24643 4589
rect 15101 4584 17050 4586
rect 15101 4528 15106 4584
rect 15162 4528 17050 4584
rect 15101 4526 17050 4528
rect 17174 4584 24643 4586
rect 17174 4528 24582 4584
rect 24638 4528 24643 4584
rect 17174 4526 24643 4528
rect 15101 4523 15167 4526
rect 7741 4452 7807 4453
rect 7741 4450 7788 4452
rect 7696 4448 7788 4450
rect 7696 4392 7746 4448
rect 7696 4390 7788 4392
rect 7741 4388 7788 4390
rect 7852 4388 7858 4452
rect 8109 4450 8175 4453
rect 11145 4450 11211 4453
rect 8109 4448 11211 4450
rect 8109 4392 8114 4448
rect 8170 4392 11150 4448
rect 11206 4392 11211 4448
rect 8109 4390 11211 4392
rect 16990 4450 17050 4526
rect 24577 4523 24643 4526
rect 18873 4450 18939 4453
rect 16990 4448 18939 4450
rect 16990 4392 18878 4448
rect 18934 4392 18939 4448
rect 16990 4390 18939 4392
rect 7741 4387 7807 4388
rect 8109 4387 8175 4390
rect 11145 4387 11211 4390
rect 18873 4387 18939 4390
rect 20662 4388 20668 4452
rect 20732 4450 20738 4452
rect 22369 4450 22435 4453
rect 20732 4448 22435 4450
rect 20732 4392 22374 4448
rect 22430 4392 22435 4448
rect 20732 4390 22435 4392
rect 20732 4388 20738 4390
rect 22369 4387 22435 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 2129 4314 2195 4317
rect 7925 4314 7991 4317
rect 8150 4314 8156 4316
rect 2129 4312 5458 4314
rect 2129 4256 2134 4312
rect 2190 4256 5458 4312
rect 2129 4254 5458 4256
rect 2129 4251 2195 4254
rect 0 4178 480 4208
rect 5398 4181 5458 4254
rect 7925 4312 8156 4314
rect 7925 4256 7930 4312
rect 7986 4256 8156 4312
rect 7925 4254 8156 4256
rect 7925 4251 7991 4254
rect 8150 4252 8156 4254
rect 8220 4252 8226 4316
rect 8569 4314 8635 4317
rect 14365 4314 14431 4317
rect 8569 4312 14431 4314
rect 8569 4256 8574 4312
rect 8630 4256 14370 4312
rect 14426 4256 14431 4312
rect 8569 4254 14431 4256
rect 8569 4251 8635 4254
rect 14365 4251 14431 4254
rect 20161 4314 20227 4317
rect 22921 4314 22987 4317
rect 20161 4312 22987 4314
rect 20161 4256 20166 4312
rect 20222 4256 22926 4312
rect 22982 4256 22987 4312
rect 20161 4254 22987 4256
rect 24718 4314 24778 4662
rect 27520 4314 28000 4344
rect 24718 4254 28000 4314
rect 20161 4251 20227 4254
rect 22921 4251 22987 4254
rect 27520 4224 28000 4254
rect 3785 4178 3851 4181
rect 0 4176 3851 4178
rect 0 4120 3790 4176
rect 3846 4120 3851 4176
rect 0 4118 3851 4120
rect 5398 4178 5507 4181
rect 11697 4178 11763 4181
rect 5398 4176 11763 4178
rect 5398 4120 5446 4176
rect 5502 4120 11702 4176
rect 11758 4120 11763 4176
rect 5398 4118 11763 4120
rect 0 4088 480 4118
rect 3785 4115 3851 4118
rect 5441 4115 5507 4118
rect 11697 4115 11763 4118
rect 19149 4178 19215 4181
rect 23657 4178 23723 4181
rect 19149 4176 23723 4178
rect 19149 4120 19154 4176
rect 19210 4120 23662 4176
rect 23718 4120 23723 4176
rect 19149 4118 23723 4120
rect 19149 4115 19215 4118
rect 23657 4115 23723 4118
rect 6085 4042 6151 4045
rect 9581 4042 9647 4045
rect 15653 4042 15719 4045
rect 6085 4040 15719 4042
rect 6085 3984 6090 4040
rect 6146 3984 9586 4040
rect 9642 3984 15658 4040
rect 15714 3984 15719 4040
rect 6085 3982 15719 3984
rect 6085 3979 6151 3982
rect 9581 3979 9647 3982
rect 15653 3979 15719 3982
rect 18321 4042 18387 4045
rect 19517 4042 19583 4045
rect 18321 4040 19583 4042
rect 18321 3984 18326 4040
rect 18382 3984 19522 4040
rect 19578 3984 19583 4040
rect 18321 3982 19583 3984
rect 18321 3979 18387 3982
rect 19517 3979 19583 3982
rect 22870 3980 22876 4044
rect 22940 4042 22946 4044
rect 23013 4042 23079 4045
rect 22940 4040 23079 4042
rect 22940 3984 23018 4040
rect 23074 3984 23079 4040
rect 22940 3982 23079 3984
rect 22940 3980 22946 3982
rect 23013 3979 23079 3982
rect 23422 3980 23428 4044
rect 23492 4042 23498 4044
rect 23492 3982 26434 4042
rect 23492 3980 23498 3982
rect 1485 3906 1551 3909
rect 6494 3906 6500 3908
rect 1485 3904 6500 3906
rect 1485 3848 1490 3904
rect 1546 3848 6500 3904
rect 1485 3846 6500 3848
rect 1485 3843 1551 3846
rect 6494 3844 6500 3846
rect 6564 3844 6570 3908
rect 6729 3906 6795 3909
rect 8293 3906 8359 3909
rect 6729 3904 8359 3906
rect 6729 3848 6734 3904
rect 6790 3848 8298 3904
rect 8354 3848 8359 3904
rect 6729 3846 8359 3848
rect 6729 3843 6795 3846
rect 8293 3843 8359 3846
rect 20253 3906 20319 3909
rect 23473 3906 23539 3909
rect 20253 3904 23539 3906
rect 20253 3848 20258 3904
rect 20314 3848 23478 3904
rect 23534 3848 23539 3904
rect 20253 3846 23539 3848
rect 20253 3843 20319 3846
rect 23473 3843 23539 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 2497 3770 2563 3773
rect 4613 3770 4679 3773
rect 2497 3768 4679 3770
rect 2497 3712 2502 3768
rect 2558 3712 4618 3768
rect 4674 3712 4679 3768
rect 2497 3710 4679 3712
rect 2497 3707 2563 3710
rect 4613 3707 4679 3710
rect 6453 3770 6519 3773
rect 9581 3770 9647 3773
rect 6453 3768 9647 3770
rect 6453 3712 6458 3768
rect 6514 3712 9586 3768
rect 9642 3712 9647 3768
rect 6453 3710 9647 3712
rect 6453 3707 6519 3710
rect 9581 3707 9647 3710
rect 16481 3770 16547 3773
rect 19425 3770 19491 3773
rect 16481 3768 19491 3770
rect 16481 3712 16486 3768
rect 16542 3712 19430 3768
rect 19486 3712 19491 3768
rect 16481 3710 19491 3712
rect 16481 3707 16547 3710
rect 19425 3707 19491 3710
rect 22134 3708 22140 3772
rect 22204 3770 22210 3772
rect 22277 3770 22343 3773
rect 22204 3768 22343 3770
rect 22204 3712 22282 3768
rect 22338 3712 22343 3768
rect 22204 3710 22343 3712
rect 22204 3708 22210 3710
rect 22277 3707 22343 3710
rect 23289 3770 23355 3773
rect 24945 3770 25011 3773
rect 23289 3768 25011 3770
rect 23289 3712 23294 3768
rect 23350 3712 24950 3768
rect 25006 3712 25011 3768
rect 23289 3710 25011 3712
rect 23289 3707 23355 3710
rect 24945 3707 25011 3710
rect 7281 3634 7347 3637
rect 12341 3634 12407 3637
rect 7281 3632 12407 3634
rect 7281 3576 7286 3632
rect 7342 3576 12346 3632
rect 12402 3576 12407 3632
rect 7281 3574 12407 3576
rect 7281 3571 7347 3574
rect 12341 3571 12407 3574
rect 14365 3634 14431 3637
rect 26233 3634 26299 3637
rect 14365 3632 26299 3634
rect 14365 3576 14370 3632
rect 14426 3576 26238 3632
rect 26294 3576 26299 3632
rect 14365 3574 26299 3576
rect 26374 3634 26434 3982
rect 27520 3634 28000 3664
rect 26374 3574 28000 3634
rect 14365 3571 14431 3574
rect 26233 3571 26299 3574
rect 27520 3544 28000 3574
rect 0 3498 480 3528
rect 3417 3498 3483 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3408 480 3438
rect 3417 3435 3483 3438
rect 3969 3498 4035 3501
rect 10777 3498 10843 3501
rect 3969 3496 10843 3498
rect 3969 3440 3974 3496
rect 4030 3440 10782 3496
rect 10838 3440 10843 3496
rect 3969 3438 10843 3440
rect 3969 3435 4035 3438
rect 10777 3435 10843 3438
rect 22001 3498 22067 3501
rect 23289 3498 23355 3501
rect 24853 3498 24919 3501
rect 22001 3496 23355 3498
rect 22001 3440 22006 3496
rect 22062 3440 23294 3496
rect 23350 3440 23355 3496
rect 22001 3438 23355 3440
rect 22001 3435 22067 3438
rect 23289 3435 23355 3438
rect 23430 3496 24919 3498
rect 23430 3440 24858 3496
rect 24914 3440 24919 3496
rect 23430 3438 24919 3440
rect 6269 3362 6335 3365
rect 8477 3362 8543 3365
rect 11237 3362 11303 3365
rect 6269 3360 11303 3362
rect 6269 3304 6274 3360
rect 6330 3304 8482 3360
rect 8538 3304 11242 3360
rect 11298 3304 11303 3360
rect 6269 3302 11303 3304
rect 6269 3299 6335 3302
rect 8477 3299 8543 3302
rect 11237 3299 11303 3302
rect 18137 3362 18203 3365
rect 23430 3362 23490 3438
rect 24853 3435 24919 3438
rect 18137 3360 23490 3362
rect 18137 3304 18142 3360
rect 18198 3304 23490 3360
rect 18137 3302 23490 3304
rect 18137 3299 18203 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 15745 3226 15811 3229
rect 17769 3226 17835 3229
rect 15745 3224 17835 3226
rect 15745 3168 15750 3224
rect 15806 3168 17774 3224
rect 17830 3168 17835 3224
rect 15745 3166 17835 3168
rect 15745 3163 15811 3166
rect 17769 3163 17835 3166
rect 18413 3226 18479 3229
rect 24025 3226 24091 3229
rect 18413 3224 24091 3226
rect 18413 3168 18418 3224
rect 18474 3168 24030 3224
rect 24086 3168 24091 3224
rect 18413 3166 24091 3168
rect 18413 3163 18479 3166
rect 24025 3163 24091 3166
rect 3049 3090 3115 3093
rect 5717 3090 5783 3093
rect 8109 3092 8175 3093
rect 8109 3090 8156 3092
rect 3049 3088 3250 3090
rect 3049 3032 3054 3088
rect 3110 3032 3250 3088
rect 3049 3030 3250 3032
rect 3049 3027 3115 3030
rect 0 2954 480 2984
rect 1669 2954 1735 2957
rect 3190 2954 3250 3030
rect 5717 3088 8156 3090
rect 5717 3032 5722 3088
rect 5778 3032 8114 3088
rect 5717 3030 8156 3032
rect 5717 3027 5783 3030
rect 8109 3028 8156 3030
rect 8220 3028 8226 3092
rect 12893 3090 12959 3093
rect 16430 3090 16436 3092
rect 12893 3088 16436 3090
rect 12893 3032 12898 3088
rect 12954 3032 16436 3088
rect 12893 3030 16436 3032
rect 8109 3027 8175 3028
rect 12893 3027 12959 3030
rect 16430 3028 16436 3030
rect 16500 3028 16506 3092
rect 19701 3090 19767 3093
rect 24485 3090 24551 3093
rect 19701 3088 24551 3090
rect 19701 3032 19706 3088
rect 19762 3032 24490 3088
rect 24546 3032 24551 3088
rect 19701 3030 24551 3032
rect 19701 3027 19767 3030
rect 24485 3027 24551 3030
rect 11145 2954 11211 2957
rect 0 2894 1410 2954
rect 0 2864 480 2894
rect 1350 2818 1410 2894
rect 1669 2952 3020 2954
rect 1669 2896 1674 2952
rect 1730 2896 3020 2952
rect 1669 2894 3020 2896
rect 3190 2952 11211 2954
rect 3190 2896 11150 2952
rect 11206 2896 11211 2952
rect 3190 2894 11211 2896
rect 1669 2891 1735 2894
rect 2960 2818 3020 2894
rect 11145 2891 11211 2894
rect 17769 2954 17835 2957
rect 22645 2954 22711 2957
rect 17769 2952 22711 2954
rect 17769 2896 17774 2952
rect 17830 2896 22650 2952
rect 22706 2896 22711 2952
rect 17769 2894 22711 2896
rect 17769 2891 17835 2894
rect 22645 2891 22711 2894
rect 23606 2892 23612 2956
rect 23676 2954 23682 2956
rect 23749 2954 23815 2957
rect 26233 2954 26299 2957
rect 23676 2952 26299 2954
rect 23676 2896 23754 2952
rect 23810 2896 26238 2952
rect 26294 2896 26299 2952
rect 23676 2894 26299 2896
rect 23676 2892 23682 2894
rect 23749 2891 23815 2894
rect 26233 2891 26299 2894
rect 26417 2954 26483 2957
rect 27520 2954 28000 2984
rect 26417 2952 28000 2954
rect 26417 2896 26422 2952
rect 26478 2896 28000 2952
rect 26417 2894 28000 2896
rect 26417 2891 26483 2894
rect 27520 2864 28000 2894
rect 9305 2818 9371 2821
rect 1350 2758 2882 2818
rect 2960 2816 9371 2818
rect 2960 2760 9310 2816
rect 9366 2760 9371 2816
rect 2960 2758 9371 2760
rect 2822 2682 2882 2758
rect 9305 2755 9371 2758
rect 16573 2818 16639 2821
rect 19333 2818 19399 2821
rect 16573 2816 19399 2818
rect 16573 2760 16578 2816
rect 16634 2760 19338 2816
rect 19394 2760 19399 2816
rect 16573 2758 19399 2760
rect 16573 2755 16639 2758
rect 19333 2755 19399 2758
rect 22369 2818 22435 2821
rect 22502 2818 22508 2820
rect 22369 2816 22508 2818
rect 22369 2760 22374 2816
rect 22430 2760 22508 2816
rect 22369 2758 22508 2760
rect 22369 2755 22435 2758
rect 22502 2756 22508 2758
rect 22572 2756 22578 2820
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 4061 2682 4127 2685
rect 2822 2680 4127 2682
rect 2822 2624 4066 2680
rect 4122 2624 4127 2680
rect 2822 2622 4127 2624
rect 4061 2619 4127 2622
rect 5349 2682 5415 2685
rect 9121 2682 9187 2685
rect 5349 2680 9187 2682
rect 5349 2624 5354 2680
rect 5410 2624 9126 2680
rect 9182 2624 9187 2680
rect 5349 2622 9187 2624
rect 5349 2619 5415 2622
rect 9121 2619 9187 2622
rect 11094 2620 11100 2684
rect 11164 2682 11170 2684
rect 18229 2682 18295 2685
rect 11164 2680 18295 2682
rect 11164 2624 18234 2680
rect 18290 2624 18295 2680
rect 11164 2622 18295 2624
rect 11164 2620 11170 2622
rect 18229 2619 18295 2622
rect 2129 2546 2195 2549
rect 6637 2546 6703 2549
rect 2129 2544 6703 2546
rect 2129 2488 2134 2544
rect 2190 2488 6642 2544
rect 6698 2488 6703 2544
rect 2129 2486 6703 2488
rect 2129 2483 2195 2486
rect 6637 2483 6703 2486
rect 10133 2546 10199 2549
rect 16021 2546 16087 2549
rect 10133 2544 16087 2546
rect 10133 2488 10138 2544
rect 10194 2488 16026 2544
rect 16082 2488 16087 2544
rect 10133 2486 16087 2488
rect 10133 2483 10199 2486
rect 16021 2483 16087 2486
rect 19425 2546 19491 2549
rect 25129 2546 25195 2549
rect 19425 2544 25195 2546
rect 19425 2488 19430 2544
rect 19486 2488 25134 2544
rect 25190 2488 25195 2544
rect 19425 2486 25195 2488
rect 19425 2483 19491 2486
rect 25129 2483 25195 2486
rect 12801 2410 12867 2413
rect 1350 2408 12867 2410
rect 1350 2352 12806 2408
rect 12862 2352 12867 2408
rect 1350 2350 12867 2352
rect 0 2274 480 2304
rect 1350 2274 1410 2350
rect 12801 2347 12867 2350
rect 13905 2410 13971 2413
rect 18781 2410 18847 2413
rect 23657 2410 23723 2413
rect 25037 2410 25103 2413
rect 13905 2408 23723 2410
rect 13905 2352 13910 2408
rect 13966 2352 18786 2408
rect 18842 2352 23662 2408
rect 23718 2352 23723 2408
rect 13905 2350 23723 2352
rect 13905 2347 13971 2350
rect 18781 2347 18847 2350
rect 23657 2347 23723 2350
rect 23982 2408 25103 2410
rect 23982 2352 25042 2408
rect 25098 2352 25103 2408
rect 23982 2350 25103 2352
rect 0 2214 1410 2274
rect 2497 2274 2563 2277
rect 4797 2274 4863 2277
rect 2497 2272 4863 2274
rect 2497 2216 2502 2272
rect 2558 2216 4802 2272
rect 4858 2216 4863 2272
rect 2497 2214 4863 2216
rect 0 2184 480 2214
rect 2497 2211 2563 2214
rect 4797 2211 4863 2214
rect 5993 2274 6059 2277
rect 6637 2274 6703 2277
rect 9121 2274 9187 2277
rect 5993 2272 9187 2274
rect 5993 2216 5998 2272
rect 6054 2216 6642 2272
rect 6698 2216 9126 2272
rect 9182 2216 9187 2272
rect 5993 2214 9187 2216
rect 5993 2211 6059 2214
rect 6637 2211 6703 2214
rect 9121 2211 9187 2214
rect 10777 2274 10843 2277
rect 13629 2274 13695 2277
rect 10777 2272 13695 2274
rect 10777 2216 10782 2272
rect 10838 2216 13634 2272
rect 13690 2216 13695 2272
rect 10777 2214 13695 2216
rect 10777 2211 10843 2214
rect 13629 2211 13695 2214
rect 21173 2274 21239 2277
rect 23982 2274 24042 2350
rect 25037 2347 25103 2350
rect 21173 2272 24042 2274
rect 21173 2216 21178 2272
rect 21234 2216 24042 2272
rect 21173 2214 24042 2216
rect 26785 2274 26851 2277
rect 27520 2274 28000 2304
rect 26785 2272 28000 2274
rect 26785 2216 26790 2272
rect 26846 2216 28000 2272
rect 26785 2214 28000 2216
rect 21173 2211 21239 2214
rect 26785 2211 26851 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 27520 2184 28000 2214
rect 24277 2143 24597 2144
rect 3693 2140 3759 2141
rect 3693 2138 3740 2140
rect 3648 2136 3740 2138
rect 3648 2080 3698 2136
rect 3648 2078 3740 2080
rect 3693 2076 3740 2078
rect 3804 2076 3810 2140
rect 5993 2138 6059 2141
rect 9857 2138 9923 2141
rect 5993 2136 9923 2138
rect 5993 2080 5998 2136
rect 6054 2080 9862 2136
rect 9918 2080 9923 2136
rect 5993 2078 9923 2080
rect 3693 2075 3759 2076
rect 5993 2075 6059 2078
rect 9857 2075 9923 2078
rect 16941 2138 17007 2141
rect 20989 2138 21055 2141
rect 16941 2136 21055 2138
rect 16941 2080 16946 2136
rect 17002 2080 20994 2136
rect 21050 2080 21055 2136
rect 16941 2078 21055 2080
rect 16941 2075 17007 2078
rect 20989 2075 21055 2078
rect 4061 2002 4127 2005
rect 8661 2002 8727 2005
rect 17309 2002 17375 2005
rect 4061 2000 8727 2002
rect 4061 1944 4066 2000
rect 4122 1944 8666 2000
rect 8722 1944 8727 2000
rect 4061 1942 8727 1944
rect 4061 1939 4127 1942
rect 8661 1939 8727 1942
rect 8894 2000 17375 2002
rect 8894 1944 17314 2000
rect 17370 1944 17375 2000
rect 8894 1942 17375 1944
rect 5257 1866 5323 1869
rect 8894 1866 8954 1942
rect 17309 1939 17375 1942
rect 5257 1864 8954 1866
rect 5257 1808 5262 1864
rect 5318 1808 8954 1864
rect 5257 1806 8954 1808
rect 9121 1866 9187 1869
rect 20897 1866 20963 1869
rect 25221 1866 25287 1869
rect 9121 1864 20963 1866
rect 9121 1808 9126 1864
rect 9182 1808 20902 1864
rect 20958 1808 20963 1864
rect 9121 1806 20963 1808
rect 5257 1803 5323 1806
rect 9121 1803 9187 1806
rect 20897 1803 20963 1806
rect 21222 1864 25287 1866
rect 21222 1808 25226 1864
rect 25282 1808 25287 1864
rect 21222 1806 25287 1808
rect 2957 1730 3023 1733
rect 14181 1730 14247 1733
rect 2957 1728 14247 1730
rect 2957 1672 2962 1728
rect 3018 1672 14186 1728
rect 14242 1672 14247 1728
rect 2957 1670 14247 1672
rect 2957 1667 3023 1670
rect 14181 1667 14247 1670
rect 15377 1730 15443 1733
rect 21222 1730 21282 1806
rect 25221 1803 25287 1806
rect 15377 1728 21282 1730
rect 15377 1672 15382 1728
rect 15438 1672 21282 1728
rect 15377 1670 21282 1672
rect 23565 1730 23631 1733
rect 23565 1728 27538 1730
rect 23565 1672 23570 1728
rect 23626 1672 27538 1728
rect 23565 1670 27538 1672
rect 15377 1667 15443 1670
rect 23565 1667 23631 1670
rect 27478 1624 27538 1670
rect 0 1594 480 1624
rect 5993 1594 6059 1597
rect 0 1592 6059 1594
rect 0 1536 5998 1592
rect 6054 1536 6059 1592
rect 0 1534 6059 1536
rect 0 1504 480 1534
rect 5993 1531 6059 1534
rect 6361 1594 6427 1597
rect 17125 1594 17191 1597
rect 6361 1592 17191 1594
rect 6361 1536 6366 1592
rect 6422 1536 17130 1592
rect 17186 1536 17191 1592
rect 6361 1534 17191 1536
rect 6361 1531 6427 1534
rect 17125 1531 17191 1534
rect 18321 1594 18387 1597
rect 25497 1594 25563 1597
rect 18321 1592 25563 1594
rect 18321 1536 18326 1592
rect 18382 1536 25502 1592
rect 25558 1536 25563 1592
rect 18321 1534 25563 1536
rect 27478 1534 28000 1624
rect 18321 1531 18387 1534
rect 25497 1531 25563 1534
rect 27520 1504 28000 1534
rect 2221 1458 2287 1461
rect 11697 1458 11763 1461
rect 2221 1456 11763 1458
rect 2221 1400 2226 1456
rect 2282 1400 11702 1456
rect 11758 1400 11763 1456
rect 2221 1398 11763 1400
rect 2221 1395 2287 1398
rect 11697 1395 11763 1398
rect 15837 1458 15903 1461
rect 16941 1458 17007 1461
rect 15837 1456 17007 1458
rect 15837 1400 15842 1456
rect 15898 1400 16946 1456
rect 17002 1400 17007 1456
rect 15837 1398 17007 1400
rect 15837 1395 15903 1398
rect 16941 1395 17007 1398
rect 17125 1458 17191 1461
rect 22921 1458 22987 1461
rect 17125 1456 22987 1458
rect 17125 1400 17130 1456
rect 17186 1400 22926 1456
rect 22982 1400 22987 1456
rect 17125 1398 22987 1400
rect 17125 1395 17191 1398
rect 22921 1395 22987 1398
rect 12985 1322 13051 1325
rect 25773 1322 25839 1325
rect 12985 1320 25839 1322
rect 12985 1264 12990 1320
rect 13046 1264 25778 1320
rect 25834 1264 25839 1320
rect 12985 1262 25839 1264
rect 12985 1259 13051 1262
rect 25773 1259 25839 1262
rect 17217 1186 17283 1189
rect 4800 1184 17283 1186
rect 4800 1128 17222 1184
rect 17278 1128 17283 1184
rect 4800 1126 17283 1128
rect 0 914 480 944
rect 4800 914 4860 1126
rect 17217 1123 17283 1126
rect 0 854 4860 914
rect 7557 914 7623 917
rect 13629 914 13695 917
rect 7557 912 13695 914
rect 7557 856 7562 912
rect 7618 856 13634 912
rect 13690 856 13695 912
rect 7557 854 13695 856
rect 0 824 480 854
rect 7557 851 7623 854
rect 13629 851 13695 854
rect 19057 914 19123 917
rect 27520 914 28000 944
rect 19057 912 28000 914
rect 19057 856 19062 912
rect 19118 856 28000 912
rect 19057 854 28000 856
rect 19057 851 19123 854
rect 27520 824 28000 854
rect 21766 580 21772 644
rect 21836 642 21842 644
rect 21836 611 21880 642
rect 21836 608 21883 611
rect 21836 606 21894 608
rect 21817 550 21822 580
rect 21878 550 21894 606
rect 21817 548 21894 550
rect 21817 545 21883 548
rect 0 370 480 400
rect 9949 370 10015 373
rect 0 368 10015 370
rect 0 312 9954 368
rect 10010 312 10015 368
rect 0 310 10015 312
rect 0 280 480 310
rect 9949 307 10015 310
rect 26325 370 26391 373
rect 27520 370 28000 400
rect 26325 368 28000 370
rect 26325 312 26330 368
rect 26386 312 28000 368
rect 26325 310 28000 312
rect 26325 307 26391 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 19380 25196 19444 25260
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 9628 21388 9692 21452
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 9628 20300 9692 20364
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 2084 18048 2148 18052
rect 2084 17992 2098 18048
rect 2098 17992 2148 18048
rect 2084 17988 2148 17992
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 23980 17096 24044 17100
rect 23980 17040 23994 17096
rect 23994 17040 24044 17096
rect 23980 17036 24044 17040
rect 6316 16900 6380 16964
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 2452 16220 2516 16284
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5212 15464 5276 15468
rect 5212 15408 5262 15464
rect 5262 15408 5276 15464
rect 5212 15404 5276 15408
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 6684 14996 6748 15060
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 21588 14588 21652 14652
rect 2636 14512 2700 14516
rect 2636 14456 2650 14512
rect 2650 14456 2700 14512
rect 2636 14452 2700 14456
rect 23244 14240 23308 14244
rect 23244 14184 23258 14240
rect 23258 14184 23308 14240
rect 23244 14180 23308 14184
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 2268 13364 2332 13428
rect 18644 13908 18708 13972
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 23980 13500 24044 13564
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 23428 12820 23492 12884
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 6132 12336 6196 12340
rect 6132 12280 6182 12336
rect 6182 12280 6196 12336
rect 6132 12276 6196 12280
rect 6684 12336 6748 12340
rect 6684 12280 6698 12336
rect 6698 12280 6748 12336
rect 6684 12276 6748 12280
rect 2268 12140 2332 12204
rect 23244 12200 23308 12204
rect 23244 12144 23258 12200
rect 23258 12144 23308 12200
rect 2636 12004 2700 12068
rect 23244 12140 23308 12144
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 11100 11868 11164 11932
rect 19196 11868 19260 11932
rect 6132 11460 6196 11524
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 23060 11324 23124 11388
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 2452 10372 2516 10436
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 20300 10236 20364 10300
rect 23612 10296 23676 10300
rect 23612 10240 23626 10296
rect 23626 10240 23676 10296
rect 23612 10236 23676 10240
rect 21588 9964 21652 10028
rect 5212 9888 5276 9892
rect 5212 9832 5262 9888
rect 5262 9832 5276 9888
rect 5212 9828 5276 9832
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 20116 9692 20180 9756
rect 18644 9556 18708 9620
rect 19012 9556 19076 9620
rect 18828 9284 18892 9348
rect 22508 9344 22572 9348
rect 22508 9288 22522 9344
rect 22522 9288 22572 9344
rect 22508 9284 22572 9288
rect 23060 9284 23124 9348
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 11100 9148 11164 9212
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 6500 8876 6564 8940
rect 6132 8740 6196 8804
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 3740 8528 3804 8532
rect 3740 8472 3754 8528
rect 3754 8472 3804 8528
rect 3740 8468 3804 8472
rect 10916 8332 10980 8396
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 22876 8060 22940 8124
rect 18092 7788 18156 7852
rect 19380 7788 19444 7852
rect 20116 7712 20180 7716
rect 20116 7656 20130 7712
rect 20130 7656 20180 7712
rect 20116 7652 20180 7656
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10916 7380 10980 7444
rect 20116 7168 20180 7172
rect 20116 7112 20166 7168
rect 20166 7112 20180 7168
rect 20116 7108 20180 7112
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 21772 6972 21836 7036
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 5396 6428 5460 6492
rect 3372 6156 3436 6220
rect 15516 6488 15580 6492
rect 15516 6432 15530 6488
rect 15530 6432 15580 6488
rect 15516 6428 15580 6432
rect 20116 6292 20180 6356
rect 23060 6352 23124 6356
rect 23060 6296 23110 6352
rect 23110 6296 23124 6352
rect 23060 6292 23124 6296
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 6316 5884 6380 5948
rect 6868 5884 6932 5948
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 14228 5536 14292 5540
rect 14228 5480 14278 5536
rect 14278 5480 14292 5536
rect 14228 5476 14292 5480
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 3004 5128 3068 5132
rect 3004 5072 3018 5128
rect 3018 5072 3068 5128
rect 3004 5068 3068 5072
rect 17908 5068 17972 5132
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 2084 4796 2148 4860
rect 14228 4796 14292 4860
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 20300 4796 20364 4860
rect 19196 4660 19260 4724
rect 23612 4660 23676 4724
rect 7788 4448 7852 4452
rect 7788 4392 7802 4448
rect 7802 4392 7852 4448
rect 7788 4388 7852 4392
rect 20668 4388 20732 4452
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 8156 4252 8220 4316
rect 22876 3980 22940 4044
rect 23428 3980 23492 4044
rect 6500 3844 6564 3908
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 22140 3708 22204 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 8156 3088 8220 3092
rect 8156 3032 8170 3088
rect 8170 3032 8220 3088
rect 8156 3028 8220 3032
rect 16436 3028 16500 3092
rect 23612 2892 23676 2956
rect 22508 2756 22572 2820
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 11100 2620 11164 2684
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 3740 2136 3804 2140
rect 3740 2080 3754 2136
rect 3754 2080 3804 2136
rect 3740 2076 3804 2080
rect 21772 606 21836 644
rect 21772 580 21822 606
rect 21822 580 21836 606
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 9627 21452 9693 21453
rect 9627 21388 9628 21452
rect 9692 21388 9693 21452
rect 9627 21387 9693 21388
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 9630 20365 9690 21387
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 9627 20364 9693 20365
rect 9627 20300 9628 20364
rect 9692 20300 9693 20364
rect 9627 20299 9693 20300
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 2083 18052 2149 18053
rect 2083 17988 2084 18052
rect 2148 17988 2149 18052
rect 2083 17987 2149 17988
rect 2086 7938 2146 17987
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 6315 16964 6381 16965
rect 6315 16900 6316 16964
rect 6380 16900 6381 16964
rect 6315 16899 6381 16900
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 2451 16284 2517 16285
rect 2451 16220 2452 16284
rect 2516 16220 2517 16284
rect 2451 16219 2517 16220
rect 2267 13428 2333 13429
rect 2267 13364 2268 13428
rect 2332 13364 2333 13428
rect 2267 13363 2333 13364
rect 2270 12205 2330 13363
rect 2267 12204 2333 12205
rect 2267 12140 2268 12204
rect 2332 12140 2333 12204
rect 2267 12139 2333 12140
rect 2454 10437 2514 16219
rect 5211 15468 5277 15469
rect 5211 15404 5212 15468
rect 5276 15404 5277 15468
rect 5211 15403 5277 15404
rect 2635 14516 2701 14517
rect 2635 14452 2636 14516
rect 2700 14452 2701 14516
rect 2635 14451 2701 14452
rect 2638 12069 2698 14451
rect 2635 12068 2701 12069
rect 2635 12004 2636 12068
rect 2700 12004 2701 12068
rect 2635 12003 2701 12004
rect 2451 10436 2517 10437
rect 2451 10372 2452 10436
rect 2516 10372 2517 10436
rect 2451 10371 2517 10372
rect 5214 9893 5274 15403
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 6131 12340 6197 12341
rect 6131 12276 6132 12340
rect 6196 12276 6197 12340
rect 6131 12275 6197 12276
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 6134 11525 6194 12275
rect 6131 11524 6197 11525
rect 6131 11460 6132 11524
rect 6196 11460 6197 11524
rect 6131 11459 6197 11460
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5211 9892 5277 9893
rect 5211 9828 5212 9892
rect 5276 9828 5277 9892
rect 5211 9827 5277 9828
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 6134 8805 6194 11459
rect 6131 8804 6197 8805
rect 6131 8740 6132 8804
rect 6196 8740 6197 8804
rect 6131 8739 6197 8740
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 3739 8532 3805 8533
rect 3739 8468 3740 8532
rect 3804 8468 3805 8532
rect 3739 8467 3805 8468
rect 2086 4861 2146 7702
rect 3371 6220 3437 6221
rect 3371 6156 3372 6220
rect 3436 6156 3437 6220
rect 3371 6155 3437 6156
rect 2083 4860 2149 4861
rect 2083 4796 2084 4860
rect 2148 4796 2149 4860
rect 2083 4795 2149 4796
rect 3374 2498 3434 6155
rect 3742 2141 3802 8467
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 6318 5949 6378 16899
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 6683 15060 6749 15061
rect 6683 14996 6684 15060
rect 6748 14996 6749 15060
rect 6683 14995 6749 14996
rect 6686 12341 6746 14995
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 6683 12340 6749 12341
rect 6683 12276 6684 12340
rect 6748 12276 6749 12340
rect 6683 12275 6749 12276
rect 10277 11456 10597 12480
rect 14944 25056 15264 25616
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19379 25260 19445 25261
rect 19379 25196 19380 25260
rect 19444 25196 19445 25260
rect 19379 25195 19445 25196
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 18643 13972 18709 13973
rect 18643 13908 18644 13972
rect 18708 13908 18709 13972
rect 18643 13907 18709 13908
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 11099 11932 11165 11933
rect 11099 11868 11100 11932
rect 11164 11868 11165 11932
rect 11099 11867 11165 11868
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 6499 8940 6565 8941
rect 6499 8876 6500 8940
rect 6564 8876 6565 8940
rect 6499 8875 6565 8876
rect 6315 5948 6381 5949
rect 6315 5884 6316 5948
rect 6380 5884 6381 5948
rect 6315 5883 6381 5884
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 6502 3909 6562 8875
rect 10277 8192 10597 9216
rect 11102 9213 11162 11867
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 11099 9212 11165 9213
rect 11099 9148 11100 9212
rect 11164 9148 11165 9212
rect 11099 9147 11165 9148
rect 14944 8736 15264 9760
rect 18646 9621 18706 13907
rect 19195 11932 19261 11933
rect 19195 11868 19196 11932
rect 19260 11868 19261 11932
rect 19195 11867 19261 11868
rect 18643 9620 18709 9621
rect 18643 9556 18644 9620
rect 18708 9556 18709 9620
rect 18643 9555 18709 9556
rect 19011 9620 19077 9621
rect 19011 9556 19012 9620
rect 19076 9556 19077 9620
rect 19011 9555 19077 9556
rect 18827 9348 18893 9349
rect 18827 9284 18828 9348
rect 18892 9284 18893 9348
rect 18827 9283 18893 9284
rect 18830 9210 18890 9283
rect 19014 9210 19074 9555
rect 18830 9150 19074 9210
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 10915 8396 10981 8397
rect 10915 8332 10916 8396
rect 10980 8332 10981 8396
rect 10915 8331 10981 8332
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10918 7445 10978 8331
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 10915 7444 10981 7445
rect 10915 7380 10916 7444
rect 10980 7380 10981 7444
rect 10915 7379 10981 7380
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 6867 5948 6933 5949
rect 6867 5898 6868 5948
rect 6932 5898 6933 5948
rect 10277 4928 10597 5952
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14227 5540 14293 5541
rect 14227 5476 14228 5540
rect 14292 5476 14293 5540
rect 14227 5475 14293 5476
rect 14230 5218 14290 5475
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 8155 4316 8221 4317
rect 8155 4252 8156 4316
rect 8220 4252 8221 4316
rect 8155 4251 8221 4252
rect 6499 3908 6565 3909
rect 6499 3844 6500 3908
rect 6564 3844 6565 3908
rect 8158 3858 8218 4251
rect 6499 3843 6565 3844
rect 10277 3840 10597 4864
rect 14227 4860 14293 4861
rect 14227 4796 14228 4860
rect 14292 4796 14293 4860
rect 14227 4795 14293 4796
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 3739 2140 3805 2141
rect 3739 2076 3740 2140
rect 3804 2076 3805 2140
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 14230 3178 14290 4795
rect 14944 4384 15264 5408
rect 19198 4725 19258 11867
rect 19382 7853 19442 25195
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 23979 17100 24045 17101
rect 23979 17036 23980 17100
rect 24044 17036 24045 17100
rect 23979 17035 24045 17036
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 21587 14652 21653 14653
rect 21587 14588 21588 14652
rect 21652 14588 21653 14652
rect 21587 14587 21653 14588
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 20299 10300 20365 10301
rect 20299 10236 20300 10300
rect 20364 10236 20365 10300
rect 20299 10235 20365 10236
rect 20115 9756 20181 9757
rect 20115 9692 20116 9756
rect 20180 9692 20181 9756
rect 20115 9691 20181 9692
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19379 7852 19445 7853
rect 19379 7788 19380 7852
rect 19444 7788 19445 7852
rect 19379 7787 19445 7788
rect 19610 7104 19930 8128
rect 20118 7717 20178 9691
rect 20115 7716 20181 7717
rect 20115 7652 20116 7716
rect 20180 7652 20181 7716
rect 20115 7651 20181 7652
rect 20115 7172 20181 7173
rect 20115 7108 20116 7172
rect 20180 7108 20181 7172
rect 20115 7107 20181 7108
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 20118 6357 20178 7107
rect 20115 6356 20181 6357
rect 20115 6292 20116 6356
rect 20180 6292 20181 6356
rect 20115 6291 20181 6292
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 20302 5898 20362 10235
rect 21590 10029 21650 14587
rect 23243 14244 23309 14245
rect 23243 14180 23244 14244
rect 23308 14180 23309 14244
rect 23243 14179 23309 14180
rect 23246 12205 23306 14179
rect 23982 13565 24042 17035
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 23979 13564 24045 13565
rect 23979 13500 23980 13564
rect 24044 13500 24045 13564
rect 23979 13499 24045 13500
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 23427 12884 23493 12885
rect 23427 12820 23428 12884
rect 23492 12820 23493 12884
rect 23427 12819 23493 12820
rect 23243 12204 23309 12205
rect 23243 12140 23244 12204
rect 23308 12140 23309 12204
rect 23243 12139 23309 12140
rect 23059 11388 23125 11389
rect 23059 11324 23060 11388
rect 23124 11324 23125 11388
rect 23059 11323 23125 11324
rect 21587 10028 21653 10029
rect 21587 9964 21588 10028
rect 21652 9964 21653 10028
rect 21587 9963 21653 9964
rect 23062 9349 23122 11323
rect 22507 9348 22573 9349
rect 22507 9284 22508 9348
rect 22572 9284 22573 9348
rect 22507 9283 22573 9284
rect 23059 9348 23125 9349
rect 23059 9284 23060 9348
rect 23124 9284 23125 9348
rect 23059 9283 23125 9284
rect 21771 7036 21837 7037
rect 21771 6972 21772 7036
rect 21836 6972 21837 7036
rect 21771 6971 21837 6972
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19195 4724 19261 4725
rect 19195 4660 19196 4724
rect 19260 4660 19261 4724
rect 19195 4659 19261 4660
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 11099 2684 11165 2685
rect 11099 2620 11100 2684
rect 11164 2620 11165 2684
rect 11099 2619 11165 2620
rect 11102 2498 11162 2619
rect 14944 2208 15264 3232
rect 19610 3840 19930 4864
rect 20302 4861 20362 5662
rect 20299 4860 20365 4861
rect 20299 4796 20300 4860
rect 20364 4796 20365 4860
rect 20299 4795 20365 4796
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 3739 2075 3805 2076
rect 21774 645 21834 6971
rect 22510 2821 22570 9283
rect 22875 8124 22941 8125
rect 22875 8060 22876 8124
rect 22940 8060 22941 8124
rect 22875 8059 22941 8060
rect 22878 4045 22938 8059
rect 23062 6357 23122 9283
rect 23059 6356 23125 6357
rect 23059 6292 23060 6356
rect 23124 6292 23125 6356
rect 23059 6291 23125 6292
rect 23430 4045 23490 12819
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 23611 10300 23677 10301
rect 23611 10236 23612 10300
rect 23676 10236 23677 10300
rect 23611 10235 23677 10236
rect 23614 4725 23674 10235
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 23611 4724 23677 4725
rect 23611 4660 23612 4724
rect 23676 4660 23677 4724
rect 23611 4659 23677 4660
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 22875 4044 22941 4045
rect 22875 3980 22876 4044
rect 22940 3980 22941 4044
rect 22875 3979 22941 3980
rect 23427 4044 23493 4045
rect 23427 3980 23428 4044
rect 23492 3980 23493 4044
rect 23427 3979 23493 3980
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 23611 2892 23612 2942
rect 23676 2892 23677 2942
rect 23611 2891 23677 2892
rect 22507 2820 22573 2821
rect 22507 2756 22508 2820
rect 22572 2756 22573 2820
rect 22507 2755 22573 2756
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 21771 644 21837 645
rect 21771 580 21772 644
rect 21836 580 21837 644
rect 21771 579 21837 580
<< via4 >>
rect 1998 7702 2234 7938
rect 2918 5132 3154 5218
rect 2918 5068 3004 5132
rect 3004 5068 3068 5132
rect 3068 5068 3154 5132
rect 2918 4982 3154 5068
rect 3286 2262 3522 2498
rect 5310 6492 5546 6578
rect 5310 6428 5396 6492
rect 5396 6428 5460 6492
rect 5460 6428 5546 6492
rect 5310 6342 5546 6428
rect 18006 7852 18242 7938
rect 18006 7788 18092 7852
rect 18092 7788 18156 7852
rect 18156 7788 18242 7852
rect 18006 7702 18242 7788
rect 6782 5884 6868 5898
rect 6868 5884 6932 5898
rect 6932 5884 7018 5898
rect 6782 5662 7018 5884
rect 15430 6492 15666 6578
rect 15430 6428 15516 6492
rect 15516 6428 15580 6492
rect 15580 6428 15666 6492
rect 15430 6342 15666 6428
rect 14142 4982 14378 5218
rect 7702 4452 7938 4538
rect 7702 4388 7788 4452
rect 7788 4388 7852 4452
rect 7852 4388 7938 4452
rect 7702 4302 7938 4388
rect 8070 3622 8306 3858
rect 8070 3092 8306 3178
rect 8070 3028 8156 3092
rect 8156 3028 8220 3092
rect 8220 3028 8306 3092
rect 8070 2942 8306 3028
rect 17822 5132 18058 5218
rect 17822 5068 17908 5132
rect 17908 5068 17972 5132
rect 17972 5068 18058 5132
rect 17822 4982 18058 5068
rect 20214 5662 20450 5898
rect 14142 2942 14378 3178
rect 11014 2262 11250 2498
rect 20582 4452 20818 4538
rect 20582 4388 20668 4452
rect 20668 4388 20732 4452
rect 20732 4388 20818 4452
rect 20582 4302 20818 4388
rect 16350 3092 16586 3178
rect 16350 3028 16436 3092
rect 16436 3028 16500 3092
rect 16500 3028 16586 3092
rect 16350 2942 16586 3028
rect 22054 3772 22290 3858
rect 22054 3708 22140 3772
rect 22140 3708 22204 3772
rect 22204 3708 22290 3772
rect 22054 3622 22290 3708
rect 23526 2956 23762 3178
rect 23526 2942 23612 2956
rect 23612 2942 23676 2956
rect 23676 2942 23762 2956
<< metal5 >>
rect 1956 7938 18284 7980
rect 1956 7702 1998 7938
rect 2234 7702 18006 7938
rect 18242 7702 18284 7938
rect 1956 7660 18284 7702
rect 5268 6578 15708 6620
rect 5268 6342 5310 6578
rect 5546 6342 15430 6578
rect 15666 6342 15708 6578
rect 5268 6300 15708 6342
rect 6740 5898 20492 5940
rect 6740 5662 6782 5898
rect 7018 5662 20214 5898
rect 20450 5662 20492 5898
rect 6740 5620 20492 5662
rect 2876 5218 18100 5260
rect 2876 4982 2918 5218
rect 3154 4982 14142 5218
rect 14378 4982 17822 5218
rect 18058 4982 18100 5218
rect 2876 4940 18100 4982
rect 7660 4538 20860 4580
rect 7660 4302 7702 4538
rect 7938 4302 20582 4538
rect 20818 4302 20860 4538
rect 7660 4260 20860 4302
rect 8028 3858 22332 3900
rect 8028 3622 8070 3858
rect 8306 3622 22054 3858
rect 22290 3622 22332 3858
rect 8028 3580 22332 3622
rect 8028 3178 14420 3220
rect 8028 2942 8070 3178
rect 8306 2942 14142 3178
rect 14378 2942 14420 3178
rect 8028 2900 14420 2942
rect 16308 3178 23804 3220
rect 16308 2942 16350 3178
rect 16586 2942 23526 3178
rect 23762 2942 23804 3178
rect 16308 2900 23804 2942
rect 3244 2498 11292 2540
rect 3244 2262 3286 2498
rect 3522 2262 11014 2498
rect 11250 2262 11292 2498
rect 3244 2220 11292 2262
use scs8hd_fill_2  FILLER_1_9 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_5.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use scs8hd_conb_1  _047_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_13
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l2_in_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_2_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_55 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6164 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_51
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_85
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_81
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _083_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_116
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_121
timestamp 1586364061
transform 1 0 12236 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_152
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 1786 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_177
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_181
timestamp 1586364061
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _127_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_39.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_224
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_228
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _125_
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _126_
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_243
timestamp 1586364061
transform 1 0 23460 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_239
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23644 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_4  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23736 0 1 2720
box -38 -48 590 592
use scs8hd_buf_4  mux_bottom_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_256
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_252
timestamp 1586364061
transform 1 0 24288 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_255
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_19.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 590 592
use scs8hd_buf_2  _124_
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_270
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_271 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_267
timestamp 1586364061
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_274
timestamp 1586364061
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_38
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_42
timestamp 1586364061
transform 1 0 4968 0 -1 3808
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_191
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_195
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 590 592
use scs8hd_buf_4  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_21.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22540 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_221
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_225
timestamp 1586364061
transform 1 0 21804 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24472 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_252
timestamp 1586364061
transform 1 0 24288 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_256
timestamp 1586364061
transform 1 0 24656 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 25024 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_264
timestamp 1586364061
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25576 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_272
timestamp 1586364061
transform 1 0 26128 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_268
timestamp 1586364061
transform 1 0 25760 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5244 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_78
timestamp 1586364061
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_82
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_134
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_151
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_155
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_158
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_track_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_190
timestamp 1586364061
transform 1 0 18584 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_21.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_212
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_19.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_222
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_23.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_251
timestamp 1586364061
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_255
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 24932 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 26220 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_263
timestamp 1586364061
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_267
timestamp 1586364061
transform 1 0 25668 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_271
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_275
timestamp 1586364061
transform 1 0 26404 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_58
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_62
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_75
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_79
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9752 0 -1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_137
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_148
timestamp 1586364061
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14904 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_21.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_179
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_183
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_189
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_193
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_21.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_19.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22356 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_229
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_252
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_257
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 314 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 25024 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_264
timestamp 1586364061
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_268
timestamp 1586364061
transform 1 0 25760 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_108
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_134
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_151
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_172
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_176
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_21.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_180
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_188
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_192
timestamp 1586364061
transform 1 0 18768 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_216
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_19.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_223
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 24564 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23828 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24196 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_249
timestamp 1586364061
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_253
timestamp 1586364061
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_259
timestamp 1586364061
transform 1 0 24932 0 1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_265 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_13
timestamp 1586364061
transform 1 0 2300 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_49
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_67
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_79
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_96
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_100
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_100
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_164
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_162
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16192 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_buf_4  mux_right_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_190
timestamp 1586364061
transform 1 0 18584 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_23.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_23.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 1786 592
use scs8hd_buf_4  mux_bottom_track_21.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_204
timestamp 1586364061
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_208
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_218
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_222
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_225
timestamp 1586364061
transform 1 0 21804 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_221
timestamp 1586364061
transform 1 0 21436 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_19.mux_l1_in_1_
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_19.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1786 592
use scs8hd_buf_4  mux_right_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_241
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_255 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_264
timestamp 1586364061
transform 1 0 25392 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_7_268
timestamp 1586364061
transform 1 0 25760 0 1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_6_267
timestamp 1586364061
transform 1 0 25668 0 -1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_276
timestamp 1586364061
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1472 0 -1 7072
box -38 -48 1786 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_29
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_53
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_57
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_61
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_77
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10304 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_126
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_132
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_23.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18124 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_179
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_183
timestamp 1586364061
transform 1 0 17940 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_187
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _121_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22632 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21620 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_219
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_225
timestamp 1586364061
transform 1 0 21804 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_229
timestamp 1586364061
transform 1 0 22172 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_233
timestamp 1586364061
transform 1 0 22540 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_253
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 25116 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_265
timestamp 1586364061
transform 1 0 25484 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_273
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _049_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_65
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_69
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_131
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_154
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_158
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 314 592
use scs8hd_buf_2  _122_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_23.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_216
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_266
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_270
timestamp 1586364061
transform 1 0 25944 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_276
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_12
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_29
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_4  mux_left_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_87
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_115
timestamp 1586364061
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_139
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_13.mux_l1_in_1_
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_171
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_175
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_23.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_187
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_191
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_212
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_219
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_4  mux_bottom_track_37.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24288 0 -1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_243
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_43
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_68
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_72
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_85
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_89
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_131
timestamp 1586364061
transform 1 0 13156 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_201
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_218
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21528 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_235
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 590 592
use scs8hd_buf_4  mux_bottom_track_35.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_251
timestamp 1586364061
transform 1 0 24196 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_255
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_263
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_267
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_275
timestamp 1586364061
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_16
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_22
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_26
timestamp 1586364061
transform 1 0 3496 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_32.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_69
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_118
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_122
timestamp 1586364061
transform 1 0 12328 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_39.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_167
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_171
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_175
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20332 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_207
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_234
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_track_37.mux_l1_in_0_
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_242
timestamp 1586364061
transform 1 0 23368 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_261
timestamp 1586364061
transform 1 0 25116 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_273
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_16
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_28
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_24
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_20
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_25
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5980 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_52
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_49
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 7912 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_72
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_76
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_116
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_124
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_134
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_139
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_152
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_39.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15364 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_174
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_188
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_195
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_191
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_192
timestamp 1586364061
transform 1 0 18768 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_14_204
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_199
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _120_
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_216
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_39.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21436 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_15.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21252 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_233
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_237
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_244
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_240
timestamp 1586364061
transform 1 0 23184 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_241
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_37.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24012 0 1 9248
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_37.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_13_262
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 25576 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_267
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_3_
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_9
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_44
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 1786 592
use scs8hd_buf_4  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_70
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_39.mux_l1_in_0_
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _119_
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_203
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_207
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_211
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_218
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_35.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_222
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_37.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_264
timestamp 1586364061
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_268
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4968 0 -1 11424
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_16_40
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_109
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_135
timestamp 1586364061
transform 1 0 13524 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_139
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_147
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_160
timestamp 1586364061
transform 1 0 15824 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_177
timestamp 1586364061
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18124 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17572 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_181
timestamp 1586364061
transform 1 0 17756 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_195
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _118_
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_35.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22724 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22540 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21620 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_221
timestamp 1586364061
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_225
timestamp 1586364061
transform 1 0 21804 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_229
timestamp 1586364061
transform 1 0 22172 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_254
timestamp 1586364061
transform 1 0 24472 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 25208 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25024 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_258
timestamp 1586364061
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_266
timestamp 1586364061
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_50
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_54
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_58
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_76
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_80
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_33.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_129
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_11.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_163
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _123_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_188
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_192
timestamp 1586364061
transform 1 0 18768 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_195
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_199
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _117_
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_222
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_226
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_35.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_266
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_270
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1786 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_26
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_75
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_87
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_99
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_103
timestamp 1586364061
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_track_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_11.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_160
timestamp 1586364061
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_164
timestamp 1586364061
transform 1 0 16192 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_168
timestamp 1586364061
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_189
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_193
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 22264 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_232
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_237
timestamp 1586364061
transform 1 0 22908 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23368 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24380 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23184 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_255
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_265
timestamp 1586364061
transform 1 0 25484 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_273
timestamp 1586364061
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_9
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_17
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_25
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_21
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_3_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_58
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 866 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_79
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_70
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_19_102
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_116
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_112
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_33.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_152
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_11.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_170
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_176
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_193
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_201
timestamp 1586364061
transform 1 0 19596 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_200
timestamp 1586364061
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_227
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_223
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_229
timestamp 1586364061
transform 1 0 22172 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_235
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22540 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22172 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _116_
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_35.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22724 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_31.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23920 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24656 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_239
timestamp 1586364061
transform 1 0 23092 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_254
timestamp 1586364061
transform 1 0 24472 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_266
timestamp 1586364061
transform 1 0 25576 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_258
timestamp 1586364061
transform 1 0 24840 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_264
timestamp 1586364061
transform 1 0 25392 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_261
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25024 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 25208 0 -1 13600
box -38 -48 406 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_273
timestamp 1586364061
transform 1 0 26220 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 26036 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 1786 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_26
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_43
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_47
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_96
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_100
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_146
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_169
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_173
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 774 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_181
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_191
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_195
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_21_218
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_222
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24104 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_conb_1  _055_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_58
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_3_
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_75
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_79
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10580 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_112
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_116
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 13708 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12144 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_133
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 406 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_157
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 15732 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_161
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_184
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_188
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_191
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 590 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_27.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_199
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22540 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_230
timestamp 1586364061
transform 1 0 22264 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 24472 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_252
timestamp 1586364061
transform 1 0 24288 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_256
timestamp 1586364061
transform 1 0 24656 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_track_31.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25024 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_266
timestamp 1586364061
transform 1 0 25576 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5244 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_43
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l1_in_3_
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_104
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_108
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 774 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_140
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_148
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 590 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_27.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_23_199
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_27.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_224
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_234
timestamp 1586364061
transform 1 0 22632 0 1 14688
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_31.mux_l1_in_0_
timestamp 1586364061
transform 1 0 24380 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 24196 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23828 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_249
timestamp 1586364061
transform 1 0 24012 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_262
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_23_274
timestamp 1586364061
transform 1 0 26312 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_24_9
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4324 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use scs8hd_conb_1  _066_
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_48
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_55
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_63
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_79
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 130 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_24_101
timestamp 1586364061
transform 1 0 10396 0 -1 15776
box -38 -48 130 592
use scs8hd_conb_1  _054_
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_140
timestamp 1586364061
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_conb_1  _062_
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_171
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_177
timestamp 1586364061
transform 1 0 17388 0 -1 15776
box -38 -48 774 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_27.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_189
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_track_27.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22816 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_234
timestamp 1586364061
transform 1 0 22632 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_238
timestamp 1586364061
transform 1 0 23000 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_31.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23920 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_242
timestamp 1586364061
transform 1 0 23368 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_247
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_267
timestamp 1586364061
transform 1 0 25668 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 406 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_19
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 3036 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_23
timestamp 1586364061
transform 1 0 3220 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_28
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_41
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_45
timestamp 1586364061
transform 1 0 5244 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_49
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_25_94
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_97
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_139
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_151
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _056_
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_163
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_168
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _059_
timestamp 1586364061
transform 1 0 18952 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_180
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_192
timestamp 1586364061
transform 1 0 18768 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 774 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_29.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_209
timestamp 1586364061
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_213
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_31.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_264
timestamp 1586364061
transform 1 0 25392 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_268
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_11
timestamp 1586364061
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2300 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_23
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_35
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_53
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_65
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_77
timestamp 1586364061
transform 1 0 8188 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_99
timestamp 1586364061
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_103
timestamp 1586364061
transform 1 0 10580 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_115
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_127
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_139
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_152
timestamp 1586364061
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_162
timestamp 1586364061
transform 1 0 16008 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_168
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_176
timestamp 1586364061
transform 1 0 17296 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_conb_1  _057_
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 314 592
use scs8hd_conb_1  _063_
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_182
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_195
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 774 592
use scs8hd_conb_1  _064_
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 314 592
use scs8hd_conb_1  _065_
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21068 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_207
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_225
timestamp 1586364061
transform 1 0 21804 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_219
timestamp 1586364061
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_29.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 866 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 21436 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_229
timestamp 1586364061
transform 1 0 22172 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22356 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_29.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22540 0 -1 16864
box -38 -48 1786 592
use scs8hd_buf_4  mux_bottom_track_29.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_252
timestamp 1586364061
transform 1 0 24288 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_251
timestamp 1586364061
transform 1 0 24196 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_263
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_264
timestamp 1586364061
transform 1 0 25392 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 25484 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 25024 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_275
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_267
timestamp 1586364061
transform 1 0 25668 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_272
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 406 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_198
timestamp 1586364061
transform 1 0 19320 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _061_
timestamp 1586364061
transform 1 0 19504 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_203
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_211
timestamp 1586364061
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 21344 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_29.mux_l1_in_0_
timestamp 1586364061
transform 1 0 22356 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_219
timestamp 1586364061
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_223
timestamp 1586364061
transform 1 0 21620 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_229
timestamp 1586364061
transform 1 0 22172 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_240
timestamp 1586364061
transform 1 0 23184 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_28_252
timestamp 1586364061
transform 1 0 24288 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_259
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 774 592
use scs8hd_conb_1  _058_
timestamp 1586364061
transform 1 0 20148 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_204
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_210
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 1142 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 22540 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_222
timestamp 1586364061
transform 1 0 21528 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_29_230
timestamp 1586364061
transform 1 0 22264 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 774 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 23828 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_249
timestamp 1586364061
transform 1 0 24012 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_259
timestamp 1586364061
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_263
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_29_275
timestamp 1586364061
transform 1 0 26404 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_conb_1  _060_
timestamp 1586364061
transform 1 0 22448 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_231
timestamp 1586364061
transform 1 0 22356 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_235
timestamp 1586364061
transform 1 0 22724 0 -1 19040
box -38 -48 774 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 23460 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_247
timestamp 1586364061
transform 1 0 23828 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_259
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_271
timestamp 1586364061
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_259
timestamp 1586364061
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_263
timestamp 1586364061
transform 1 0 25300 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_31_275
timestamp 1586364061
transform 1 0 26404 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_conb_1  _067_
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_258
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_270
timestamp 1586364061
transform 1 0 25944 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2594 0 2650 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 3146 0 3202 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3790 0 3846 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 4342 0 4398 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal3 s 0 26936 480 27056 6 ccff_head
port 8 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 19728 480 19848 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 20408 480 20528 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 21088 480 21208 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 23672 480 23792 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 24352 480 24472 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 25032 480 25152 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 25576 480 25696 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 16464 480 16584 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 17144 480 17264 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 17824 480 17944 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 18504 480 18624 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 6672 480 6792 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 8712 480 8832 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 9392 480 9512 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 9936 480 10056 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 10616 480 10736 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 11296 480 11416 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 12656 480 12776 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 1504 480 1624 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 2864 480 2984 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 4088 480 4208 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 5448 480 5568 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 6128 480 6248 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 27520 20952 28000 21072 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 27520 21496 28000 21616 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 27520 22176 28000 22296 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 27520 22856 28000 22976 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 27520 23536 28000 23656 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 27520 24896 28000 25016 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 27520 25576 28000 25696 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 27520 26256 28000 26376 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 27520 15512 28000 15632 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 27520 16192 28000 16312 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 27520 16872 28000 16992 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 27520 17552 28000 17672 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 27520 18232 28000 18352 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 27520 18912 28000 19032 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 27520 280 28000 400 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 27520 6944 28000 7064 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 27520 7488 28000 7608 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 27520 10208 28000 10328 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 27520 10888 28000 11008 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 27520 11568 28000 11688 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 27520 12928 28000 13048 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 27520 824 28000 944 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 27520 1504 28000 1624 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 27520 2184 28000 2304 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 27520 2864 28000 2984 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 27520 3544 28000 3664 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 27520 4224 28000 4344 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 27520 5584 28000 5704 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 27520 6264 28000 6384 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 14830 0 14886 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 22374 0 22430 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 23018 0 23074 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 23570 0 23626 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 24122 0 24178 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 25318 0 25374 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 25870 0 25926 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 27618 0 27674 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 18878 0 18934 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 19522 0 19578 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 21270 0 21326 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 21822 0 21878 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal3 s 0 26256 480 26376 6 left_top_grid_pin_1_
port 130 nsew default input
rlabel metal3 s 0 27616 480 27736 6 prog_clk
port 131 nsew default input
rlabel metal3 s 27520 26936 28000 27056 6 right_top_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 133 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 27736
<< end >>
