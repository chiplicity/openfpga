magic
tech EFS8A
magscale 1 2
timestamp 1602525323
<< locali >>
rect 9643 35785 9781 35819
rect 7015 34153 7021 34187
rect 7015 34085 7049 34153
rect 11287 34017 11322 34051
rect 9131 33303 9165 33371
rect 9131 33269 9137 33303
rect 4905 32827 4939 32929
rect 4715 32215 4749 32283
rect 4715 32181 4721 32215
rect 8435 31841 8470 31875
rect 3433 29087 3467 29257
rect 4307 28985 4445 29019
rect 3111 28713 3157 28747
rect 6555 28713 6561 28747
rect 6555 28645 6589 28713
rect 2915 28577 3042 28611
rect 11287 28577 11322 28611
rect 2283 28169 2421 28203
rect 3295 28169 3433 28203
rect 4755 27557 4800 27591
rect 10051 25449 10057 25483
rect 10051 25381 10085 25449
rect 11287 24225 11322 24259
rect 4169 23545 4261 23579
rect 5359 23511 5393 23579
rect 5359 23477 5365 23511
rect 8159 23137 8194 23171
rect 10735 23137 10770 23171
rect 4813 22491 4847 22661
rect 11287 22049 11322 22083
rect 4439 20009 4445 20043
rect 4439 19941 4473 20009
rect 7751 18921 7757 18955
rect 7751 18853 7785 18921
rect 3709 18139 3743 18377
rect 4905 16983 4939 17085
rect 5543 16745 5549 16779
rect 5543 16677 5577 16745
rect 9631 16609 9758 16643
rect 10735 16609 10770 16643
rect 5641 15963 5675 16133
rect 6279 15657 6285 15691
rect 6279 15589 6313 15657
rect 6469 15011 6503 15113
rect 2915 14433 3042 14467
rect 11471 14433 11506 14467
rect 2915 13345 3042 13379
rect 5089 13175 5123 13345
rect 10735 10081 10862 10115
rect 11287 8993 11322 9027
rect 8619 7905 8654 7939
rect 11287 7905 11322 7939
rect 3157 7191 3191 7293
rect 12851 3553 12886 3587
<< viali >>
rect 9781 35785 9815 35819
rect 8493 35649 8527 35683
rect 6904 35581 6938 35615
rect 9540 35581 9574 35615
rect 9965 35581 9999 35615
rect 7849 35513 7883 35547
rect 8033 35513 8067 35547
rect 8125 35513 8159 35547
rect 4905 35445 4939 35479
rect 6975 35445 7009 35479
rect 7389 35445 7423 35479
rect 4215 35241 4249 35275
rect 8033 35241 8067 35275
rect 9873 35241 9907 35275
rect 5273 35173 5307 35207
rect 7113 35173 7147 35207
rect 4123 35105 4157 35139
rect 8493 35105 8527 35139
rect 9689 35105 9723 35139
rect 5181 35037 5215 35071
rect 7021 35037 7055 35071
rect 7665 35037 7699 35071
rect 5733 34969 5767 35003
rect 8677 34969 8711 35003
rect 4813 34901 4847 34935
rect 6837 34901 6871 34935
rect 9045 34901 9079 34935
rect 3893 34697 3927 34731
rect 5733 34697 5767 34731
rect 6009 34697 6043 34731
rect 7757 34697 7791 34731
rect 9689 34697 9723 34731
rect 12725 34697 12759 34731
rect 3617 34629 3651 34663
rect 9229 34629 9263 34663
rect 4813 34561 4847 34595
rect 10149 34561 10183 34595
rect 3709 34493 3743 34527
rect 6837 34493 6871 34527
rect 12541 34493 12575 34527
rect 13093 34493 13127 34527
rect 4721 34425 4755 34459
rect 5134 34425 5168 34459
rect 6561 34425 6595 34459
rect 7158 34425 7192 34459
rect 8677 34425 8711 34459
rect 8769 34425 8803 34459
rect 4261 34357 4295 34391
rect 8033 34357 8067 34391
rect 8401 34357 8435 34391
rect 4905 34153 4939 34187
rect 5641 34153 5675 34187
rect 6561 34153 6595 34187
rect 7021 34153 7055 34187
rect 7573 34153 7607 34187
rect 9781 34153 9815 34187
rect 9321 34085 9355 34119
rect 4721 34017 4755 34051
rect 5089 34017 5123 34051
rect 8401 34017 8435 34051
rect 9965 34017 9999 34051
rect 10149 34017 10183 34051
rect 10701 34017 10735 34051
rect 11253 34017 11287 34051
rect 3341 33949 3375 33983
rect 6653 33949 6687 33983
rect 8585 33881 8619 33915
rect 8953 33813 8987 33847
rect 11391 33813 11425 33847
rect 4629 33609 4663 33643
rect 8493 33609 8527 33643
rect 9965 33609 9999 33643
rect 10425 33541 10459 33575
rect 4353 33473 4387 33507
rect 8769 33473 8803 33507
rect 11529 33473 11563 33507
rect 3157 33405 3191 33439
rect 3525 33405 3559 33439
rect 3709 33405 3743 33439
rect 3985 33405 4019 33439
rect 4813 33405 4847 33439
rect 6837 33405 6871 33439
rect 8033 33405 8067 33439
rect 10609 33405 10643 33439
rect 10977 33405 11011 33439
rect 5134 33337 5168 33371
rect 6193 33337 6227 33371
rect 6561 33337 6595 33371
rect 7158 33337 7192 33371
rect 5733 33269 5767 33303
rect 7757 33269 7791 33303
rect 9137 33269 9171 33303
rect 9689 33269 9723 33303
rect 10609 33269 10643 33303
rect 4997 33065 5031 33099
rect 6653 33065 6687 33099
rect 11437 33065 11471 33099
rect 3157 32997 3191 33031
rect 5365 32997 5399 33031
rect 7066 32997 7100 33031
rect 9965 32997 9999 33031
rect 2697 32929 2731 32963
rect 2973 32929 3007 32963
rect 4905 32929 4939 32963
rect 8560 32929 8594 32963
rect 9413 32929 9447 32963
rect 11345 32929 11379 32963
rect 11805 32929 11839 32963
rect 4353 32861 4387 32895
rect 5273 32861 5307 32895
rect 5641 32861 5675 32895
rect 6745 32861 6779 32895
rect 9873 32861 9907 32895
rect 10333 32861 10367 32895
rect 12909 32861 12943 32895
rect 4629 32793 4663 32827
rect 4905 32793 4939 32827
rect 7665 32725 7699 32759
rect 8631 32725 8665 32759
rect 9045 32725 9079 32759
rect 11253 32725 11287 32759
rect 2881 32521 2915 32555
rect 9965 32521 9999 32555
rect 11621 32521 11655 32555
rect 12173 32521 12207 32555
rect 8125 32453 8159 32487
rect 7849 32385 7883 32419
rect 8677 32385 8711 32419
rect 13001 32385 13035 32419
rect 3893 32317 3927 32351
rect 4353 32317 4387 32351
rect 9597 32317 9631 32351
rect 10425 32317 10459 32351
rect 12449 32317 12483 32351
rect 12909 32317 12943 32351
rect 6285 32249 6319 32283
rect 7205 32249 7239 32283
rect 7297 32249 7331 32283
rect 8998 32249 9032 32283
rect 10241 32249 10275 32283
rect 10746 32249 10780 32283
rect 2513 32181 2547 32215
rect 4261 32181 4295 32215
rect 4721 32181 4755 32215
rect 5273 32181 5307 32215
rect 5917 32181 5951 32215
rect 6653 32181 6687 32215
rect 8585 32181 8619 32215
rect 11345 32181 11379 32215
rect 2789 31977 2823 32011
rect 5457 31977 5491 32011
rect 5825 31977 5859 32011
rect 8953 31977 8987 32011
rect 9505 31977 9539 32011
rect 10701 31977 10735 32011
rect 11345 31977 11379 32011
rect 4623 31909 4657 31943
rect 7021 31909 7055 31943
rect 9873 31909 9907 31943
rect 2605 31841 2639 31875
rect 8401 31841 8435 31875
rect 11529 31841 11563 31875
rect 11713 31841 11747 31875
rect 12449 31841 12483 31875
rect 4261 31773 4295 31807
rect 6929 31773 6963 31807
rect 9781 31773 9815 31807
rect 7481 31705 7515 31739
rect 10333 31705 10367 31739
rect 5181 31637 5215 31671
rect 7849 31637 7883 31671
rect 8539 31637 8573 31671
rect 2605 31433 2639 31467
rect 4537 31433 4571 31467
rect 6653 31433 6687 31467
rect 7941 31433 7975 31467
rect 9045 31433 9079 31467
rect 9597 31433 9631 31467
rect 11621 31433 11655 31467
rect 5641 31365 5675 31399
rect 10333 31365 10367 31399
rect 4169 31297 4203 31331
rect 4813 31297 4847 31331
rect 6193 31297 6227 31331
rect 6929 31297 6963 31331
rect 3433 31229 3467 31263
rect 3893 31229 3927 31263
rect 8620 31229 8654 31263
rect 5089 31161 5123 31195
rect 5181 31161 5215 31195
rect 7021 31161 7055 31195
rect 7573 31161 7607 31195
rect 9781 31161 9815 31195
rect 9873 31161 9907 31195
rect 10701 31161 10735 31195
rect 3249 31093 3283 31127
rect 8401 31093 8435 31127
rect 8723 31093 8757 31127
rect 11253 31093 11287 31127
rect 3525 30889 3559 30923
rect 4445 30889 4479 30923
rect 6561 30889 6595 30923
rect 7573 30889 7607 30923
rect 5089 30821 5123 30855
rect 8217 30821 8251 30855
rect 9781 30821 9815 30855
rect 9873 30821 9907 30855
rect 6745 30753 6779 30787
rect 7021 30753 7055 30787
rect 9137 30753 9171 30787
rect 11288 30753 11322 30787
rect 4813 30685 4847 30719
rect 4997 30685 5031 30719
rect 8125 30685 8159 30719
rect 10057 30685 10091 30719
rect 5549 30617 5583 30651
rect 8677 30617 8711 30651
rect 9413 30549 9447 30583
rect 11391 30549 11425 30583
rect 4353 30345 4387 30379
rect 6561 30345 6595 30379
rect 9505 30345 9539 30379
rect 10517 30345 10551 30379
rect 11253 30345 11287 30379
rect 9229 30277 9263 30311
rect 4721 30209 4755 30243
rect 5181 30141 5215 30175
rect 5733 30141 5767 30175
rect 6872 30141 6906 30175
rect 7297 30141 7331 30175
rect 7941 30141 7975 30175
rect 9724 30141 9758 30175
rect 10149 30141 10183 30175
rect 5917 30073 5951 30107
rect 8262 30073 8296 30107
rect 4997 30005 5031 30039
rect 6975 30005 7009 30039
rect 7757 30005 7791 30039
rect 8861 30005 8895 30039
rect 9827 30005 9861 30039
rect 1593 29801 1627 29835
rect 6837 29801 6871 29835
rect 8125 29801 8159 29835
rect 12265 29801 12299 29835
rect 5089 29733 5123 29767
rect 5641 29733 5675 29767
rect 6561 29733 6595 29767
rect 7205 29733 7239 29767
rect 7757 29733 7791 29767
rect 9873 29733 9907 29767
rect 1409 29665 1443 29699
rect 8620 29665 8654 29699
rect 12081 29665 12115 29699
rect 4997 29597 5031 29631
rect 7113 29597 7147 29631
rect 8723 29597 8757 29631
rect 9781 29597 9815 29631
rect 10333 29529 10367 29563
rect 4721 29461 4755 29495
rect 8493 29461 8527 29495
rect 3433 29257 3467 29291
rect 3709 29257 3743 29291
rect 9689 29257 9723 29291
rect 11161 29257 11195 29291
rect 5825 29189 5859 29223
rect 9229 29189 9263 29223
rect 6837 29121 6871 29155
rect 8677 29121 8711 29155
rect 10241 29121 10275 29155
rect 10517 29121 10551 29155
rect 3224 29053 3258 29087
rect 3433 29053 3467 29087
rect 4236 29053 4270 29087
rect 4629 29053 4663 29087
rect 7757 29053 7791 29087
rect 8033 29053 8067 29087
rect 4445 28985 4479 29019
rect 5273 28985 5307 29019
rect 5365 28985 5399 29019
rect 6285 28985 6319 29019
rect 7158 28985 7192 29019
rect 8769 28985 8803 29019
rect 10333 28985 10367 29019
rect 1593 28917 1627 28951
rect 3295 28917 3329 28951
rect 3985 28917 4019 28951
rect 5089 28917 5123 28951
rect 6653 28917 6687 28951
rect 8401 28917 8435 28951
rect 9965 28917 9999 28951
rect 12173 28917 12207 28951
rect 3157 28713 3191 28747
rect 5641 28713 5675 28747
rect 6561 28713 6595 28747
rect 7113 28713 7147 28747
rect 7481 28713 7515 28747
rect 8953 28713 8987 28747
rect 10701 28713 10735 28747
rect 12403 28713 12437 28747
rect 4813 28645 4847 28679
rect 7757 28645 7791 28679
rect 8125 28645 8159 28679
rect 9873 28645 9907 28679
rect 10425 28645 10459 28679
rect 2881 28577 2915 28611
rect 11253 28577 11287 28611
rect 12332 28577 12366 28611
rect 4721 28509 4755 28543
rect 6193 28509 6227 28543
rect 8033 28509 8067 28543
rect 8309 28509 8343 28543
rect 9505 28509 9539 28543
rect 9781 28509 9815 28543
rect 11391 28509 11425 28543
rect 5273 28441 5307 28475
rect 2421 28169 2455 28203
rect 3433 28169 3467 28203
rect 5733 28169 5767 28203
rect 9045 28169 9079 28203
rect 3617 28101 3651 28135
rect 11253 28101 11287 28135
rect 2697 28033 2731 28067
rect 9689 28033 9723 28067
rect 2212 27965 2246 27999
rect 3224 27965 3258 27999
rect 4169 27965 4203 27999
rect 6888 27965 6922 27999
rect 7297 27965 7331 27999
rect 8125 27965 8159 27999
rect 9873 27965 9907 27999
rect 4531 27897 4565 27931
rect 6193 27897 6227 27931
rect 6975 27897 7009 27931
rect 8446 27897 8480 27931
rect 10194 27897 10228 27931
rect 3065 27829 3099 27863
rect 4077 27829 4111 27863
rect 5089 27829 5123 27863
rect 5365 27829 5399 27863
rect 6653 27829 6687 27863
rect 7941 27829 7975 27863
rect 9321 27829 9355 27863
rect 10793 27829 10827 27863
rect 12633 27829 12667 27863
rect 7665 27625 7699 27659
rect 9505 27625 9539 27659
rect 4721 27557 4755 27591
rect 6377 27557 6411 27591
rect 6929 27557 6963 27591
rect 8493 27557 8527 27591
rect 9873 27557 9907 27591
rect 2697 27489 2731 27523
rect 2973 27489 3007 27523
rect 5365 27489 5399 27523
rect 7757 27489 7791 27523
rect 8217 27489 8251 27523
rect 3157 27421 3191 27455
rect 4445 27421 4479 27455
rect 6285 27421 6319 27455
rect 9781 27421 9815 27455
rect 10333 27353 10367 27387
rect 4261 27285 4295 27319
rect 8861 27285 8895 27319
rect 2697 27081 2731 27115
rect 6285 27081 6319 27115
rect 8677 27081 8711 27115
rect 9873 27081 9907 27115
rect 10241 27081 10275 27115
rect 10563 27081 10597 27115
rect 6561 27013 6595 27047
rect 8309 27013 8343 27047
rect 3893 26945 3927 26979
rect 5089 26945 5123 26979
rect 8033 26945 8067 26979
rect 2145 26877 2179 26911
rect 3065 26877 3099 26911
rect 3433 26877 3467 26911
rect 3617 26877 3651 26911
rect 7297 26877 7331 26911
rect 7757 26877 7791 26911
rect 8861 26877 8895 26911
rect 9321 26877 9355 26911
rect 10460 26877 10494 26911
rect 10885 26877 10919 26911
rect 4813 26809 4847 26843
rect 4905 26809 4939 26843
rect 5733 26809 5767 26843
rect 1961 26741 1995 26775
rect 2329 26741 2363 26775
rect 4537 26741 4571 26775
rect 7113 26741 7147 26775
rect 8953 26741 8987 26775
rect 3157 26537 3191 26571
rect 5089 26537 5123 26571
rect 7297 26537 7331 26571
rect 7665 26537 7699 26571
rect 9781 26537 9815 26571
rect 2513 26469 2547 26503
rect 3525 26469 3559 26503
rect 4813 26469 4847 26503
rect 6377 26469 6411 26503
rect 2973 26401 3007 26435
rect 4353 26401 4387 26435
rect 4537 26401 4571 26435
rect 5733 26401 5767 26435
rect 6101 26401 6135 26435
rect 8033 26401 8067 26435
rect 8309 26401 8343 26435
rect 9689 26401 9723 26435
rect 10149 26401 10183 26435
rect 11320 26401 11354 26435
rect 8585 26333 8619 26367
rect 5457 26265 5491 26299
rect 8861 26265 8895 26299
rect 10793 26197 10827 26231
rect 11391 26197 11425 26231
rect 4215 25993 4249 26027
rect 4905 25993 4939 26027
rect 6101 25993 6135 26027
rect 9965 25993 9999 26027
rect 10333 25993 10367 26027
rect 5273 25925 5307 25959
rect 8217 25857 8251 25891
rect 10609 25857 10643 25891
rect 12449 25857 12483 25891
rect 4112 25789 4146 25823
rect 4537 25789 4571 25823
rect 5089 25789 5123 25823
rect 7205 25789 7239 25823
rect 7665 25789 7699 25823
rect 7941 25789 7975 25823
rect 8769 25789 8803 25823
rect 9689 25789 9723 25823
rect 3985 25721 4019 25755
rect 9090 25721 9124 25755
rect 10701 25721 10735 25755
rect 11253 25721 11287 25755
rect 3065 25653 3099 25687
rect 5733 25653 5767 25687
rect 7113 25653 7147 25687
rect 8585 25653 8619 25687
rect 11529 25653 11563 25687
rect 4629 25449 4663 25483
rect 8401 25449 8435 25483
rect 8769 25449 8803 25483
rect 10057 25449 10091 25483
rect 10609 25449 10643 25483
rect 10885 25449 10919 25483
rect 6009 25381 6043 25415
rect 7205 25381 7239 25415
rect 7573 25381 7607 25415
rect 11621 25381 11655 25415
rect 4445 25313 4479 25347
rect 9689 25313 9723 25347
rect 5917 25245 5951 25279
rect 6561 25245 6595 25279
rect 7481 25245 7515 25279
rect 8125 25245 8159 25279
rect 11529 25245 11563 25279
rect 11805 25245 11839 25279
rect 5089 25109 5123 25143
rect 5457 25109 5491 25143
rect 6929 25109 6963 25143
rect 3295 24905 3329 24939
rect 4997 24905 5031 24939
rect 8677 24905 8711 24939
rect 10057 24905 10091 24939
rect 11621 24905 11655 24939
rect 3617 24837 3651 24871
rect 11989 24837 12023 24871
rect 6561 24769 6595 24803
rect 7205 24769 7239 24803
rect 8217 24769 8251 24803
rect 8861 24769 8895 24803
rect 11345 24769 11379 24803
rect 3224 24701 3258 24735
rect 4220 24701 4254 24735
rect 4629 24701 4663 24735
rect 9781 24701 9815 24735
rect 10425 24701 10459 24735
rect 4077 24633 4111 24667
rect 4307 24633 4341 24667
rect 5273 24633 5307 24667
rect 5365 24633 5399 24667
rect 5917 24633 5951 24667
rect 6929 24633 6963 24667
rect 7021 24633 7055 24667
rect 9182 24633 9216 24667
rect 10701 24633 10735 24667
rect 10793 24633 10827 24667
rect 6193 24565 6227 24599
rect 7849 24565 7883 24599
rect 3111 24361 3145 24395
rect 8861 24361 8895 24395
rect 9413 24361 9447 24395
rect 11391 24361 11425 24395
rect 5226 24293 5260 24327
rect 6837 24293 6871 24327
rect 9873 24293 9907 24327
rect 3040 24225 3074 24259
rect 6101 24225 6135 24259
rect 8252 24225 8286 24259
rect 11253 24225 11287 24259
rect 4905 24157 4939 24191
rect 6561 24157 6595 24191
rect 6745 24157 6779 24191
rect 9781 24157 9815 24191
rect 10057 24157 10091 24191
rect 7297 24089 7331 24123
rect 3525 24021 3559 24055
rect 4721 24021 4755 24055
rect 5825 24021 5859 24055
rect 8355 24021 8389 24055
rect 10701 24021 10735 24055
rect 2329 23817 2363 23851
rect 6193 23817 6227 23851
rect 7849 23817 7883 23851
rect 9505 23817 9539 23851
rect 3065 23749 3099 23783
rect 5917 23749 5951 23783
rect 10977 23749 11011 23783
rect 2559 23681 2593 23715
rect 6929 23681 6963 23715
rect 7297 23681 7331 23715
rect 8493 23681 8527 23715
rect 8769 23681 8803 23715
rect 10333 23681 10367 23715
rect 11345 23681 11379 23715
rect 2456 23613 2490 23647
rect 3433 23613 3467 23647
rect 3893 23613 3927 23647
rect 4997 23613 5031 23647
rect 4261 23545 4295 23579
rect 7021 23545 7055 23579
rect 8585 23545 8619 23579
rect 10057 23545 10091 23579
rect 10149 23545 10183 23579
rect 4445 23477 4479 23511
rect 4813 23477 4847 23511
rect 5365 23477 5399 23511
rect 6561 23477 6595 23511
rect 8217 23477 8251 23511
rect 9781 23477 9815 23511
rect 3065 23273 3099 23307
rect 5549 23273 5583 23307
rect 5825 23273 5859 23307
rect 7665 23273 7699 23307
rect 8263 23273 8297 23307
rect 8585 23273 8619 23307
rect 9689 23273 9723 23307
rect 3525 23205 3559 23239
rect 4991 23205 5025 23239
rect 6698 23205 6732 23239
rect 2881 23137 2915 23171
rect 8125 23137 8159 23171
rect 10701 23137 10735 23171
rect 4629 23069 4663 23103
rect 6377 23069 6411 23103
rect 7297 23001 7331 23035
rect 4537 22933 4571 22967
rect 6193 22933 6227 22967
rect 10149 22933 10183 22967
rect 10839 22933 10873 22967
rect 2881 22729 2915 22763
rect 3525 22729 3559 22763
rect 7757 22729 7791 22763
rect 10701 22729 10735 22763
rect 4813 22661 4847 22695
rect 4353 22593 4387 22627
rect 4721 22593 4755 22627
rect 3893 22525 3927 22559
rect 4169 22525 4203 22559
rect 5917 22593 5951 22627
rect 9413 22593 9447 22627
rect 5273 22525 5307 22559
rect 5641 22525 5675 22559
rect 6837 22525 6871 22559
rect 10920 22525 10954 22559
rect 11345 22525 11379 22559
rect 4813 22457 4847 22491
rect 6285 22457 6319 22491
rect 6653 22457 6687 22491
rect 7199 22457 7233 22491
rect 9505 22457 9539 22491
rect 10057 22457 10091 22491
rect 5089 22389 5123 22423
rect 8125 22389 8159 22423
rect 9229 22389 9263 22423
rect 11023 22389 11057 22423
rect 4261 22185 4295 22219
rect 4537 22185 4571 22219
rect 5457 22185 5491 22219
rect 9413 22185 9447 22219
rect 8211 22117 8245 22151
rect 9873 22117 9907 22151
rect 10425 22117 10459 22151
rect 4445 22049 4479 22083
rect 4997 22049 5031 22083
rect 6285 22049 6319 22083
rect 6837 22049 6871 22083
rect 8769 22049 8803 22083
rect 11253 22049 11287 22083
rect 7021 21981 7055 22015
rect 7849 21981 7883 22015
rect 9781 21981 9815 22015
rect 3709 21913 3743 21947
rect 7297 21845 7331 21879
rect 10793 21845 10827 21879
rect 11391 21845 11425 21879
rect 6285 21641 6319 21675
rect 7021 21641 7055 21675
rect 9781 21641 9815 21675
rect 10609 21573 10643 21607
rect 5917 21505 5951 21539
rect 10057 21505 10091 21539
rect 3560 21437 3594 21471
rect 3985 21437 4019 21471
rect 5089 21437 5123 21471
rect 5457 21437 5491 21471
rect 5641 21437 5675 21471
rect 6837 21437 6871 21471
rect 8217 21437 8251 21471
rect 4537 21369 4571 21403
rect 7297 21369 7331 21403
rect 7757 21369 7791 21403
rect 8033 21369 8067 21403
rect 8538 21369 8572 21403
rect 10149 21369 10183 21403
rect 3663 21301 3697 21335
rect 9137 21301 9171 21335
rect 11253 21301 11287 21335
rect 3617 21097 3651 21131
rect 7849 21097 7883 21131
rect 9045 21097 9079 21131
rect 9505 21097 9539 21131
rect 10701 21097 10735 21131
rect 11391 21097 11425 21131
rect 4261 21029 4295 21063
rect 6377 21029 6411 21063
rect 7205 21029 7239 21063
rect 8217 21029 8251 21063
rect 9873 21029 9907 21063
rect 10425 21029 10459 21063
rect 6653 20961 6687 20995
rect 7021 20961 7055 20995
rect 11288 20961 11322 20995
rect 4169 20893 4203 20927
rect 7573 20893 7607 20927
rect 8125 20893 8159 20927
rect 8769 20893 8803 20927
rect 9781 20893 9815 20927
rect 4721 20825 4755 20859
rect 5181 20757 5215 20791
rect 5549 20757 5583 20791
rect 6561 20553 6595 20587
rect 7941 20553 7975 20587
rect 9689 20553 9723 20587
rect 2743 20485 2777 20519
rect 3709 20417 3743 20451
rect 5273 20417 5307 20451
rect 10517 20417 10551 20451
rect 2672 20349 2706 20383
rect 3065 20349 3099 20383
rect 6837 20349 6871 20383
rect 7297 20349 7331 20383
rect 7573 20349 7607 20383
rect 8401 20349 8435 20383
rect 3525 20281 3559 20315
rect 3801 20281 3835 20315
rect 4353 20281 4387 20315
rect 5365 20281 5399 20315
rect 5917 20281 5951 20315
rect 8722 20281 8756 20315
rect 10241 20281 10275 20315
rect 10333 20281 10367 20315
rect 4721 20213 4755 20247
rect 5089 20213 5123 20247
rect 6285 20213 6319 20247
rect 8217 20213 8251 20247
rect 9321 20213 9355 20247
rect 11253 20213 11287 20247
rect 3893 20009 3927 20043
rect 4445 20009 4479 20043
rect 4997 20009 5031 20043
rect 6929 20009 6963 20043
rect 7205 20009 7239 20043
rect 7481 20009 7515 20043
rect 8953 20009 8987 20043
rect 9505 20009 9539 20043
rect 9827 20009 9861 20043
rect 10517 20009 10551 20043
rect 10839 20009 10873 20043
rect 5917 19941 5951 19975
rect 6009 19941 6043 19975
rect 8585 19941 8619 19975
rect 2697 19873 2731 19907
rect 2973 19873 3007 19907
rect 3157 19873 3191 19907
rect 5273 19873 5307 19907
rect 7389 19873 7423 19907
rect 7941 19873 7975 19907
rect 9724 19873 9758 19907
rect 10241 19873 10275 19907
rect 10736 19873 10770 19907
rect 4077 19805 4111 19839
rect 6193 19805 6227 19839
rect 3525 19669 3559 19703
rect 2973 19465 3007 19499
rect 5917 19465 5951 19499
rect 7757 19465 7791 19499
rect 8033 19465 8067 19499
rect 10287 19465 10321 19499
rect 4077 19397 4111 19431
rect 2605 19329 2639 19363
rect 4997 19329 5031 19363
rect 9597 19329 9631 19363
rect 1777 19261 1811 19295
rect 1869 19261 1903 19295
rect 2329 19261 2363 19295
rect 6837 19261 6871 19295
rect 8585 19261 8619 19295
rect 9045 19261 9079 19295
rect 10184 19261 10218 19295
rect 3249 19193 3283 19227
rect 3525 19193 3559 19227
rect 3617 19193 3651 19227
rect 4537 19193 4571 19227
rect 4905 19193 4939 19227
rect 5318 19193 5352 19227
rect 7158 19193 7192 19227
rect 6193 19125 6227 19159
rect 6653 19125 6687 19159
rect 8493 19125 8527 19159
rect 8677 19125 8711 19159
rect 9965 19125 9999 19159
rect 10701 19125 10735 19159
rect 4261 18921 4295 18955
rect 5733 18921 5767 18955
rect 7757 18921 7791 18955
rect 2605 18853 2639 18887
rect 5175 18853 5209 18887
rect 6009 18853 6043 18887
rect 1444 18785 1478 18819
rect 3157 18785 3191 18819
rect 7389 18785 7423 18819
rect 2513 18717 2547 18751
rect 4721 18717 4755 18751
rect 4813 18717 4847 18751
rect 1547 18649 1581 18683
rect 1961 18581 1995 18615
rect 3525 18581 3559 18615
rect 6837 18581 6871 18615
rect 7205 18581 7239 18615
rect 8309 18581 8343 18615
rect 8585 18581 8619 18615
rect 2421 18377 2455 18411
rect 2789 18377 2823 18411
rect 3709 18377 3743 18411
rect 3801 18377 3835 18411
rect 6653 18377 6687 18411
rect 2028 18173 2062 18207
rect 3024 18173 3058 18207
rect 5733 18309 5767 18343
rect 4077 18241 4111 18275
rect 4721 18241 4755 18275
rect 8677 18241 8711 18275
rect 5549 18173 5583 18207
rect 6009 18173 6043 18207
rect 10460 18173 10494 18207
rect 10885 18173 10919 18207
rect 3111 18105 3145 18139
rect 3709 18105 3743 18139
rect 4169 18105 4203 18139
rect 5089 18105 5123 18139
rect 7205 18105 7239 18139
rect 7297 18105 7331 18139
rect 7849 18105 7883 18139
rect 8998 18105 9032 18139
rect 1593 18037 1627 18071
rect 2099 18037 2133 18071
rect 3525 18037 3559 18071
rect 5365 18037 5399 18071
rect 8125 18037 8159 18071
rect 8493 18037 8527 18071
rect 9597 18037 9631 18071
rect 10563 18037 10597 18071
rect 2513 17833 2547 17867
rect 3111 17833 3145 17867
rect 8769 17833 8803 17867
rect 4261 17765 4295 17799
rect 4813 17765 4847 17799
rect 6101 17765 6135 17799
rect 7894 17765 7928 17799
rect 9781 17765 9815 17799
rect 9873 17765 9907 17799
rect 3040 17697 3074 17731
rect 4169 17629 4203 17663
rect 6009 17629 6043 17663
rect 6285 17629 6319 17663
rect 7573 17629 7607 17663
rect 10057 17629 10091 17663
rect 5273 17493 5307 17527
rect 7205 17493 7239 17527
rect 8493 17493 8527 17527
rect 3157 17289 3191 17323
rect 4629 17289 4663 17323
rect 6561 17289 6595 17323
rect 7481 17289 7515 17323
rect 9413 17289 9447 17323
rect 10517 17289 10551 17323
rect 11529 17289 11563 17323
rect 8585 17221 8619 17255
rect 3525 17153 3559 17187
rect 4353 17153 4387 17187
rect 5917 17153 5951 17187
rect 9597 17153 9631 17187
rect 10885 17153 10919 17187
rect 3617 17085 3651 17119
rect 4077 17085 4111 17119
rect 4905 17085 4939 17119
rect 5181 17085 5215 17119
rect 5641 17085 5675 17119
rect 6996 17085 7030 17119
rect 11136 17085 11170 17119
rect 2605 17017 2639 17051
rect 6193 17017 6227 17051
rect 8033 17017 8067 17051
rect 8125 17017 8159 17051
rect 9689 17017 9723 17051
rect 10241 17017 10275 17051
rect 4905 16949 4939 16983
rect 4997 16949 5031 16983
rect 7067 16949 7101 16983
rect 7757 16949 7791 16983
rect 8953 16949 8987 16983
rect 11207 16949 11241 16983
rect 3617 16745 3651 16779
rect 4629 16745 4663 16779
rect 5549 16745 5583 16779
rect 6101 16745 6135 16779
rect 7067 16745 7101 16779
rect 7573 16745 7607 16779
rect 10149 16745 10183 16779
rect 8125 16677 8159 16711
rect 8217 16677 8251 16711
rect 9137 16677 9171 16711
rect 2973 16609 3007 16643
rect 4169 16609 4203 16643
rect 6964 16609 6998 16643
rect 9597 16609 9631 16643
rect 10701 16609 10735 16643
rect 5181 16541 5215 16575
rect 8401 16541 8435 16575
rect 3157 16473 3191 16507
rect 4353 16473 4387 16507
rect 10839 16473 10873 16507
rect 9827 16405 9861 16439
rect 3065 16201 3099 16235
rect 4445 16201 4479 16235
rect 5457 16201 5491 16235
rect 8401 16201 8435 16235
rect 10609 16201 10643 16235
rect 5641 16133 5675 16167
rect 10885 16133 10919 16167
rect 2697 15997 2731 16031
rect 3525 15997 3559 16031
rect 5273 15997 5307 16031
rect 6561 16065 6595 16099
rect 7573 16065 7607 16099
rect 8125 16065 8159 16099
rect 9229 16065 9263 16099
rect 9505 16065 9539 16099
rect 7021 15997 7055 16031
rect 7481 15997 7515 16031
rect 10701 15997 10735 16031
rect 11253 15997 11287 16031
rect 3846 15929 3880 15963
rect 5089 15929 5123 15963
rect 5641 15929 5675 15963
rect 6285 15929 6319 15963
rect 9045 15929 9079 15963
rect 9321 15929 9355 15963
rect 3341 15861 3375 15895
rect 4721 15861 4755 15895
rect 5825 15861 5859 15895
rect 10149 15861 10183 15895
rect 4169 15657 4203 15691
rect 5181 15657 5215 15691
rect 6285 15657 6319 15691
rect 9229 15657 9263 15691
rect 11345 15657 11379 15691
rect 3157 15589 3191 15623
rect 7849 15589 7883 15623
rect 9873 15589 9907 15623
rect 2605 15521 2639 15555
rect 2881 15521 2915 15555
rect 4077 15521 4111 15555
rect 4629 15521 4663 15555
rect 6837 15521 6871 15555
rect 11253 15521 11287 15555
rect 11713 15521 11747 15555
rect 5917 15453 5951 15487
rect 7757 15453 7791 15487
rect 8033 15453 8067 15487
rect 9781 15453 9815 15487
rect 10057 15453 10091 15487
rect 7481 15385 7515 15419
rect 3617 15317 3651 15351
rect 7113 15317 7147 15351
rect 10701 15317 10735 15351
rect 2145 15113 2179 15147
rect 2789 15113 2823 15147
rect 4537 15113 4571 15147
rect 5549 15113 5583 15147
rect 6469 15113 6503 15147
rect 6653 15113 6687 15147
rect 7849 15113 7883 15147
rect 9321 15113 9355 15147
rect 9689 15113 9723 15147
rect 11345 15113 11379 15147
rect 11713 15113 11747 15147
rect 2513 15045 2547 15079
rect 6469 14977 6503 15011
rect 8401 14977 8435 15011
rect 10517 14977 10551 15011
rect 2605 14909 2639 14943
rect 3065 14909 3099 14943
rect 3617 14909 3651 14943
rect 5365 14909 5399 14943
rect 7573 14909 7607 14943
rect 3433 14841 3467 14875
rect 3979 14841 4013 14875
rect 6929 14841 6963 14875
rect 7021 14841 7055 14875
rect 8722 14841 8756 14875
rect 10241 14841 10275 14875
rect 10333 14841 10367 14875
rect 4813 14773 4847 14807
rect 5273 14773 5307 14807
rect 6009 14773 6043 14807
rect 8217 14773 8251 14807
rect 3111 14569 3145 14603
rect 4353 14569 4387 14603
rect 7941 14569 7975 14603
rect 8493 14569 8527 14603
rect 10609 14569 10643 14603
rect 3617 14501 3651 14535
rect 7113 14501 7147 14535
rect 10010 14501 10044 14535
rect 10885 14501 10919 14535
rect 2881 14433 2915 14467
rect 4169 14433 4203 14467
rect 4721 14433 4755 14467
rect 5365 14433 5399 14467
rect 5641 14433 5675 14467
rect 8652 14433 8686 14467
rect 9045 14433 9079 14467
rect 11437 14433 11471 14467
rect 5825 14365 5859 14399
rect 7021 14365 7055 14399
rect 7665 14365 7699 14399
rect 9689 14365 9723 14399
rect 8723 14297 8757 14331
rect 9505 14297 9539 14331
rect 11575 14297 11609 14331
rect 6193 14229 6227 14263
rect 6837 14229 6871 14263
rect 5089 14025 5123 14059
rect 6193 14025 6227 14059
rect 9781 14025 9815 14059
rect 9321 13957 9355 13991
rect 3065 13889 3099 13923
rect 5917 13889 5951 13923
rect 8769 13889 8803 13923
rect 3893 13821 3927 13855
rect 4169 13821 4203 13855
rect 5181 13821 5215 13855
rect 5641 13821 5675 13855
rect 6929 13821 6963 13855
rect 8125 13821 8159 13855
rect 10517 13821 10551 13855
rect 10793 13821 10827 13855
rect 2697 13753 2731 13787
rect 7250 13753 7284 13787
rect 8861 13753 8895 13787
rect 10149 13753 10183 13787
rect 3433 13685 3467 13719
rect 3709 13685 3743 13719
rect 4721 13685 4755 13719
rect 6653 13685 6687 13719
rect 7849 13685 7883 13719
rect 8493 13685 8527 13719
rect 10333 13685 10367 13719
rect 11529 13685 11563 13719
rect 1593 13481 1627 13515
rect 6745 13481 6779 13515
rect 7113 13481 7147 13515
rect 8861 13481 8895 13515
rect 9505 13481 9539 13515
rect 10701 13481 10735 13515
rect 4997 13413 5031 13447
rect 6187 13413 6221 13447
rect 7894 13413 7928 13447
rect 9873 13413 9907 13447
rect 1409 13345 1443 13379
rect 2881 13345 2915 13379
rect 4261 13345 4295 13379
rect 4813 13345 4847 13379
rect 5089 13345 5123 13379
rect 5825 13345 5859 13379
rect 7389 13345 7423 13379
rect 3111 13209 3145 13243
rect 7573 13277 7607 13311
rect 9781 13277 9815 13311
rect 10057 13277 10091 13311
rect 3709 13141 3743 13175
rect 5089 13141 5123 13175
rect 5365 13141 5399 13175
rect 5733 13141 5767 13175
rect 8493 13141 8527 13175
rect 1593 12937 1627 12971
rect 3065 12937 3099 12971
rect 3433 12937 3467 12971
rect 3755 12937 3789 12971
rect 6975 12937 7009 12971
rect 9229 12937 9263 12971
rect 10563 12937 10597 12971
rect 3893 12869 3927 12903
rect 10241 12869 10275 12903
rect 3985 12801 4019 12835
rect 6561 12801 6595 12835
rect 7941 12801 7975 12835
rect 3617 12733 3651 12767
rect 5181 12733 5215 12767
rect 5733 12733 5767 12767
rect 6872 12733 6906 12767
rect 7297 12733 7331 12767
rect 8585 12733 8619 12767
rect 9448 12733 9482 12767
rect 9873 12733 9907 12767
rect 10492 12733 10526 12767
rect 5089 12665 5123 12699
rect 5917 12665 5951 12699
rect 8033 12665 8067 12699
rect 9551 12665 9585 12699
rect 2697 12597 2731 12631
rect 4261 12597 4295 12631
rect 4721 12597 4755 12631
rect 6285 12597 6319 12631
rect 7665 12597 7699 12631
rect 8861 12597 8895 12631
rect 10977 12597 11011 12631
rect 4813 12393 4847 12427
rect 7573 12393 7607 12427
rect 8769 12393 8803 12427
rect 9781 12393 9815 12427
rect 13645 12393 13679 12427
rect 3157 12325 3191 12359
rect 7941 12325 7975 12359
rect 2605 12257 2639 12291
rect 2789 12257 2823 12291
rect 4169 12257 4203 12291
rect 5733 12257 5767 12291
rect 6193 12257 6227 12291
rect 9689 12257 9723 12291
rect 10149 12257 10183 12291
rect 13461 12257 13495 12291
rect 2513 12189 2547 12223
rect 3709 12189 3743 12223
rect 4537 12189 4571 12223
rect 5181 12189 5215 12223
rect 6469 12189 6503 12223
rect 7849 12189 7883 12223
rect 8493 12189 8527 12223
rect 5549 12121 5583 12155
rect 4307 12053 4341 12087
rect 4445 12053 4479 12087
rect 7113 12053 7147 12087
rect 1685 11849 1719 11883
rect 1961 11849 1995 11883
rect 2329 11849 2363 11883
rect 3893 11849 3927 11883
rect 4261 11849 4295 11883
rect 4813 11849 4847 11883
rect 6469 11849 6503 11883
rect 8677 11849 8711 11883
rect 10057 11849 10091 11883
rect 10425 11849 10459 11883
rect 13461 11849 13495 11883
rect 2697 11781 2731 11815
rect 4629 11781 4663 11815
rect 7665 11781 7699 11815
rect 4721 11713 4755 11747
rect 7113 11713 7147 11747
rect 8861 11713 8895 11747
rect 1777 11645 1811 11679
rect 3433 11645 3467 11679
rect 3525 11645 3559 11679
rect 4500 11645 4534 11679
rect 5457 11645 5491 11679
rect 5733 11645 5767 11679
rect 4353 11577 4387 11611
rect 7205 11577 7239 11611
rect 9182 11577 9216 11611
rect 6193 11509 6227 11543
rect 8033 11509 8067 11543
rect 9781 11509 9815 11543
rect 10609 11509 10643 11543
rect 1593 11305 1627 11339
rect 4537 11305 4571 11339
rect 5457 11305 5491 11339
rect 7573 11305 7607 11339
rect 7941 11305 7975 11339
rect 8953 11305 8987 11339
rect 1961 11237 1995 11271
rect 6974 11237 7008 11271
rect 8217 11237 8251 11271
rect 9873 11237 9907 11271
rect 10425 11237 10459 11271
rect 1409 11169 1443 11203
rect 2421 11169 2455 11203
rect 2697 11169 2731 11203
rect 4077 11169 4111 11203
rect 4307 11169 4341 11203
rect 5641 11169 5675 11203
rect 6653 11169 6687 11203
rect 2973 11101 3007 11135
rect 8401 11101 8435 11135
rect 9781 11101 9815 11135
rect 2329 11033 2363 11067
rect 2513 11033 2547 11067
rect 4169 11033 4203 11067
rect 5089 11033 5123 11067
rect 5825 11033 5859 11067
rect 3525 10965 3559 10999
rect 3801 10965 3835 10999
rect 1685 10761 1719 10795
rect 2513 10761 2547 10795
rect 4169 10761 4203 10795
rect 4491 10761 4525 10795
rect 4813 10761 4847 10795
rect 8493 10761 8527 10795
rect 9689 10761 9723 10795
rect 10057 10761 10091 10795
rect 4629 10693 4663 10727
rect 5365 10693 5399 10727
rect 3801 10625 3835 10659
rect 4721 10625 4755 10659
rect 5733 10625 5767 10659
rect 8769 10625 8803 10659
rect 9045 10625 9079 10659
rect 1777 10557 1811 10591
rect 2881 10557 2915 10591
rect 3525 10557 3559 10591
rect 6929 10557 6963 10591
rect 4353 10489 4387 10523
rect 7250 10489 7284 10523
rect 8861 10489 8895 10523
rect 1961 10421 1995 10455
rect 6285 10421 6319 10455
rect 6653 10421 6687 10455
rect 7849 10421 7883 10455
rect 1593 10217 1627 10251
rect 3157 10217 3191 10251
rect 3893 10217 3927 10251
rect 4905 10217 4939 10251
rect 5641 10217 5675 10251
rect 6837 10217 6871 10251
rect 7665 10217 7699 10251
rect 8677 10217 8711 10251
rect 6561 10149 6595 10183
rect 7205 10149 7239 10183
rect 1409 10081 1443 10115
rect 2973 10081 3007 10115
rect 4261 10081 4295 10115
rect 6101 10081 6135 10115
rect 6285 10081 6319 10115
rect 7389 10081 7423 10115
rect 7573 10081 7607 10115
rect 9756 10081 9790 10115
rect 10701 10081 10735 10115
rect 4629 10013 4663 10047
rect 4426 9945 4460 9979
rect 4537 9945 4571 9979
rect 2421 9877 2455 9911
rect 2789 9877 2823 9911
rect 5365 9877 5399 9911
rect 8309 9877 8343 9911
rect 9827 9877 9861 9911
rect 10931 9877 10965 9911
rect 2973 9673 3007 9707
rect 3709 9673 3743 9707
rect 4997 9673 5031 9707
rect 6285 9673 6319 9707
rect 7941 9673 7975 9707
rect 10149 9673 10183 9707
rect 10885 9673 10919 9707
rect 3249 9605 3283 9639
rect 4629 9605 4663 9639
rect 7251 9605 7285 9639
rect 10609 9605 10643 9639
rect 4261 9537 4295 9571
rect 8217 9537 8251 9571
rect 9137 9537 9171 9571
rect 3801 9469 3835 9503
rect 3985 9469 4019 9503
rect 5181 9469 5215 9503
rect 5641 9469 5675 9503
rect 7180 9469 7214 9503
rect 7573 9469 7607 9503
rect 9756 9469 9790 9503
rect 5917 9401 5951 9435
rect 8309 9401 8343 9435
rect 8861 9401 8895 9435
rect 1685 9333 1719 9367
rect 6653 9333 6687 9367
rect 9827 9333 9861 9367
rect 3157 9129 3191 9163
rect 5365 9129 5399 9163
rect 7481 9129 7515 9163
rect 3525 9061 3559 9095
rect 3893 9061 3927 9095
rect 8125 9061 8159 9095
rect 8677 9061 8711 9095
rect 9781 9061 9815 9095
rect 9873 9061 9907 9095
rect 2973 8993 3007 9027
rect 4353 8993 4387 9027
rect 4905 8993 4939 9027
rect 5733 8993 5767 9027
rect 5917 8993 5951 9027
rect 6377 8993 6411 9027
rect 11253 8993 11287 9027
rect 5089 8925 5123 8959
rect 6653 8925 6687 8959
rect 8033 8925 8067 8959
rect 10057 8925 10091 8959
rect 6929 8789 6963 8823
rect 8953 8789 8987 8823
rect 11391 8789 11425 8823
rect 3249 8585 3283 8619
rect 4077 8585 4111 8619
rect 7757 8585 7791 8619
rect 8125 8585 8159 8619
rect 9689 8585 9723 8619
rect 11253 8585 11287 8619
rect 9229 8517 9263 8551
rect 10793 8517 10827 8551
rect 5917 8449 5951 8483
rect 6837 8449 6871 8483
rect 8677 8449 8711 8483
rect 10241 8449 10275 8483
rect 2789 8381 2823 8415
rect 3985 8381 4019 8415
rect 5181 8381 5215 8415
rect 5641 8381 5675 8415
rect 3801 8313 3835 8347
rect 7199 8313 7233 8347
rect 8769 8313 8803 8347
rect 10333 8313 10367 8347
rect 2697 8245 2731 8279
rect 2973 8245 3007 8279
rect 3617 8245 3651 8279
rect 4629 8245 4663 8279
rect 5089 8245 5123 8279
rect 6193 8245 6227 8279
rect 6653 8245 6687 8279
rect 8401 8245 8435 8279
rect 9965 8245 9999 8279
rect 2145 8041 2179 8075
rect 2789 8041 2823 8075
rect 3157 8041 3191 8075
rect 5825 8041 5859 8075
rect 6653 8041 6687 8075
rect 8033 8041 8067 8075
rect 9505 8041 9539 8075
rect 10793 8041 10827 8075
rect 7199 7973 7233 8007
rect 8723 7973 8757 8007
rect 9873 7973 9907 8007
rect 11391 7973 11425 8007
rect 1961 7905 1995 7939
rect 2973 7905 3007 7939
rect 3893 7905 3927 7939
rect 4077 7905 4111 7939
rect 4353 7905 4387 7939
rect 5641 7905 5675 7939
rect 6101 7905 6135 7939
rect 6837 7905 6871 7939
rect 8585 7905 8619 7939
rect 11253 7905 11287 7939
rect 2513 7837 2547 7871
rect 4537 7837 4571 7871
rect 9781 7837 9815 7871
rect 10057 7837 10091 7871
rect 4169 7769 4203 7803
rect 7757 7769 7791 7803
rect 3433 7701 3467 7735
rect 5273 7701 5307 7735
rect 1593 7497 1627 7531
rect 2605 7497 2639 7531
rect 2973 7497 3007 7531
rect 6193 7497 6227 7531
rect 7757 7497 7791 7531
rect 8493 7497 8527 7531
rect 9781 7497 9815 7531
rect 3525 7361 3559 7395
rect 4445 7361 4479 7395
rect 5917 7361 5951 7395
rect 8585 7361 8619 7395
rect 10425 7361 10459 7395
rect 10701 7361 10735 7395
rect 1409 7293 1443 7327
rect 2421 7293 2455 7327
rect 3157 7293 3191 7327
rect 3433 7293 3467 7327
rect 3709 7293 3743 7327
rect 5089 7293 5123 7327
rect 5365 7293 5399 7327
rect 5641 7293 5675 7327
rect 6837 7293 6871 7327
rect 8033 7293 8067 7327
rect 9505 7293 9539 7327
rect 10149 7293 10183 7327
rect 2329 7225 2363 7259
rect 6653 7225 6687 7259
rect 7199 7225 7233 7259
rect 8906 7225 8940 7259
rect 10517 7225 10551 7259
rect 1961 7157 1995 7191
rect 3157 7157 3191 7191
rect 3249 7157 3283 7191
rect 3893 7157 3927 7191
rect 11345 7157 11379 7191
rect 2881 6953 2915 6987
rect 3525 6953 3559 6987
rect 4537 6953 4571 6987
rect 6101 6953 6135 6987
rect 8125 6953 8159 6987
rect 10701 6953 10735 6987
rect 6929 6885 6963 6919
rect 7526 6885 7560 6919
rect 8585 6885 8619 6919
rect 8953 6885 8987 6919
rect 9505 6885 9539 6919
rect 9781 6885 9815 6919
rect 9873 6885 9907 6919
rect 2421 6817 2455 6851
rect 2697 6817 2731 6851
rect 3801 6817 3835 6851
rect 4077 6817 4111 6851
rect 4353 6817 4387 6851
rect 5641 6817 5675 6851
rect 5917 6817 5951 6851
rect 7205 6817 7239 6851
rect 5273 6749 5307 6783
rect 10057 6749 10091 6783
rect 2513 6681 2547 6715
rect 4169 6681 4203 6715
rect 5733 6681 5767 6715
rect 2145 6409 2179 6443
rect 9689 6409 9723 6443
rect 10425 6409 10459 6443
rect 9045 6341 9079 6375
rect 4997 6273 5031 6307
rect 8493 6273 8527 6307
rect 9965 6273 9999 6307
rect 3525 6205 3559 6239
rect 5089 6205 5123 6239
rect 6377 6205 6411 6239
rect 6837 6205 6871 6239
rect 7297 6205 7331 6239
rect 2513 6137 2547 6171
rect 4169 6137 4203 6171
rect 8217 6137 8251 6171
rect 8585 6137 8619 6171
rect 2789 6069 2823 6103
rect 3249 6069 3283 6103
rect 4537 6069 4571 6103
rect 4813 6069 4847 6103
rect 6009 6069 6043 6103
rect 7113 6069 7147 6103
rect 7849 6069 7883 6103
rect 3525 5865 3559 5899
rect 6469 5865 6503 5899
rect 6929 5865 6963 5899
rect 8033 5865 8067 5899
rect 9137 5865 9171 5899
rect 7434 5797 7468 5831
rect 8493 5797 8527 5831
rect 8769 5797 8803 5831
rect 3893 5729 3927 5763
rect 4065 5729 4099 5763
rect 4353 5729 4387 5763
rect 5641 5729 5675 5763
rect 5825 5729 5859 5763
rect 7113 5729 7147 5763
rect 9724 5729 9758 5763
rect 4537 5661 4571 5695
rect 5181 5661 5215 5695
rect 4169 5593 4203 5627
rect 5549 5525 5583 5559
rect 5917 5525 5951 5559
rect 9827 5525 9861 5559
rect 2697 5321 2731 5355
rect 3065 5321 3099 5355
rect 9597 5321 9631 5355
rect 4905 5253 4939 5287
rect 5181 5253 5215 5287
rect 9873 5253 9907 5287
rect 7389 5185 7423 5219
rect 10241 5185 10275 5219
rect 2513 5117 2547 5151
rect 3433 5117 3467 5151
rect 4077 5117 4111 5151
rect 4261 5117 4295 5151
rect 5365 5117 5399 5151
rect 5825 5117 5859 5151
rect 6837 5117 6871 5151
rect 9045 5117 9079 5151
rect 9689 5117 9723 5151
rect 10828 5117 10862 5151
rect 11253 5117 11287 5151
rect 6469 5049 6503 5083
rect 7757 5049 7791 5083
rect 8033 5049 8067 5083
rect 8125 5049 8159 5083
rect 8677 5049 8711 5083
rect 10931 5049 10965 5083
rect 4537 4981 4571 5015
rect 6193 4981 6227 5015
rect 7021 4981 7055 5015
rect 2881 4777 2915 4811
rect 4261 4777 4295 4811
rect 4721 4777 4755 4811
rect 7389 4777 7423 4811
rect 8953 4777 8987 4811
rect 9413 4777 9447 4811
rect 2605 4709 2639 4743
rect 6561 4709 6595 4743
rect 7113 4709 7147 4743
rect 8125 4709 8159 4743
rect 2789 4641 2823 4675
rect 5457 4641 5491 4675
rect 5825 4641 5859 4675
rect 9873 4641 9907 4675
rect 11288 4641 11322 4675
rect 5549 4573 5583 4607
rect 6469 4573 6503 4607
rect 7757 4573 7791 4607
rect 8033 4573 8067 4607
rect 8677 4573 8711 4607
rect 9689 4573 9723 4607
rect 6193 4437 6227 4471
rect 11391 4437 11425 4471
rect 2789 4233 2823 4267
rect 4261 4233 4295 4267
rect 6193 4233 6227 4267
rect 7757 4233 7791 4267
rect 11253 4233 11287 4267
rect 9229 4165 9263 4199
rect 3985 4097 4019 4131
rect 8677 4097 8711 4131
rect 2145 4029 2179 4063
rect 2304 4029 2338 4063
rect 3341 4029 3375 4063
rect 5089 4029 5123 4063
rect 5273 4029 5307 4063
rect 5641 4029 5675 4063
rect 6837 4029 6871 4063
rect 10057 4029 10091 4063
rect 10241 4029 10275 4063
rect 3157 3961 3191 3995
rect 4721 3961 4755 3995
rect 5917 3961 5951 3995
rect 7158 3961 7192 3995
rect 8493 3961 8527 3995
rect 8769 3961 8803 3995
rect 10149 3961 10183 3995
rect 2375 3893 2409 3927
rect 6653 3893 6687 3927
rect 8125 3893 8159 3927
rect 9689 3893 9723 3927
rect 2697 3689 2731 3723
rect 3111 3689 3145 3723
rect 6009 3689 6043 3723
rect 8125 3689 8159 3723
rect 6653 3621 6687 3655
rect 7158 3621 7192 3655
rect 9873 3621 9907 3655
rect 11253 3621 11287 3655
rect 3040 3553 3074 3587
rect 4353 3553 4387 3587
rect 4721 3553 4755 3587
rect 5089 3553 5123 3587
rect 5733 3553 5767 3587
rect 6285 3553 6319 3587
rect 7757 3553 7791 3587
rect 11805 3553 11839 3587
rect 12817 3553 12851 3587
rect 5641 3485 5675 3519
rect 6837 3485 6871 3519
rect 8585 3485 8619 3519
rect 9781 3485 9815 3519
rect 10333 3417 10367 3451
rect 9413 3349 9447 3383
rect 12955 3349 12989 3383
rect 2605 3145 2639 3179
rect 3065 3145 3099 3179
rect 4629 3145 4663 3179
rect 8401 3145 8435 3179
rect 8861 3145 8895 3179
rect 10333 3145 10367 3179
rect 11805 3145 11839 3179
rect 12909 3145 12943 3179
rect 4353 3077 4387 3111
rect 7757 3077 7791 3111
rect 11069 3077 11103 3111
rect 3341 3009 3375 3043
rect 3985 3009 4019 3043
rect 9413 3009 9447 3043
rect 10057 3009 10091 3043
rect 4813 2941 4847 2975
rect 5457 2941 5491 2975
rect 5641 2941 5675 2975
rect 6837 2941 6871 2975
rect 8033 2941 8067 2975
rect 10885 2941 10919 2975
rect 11437 2941 11471 2975
rect 12500 2941 12534 2975
rect 13277 2941 13311 2975
rect 3433 2873 3467 2907
rect 7158 2873 7192 2907
rect 9229 2873 9263 2907
rect 9505 2873 9539 2907
rect 12587 2873 12621 2907
rect 5917 2805 5951 2839
rect 6285 2805 6319 2839
rect 6653 2805 6687 2839
rect 3341 2601 3375 2635
rect 3893 2601 3927 2635
rect 5825 2601 5859 2635
rect 7849 2601 7883 2635
rect 8677 2601 8711 2635
rect 9597 2601 9631 2635
rect 1961 2533 1995 2567
rect 7250 2533 7284 2567
rect 9137 2533 9171 2567
rect 9873 2533 9907 2567
rect 9965 2533 9999 2567
rect 2053 2465 2087 2499
rect 4721 2465 4755 2499
rect 5549 2465 5583 2499
rect 6929 2465 6963 2499
rect 8125 2465 8159 2499
rect 11345 2465 11379 2499
rect 11897 2465 11931 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 5457 2397 5491 2431
rect 6101 2397 6135 2431
rect 10149 2397 10183 2431
rect 1777 2261 1811 2295
rect 4537 2261 4571 2295
rect 6653 2261 6687 2295
rect 11529 2261 11563 2295
rect 12817 2261 12851 2295
<< metal1 >>
rect 658 39584 664 39636
rect 716 39624 722 39636
rect 2498 39624 2504 39636
rect 716 39596 2504 39624
rect 716 39584 722 39596
rect 2498 39584 2504 39596
rect 2556 39584 2562 39636
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 9766 35980 9772 36032
rect 9824 36020 9830 36032
rect 15470 36020 15476 36032
rect 9824 35992 15476 36020
rect 9824 35980 9830 35992
rect 15470 35980 15476 35992
rect 15528 35980 15534 36032
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 9766 35816 9772 35828
rect 9727 35788 9772 35816
rect 9766 35776 9772 35788
rect 9824 35776 9830 35828
rect 8478 35680 8484 35692
rect 8439 35652 8484 35680
rect 8478 35640 8484 35652
rect 8536 35680 8542 35692
rect 8536 35652 9076 35680
rect 8536 35640 8542 35652
rect 4154 35572 4160 35624
rect 4212 35612 4218 35624
rect 6892 35615 6950 35621
rect 6892 35612 6904 35615
rect 4212 35584 6904 35612
rect 4212 35572 4218 35584
rect 6892 35581 6904 35584
rect 6938 35612 6950 35615
rect 9048 35612 9076 35652
rect 9528 35615 9586 35621
rect 9528 35612 9540 35615
rect 6938 35584 7420 35612
rect 9048 35584 9540 35612
rect 6938 35581 6950 35584
rect 6892 35575 6950 35581
rect 4890 35476 4896 35488
rect 4851 35448 4896 35476
rect 4890 35436 4896 35448
rect 4948 35436 4954 35488
rect 6730 35436 6736 35488
rect 6788 35476 6794 35488
rect 7392 35485 7420 35584
rect 9528 35581 9540 35584
rect 9574 35612 9586 35615
rect 9953 35615 10011 35621
rect 9953 35612 9965 35615
rect 9574 35584 9965 35612
rect 9574 35581 9586 35584
rect 9528 35575 9586 35581
rect 9953 35581 9965 35584
rect 9999 35581 10011 35615
rect 9953 35575 10011 35581
rect 7837 35547 7895 35553
rect 7837 35513 7849 35547
rect 7883 35544 7895 35547
rect 8018 35544 8024 35556
rect 7883 35516 8024 35544
rect 7883 35513 7895 35516
rect 7837 35507 7895 35513
rect 8018 35504 8024 35516
rect 8076 35504 8082 35556
rect 8110 35504 8116 35556
rect 8168 35544 8174 35556
rect 8168 35516 8213 35544
rect 8168 35504 8174 35516
rect 6963 35479 7021 35485
rect 6963 35476 6975 35479
rect 6788 35448 6975 35476
rect 6788 35436 6794 35448
rect 6963 35445 6975 35448
rect 7009 35445 7021 35479
rect 6963 35439 7021 35445
rect 7377 35479 7435 35485
rect 7377 35445 7389 35479
rect 7423 35476 7435 35479
rect 9674 35476 9680 35488
rect 7423 35448 9680 35476
rect 7423 35445 7435 35448
rect 7377 35439 7435 35445
rect 9674 35436 9680 35448
rect 9732 35436 9738 35488
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 106 35232 112 35284
rect 164 35272 170 35284
rect 4203 35275 4261 35281
rect 4203 35272 4215 35275
rect 164 35244 4215 35272
rect 164 35232 170 35244
rect 4203 35241 4215 35244
rect 4249 35241 4261 35275
rect 4203 35235 4261 35241
rect 8021 35275 8079 35281
rect 8021 35241 8033 35275
rect 8067 35272 8079 35275
rect 8110 35272 8116 35284
rect 8067 35244 8116 35272
rect 8067 35241 8079 35244
rect 8021 35235 8079 35241
rect 8110 35232 8116 35244
rect 8168 35232 8174 35284
rect 8846 35232 8852 35284
rect 8904 35272 8910 35284
rect 9861 35275 9919 35281
rect 9861 35272 9873 35275
rect 8904 35244 9873 35272
rect 8904 35232 8910 35244
rect 9861 35241 9873 35244
rect 9907 35241 9919 35275
rect 9861 35235 9919 35241
rect 5258 35204 5264 35216
rect 5219 35176 5264 35204
rect 5258 35164 5264 35176
rect 5316 35164 5322 35216
rect 7101 35207 7159 35213
rect 7101 35173 7113 35207
rect 7147 35204 7159 35207
rect 7742 35204 7748 35216
rect 7147 35176 7748 35204
rect 7147 35173 7159 35176
rect 7101 35167 7159 35173
rect 7742 35164 7748 35176
rect 7800 35164 7806 35216
rect 3970 35096 3976 35148
rect 4028 35136 4034 35148
rect 4111 35139 4169 35145
rect 4111 35136 4123 35139
rect 4028 35108 4123 35136
rect 4028 35096 4034 35108
rect 4111 35105 4123 35108
rect 4157 35105 4169 35139
rect 4111 35099 4169 35105
rect 4126 35000 4154 35099
rect 8386 35096 8392 35148
rect 8444 35136 8450 35148
rect 8481 35139 8539 35145
rect 8481 35136 8493 35139
rect 8444 35108 8493 35136
rect 8444 35096 8450 35108
rect 8481 35105 8493 35108
rect 8527 35105 8539 35139
rect 9674 35136 9680 35148
rect 9587 35108 9680 35136
rect 8481 35099 8539 35105
rect 9674 35096 9680 35108
rect 9732 35136 9738 35148
rect 11422 35136 11428 35148
rect 9732 35108 11428 35136
rect 9732 35096 9738 35108
rect 11422 35096 11428 35108
rect 11480 35096 11486 35148
rect 4890 35028 4896 35080
rect 4948 35068 4954 35080
rect 5169 35071 5227 35077
rect 5169 35068 5181 35071
rect 4948 35040 5181 35068
rect 4948 35028 4954 35040
rect 5169 35037 5181 35040
rect 5215 35068 5227 35071
rect 5994 35068 6000 35080
rect 5215 35040 6000 35068
rect 5215 35037 5227 35040
rect 5169 35031 5227 35037
rect 5994 35028 6000 35040
rect 6052 35028 6058 35080
rect 6730 35028 6736 35080
rect 6788 35068 6794 35080
rect 7009 35071 7067 35077
rect 7009 35068 7021 35071
rect 6788 35040 7021 35068
rect 6788 35028 6794 35040
rect 7009 35037 7021 35040
rect 7055 35037 7067 35071
rect 7009 35031 7067 35037
rect 7653 35071 7711 35077
rect 7653 35037 7665 35071
rect 7699 35068 7711 35071
rect 8570 35068 8576 35080
rect 7699 35040 8576 35068
rect 7699 35037 7711 35040
rect 7653 35031 7711 35037
rect 8570 35028 8576 35040
rect 8628 35028 8634 35080
rect 5718 35000 5724 35012
rect 4126 34972 5724 35000
rect 5718 34960 5724 34972
rect 5776 34960 5782 35012
rect 8665 35003 8723 35009
rect 8665 34969 8677 35003
rect 8711 35000 8723 35003
rect 9766 35000 9772 35012
rect 8711 34972 9772 35000
rect 8711 34969 8723 34972
rect 8665 34963 8723 34969
rect 9766 34960 9772 34972
rect 9824 34960 9830 35012
rect 4798 34932 4804 34944
rect 4759 34904 4804 34932
rect 4798 34892 4804 34904
rect 4856 34892 4862 34944
rect 6822 34932 6828 34944
rect 6783 34904 6828 34932
rect 6822 34892 6828 34904
rect 6880 34892 6886 34944
rect 8754 34892 8760 34944
rect 8812 34932 8818 34944
rect 9033 34935 9091 34941
rect 9033 34932 9045 34935
rect 8812 34904 9045 34932
rect 8812 34892 8818 34904
rect 9033 34901 9045 34904
rect 9079 34901 9091 34935
rect 9033 34895 9091 34901
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 3510 34688 3516 34740
rect 3568 34728 3574 34740
rect 3881 34731 3939 34737
rect 3881 34728 3893 34731
rect 3568 34700 3893 34728
rect 3568 34688 3574 34700
rect 3881 34697 3893 34700
rect 3927 34697 3939 34731
rect 3881 34691 3939 34697
rect 5258 34688 5264 34740
rect 5316 34728 5322 34740
rect 5626 34728 5632 34740
rect 5316 34700 5632 34728
rect 5316 34688 5322 34700
rect 5626 34688 5632 34700
rect 5684 34728 5690 34740
rect 5721 34731 5779 34737
rect 5721 34728 5733 34731
rect 5684 34700 5733 34728
rect 5684 34688 5690 34700
rect 5721 34697 5733 34700
rect 5767 34697 5779 34731
rect 5994 34728 6000 34740
rect 5955 34700 6000 34728
rect 5721 34691 5779 34697
rect 5994 34688 6000 34700
rect 6052 34688 6058 34740
rect 7745 34731 7803 34737
rect 7745 34697 7757 34731
rect 7791 34728 7803 34731
rect 8110 34728 8116 34740
rect 7791 34700 8116 34728
rect 7791 34697 7803 34700
rect 7745 34691 7803 34697
rect 8110 34688 8116 34700
rect 8168 34688 8174 34740
rect 9674 34728 9680 34740
rect 9635 34700 9680 34728
rect 9674 34688 9680 34700
rect 9732 34688 9738 34740
rect 12713 34731 12771 34737
rect 12713 34697 12725 34731
rect 12759 34728 12771 34731
rect 13722 34728 13728 34740
rect 12759 34700 13728 34728
rect 12759 34697 12771 34700
rect 12713 34691 12771 34697
rect 13722 34688 13728 34700
rect 13780 34688 13786 34740
rect 3605 34663 3663 34669
rect 3605 34629 3617 34663
rect 3651 34660 3663 34663
rect 3970 34660 3976 34672
rect 3651 34632 3976 34660
rect 3651 34629 3663 34632
rect 3605 34623 3663 34629
rect 3970 34620 3976 34632
rect 4028 34620 4034 34672
rect 7834 34620 7840 34672
rect 7892 34660 7898 34672
rect 8478 34660 8484 34672
rect 7892 34632 8484 34660
rect 7892 34620 7898 34632
rect 8478 34620 8484 34632
rect 8536 34660 8542 34672
rect 9217 34663 9275 34669
rect 9217 34660 9229 34663
rect 8536 34632 9229 34660
rect 8536 34620 8542 34632
rect 9217 34629 9229 34632
rect 9263 34629 9275 34663
rect 9217 34623 9275 34629
rect 4798 34592 4804 34604
rect 4759 34564 4804 34592
rect 4798 34552 4804 34564
rect 4856 34552 4862 34604
rect 8018 34552 8024 34604
rect 8076 34592 8082 34604
rect 10137 34595 10195 34601
rect 10137 34592 10149 34595
rect 8076 34564 10149 34592
rect 8076 34552 8082 34564
rect 10137 34561 10149 34564
rect 10183 34561 10195 34595
rect 10137 34555 10195 34561
rect 3697 34527 3755 34533
rect 3697 34493 3709 34527
rect 3743 34524 3755 34527
rect 6822 34524 6828 34536
rect 3743 34496 4016 34524
rect 6735 34496 6828 34524
rect 3743 34493 3755 34496
rect 3697 34487 3755 34493
rect 3988 34400 4016 34496
rect 6822 34484 6828 34496
rect 6880 34524 6886 34536
rect 6880 34496 8524 34524
rect 6880 34484 6886 34496
rect 4614 34416 4620 34468
rect 4672 34456 4678 34468
rect 4709 34459 4767 34465
rect 4709 34456 4721 34459
rect 4672 34428 4721 34456
rect 4672 34416 4678 34428
rect 4709 34425 4721 34428
rect 4755 34456 4767 34459
rect 5122 34459 5180 34465
rect 5122 34456 5134 34459
rect 4755 34428 5134 34456
rect 4755 34425 4767 34428
rect 4709 34419 4767 34425
rect 5122 34425 5134 34428
rect 5168 34456 5180 34459
rect 6549 34459 6607 34465
rect 6549 34456 6561 34459
rect 5168 34428 6561 34456
rect 5168 34425 5180 34428
rect 5122 34419 5180 34425
rect 6549 34425 6561 34428
rect 6595 34456 6607 34459
rect 7006 34456 7012 34468
rect 6595 34428 7012 34456
rect 6595 34425 6607 34428
rect 6549 34419 6607 34425
rect 7006 34416 7012 34428
rect 7064 34456 7070 34468
rect 7146 34459 7204 34465
rect 7146 34456 7158 34459
rect 7064 34428 7158 34456
rect 7064 34416 7070 34428
rect 7146 34425 7158 34428
rect 7192 34425 7204 34459
rect 7146 34419 7204 34425
rect 3970 34348 3976 34400
rect 4028 34388 4034 34400
rect 4249 34391 4307 34397
rect 4249 34388 4261 34391
rect 4028 34360 4261 34388
rect 4028 34348 4034 34360
rect 4249 34357 4261 34360
rect 4295 34357 4307 34391
rect 4249 34351 4307 34357
rect 7742 34348 7748 34400
rect 7800 34388 7806 34400
rect 8021 34391 8079 34397
rect 8021 34388 8033 34391
rect 7800 34360 8033 34388
rect 7800 34348 7806 34360
rect 8021 34357 8033 34360
rect 8067 34357 8079 34391
rect 8386 34388 8392 34400
rect 8347 34360 8392 34388
rect 8021 34351 8079 34357
rect 8386 34348 8392 34360
rect 8444 34348 8450 34400
rect 8496 34388 8524 34496
rect 10778 34484 10784 34536
rect 10836 34524 10842 34536
rect 12529 34527 12587 34533
rect 12529 34524 12541 34527
rect 10836 34496 12541 34524
rect 10836 34484 10842 34496
rect 12529 34493 12541 34496
rect 12575 34524 12587 34527
rect 13081 34527 13139 34533
rect 13081 34524 13093 34527
rect 12575 34496 13093 34524
rect 12575 34493 12587 34496
rect 12529 34487 12587 34493
rect 13081 34493 13093 34496
rect 13127 34493 13139 34527
rect 13081 34487 13139 34493
rect 8662 34456 8668 34468
rect 8623 34428 8668 34456
rect 8662 34416 8668 34428
rect 8720 34416 8726 34468
rect 8754 34416 8760 34468
rect 8812 34456 8818 34468
rect 8812 34428 8857 34456
rect 8812 34416 8818 34428
rect 8846 34388 8852 34400
rect 8496 34360 8852 34388
rect 8846 34348 8852 34360
rect 8904 34348 8910 34400
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 4798 34144 4804 34196
rect 4856 34184 4862 34196
rect 4893 34187 4951 34193
rect 4893 34184 4905 34187
rect 4856 34156 4905 34184
rect 4856 34144 4862 34156
rect 4893 34153 4905 34156
rect 4939 34153 4951 34187
rect 5626 34184 5632 34196
rect 5587 34156 5632 34184
rect 4893 34147 4951 34153
rect 5626 34144 5632 34156
rect 5684 34144 5690 34196
rect 6549 34187 6607 34193
rect 6549 34153 6561 34187
rect 6595 34184 6607 34187
rect 6730 34184 6736 34196
rect 6595 34156 6736 34184
rect 6595 34153 6607 34156
rect 6549 34147 6607 34153
rect 6730 34144 6736 34156
rect 6788 34144 6794 34196
rect 7006 34184 7012 34196
rect 6967 34156 7012 34184
rect 7006 34144 7012 34156
rect 7064 34144 7070 34196
rect 7561 34187 7619 34193
rect 7561 34153 7573 34187
rect 7607 34184 7619 34187
rect 8754 34184 8760 34196
rect 7607 34156 8760 34184
rect 7607 34153 7619 34156
rect 7561 34147 7619 34153
rect 8754 34144 8760 34156
rect 8812 34144 8818 34196
rect 8846 34144 8852 34196
rect 8904 34184 8910 34196
rect 9769 34187 9827 34193
rect 9769 34184 9781 34187
rect 8904 34156 9781 34184
rect 8904 34144 8910 34156
rect 9769 34153 9781 34156
rect 9815 34153 9827 34187
rect 9769 34147 9827 34153
rect 8662 34076 8668 34128
rect 8720 34116 8726 34128
rect 9309 34119 9367 34125
rect 9309 34116 9321 34119
rect 8720 34088 9321 34116
rect 8720 34076 8726 34088
rect 8864 34060 8892 34088
rect 9309 34085 9321 34088
rect 9355 34085 9367 34119
rect 9309 34079 9367 34085
rect 4706 34048 4712 34060
rect 4667 34020 4712 34048
rect 4706 34008 4712 34020
rect 4764 34008 4770 34060
rect 5077 34051 5135 34057
rect 5077 34048 5089 34051
rect 4816 34020 5089 34048
rect 3329 33983 3387 33989
rect 3329 33949 3341 33983
rect 3375 33980 3387 33983
rect 3510 33980 3516 33992
rect 3375 33952 3516 33980
rect 3375 33949 3387 33952
rect 3329 33943 3387 33949
rect 3510 33940 3516 33952
rect 3568 33980 3574 33992
rect 4816 33980 4844 34020
rect 5077 34017 5089 34020
rect 5123 34017 5135 34051
rect 5077 34011 5135 34017
rect 8389 34051 8447 34057
rect 8389 34017 8401 34051
rect 8435 34048 8447 34051
rect 8478 34048 8484 34060
rect 8435 34020 8484 34048
rect 8435 34017 8447 34020
rect 8389 34011 8447 34017
rect 8478 34008 8484 34020
rect 8536 34048 8542 34060
rect 8536 34020 8800 34048
rect 8536 34008 8542 34020
rect 6638 33980 6644 33992
rect 3568 33952 4844 33980
rect 6599 33952 6644 33980
rect 3568 33940 3574 33952
rect 6638 33940 6644 33952
rect 6696 33940 6702 33992
rect 7650 33872 7656 33924
rect 7708 33912 7714 33924
rect 8573 33915 8631 33921
rect 8573 33912 8585 33915
rect 7708 33884 8585 33912
rect 7708 33872 7714 33884
rect 8573 33881 8585 33884
rect 8619 33881 8631 33915
rect 8772 33912 8800 34020
rect 8846 34008 8852 34060
rect 8904 34008 8910 34060
rect 9950 34048 9956 34060
rect 9911 34020 9956 34048
rect 9950 34008 9956 34020
rect 10008 34008 10014 34060
rect 10137 34051 10195 34057
rect 10137 34017 10149 34051
rect 10183 34048 10195 34051
rect 10689 34051 10747 34057
rect 10689 34048 10701 34051
rect 10183 34020 10701 34048
rect 10183 34017 10195 34020
rect 10137 34011 10195 34017
rect 10689 34017 10701 34020
rect 10735 34048 10747 34051
rect 10962 34048 10968 34060
rect 10735 34020 10968 34048
rect 10735 34017 10747 34020
rect 10689 34011 10747 34017
rect 9398 33940 9404 33992
rect 9456 33980 9462 33992
rect 10152 33980 10180 34011
rect 10962 34008 10968 34020
rect 11020 34008 11026 34060
rect 11238 34048 11244 34060
rect 11199 34020 11244 34048
rect 11238 34008 11244 34020
rect 11296 34008 11302 34060
rect 11422 33980 11428 33992
rect 9456 33952 10180 33980
rect 9456 33940 9462 33952
rect 11394 33940 11428 33980
rect 11480 33940 11486 33992
rect 9582 33912 9588 33924
rect 8772 33884 9588 33912
rect 8573 33875 8631 33881
rect 9582 33872 9588 33884
rect 9640 33872 9646 33924
rect 8754 33804 8760 33856
rect 8812 33844 8818 33856
rect 11394 33853 11422 33940
rect 8941 33847 8999 33853
rect 8941 33844 8953 33847
rect 8812 33816 8953 33844
rect 8812 33804 8818 33816
rect 8941 33813 8953 33816
rect 8987 33813 8999 33847
rect 8941 33807 8999 33813
rect 11379 33847 11437 33853
rect 11379 33813 11391 33847
rect 11425 33813 11437 33847
rect 11379 33807 11437 33813
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 4614 33640 4620 33652
rect 4575 33612 4620 33640
rect 4614 33600 4620 33612
rect 4672 33600 4678 33652
rect 8478 33640 8484 33652
rect 8439 33612 8484 33640
rect 8478 33600 8484 33612
rect 8536 33600 8542 33652
rect 9490 33600 9496 33652
rect 9548 33640 9554 33652
rect 9950 33640 9956 33652
rect 9548 33612 9956 33640
rect 9548 33600 9554 33612
rect 9950 33600 9956 33612
rect 10008 33600 10014 33652
rect 9674 33572 9680 33584
rect 4126 33544 9680 33572
rect 4126 33504 4154 33544
rect 9674 33532 9680 33544
rect 9732 33572 9738 33584
rect 10413 33575 10471 33581
rect 10413 33572 10425 33575
rect 9732 33544 10425 33572
rect 9732 33532 9738 33544
rect 10413 33541 10425 33544
rect 10459 33572 10471 33575
rect 10594 33572 10600 33584
rect 10459 33544 10600 33572
rect 10459 33541 10471 33544
rect 10413 33535 10471 33541
rect 10594 33532 10600 33544
rect 10652 33532 10658 33584
rect 3528 33476 4154 33504
rect 4341 33507 4399 33513
rect 3528 33445 3556 33476
rect 4341 33473 4353 33507
rect 4387 33504 4399 33507
rect 4706 33504 4712 33516
rect 4387 33476 4712 33504
rect 4387 33473 4399 33476
rect 4341 33467 4399 33473
rect 4706 33464 4712 33476
rect 4764 33504 4770 33516
rect 7650 33504 7656 33516
rect 4764 33476 7656 33504
rect 4764 33464 4770 33476
rect 7650 33464 7656 33476
rect 7708 33464 7714 33516
rect 8754 33504 8760 33516
rect 8715 33476 8760 33504
rect 8754 33464 8760 33476
rect 8812 33464 8818 33516
rect 10318 33464 10324 33516
rect 10376 33504 10382 33516
rect 11238 33504 11244 33516
rect 10376 33476 11244 33504
rect 10376 33464 10382 33476
rect 11238 33464 11244 33476
rect 11296 33504 11302 33516
rect 11517 33507 11575 33513
rect 11517 33504 11529 33507
rect 11296 33476 11529 33504
rect 11296 33464 11302 33476
rect 11517 33473 11529 33476
rect 11563 33473 11575 33507
rect 11517 33467 11575 33473
rect 3145 33439 3203 33445
rect 3145 33405 3157 33439
rect 3191 33436 3203 33439
rect 3513 33439 3571 33445
rect 3513 33436 3525 33439
rect 3191 33408 3525 33436
rect 3191 33405 3203 33408
rect 3145 33399 3203 33405
rect 3513 33405 3525 33408
rect 3559 33405 3571 33439
rect 3513 33399 3571 33405
rect 3602 33396 3608 33448
rect 3660 33436 3666 33448
rect 3697 33439 3755 33445
rect 3697 33436 3709 33439
rect 3660 33408 3709 33436
rect 3660 33396 3666 33408
rect 3697 33405 3709 33408
rect 3743 33405 3755 33439
rect 3697 33399 3755 33405
rect 3973 33439 4031 33445
rect 3973 33405 3985 33439
rect 4019 33436 4031 33439
rect 4801 33439 4859 33445
rect 4801 33436 4813 33439
rect 4019 33408 4813 33436
rect 4019 33405 4031 33408
rect 3973 33399 4031 33405
rect 4801 33405 4813 33408
rect 4847 33436 4859 33439
rect 4982 33436 4988 33448
rect 4847 33408 4988 33436
rect 4847 33405 4859 33408
rect 4801 33399 4859 33405
rect 4982 33396 4988 33408
rect 5040 33396 5046 33448
rect 5258 33396 5264 33448
rect 5316 33436 5322 33448
rect 6825 33439 6883 33445
rect 6825 33436 6837 33439
rect 5316 33408 6837 33436
rect 5316 33396 5322 33408
rect 6825 33405 6837 33408
rect 6871 33436 6883 33439
rect 8021 33439 8079 33445
rect 8021 33436 8033 33439
rect 6871 33408 8033 33436
rect 6871 33405 6883 33408
rect 6825 33399 6883 33405
rect 8021 33405 8033 33408
rect 8067 33405 8079 33439
rect 8021 33399 8079 33405
rect 9306 33396 9312 33448
rect 9364 33436 9370 33448
rect 10594 33436 10600 33448
rect 9364 33408 9674 33436
rect 10555 33408 10600 33436
rect 9364 33396 9370 33408
rect 4614 33328 4620 33380
rect 4672 33368 4678 33380
rect 5122 33371 5180 33377
rect 5122 33368 5134 33371
rect 4672 33340 5134 33368
rect 4672 33328 4678 33340
rect 5122 33337 5134 33340
rect 5168 33368 5180 33371
rect 6181 33371 6239 33377
rect 6181 33368 6193 33371
rect 5168 33340 6193 33368
rect 5168 33337 5180 33340
rect 5122 33331 5180 33337
rect 6181 33337 6193 33340
rect 6227 33368 6239 33371
rect 6549 33371 6607 33377
rect 6549 33368 6561 33371
rect 6227 33340 6561 33368
rect 6227 33337 6239 33340
rect 6181 33331 6239 33337
rect 6549 33337 6561 33340
rect 6595 33368 6607 33371
rect 6730 33368 6736 33380
rect 6595 33340 6736 33368
rect 6595 33337 6607 33340
rect 6549 33331 6607 33337
rect 6730 33328 6736 33340
rect 6788 33368 6794 33380
rect 7146 33371 7204 33377
rect 7146 33368 7158 33371
rect 6788 33340 7158 33368
rect 6788 33328 6794 33340
rect 7146 33337 7158 33340
rect 7192 33337 7204 33371
rect 9646 33368 9674 33408
rect 10594 33396 10600 33408
rect 10652 33396 10658 33448
rect 10962 33436 10968 33448
rect 10923 33408 10968 33436
rect 10962 33396 10968 33408
rect 11020 33396 11026 33448
rect 9646 33340 10456 33368
rect 7146 33331 7204 33337
rect 5718 33300 5724 33312
rect 5679 33272 5724 33300
rect 5718 33260 5724 33272
rect 5776 33260 5782 33312
rect 7006 33260 7012 33312
rect 7064 33300 7070 33312
rect 7742 33300 7748 33312
rect 7064 33272 7748 33300
rect 7064 33260 7070 33272
rect 7742 33260 7748 33272
rect 7800 33260 7806 33312
rect 9122 33300 9128 33312
rect 9083 33272 9128 33300
rect 9122 33260 9128 33272
rect 9180 33260 9186 33312
rect 9582 33260 9588 33312
rect 9640 33300 9646 33312
rect 9677 33303 9735 33309
rect 9677 33300 9689 33303
rect 9640 33272 9689 33300
rect 9640 33260 9646 33272
rect 9677 33269 9689 33272
rect 9723 33269 9735 33303
rect 10428 33300 10456 33340
rect 10597 33303 10655 33309
rect 10597 33300 10609 33303
rect 10428 33272 10609 33300
rect 9677 33263 9735 33269
rect 10597 33269 10609 33272
rect 10643 33269 10655 33303
rect 10597 33263 10655 33269
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 4982 33096 4988 33108
rect 4943 33068 4988 33096
rect 4982 33056 4988 33068
rect 5040 33056 5046 33108
rect 6638 33096 6644 33108
rect 6551 33068 6644 33096
rect 6638 33056 6644 33068
rect 6696 33096 6702 33108
rect 9306 33096 9312 33108
rect 6696 33068 9312 33096
rect 6696 33056 6702 33068
rect 9306 33056 9312 33068
rect 9364 33056 9370 33108
rect 10778 33096 10784 33108
rect 9416 33068 10784 33096
rect 3145 33031 3203 33037
rect 3145 32997 3157 33031
rect 3191 33028 3203 33031
rect 5258 33028 5264 33040
rect 3191 33000 5264 33028
rect 3191 32997 3203 33000
rect 3145 32991 3203 32997
rect 5258 32988 5264 33000
rect 5316 32988 5322 33040
rect 5353 33031 5411 33037
rect 5353 32997 5365 33031
rect 5399 33028 5411 33031
rect 5534 33028 5540 33040
rect 5399 33000 5540 33028
rect 5399 32997 5411 33000
rect 5353 32991 5411 32997
rect 5534 32988 5540 33000
rect 5592 33028 5598 33040
rect 5718 33028 5724 33040
rect 5592 33000 5724 33028
rect 5592 32988 5598 33000
rect 5718 32988 5724 33000
rect 5776 32988 5782 33040
rect 6730 32988 6736 33040
rect 6788 33028 6794 33040
rect 7054 33031 7112 33037
rect 7054 33028 7066 33031
rect 6788 33000 7066 33028
rect 6788 32988 6794 33000
rect 7054 32997 7066 33000
rect 7100 32997 7112 33031
rect 9416 33028 9444 33068
rect 10778 33056 10784 33068
rect 10836 33056 10842 33108
rect 11422 33096 11428 33108
rect 11383 33068 11428 33096
rect 11422 33056 11428 33068
rect 11480 33056 11486 33108
rect 7054 32991 7112 32997
rect 8680 33000 9444 33028
rect 8680 32972 8708 33000
rect 9490 32988 9496 33040
rect 9548 33028 9554 33040
rect 9953 33031 10011 33037
rect 9953 33028 9965 33031
rect 9548 33000 9965 33028
rect 9548 32988 9554 33000
rect 9953 32997 9965 33000
rect 9999 32997 10011 33031
rect 9953 32991 10011 32997
rect 10042 32988 10048 33040
rect 10100 33028 10106 33040
rect 12158 33028 12164 33040
rect 10100 33000 12164 33028
rect 10100 32988 10106 33000
rect 12158 32988 12164 33000
rect 12216 32988 12222 33040
rect 2682 32960 2688 32972
rect 2643 32932 2688 32960
rect 2682 32920 2688 32932
rect 2740 32920 2746 32972
rect 2866 32920 2872 32972
rect 2924 32960 2930 32972
rect 2961 32963 3019 32969
rect 2961 32960 2973 32963
rect 2924 32932 2973 32960
rect 2924 32920 2930 32932
rect 2961 32929 2973 32932
rect 3007 32960 3019 32963
rect 4893 32963 4951 32969
rect 4893 32960 4905 32963
rect 3007 32932 4905 32960
rect 3007 32929 3019 32932
rect 2961 32923 3019 32929
rect 4893 32929 4905 32932
rect 4939 32929 4951 32963
rect 4893 32923 4951 32929
rect 8548 32963 8606 32969
rect 8548 32929 8560 32963
rect 8594 32960 8606 32963
rect 8662 32960 8668 32972
rect 8594 32932 8668 32960
rect 8594 32929 8606 32932
rect 8548 32923 8606 32929
rect 8662 32920 8668 32932
rect 8720 32920 8726 32972
rect 9398 32960 9404 32972
rect 9359 32932 9404 32960
rect 9398 32920 9404 32932
rect 9456 32920 9462 32972
rect 10594 32920 10600 32972
rect 10652 32960 10658 32972
rect 11333 32963 11391 32969
rect 11333 32960 11345 32963
rect 10652 32932 11345 32960
rect 10652 32920 10658 32932
rect 11333 32929 11345 32932
rect 11379 32960 11391 32963
rect 11606 32960 11612 32972
rect 11379 32932 11612 32960
rect 11379 32929 11391 32932
rect 11333 32923 11391 32929
rect 11606 32920 11612 32932
rect 11664 32920 11670 32972
rect 11793 32963 11851 32969
rect 11793 32929 11805 32963
rect 11839 32929 11851 32963
rect 11793 32923 11851 32929
rect 4341 32895 4399 32901
rect 4341 32861 4353 32895
rect 4387 32892 4399 32895
rect 5261 32895 5319 32901
rect 5261 32892 5273 32895
rect 4387 32864 5273 32892
rect 4387 32861 4399 32864
rect 4341 32855 4399 32861
rect 5261 32861 5273 32864
rect 5307 32892 5319 32895
rect 5442 32892 5448 32904
rect 5307 32864 5448 32892
rect 5307 32861 5319 32864
rect 5261 32855 5319 32861
rect 5442 32852 5448 32864
rect 5500 32852 5506 32904
rect 5626 32892 5632 32904
rect 5587 32864 5632 32892
rect 5626 32852 5632 32864
rect 5684 32852 5690 32904
rect 5902 32852 5908 32904
rect 5960 32892 5966 32904
rect 6733 32895 6791 32901
rect 6733 32892 6745 32895
rect 5960 32864 6745 32892
rect 5960 32852 5966 32864
rect 6733 32861 6745 32864
rect 6779 32861 6791 32895
rect 6733 32855 6791 32861
rect 7098 32852 7104 32904
rect 7156 32892 7162 32904
rect 9416 32892 9444 32920
rect 7156 32864 9444 32892
rect 9861 32895 9919 32901
rect 7156 32852 7162 32864
rect 9861 32861 9873 32895
rect 9907 32861 9919 32895
rect 10318 32892 10324 32904
rect 10279 32864 10324 32892
rect 9861 32855 9919 32861
rect 4617 32827 4675 32833
rect 4617 32824 4629 32827
rect 4126 32796 4629 32824
rect 3510 32716 3516 32768
rect 3568 32756 3574 32768
rect 4126 32756 4154 32796
rect 4617 32793 4629 32796
rect 4663 32793 4675 32827
rect 4617 32787 4675 32793
rect 4893 32827 4951 32833
rect 4893 32793 4905 32827
rect 4939 32824 4951 32827
rect 7116 32824 7144 32852
rect 4939 32796 7144 32824
rect 4939 32793 4951 32796
rect 4893 32787 4951 32793
rect 9122 32784 9128 32836
rect 9180 32784 9186 32836
rect 9876 32824 9904 32855
rect 10318 32852 10324 32864
rect 10376 32852 10382 32904
rect 11514 32852 11520 32904
rect 11572 32892 11578 32904
rect 11808 32892 11836 32923
rect 12897 32895 12955 32901
rect 12897 32892 12909 32895
rect 11572 32864 11836 32892
rect 12319 32864 12909 32892
rect 11572 32852 11578 32864
rect 9950 32824 9956 32836
rect 9863 32796 9956 32824
rect 9950 32784 9956 32796
rect 10008 32824 10014 32836
rect 12319 32824 12347 32864
rect 12897 32861 12909 32864
rect 12943 32861 12955 32895
rect 12897 32855 12955 32861
rect 10008 32796 12347 32824
rect 10008 32784 10014 32796
rect 7650 32756 7656 32768
rect 3568 32728 4154 32756
rect 7611 32728 7656 32756
rect 3568 32716 3574 32728
rect 7650 32716 7656 32728
rect 7708 32716 7714 32768
rect 8018 32716 8024 32768
rect 8076 32756 8082 32768
rect 8619 32759 8677 32765
rect 8619 32756 8631 32759
rect 8076 32728 8631 32756
rect 8076 32716 8082 32728
rect 8619 32725 8631 32728
rect 8665 32725 8677 32759
rect 8619 32719 8677 32725
rect 9033 32759 9091 32765
rect 9033 32725 9045 32759
rect 9079 32756 9091 32759
rect 9140 32756 9168 32784
rect 9306 32756 9312 32768
rect 9079 32728 9312 32756
rect 9079 32725 9091 32728
rect 9033 32719 9091 32725
rect 9306 32716 9312 32728
rect 9364 32716 9370 32768
rect 11241 32759 11299 32765
rect 11241 32725 11253 32759
rect 11287 32756 11299 32759
rect 11514 32756 11520 32768
rect 11287 32728 11520 32756
rect 11287 32725 11299 32728
rect 11241 32719 11299 32725
rect 11514 32716 11520 32728
rect 11572 32716 11578 32768
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 2866 32552 2872 32564
rect 2827 32524 2872 32552
rect 2866 32512 2872 32524
rect 2924 32512 2930 32564
rect 9950 32552 9956 32564
rect 9911 32524 9956 32552
rect 9950 32512 9956 32524
rect 10008 32512 10014 32564
rect 11606 32552 11612 32564
rect 11567 32524 11612 32552
rect 11606 32512 11612 32524
rect 11664 32512 11670 32564
rect 12158 32552 12164 32564
rect 12119 32524 12164 32552
rect 12158 32512 12164 32524
rect 12216 32512 12222 32564
rect 6638 32444 6644 32496
rect 6696 32484 6702 32496
rect 8113 32487 8171 32493
rect 8113 32484 8125 32487
rect 6696 32456 8125 32484
rect 6696 32444 6702 32456
rect 8113 32453 8125 32456
rect 8159 32453 8171 32487
rect 8113 32447 8171 32453
rect 7834 32416 7840 32428
rect 7795 32388 7840 32416
rect 7834 32376 7840 32388
rect 7892 32376 7898 32428
rect 3881 32351 3939 32357
rect 3881 32317 3893 32351
rect 3927 32348 3939 32351
rect 4341 32351 4399 32357
rect 4341 32348 4353 32351
rect 3927 32320 4353 32348
rect 3927 32317 3939 32320
rect 3881 32311 3939 32317
rect 4341 32317 4353 32320
rect 4387 32348 4399 32351
rect 4798 32348 4804 32360
rect 4387 32320 4804 32348
rect 4387 32317 4399 32320
rect 4341 32311 4399 32317
rect 4798 32308 4804 32320
rect 4856 32308 4862 32360
rect 6273 32283 6331 32289
rect 6273 32249 6285 32283
rect 6319 32280 6331 32283
rect 7190 32280 7196 32292
rect 6319 32252 7097 32280
rect 7151 32252 7196 32280
rect 6319 32249 6331 32252
rect 6273 32243 6331 32249
rect 2501 32215 2559 32221
rect 2501 32181 2513 32215
rect 2547 32212 2559 32215
rect 2682 32212 2688 32224
rect 2547 32184 2688 32212
rect 2547 32181 2559 32184
rect 2501 32175 2559 32181
rect 2682 32172 2688 32184
rect 2740 32212 2746 32224
rect 3234 32212 3240 32224
rect 2740 32184 3240 32212
rect 2740 32172 2746 32184
rect 3234 32172 3240 32184
rect 3292 32172 3298 32224
rect 4249 32215 4307 32221
rect 4249 32181 4261 32215
rect 4295 32212 4307 32215
rect 4706 32212 4712 32224
rect 4295 32184 4712 32212
rect 4295 32181 4307 32184
rect 4249 32175 4307 32181
rect 4706 32172 4712 32184
rect 4764 32172 4770 32224
rect 5258 32212 5264 32224
rect 5219 32184 5264 32212
rect 5258 32172 5264 32184
rect 5316 32172 5322 32224
rect 5902 32212 5908 32224
rect 5863 32184 5908 32212
rect 5902 32172 5908 32184
rect 5960 32172 5966 32224
rect 6638 32212 6644 32224
rect 6599 32184 6644 32212
rect 6638 32172 6644 32184
rect 6696 32172 6702 32224
rect 7069 32212 7097 32252
rect 7190 32240 7196 32252
rect 7248 32240 7254 32292
rect 7285 32283 7343 32289
rect 7285 32249 7297 32283
rect 7331 32280 7343 32283
rect 7650 32280 7656 32292
rect 7331 32252 7656 32280
rect 7331 32249 7343 32252
rect 7285 32243 7343 32249
rect 7300 32212 7328 32243
rect 7650 32240 7656 32252
rect 7708 32240 7714 32292
rect 8128 32280 8156 32447
rect 8754 32444 8760 32496
rect 8812 32484 8818 32496
rect 8812 32456 12347 32484
rect 8812 32444 8818 32456
rect 8665 32419 8723 32425
rect 8665 32385 8677 32419
rect 8711 32416 8723 32419
rect 8938 32416 8944 32428
rect 8711 32388 8944 32416
rect 8711 32385 8723 32388
rect 8665 32379 8723 32385
rect 8938 32376 8944 32388
rect 8996 32416 9002 32428
rect 11422 32416 11428 32428
rect 8996 32388 11428 32416
rect 8996 32376 9002 32388
rect 11422 32376 11428 32388
rect 11480 32376 11486 32428
rect 12319 32416 12347 32456
rect 12989 32419 13047 32425
rect 12989 32416 13001 32419
rect 12319 32388 13001 32416
rect 12989 32385 13001 32388
rect 13035 32385 13047 32419
rect 12989 32379 13047 32385
rect 9585 32351 9643 32357
rect 9585 32317 9597 32351
rect 9631 32348 9643 32351
rect 9858 32348 9864 32360
rect 9631 32320 9864 32348
rect 9631 32317 9643 32320
rect 9585 32311 9643 32317
rect 9858 32308 9864 32320
rect 9916 32308 9922 32360
rect 10410 32348 10416 32360
rect 10371 32320 10416 32348
rect 10410 32308 10416 32320
rect 10468 32308 10474 32360
rect 12158 32308 12164 32360
rect 12216 32348 12222 32360
rect 12437 32351 12495 32357
rect 12437 32348 12449 32351
rect 12216 32320 12449 32348
rect 12216 32308 12222 32320
rect 12437 32317 12449 32320
rect 12483 32317 12495 32351
rect 12894 32348 12900 32360
rect 12855 32320 12900 32348
rect 12437 32311 12495 32317
rect 12894 32308 12900 32320
rect 12952 32308 12958 32360
rect 8986 32283 9044 32289
rect 8986 32280 8998 32283
rect 8128 32252 8998 32280
rect 8986 32249 8998 32252
rect 9032 32280 9044 32283
rect 9306 32280 9312 32292
rect 9032 32252 9312 32280
rect 9032 32249 9044 32252
rect 8986 32243 9044 32249
rect 9306 32240 9312 32252
rect 9364 32280 9370 32292
rect 10229 32283 10287 32289
rect 10229 32280 10241 32283
rect 9364 32252 10241 32280
rect 9364 32240 9370 32252
rect 10229 32249 10241 32252
rect 10275 32280 10287 32283
rect 10734 32283 10792 32289
rect 10734 32280 10746 32283
rect 10275 32252 10746 32280
rect 10275 32249 10287 32252
rect 10229 32243 10287 32249
rect 10734 32249 10746 32252
rect 10780 32249 10792 32283
rect 10734 32243 10792 32249
rect 7069 32184 7328 32212
rect 8573 32215 8631 32221
rect 8573 32181 8585 32215
rect 8619 32212 8631 32215
rect 8662 32212 8668 32224
rect 8619 32184 8668 32212
rect 8619 32181 8631 32184
rect 8573 32175 8631 32181
rect 8662 32172 8668 32184
rect 8720 32172 8726 32224
rect 10502 32172 10508 32224
rect 10560 32212 10566 32224
rect 11333 32215 11391 32221
rect 11333 32212 11345 32215
rect 10560 32184 11345 32212
rect 10560 32172 10566 32184
rect 11333 32181 11345 32184
rect 11379 32181 11391 32215
rect 11333 32175 11391 32181
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 2774 32008 2780 32020
rect 2735 31980 2780 32008
rect 2774 31968 2780 31980
rect 2832 31968 2838 32020
rect 5258 31968 5264 32020
rect 5316 32008 5322 32020
rect 5445 32011 5503 32017
rect 5445 32008 5457 32011
rect 5316 31980 5457 32008
rect 5316 31968 5322 31980
rect 5445 31977 5457 31980
rect 5491 31977 5503 32011
rect 5445 31971 5503 31977
rect 5534 31968 5540 32020
rect 5592 32008 5598 32020
rect 5813 32011 5871 32017
rect 5813 32008 5825 32011
rect 5592 31980 5825 32008
rect 5592 31968 5598 31980
rect 5813 31977 5825 31980
rect 5859 31977 5871 32011
rect 8938 32008 8944 32020
rect 8899 31980 8944 32008
rect 5813 31971 5871 31977
rect 8938 31968 8944 31980
rect 8996 31968 9002 32020
rect 9490 32008 9496 32020
rect 9451 31980 9496 32008
rect 9490 31968 9496 31980
rect 9548 31968 9554 32020
rect 10410 31968 10416 32020
rect 10468 32008 10474 32020
rect 10689 32011 10747 32017
rect 10689 32008 10701 32011
rect 10468 31980 10701 32008
rect 10468 31968 10474 31980
rect 10689 31977 10701 31980
rect 10735 32008 10747 32011
rect 11333 32011 11391 32017
rect 11333 32008 11345 32011
rect 10735 31980 11345 32008
rect 10735 31977 10747 31980
rect 10689 31971 10747 31977
rect 11333 31977 11345 31980
rect 11379 31977 11391 32011
rect 11333 31971 11391 31977
rect 4611 31943 4669 31949
rect 4611 31909 4623 31943
rect 4657 31940 4669 31943
rect 4706 31940 4712 31952
rect 4657 31912 4712 31940
rect 4657 31909 4669 31912
rect 4611 31903 4669 31909
rect 4706 31900 4712 31912
rect 4764 31900 4770 31952
rect 7006 31940 7012 31952
rect 6967 31912 7012 31940
rect 7006 31900 7012 31912
rect 7064 31900 7070 31952
rect 9582 31900 9588 31952
rect 9640 31940 9646 31952
rect 9861 31943 9919 31949
rect 9861 31940 9873 31943
rect 9640 31912 9873 31940
rect 9640 31900 9646 31912
rect 9861 31909 9873 31912
rect 9907 31940 9919 31943
rect 10502 31940 10508 31952
rect 9907 31912 10508 31940
rect 9907 31909 9919 31912
rect 9861 31903 9919 31909
rect 10502 31900 10508 31912
rect 10560 31900 10566 31952
rect 2590 31872 2596 31884
rect 2551 31844 2596 31872
rect 2590 31832 2596 31844
rect 2648 31832 2654 31884
rect 8386 31872 8392 31884
rect 8347 31844 8392 31872
rect 8386 31832 8392 31844
rect 8444 31832 8450 31884
rect 11514 31872 11520 31884
rect 11475 31844 11520 31872
rect 11514 31832 11520 31844
rect 11572 31832 11578 31884
rect 11698 31872 11704 31884
rect 11659 31844 11704 31872
rect 11698 31832 11704 31844
rect 11756 31872 11762 31884
rect 12437 31875 12495 31881
rect 12437 31872 12449 31875
rect 11756 31844 12449 31872
rect 11756 31832 11762 31844
rect 12437 31841 12449 31844
rect 12483 31872 12495 31875
rect 12894 31872 12900 31884
rect 12483 31844 12900 31872
rect 12483 31841 12495 31844
rect 12437 31835 12495 31841
rect 12894 31832 12900 31844
rect 12952 31832 12958 31884
rect 4246 31804 4252 31816
rect 4207 31776 4252 31804
rect 4246 31764 4252 31776
rect 4304 31764 4310 31816
rect 6917 31807 6975 31813
rect 6917 31773 6929 31807
rect 6963 31804 6975 31807
rect 8018 31804 8024 31816
rect 6963 31776 8024 31804
rect 6963 31773 6975 31776
rect 6917 31767 6975 31773
rect 8018 31764 8024 31776
rect 8076 31764 8082 31816
rect 9398 31764 9404 31816
rect 9456 31804 9462 31816
rect 9769 31807 9827 31813
rect 9769 31804 9781 31807
rect 9456 31776 9781 31804
rect 9456 31764 9462 31776
rect 9769 31773 9781 31776
rect 9815 31773 9827 31807
rect 9769 31767 9827 31773
rect 7190 31696 7196 31748
rect 7248 31736 7254 31748
rect 7469 31739 7527 31745
rect 7469 31736 7481 31739
rect 7248 31708 7481 31736
rect 7248 31696 7254 31708
rect 7469 31705 7481 31708
rect 7515 31736 7527 31739
rect 10318 31736 10324 31748
rect 7515 31708 7880 31736
rect 10279 31708 10324 31736
rect 7515 31705 7527 31708
rect 7469 31699 7527 31705
rect 7852 31680 7880 31708
rect 10318 31696 10324 31708
rect 10376 31696 10382 31748
rect 5166 31668 5172 31680
rect 5127 31640 5172 31668
rect 5166 31628 5172 31640
rect 5224 31628 5230 31680
rect 7834 31668 7840 31680
rect 7795 31640 7840 31668
rect 7834 31628 7840 31640
rect 7892 31628 7898 31680
rect 7926 31628 7932 31680
rect 7984 31668 7990 31680
rect 8527 31671 8585 31677
rect 8527 31668 8539 31671
rect 7984 31640 8539 31668
rect 7984 31628 7990 31640
rect 8527 31637 8539 31640
rect 8573 31637 8585 31671
rect 8527 31631 8585 31637
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 2590 31464 2596 31476
rect 2551 31436 2596 31464
rect 2590 31424 2596 31436
rect 2648 31424 2654 31476
rect 4525 31467 4583 31473
rect 4525 31433 4537 31467
rect 4571 31464 4583 31467
rect 4706 31464 4712 31476
rect 4571 31436 4712 31464
rect 4571 31433 4583 31436
rect 4525 31427 4583 31433
rect 4706 31424 4712 31436
rect 4764 31424 4770 31476
rect 6641 31467 6699 31473
rect 6641 31433 6653 31467
rect 6687 31464 6699 31467
rect 7006 31464 7012 31476
rect 6687 31436 7012 31464
rect 6687 31433 6699 31436
rect 6641 31427 6699 31433
rect 7006 31424 7012 31436
rect 7064 31424 7070 31476
rect 7929 31467 7987 31473
rect 7929 31433 7941 31467
rect 7975 31464 7987 31467
rect 8018 31464 8024 31476
rect 7975 31436 8024 31464
rect 7975 31433 7987 31436
rect 7929 31427 7987 31433
rect 8018 31424 8024 31436
rect 8076 31424 8082 31476
rect 8478 31424 8484 31476
rect 8536 31464 8542 31476
rect 9033 31467 9091 31473
rect 9033 31464 9045 31467
rect 8536 31436 9045 31464
rect 8536 31424 8542 31436
rect 9033 31433 9045 31436
rect 9079 31433 9091 31467
rect 9582 31464 9588 31476
rect 9543 31436 9588 31464
rect 9033 31427 9091 31433
rect 9582 31424 9588 31436
rect 9640 31424 9646 31476
rect 11514 31464 11520 31476
rect 9692 31436 11520 31464
rect 5626 31396 5632 31408
rect 5587 31368 5632 31396
rect 5626 31356 5632 31368
rect 5684 31356 5690 31408
rect 6730 31356 6736 31408
rect 6788 31396 6794 31408
rect 9692 31396 9720 31436
rect 11514 31424 11520 31436
rect 11572 31464 11578 31476
rect 11609 31467 11667 31473
rect 11609 31464 11621 31467
rect 11572 31436 11621 31464
rect 11572 31424 11578 31436
rect 11609 31433 11621 31436
rect 11655 31433 11667 31467
rect 11609 31427 11667 31433
rect 10318 31396 10324 31408
rect 6788 31368 9720 31396
rect 10279 31368 10324 31396
rect 6788 31356 6794 31368
rect 10318 31356 10324 31368
rect 10376 31356 10382 31408
rect 4157 31331 4215 31337
rect 4157 31297 4169 31331
rect 4203 31328 4215 31331
rect 4246 31328 4252 31340
rect 4203 31300 4252 31328
rect 4203 31297 4215 31300
rect 4157 31291 4215 31297
rect 4246 31288 4252 31300
rect 4304 31328 4310 31340
rect 4801 31331 4859 31337
rect 4801 31328 4813 31331
rect 4304 31300 4813 31328
rect 4304 31288 4310 31300
rect 4801 31297 4813 31300
rect 4847 31297 4859 31331
rect 4801 31291 4859 31297
rect 5166 31288 5172 31340
rect 5224 31328 5230 31340
rect 6181 31331 6239 31337
rect 6181 31328 6193 31331
rect 5224 31300 6193 31328
rect 5224 31288 5230 31300
rect 6181 31297 6193 31300
rect 6227 31297 6239 31331
rect 6181 31291 6239 31297
rect 6917 31331 6975 31337
rect 6917 31297 6929 31331
rect 6963 31328 6975 31331
rect 7926 31328 7932 31340
rect 6963 31300 7932 31328
rect 6963 31297 6975 31300
rect 6917 31291 6975 31297
rect 3421 31263 3479 31269
rect 3421 31229 3433 31263
rect 3467 31229 3479 31263
rect 3421 31223 3479 31229
rect 3234 31124 3240 31136
rect 3195 31096 3240 31124
rect 3234 31084 3240 31096
rect 3292 31124 3298 31136
rect 3436 31124 3464 31223
rect 3510 31220 3516 31272
rect 3568 31260 3574 31272
rect 3881 31263 3939 31269
rect 3881 31260 3893 31263
rect 3568 31232 3893 31260
rect 3568 31220 3574 31232
rect 3881 31229 3893 31232
rect 3927 31229 3939 31263
rect 3881 31223 3939 31229
rect 5077 31195 5135 31201
rect 5077 31161 5089 31195
rect 5123 31161 5135 31195
rect 5077 31155 5135 31161
rect 5169 31195 5227 31201
rect 5169 31161 5181 31195
rect 5215 31192 5227 31195
rect 5258 31192 5264 31204
rect 5215 31164 5264 31192
rect 5215 31161 5227 31164
rect 5169 31155 5227 31161
rect 3292 31096 3464 31124
rect 3292 31084 3298 31096
rect 4430 31084 4436 31136
rect 4488 31124 4494 31136
rect 5092 31124 5120 31155
rect 5258 31152 5264 31164
rect 5316 31152 5322 31204
rect 6196 31192 6224 31291
rect 7926 31288 7932 31300
rect 7984 31288 7990 31340
rect 8478 31220 8484 31272
rect 8536 31260 8542 31272
rect 8608 31263 8666 31269
rect 8608 31260 8620 31263
rect 8536 31232 8620 31260
rect 8536 31220 8542 31232
rect 8608 31229 8620 31232
rect 8654 31229 8666 31263
rect 8608 31223 8666 31229
rect 7009 31195 7067 31201
rect 7009 31192 7021 31195
rect 6196 31164 7021 31192
rect 7009 31161 7021 31164
rect 7055 31161 7067 31195
rect 7561 31195 7619 31201
rect 7561 31192 7573 31195
rect 7009 31155 7067 31161
rect 7202 31164 7573 31192
rect 5626 31124 5632 31136
rect 4488 31096 5632 31124
rect 4488 31084 4494 31096
rect 5626 31084 5632 31096
rect 5684 31124 5690 31136
rect 7202 31124 7230 31164
rect 7561 31161 7573 31164
rect 7607 31161 7619 31195
rect 7561 31155 7619 31161
rect 9122 31152 9128 31204
rect 9180 31192 9186 31204
rect 9766 31192 9772 31204
rect 9180 31164 9772 31192
rect 9180 31152 9186 31164
rect 9766 31152 9772 31164
rect 9824 31152 9830 31204
rect 9858 31152 9864 31204
rect 9916 31192 9922 31204
rect 10689 31195 10747 31201
rect 10689 31192 10701 31195
rect 9916 31164 10701 31192
rect 9916 31152 9922 31164
rect 10689 31161 10701 31164
rect 10735 31161 10747 31195
rect 11698 31192 11704 31204
rect 10689 31155 10747 31161
rect 11256 31164 11704 31192
rect 8386 31124 8392 31136
rect 5684 31096 7230 31124
rect 8347 31096 8392 31124
rect 5684 31084 5690 31096
rect 8386 31084 8392 31096
rect 8444 31084 8450 31136
rect 8711 31127 8769 31133
rect 8711 31093 8723 31127
rect 8757 31124 8769 31127
rect 8938 31124 8944 31136
rect 8757 31096 8944 31124
rect 8757 31093 8769 31096
rect 8711 31087 8769 31093
rect 8938 31084 8944 31096
rect 8996 31084 9002 31136
rect 9306 31084 9312 31136
rect 9364 31124 9370 31136
rect 11256 31133 11284 31164
rect 11698 31152 11704 31164
rect 11756 31152 11762 31204
rect 11241 31127 11299 31133
rect 11241 31124 11253 31127
rect 9364 31096 11253 31124
rect 9364 31084 9370 31096
rect 11241 31093 11253 31096
rect 11287 31093 11299 31127
rect 11241 31087 11299 31093
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 2958 30880 2964 30932
rect 3016 30920 3022 30932
rect 3510 30920 3516 30932
rect 3016 30892 3516 30920
rect 3016 30880 3022 30892
rect 3510 30880 3516 30892
rect 3568 30880 3574 30932
rect 4062 30880 4068 30932
rect 4120 30920 4126 30932
rect 4430 30920 4436 30932
rect 4120 30892 4436 30920
rect 4120 30880 4126 30892
rect 4430 30880 4436 30892
rect 4488 30880 4494 30932
rect 5902 30880 5908 30932
rect 5960 30920 5966 30932
rect 6549 30923 6607 30929
rect 6549 30920 6561 30923
rect 5960 30892 6561 30920
rect 5960 30880 5966 30892
rect 6549 30889 6561 30892
rect 6595 30889 6607 30923
rect 6549 30883 6607 30889
rect 7561 30923 7619 30929
rect 7561 30889 7573 30923
rect 7607 30920 7619 30923
rect 7926 30920 7932 30932
rect 7607 30892 7932 30920
rect 7607 30889 7619 30892
rect 7561 30883 7619 30889
rect 7926 30880 7932 30892
rect 7984 30880 7990 30932
rect 8220 30892 9904 30920
rect 8220 30864 8248 30892
rect 4338 30812 4344 30864
rect 4396 30852 4402 30864
rect 5077 30855 5135 30861
rect 5077 30852 5089 30855
rect 4396 30824 5089 30852
rect 4396 30812 4402 30824
rect 5077 30821 5089 30824
rect 5123 30852 5135 30855
rect 5166 30852 5172 30864
rect 5123 30824 5172 30852
rect 5123 30821 5135 30824
rect 5077 30815 5135 30821
rect 5166 30812 5172 30824
rect 5224 30812 5230 30864
rect 8202 30852 8208 30864
rect 8163 30824 8208 30852
rect 8202 30812 8208 30824
rect 8260 30812 8266 30864
rect 8938 30812 8944 30864
rect 8996 30852 9002 30864
rect 9490 30852 9496 30864
rect 8996 30824 9496 30852
rect 8996 30812 9002 30824
rect 9490 30812 9496 30824
rect 9548 30852 9554 30864
rect 9876 30861 9904 30892
rect 9769 30855 9827 30861
rect 9769 30852 9781 30855
rect 9548 30824 9781 30852
rect 9548 30812 9554 30824
rect 9769 30821 9781 30824
rect 9815 30821 9827 30855
rect 9769 30815 9827 30821
rect 9861 30855 9919 30861
rect 9861 30821 9873 30855
rect 9907 30852 9919 30855
rect 10502 30852 10508 30864
rect 9907 30824 10508 30852
rect 9907 30821 9919 30824
rect 9861 30815 9919 30821
rect 10502 30812 10508 30824
rect 10560 30812 10566 30864
rect 6730 30784 6736 30796
rect 6691 30756 6736 30784
rect 6730 30744 6736 30756
rect 6788 30744 6794 30796
rect 7009 30787 7067 30793
rect 7009 30753 7021 30787
rect 7055 30784 7067 30787
rect 7098 30784 7104 30796
rect 7055 30756 7104 30784
rect 7055 30753 7067 30756
rect 7009 30747 7067 30753
rect 7098 30744 7104 30756
rect 7156 30744 7162 30796
rect 9122 30784 9128 30796
rect 9083 30756 9128 30784
rect 9122 30744 9128 30756
rect 9180 30744 9186 30796
rect 10962 30744 10968 30796
rect 11020 30784 11026 30796
rect 11276 30787 11334 30793
rect 11276 30784 11288 30787
rect 11020 30756 11288 30784
rect 11020 30744 11026 30756
rect 11276 30753 11288 30756
rect 11322 30753 11334 30787
rect 11276 30747 11334 30753
rect 4801 30719 4859 30725
rect 4801 30716 4813 30719
rect 4126 30688 4813 30716
rect 3142 30608 3148 30660
rect 3200 30648 3206 30660
rect 4126 30648 4154 30688
rect 4801 30685 4813 30688
rect 4847 30716 4859 30719
rect 4985 30719 5043 30725
rect 4985 30716 4997 30719
rect 4847 30688 4997 30716
rect 4847 30685 4859 30688
rect 4801 30679 4859 30685
rect 4985 30685 4997 30688
rect 5031 30685 5043 30719
rect 4985 30679 5043 30685
rect 8113 30719 8171 30725
rect 8113 30685 8125 30719
rect 8159 30716 8171 30719
rect 8159 30688 9628 30716
rect 8159 30685 8171 30688
rect 8113 30679 8171 30685
rect 5534 30648 5540 30660
rect 3200 30620 4154 30648
rect 5495 30620 5540 30648
rect 3200 30608 3206 30620
rect 5534 30608 5540 30620
rect 5592 30608 5598 30660
rect 8665 30651 8723 30657
rect 8665 30617 8677 30651
rect 8711 30617 8723 30651
rect 8665 30611 8723 30617
rect 8680 30580 8708 30611
rect 9600 30592 9628 30688
rect 9766 30676 9772 30728
rect 9824 30716 9830 30728
rect 10045 30719 10103 30725
rect 10045 30716 10057 30719
rect 9824 30688 10057 30716
rect 9824 30676 9830 30688
rect 10045 30685 10057 30688
rect 10091 30716 10103 30719
rect 10410 30716 10416 30728
rect 10091 30688 10416 30716
rect 10091 30685 10103 30688
rect 10045 30679 10103 30685
rect 10410 30676 10416 30688
rect 10468 30676 10474 30728
rect 9398 30580 9404 30592
rect 8680 30552 9404 30580
rect 9398 30540 9404 30552
rect 9456 30540 9462 30592
rect 9582 30540 9588 30592
rect 9640 30580 9646 30592
rect 11379 30583 11437 30589
rect 11379 30580 11391 30583
rect 9640 30552 11391 30580
rect 9640 30540 9646 30552
rect 11379 30549 11391 30552
rect 11425 30549 11437 30583
rect 11379 30543 11437 30549
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 4338 30376 4344 30388
rect 4299 30348 4344 30376
rect 4338 30336 4344 30348
rect 4396 30336 4402 30388
rect 6549 30379 6607 30385
rect 6549 30345 6561 30379
rect 6595 30376 6607 30379
rect 7098 30376 7104 30388
rect 6595 30348 7104 30376
rect 6595 30345 6607 30348
rect 6549 30339 6607 30345
rect 4709 30243 4767 30249
rect 4709 30209 4721 30243
rect 4755 30240 4767 30243
rect 6086 30240 6092 30252
rect 4755 30212 6092 30240
rect 4755 30209 4767 30212
rect 4709 30203 4767 30209
rect 5736 30181 5764 30212
rect 6086 30200 6092 30212
rect 6144 30240 6150 30252
rect 6564 30240 6592 30339
rect 7098 30336 7104 30348
rect 7156 30336 7162 30388
rect 9490 30376 9496 30388
rect 9451 30348 9496 30376
rect 9490 30336 9496 30348
rect 9548 30336 9554 30388
rect 10502 30376 10508 30388
rect 10463 30348 10508 30376
rect 10502 30336 10508 30348
rect 10560 30336 10566 30388
rect 10962 30336 10968 30388
rect 11020 30376 11026 30388
rect 11241 30379 11299 30385
rect 11241 30376 11253 30379
rect 11020 30348 11253 30376
rect 11020 30336 11026 30348
rect 11241 30345 11253 30348
rect 11287 30345 11299 30379
rect 11241 30339 11299 30345
rect 9217 30311 9275 30317
rect 9217 30277 9229 30311
rect 9263 30308 9275 30311
rect 9582 30308 9588 30320
rect 9263 30280 9588 30308
rect 9263 30277 9275 30280
rect 9217 30271 9275 30277
rect 9582 30268 9588 30280
rect 9640 30268 9646 30320
rect 6144 30212 6592 30240
rect 6144 30200 6150 30212
rect 7374 30200 7380 30252
rect 7432 30240 7438 30252
rect 8662 30240 8668 30252
rect 7432 30212 8668 30240
rect 7432 30200 7438 30212
rect 8662 30200 8668 30212
rect 8720 30240 8726 30252
rect 8720 30212 9213 30240
rect 8720 30200 8726 30212
rect 5169 30175 5227 30181
rect 5169 30172 5181 30175
rect 5000 30144 5181 30172
rect 5000 30048 5028 30144
rect 5169 30141 5181 30144
rect 5215 30141 5227 30175
rect 5169 30135 5227 30141
rect 5721 30175 5779 30181
rect 5721 30141 5733 30175
rect 5767 30141 5779 30175
rect 5721 30135 5779 30141
rect 6178 30132 6184 30184
rect 6236 30172 6242 30184
rect 6860 30175 6918 30181
rect 6860 30172 6872 30175
rect 6236 30144 6872 30172
rect 6236 30132 6242 30144
rect 6860 30141 6872 30144
rect 6906 30172 6918 30175
rect 7285 30175 7343 30181
rect 7285 30172 7297 30175
rect 6906 30144 7297 30172
rect 6906 30141 6918 30144
rect 6860 30135 6918 30141
rect 7285 30141 7297 30144
rect 7331 30141 7343 30175
rect 7285 30135 7343 30141
rect 7929 30175 7987 30181
rect 7929 30141 7941 30175
rect 7975 30172 7987 30175
rect 8478 30172 8484 30184
rect 7975 30144 8484 30172
rect 7975 30141 7987 30144
rect 7929 30135 7987 30141
rect 8478 30132 8484 30144
rect 8536 30132 8542 30184
rect 9185 30172 9213 30212
rect 9712 30175 9770 30181
rect 9712 30172 9724 30175
rect 9185 30144 9724 30172
rect 9712 30141 9724 30144
rect 9758 30172 9770 30175
rect 10137 30175 10195 30181
rect 10137 30172 10149 30175
rect 9758 30144 10149 30172
rect 9758 30141 9770 30144
rect 9712 30135 9770 30141
rect 10137 30141 10149 30144
rect 10183 30141 10195 30175
rect 10137 30135 10195 30141
rect 5902 30104 5908 30116
rect 5863 30076 5908 30104
rect 5902 30064 5908 30076
rect 5960 30064 5966 30116
rect 8250 30107 8308 30113
rect 8250 30104 8262 30107
rect 7760 30076 8262 30104
rect 3326 29996 3332 30048
rect 3384 30036 3390 30048
rect 3970 30036 3976 30048
rect 3384 30008 3976 30036
rect 3384 29996 3390 30008
rect 3970 29996 3976 30008
rect 4028 29996 4034 30048
rect 4982 30036 4988 30048
rect 4943 30008 4988 30036
rect 4982 29996 4988 30008
rect 5040 29996 5046 30048
rect 6963 30039 7021 30045
rect 6963 30005 6975 30039
rect 7009 30036 7021 30039
rect 7190 30036 7196 30048
rect 7009 30008 7196 30036
rect 7009 30005 7021 30008
rect 6963 29999 7021 30005
rect 7190 29996 7196 30008
rect 7248 29996 7254 30048
rect 7650 29996 7656 30048
rect 7708 30036 7714 30048
rect 7760 30045 7788 30076
rect 8250 30073 8262 30076
rect 8296 30073 8308 30107
rect 8250 30067 8308 30073
rect 7745 30039 7803 30045
rect 7745 30036 7757 30039
rect 7708 30008 7757 30036
rect 7708 29996 7714 30008
rect 7745 30005 7757 30008
rect 7791 30005 7803 30039
rect 8846 30036 8852 30048
rect 8807 30008 8852 30036
rect 7745 29999 7803 30005
rect 8846 29996 8852 30008
rect 8904 29996 8910 30048
rect 9815 30039 9873 30045
rect 9815 30005 9827 30039
rect 9861 30036 9873 30039
rect 10042 30036 10048 30048
rect 9861 30008 10048 30036
rect 9861 30005 9873 30008
rect 9815 29999 9873 30005
rect 10042 29996 10048 30008
rect 10100 29996 10106 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 1578 29832 1584 29844
rect 1539 29804 1584 29832
rect 1578 29792 1584 29804
rect 1636 29792 1642 29844
rect 5902 29792 5908 29844
rect 5960 29832 5966 29844
rect 6822 29832 6828 29844
rect 5960 29804 6828 29832
rect 5960 29792 5966 29804
rect 6822 29792 6828 29804
rect 6880 29792 6886 29844
rect 8113 29835 8171 29841
rect 8113 29801 8125 29835
rect 8159 29832 8171 29835
rect 8202 29832 8208 29844
rect 8159 29804 8208 29832
rect 8159 29801 8171 29804
rect 8113 29795 8171 29801
rect 8202 29792 8208 29804
rect 8260 29832 8266 29844
rect 8846 29832 8852 29844
rect 8260 29804 8852 29832
rect 8260 29792 8266 29804
rect 8846 29792 8852 29804
rect 8904 29792 8910 29844
rect 12253 29835 12311 29841
rect 12253 29801 12265 29835
rect 12299 29832 12311 29835
rect 12434 29832 12440 29844
rect 12299 29804 12440 29832
rect 12299 29801 12311 29804
rect 12253 29795 12311 29801
rect 12434 29792 12440 29804
rect 12492 29792 12498 29844
rect 3970 29724 3976 29776
rect 4028 29764 4034 29776
rect 5077 29767 5135 29773
rect 5077 29764 5089 29767
rect 4028 29736 5089 29764
rect 4028 29724 4034 29736
rect 5077 29733 5089 29736
rect 5123 29733 5135 29767
rect 5626 29764 5632 29776
rect 5587 29736 5632 29764
rect 5077 29727 5135 29733
rect 5626 29724 5632 29736
rect 5684 29724 5690 29776
rect 6549 29767 6607 29773
rect 6549 29733 6561 29767
rect 6595 29764 6607 29767
rect 6730 29764 6736 29776
rect 6595 29736 6736 29764
rect 6595 29733 6607 29736
rect 6549 29727 6607 29733
rect 6730 29724 6736 29736
rect 6788 29724 6794 29776
rect 7098 29724 7104 29776
rect 7156 29764 7162 29776
rect 7193 29767 7251 29773
rect 7193 29764 7205 29767
rect 7156 29736 7205 29764
rect 7156 29724 7162 29736
rect 7193 29733 7205 29736
rect 7239 29733 7251 29767
rect 7193 29727 7251 29733
rect 7745 29767 7803 29773
rect 7745 29733 7757 29767
rect 7791 29764 7803 29767
rect 8754 29764 8760 29776
rect 7791 29736 8760 29764
rect 7791 29733 7803 29736
rect 7745 29727 7803 29733
rect 8754 29724 8760 29736
rect 8812 29724 8818 29776
rect 9858 29764 9864 29776
rect 9819 29736 9864 29764
rect 9858 29724 9864 29736
rect 9916 29724 9922 29776
rect 1394 29696 1400 29708
rect 1355 29668 1400 29696
rect 1394 29656 1400 29668
rect 1452 29656 1458 29708
rect 8202 29656 8208 29708
rect 8260 29696 8266 29708
rect 8386 29696 8392 29708
rect 8260 29668 8392 29696
rect 8260 29656 8266 29668
rect 8386 29656 8392 29668
rect 8444 29696 8450 29708
rect 8608 29699 8666 29705
rect 8608 29696 8620 29699
rect 8444 29668 8620 29696
rect 8444 29656 8450 29668
rect 8608 29665 8620 29668
rect 8654 29665 8666 29699
rect 12066 29696 12072 29708
rect 12027 29668 12072 29696
rect 8608 29659 8666 29665
rect 12066 29656 12072 29668
rect 12124 29656 12130 29708
rect 4985 29631 5043 29637
rect 4985 29628 4997 29631
rect 4724 29600 4997 29628
rect 3418 29452 3424 29504
rect 3476 29492 3482 29504
rect 4724 29501 4752 29600
rect 4985 29597 4997 29600
rect 5031 29597 5043 29631
rect 4985 29591 5043 29597
rect 7101 29631 7159 29637
rect 7101 29597 7113 29631
rect 7147 29628 7159 29631
rect 7466 29628 7472 29640
rect 7147 29600 7472 29628
rect 7147 29597 7159 29600
rect 7101 29591 7159 29597
rect 7466 29588 7472 29600
rect 7524 29628 7530 29640
rect 8711 29631 8769 29637
rect 8711 29628 8723 29631
rect 7524 29600 8723 29628
rect 7524 29588 7530 29600
rect 8711 29597 8723 29600
rect 8757 29597 8769 29631
rect 8711 29591 8769 29597
rect 9769 29631 9827 29637
rect 9769 29597 9781 29631
rect 9815 29628 9827 29631
rect 11146 29628 11152 29640
rect 9815 29600 11152 29628
rect 9815 29597 9827 29600
rect 9769 29591 9827 29597
rect 11146 29588 11152 29600
rect 11204 29588 11210 29640
rect 9398 29520 9404 29572
rect 9456 29560 9462 29572
rect 10318 29560 10324 29572
rect 9456 29532 10324 29560
rect 9456 29520 9462 29532
rect 10318 29520 10324 29532
rect 10376 29520 10382 29572
rect 4709 29495 4767 29501
rect 4709 29492 4721 29495
rect 3476 29464 4721 29492
rect 3476 29452 3482 29464
rect 4709 29461 4721 29464
rect 4755 29461 4767 29495
rect 8478 29492 8484 29504
rect 8439 29464 8484 29492
rect 4709 29455 4767 29461
rect 8478 29452 8484 29464
rect 8536 29452 8542 29504
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 3421 29291 3479 29297
rect 3421 29257 3433 29291
rect 3467 29288 3479 29291
rect 3697 29291 3755 29297
rect 3697 29288 3709 29291
rect 3467 29260 3709 29288
rect 3467 29257 3479 29260
rect 3421 29251 3479 29257
rect 3697 29257 3709 29260
rect 3743 29288 3755 29291
rect 4154 29288 4160 29300
rect 3743 29260 4160 29288
rect 3743 29257 3755 29260
rect 3697 29251 3755 29257
rect 4154 29248 4160 29260
rect 4212 29248 4218 29300
rect 9677 29291 9735 29297
rect 9677 29257 9689 29291
rect 9723 29288 9735 29291
rect 9858 29288 9864 29300
rect 9723 29260 9864 29288
rect 9723 29257 9735 29260
rect 9677 29251 9735 29257
rect 9858 29248 9864 29260
rect 9916 29248 9922 29300
rect 11146 29288 11152 29300
rect 11107 29260 11152 29288
rect 11146 29248 11152 29260
rect 11204 29248 11210 29300
rect 5813 29223 5871 29229
rect 5813 29189 5825 29223
rect 5859 29220 5871 29223
rect 7834 29220 7840 29232
rect 5859 29192 7840 29220
rect 5859 29189 5871 29192
rect 5813 29183 5871 29189
rect 7834 29180 7840 29192
rect 7892 29220 7898 29232
rect 8294 29220 8300 29232
rect 7892 29192 8300 29220
rect 7892 29180 7898 29192
rect 8294 29180 8300 29192
rect 8352 29180 8358 29232
rect 8754 29180 8760 29232
rect 8812 29220 8818 29232
rect 9217 29223 9275 29229
rect 9217 29220 9229 29223
rect 8812 29192 9229 29220
rect 8812 29180 8818 29192
rect 9217 29189 9229 29192
rect 9263 29189 9275 29223
rect 9217 29183 9275 29189
rect 2590 29112 2596 29164
rect 2648 29152 2654 29164
rect 3050 29152 3056 29164
rect 2648 29124 3056 29152
rect 2648 29112 2654 29124
rect 3050 29112 3056 29124
rect 3108 29152 3114 29164
rect 3108 29124 3832 29152
rect 3108 29112 3114 29124
rect 3212 29087 3270 29093
rect 3212 29053 3224 29087
rect 3258 29084 3270 29087
rect 3421 29087 3479 29093
rect 3421 29084 3433 29087
rect 3258 29056 3433 29084
rect 3258 29053 3270 29056
rect 3212 29047 3270 29053
rect 3421 29053 3433 29056
rect 3467 29053 3479 29087
rect 3804 29084 3832 29124
rect 3878 29112 3884 29164
rect 3936 29152 3942 29164
rect 4062 29152 4068 29164
rect 3936 29124 4068 29152
rect 3936 29112 3942 29124
rect 4062 29112 4068 29124
rect 4120 29112 4126 29164
rect 6822 29152 6828 29164
rect 6783 29124 6828 29152
rect 6822 29112 6828 29124
rect 6880 29112 6886 29164
rect 7190 29112 7196 29164
rect 7248 29152 7254 29164
rect 8665 29155 8723 29161
rect 8665 29152 8677 29155
rect 7248 29124 8677 29152
rect 7248 29112 7254 29124
rect 8665 29121 8677 29124
rect 8711 29152 8723 29155
rect 8938 29152 8944 29164
rect 8711 29124 8944 29152
rect 8711 29121 8723 29124
rect 8665 29115 8723 29121
rect 8938 29112 8944 29124
rect 8996 29112 9002 29164
rect 10042 29112 10048 29164
rect 10100 29152 10106 29164
rect 10229 29155 10287 29161
rect 10229 29152 10241 29155
rect 10100 29124 10241 29152
rect 10100 29112 10106 29124
rect 10229 29121 10241 29124
rect 10275 29121 10287 29155
rect 10229 29115 10287 29121
rect 10410 29112 10416 29164
rect 10468 29152 10474 29164
rect 10505 29155 10563 29161
rect 10505 29152 10517 29155
rect 10468 29124 10517 29152
rect 10468 29112 10474 29124
rect 10505 29121 10517 29124
rect 10551 29121 10563 29155
rect 10505 29115 10563 29121
rect 4224 29087 4282 29093
rect 4224 29084 4236 29087
rect 3804 29056 4236 29084
rect 3421 29047 3479 29053
rect 4224 29053 4236 29056
rect 4270 29084 4282 29087
rect 4617 29087 4675 29093
rect 4617 29084 4629 29087
rect 4270 29056 4629 29084
rect 4270 29053 4282 29056
rect 4224 29047 4282 29053
rect 4617 29053 4629 29056
rect 4663 29053 4675 29087
rect 7745 29087 7803 29093
rect 7745 29084 7757 29087
rect 4617 29047 4675 29053
rect 6104 29056 7757 29084
rect 4433 29019 4491 29025
rect 4433 28985 4445 29019
rect 4479 29016 4491 29019
rect 5258 29016 5264 29028
rect 4479 28988 5264 29016
rect 4479 28985 4491 28988
rect 4433 28979 4491 28985
rect 5258 28976 5264 28988
rect 5316 28976 5322 29028
rect 5353 29019 5411 29025
rect 5353 28985 5365 29019
rect 5399 28985 5411 29019
rect 5353 28979 5411 28985
rect 1394 28908 1400 28960
rect 1452 28948 1458 28960
rect 1581 28951 1639 28957
rect 1581 28948 1593 28951
rect 1452 28920 1593 28948
rect 1452 28908 1458 28920
rect 1581 28917 1593 28920
rect 1627 28917 1639 28951
rect 1581 28911 1639 28917
rect 3283 28951 3341 28957
rect 3283 28917 3295 28951
rect 3329 28948 3341 28951
rect 3510 28948 3516 28960
rect 3329 28920 3516 28948
rect 3329 28917 3341 28920
rect 3283 28911 3341 28917
rect 3510 28908 3516 28920
rect 3568 28908 3574 28960
rect 3970 28948 3976 28960
rect 3931 28920 3976 28948
rect 3970 28908 3976 28920
rect 4028 28908 4034 28960
rect 5077 28951 5135 28957
rect 5077 28917 5089 28951
rect 5123 28948 5135 28951
rect 5368 28948 5396 28979
rect 6104 28948 6132 29056
rect 7745 29053 7757 29056
rect 7791 29084 7803 29087
rect 8021 29087 8079 29093
rect 8021 29084 8033 29087
rect 7791 29056 8033 29084
rect 7791 29053 7803 29056
rect 7745 29047 7803 29053
rect 8021 29053 8033 29056
rect 8067 29053 8079 29087
rect 8021 29047 8079 29053
rect 6273 29019 6331 29025
rect 6273 28985 6285 29019
rect 6319 29016 6331 29019
rect 7006 29016 7012 29028
rect 6319 28988 7012 29016
rect 6319 28985 6331 28988
rect 6273 28979 6331 28985
rect 7006 28976 7012 28988
rect 7064 28976 7070 29028
rect 7146 29019 7204 29025
rect 7146 28985 7158 29019
rect 7192 29016 7204 29019
rect 7650 29016 7656 29028
rect 7192 28988 7656 29016
rect 7192 28985 7204 28988
rect 7146 28979 7204 28985
rect 6638 28948 6644 28960
rect 5123 28920 6132 28948
rect 6599 28920 6644 28948
rect 5123 28917 5135 28920
rect 5077 28911 5135 28917
rect 6638 28908 6644 28920
rect 6696 28948 6702 28960
rect 7161 28948 7189 28979
rect 7650 28976 7656 28988
rect 7708 28976 7714 29028
rect 8036 29016 8064 29047
rect 8757 29019 8815 29025
rect 8036 28988 8616 29016
rect 6696 28920 7189 28948
rect 6696 28908 6702 28920
rect 8202 28908 8208 28960
rect 8260 28948 8266 28960
rect 8389 28951 8447 28957
rect 8389 28948 8401 28951
rect 8260 28920 8401 28948
rect 8260 28908 8266 28920
rect 8389 28917 8401 28920
rect 8435 28917 8447 28951
rect 8588 28948 8616 28988
rect 8757 28985 8769 29019
rect 8803 28985 8815 29019
rect 8757 28979 8815 28985
rect 10321 29019 10379 29025
rect 10321 28985 10333 29019
rect 10367 28985 10379 29019
rect 10321 28979 10379 28985
rect 8772 28948 8800 28979
rect 9950 28948 9956 28960
rect 8588 28920 8800 28948
rect 9911 28920 9956 28948
rect 8389 28911 8447 28917
rect 9950 28908 9956 28920
rect 10008 28948 10014 28960
rect 10336 28948 10364 28979
rect 10008 28920 10364 28948
rect 10008 28908 10014 28920
rect 12066 28908 12072 28960
rect 12124 28948 12130 28960
rect 12161 28951 12219 28957
rect 12161 28948 12173 28951
rect 12124 28920 12173 28948
rect 12124 28908 12130 28920
rect 12161 28917 12173 28920
rect 12207 28948 12219 28951
rect 12618 28948 12624 28960
rect 12207 28920 12624 28948
rect 12207 28917 12219 28920
rect 12161 28911 12219 28917
rect 12618 28908 12624 28920
rect 12676 28908 12682 28960
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 3142 28744 3148 28756
rect 3103 28716 3148 28744
rect 3142 28704 3148 28716
rect 3200 28704 3206 28756
rect 5258 28704 5264 28756
rect 5316 28744 5322 28756
rect 5629 28747 5687 28753
rect 5629 28744 5641 28747
rect 5316 28716 5641 28744
rect 5316 28704 5322 28716
rect 5629 28713 5641 28716
rect 5675 28713 5687 28747
rect 5629 28707 5687 28713
rect 6549 28747 6607 28753
rect 6549 28713 6561 28747
rect 6595 28744 6607 28747
rect 6638 28744 6644 28756
rect 6595 28716 6644 28744
rect 6595 28713 6607 28716
rect 6549 28707 6607 28713
rect 6638 28704 6644 28716
rect 6696 28704 6702 28756
rect 7006 28704 7012 28756
rect 7064 28744 7070 28756
rect 7101 28747 7159 28753
rect 7101 28744 7113 28747
rect 7064 28716 7113 28744
rect 7064 28704 7070 28716
rect 7101 28713 7113 28716
rect 7147 28713 7159 28747
rect 7466 28744 7472 28756
rect 7427 28716 7472 28744
rect 7101 28707 7159 28713
rect 4801 28679 4859 28685
rect 4801 28645 4813 28679
rect 4847 28676 4859 28679
rect 5074 28676 5080 28688
rect 4847 28648 5080 28676
rect 4847 28645 4859 28648
rect 4801 28639 4859 28645
rect 5074 28636 5080 28648
rect 5132 28636 5138 28688
rect 7116 28676 7144 28707
rect 7466 28704 7472 28716
rect 7524 28704 7530 28756
rect 8938 28744 8944 28756
rect 8899 28716 8944 28744
rect 8938 28704 8944 28716
rect 8996 28704 9002 28756
rect 10042 28704 10048 28756
rect 10100 28744 10106 28756
rect 10689 28747 10747 28753
rect 10689 28744 10701 28747
rect 10100 28716 10701 28744
rect 10100 28704 10106 28716
rect 10689 28713 10701 28716
rect 10735 28713 10747 28747
rect 10689 28707 10747 28713
rect 11146 28704 11152 28756
rect 11204 28744 11210 28756
rect 12391 28747 12449 28753
rect 12391 28744 12403 28747
rect 11204 28716 12403 28744
rect 11204 28704 11210 28716
rect 12391 28713 12403 28716
rect 12437 28713 12449 28747
rect 12391 28707 12449 28713
rect 7745 28679 7803 28685
rect 7745 28676 7757 28679
rect 7116 28648 7757 28676
rect 7745 28645 7757 28648
rect 7791 28676 7803 28679
rect 8113 28679 8171 28685
rect 8113 28676 8125 28679
rect 7791 28648 8125 28676
rect 7791 28645 7803 28648
rect 7745 28639 7803 28645
rect 8113 28645 8125 28648
rect 8159 28645 8171 28679
rect 9858 28676 9864 28688
rect 9819 28648 9864 28676
rect 8113 28639 8171 28645
rect 9858 28636 9864 28648
rect 9916 28636 9922 28688
rect 10410 28676 10416 28688
rect 10371 28648 10416 28676
rect 10410 28636 10416 28648
rect 10468 28636 10474 28688
rect 106 28568 112 28620
rect 164 28608 170 28620
rect 2866 28608 2872 28620
rect 164 28580 2872 28608
rect 164 28568 170 28580
rect 2866 28568 2872 28580
rect 2924 28568 2930 28620
rect 11238 28608 11244 28620
rect 11199 28580 11244 28608
rect 11238 28568 11244 28580
rect 11296 28568 11302 28620
rect 12320 28611 12378 28617
rect 12320 28577 12332 28611
rect 12366 28608 12378 28611
rect 12618 28608 12624 28620
rect 12366 28580 12624 28608
rect 12366 28577 12378 28580
rect 12320 28571 12378 28577
rect 12618 28568 12624 28580
rect 12676 28568 12682 28620
rect 2406 28500 2412 28552
rect 2464 28540 2470 28552
rect 4706 28540 4712 28552
rect 2464 28512 4712 28540
rect 2464 28500 2470 28512
rect 4706 28500 4712 28512
rect 4764 28500 4770 28552
rect 6181 28543 6239 28549
rect 6181 28509 6193 28543
rect 6227 28540 6239 28543
rect 6638 28540 6644 28552
rect 6227 28512 6644 28540
rect 6227 28509 6239 28512
rect 6181 28503 6239 28509
rect 6638 28500 6644 28512
rect 6696 28500 6702 28552
rect 7650 28500 7656 28552
rect 7708 28540 7714 28552
rect 8021 28543 8079 28549
rect 8021 28540 8033 28543
rect 7708 28512 8033 28540
rect 7708 28500 7714 28512
rect 8021 28509 8033 28512
rect 8067 28509 8079 28543
rect 8294 28540 8300 28552
rect 8255 28512 8300 28540
rect 8021 28503 8079 28509
rect 8294 28500 8300 28512
rect 8352 28500 8358 28552
rect 9493 28543 9551 28549
rect 9493 28509 9505 28543
rect 9539 28540 9551 28543
rect 9769 28543 9827 28549
rect 9769 28540 9781 28543
rect 9539 28512 9781 28540
rect 9539 28509 9551 28512
rect 9493 28503 9551 28509
rect 9769 28509 9781 28512
rect 9815 28540 9827 28543
rect 11379 28543 11437 28549
rect 11379 28540 11391 28543
rect 9815 28512 11391 28540
rect 9815 28509 9827 28512
rect 9769 28503 9827 28509
rect 11379 28509 11391 28512
rect 11425 28509 11437 28543
rect 11379 28503 11437 28509
rect 3878 28432 3884 28484
rect 3936 28472 3942 28484
rect 4062 28472 4068 28484
rect 3936 28444 4068 28472
rect 3936 28432 3942 28444
rect 4062 28432 4068 28444
rect 4120 28432 4126 28484
rect 5261 28475 5319 28481
rect 5261 28441 5273 28475
rect 5307 28472 5319 28475
rect 5534 28472 5540 28484
rect 5307 28444 5540 28472
rect 5307 28441 5319 28444
rect 5261 28435 5319 28441
rect 5534 28432 5540 28444
rect 5592 28472 5598 28484
rect 6914 28472 6920 28484
rect 5592 28444 6920 28472
rect 5592 28432 5598 28444
rect 6914 28432 6920 28444
rect 6972 28432 6978 28484
rect 3510 28364 3516 28416
rect 3568 28404 3574 28416
rect 5994 28404 6000 28416
rect 3568 28376 6000 28404
rect 3568 28364 3574 28376
rect 5994 28364 6000 28376
rect 6052 28364 6058 28416
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 2406 28200 2412 28212
rect 2367 28172 2412 28200
rect 2406 28160 2412 28172
rect 2464 28160 2470 28212
rect 3418 28200 3424 28212
rect 3379 28172 3424 28200
rect 3418 28160 3424 28172
rect 3476 28160 3482 28212
rect 4706 28160 4712 28212
rect 4764 28200 4770 28212
rect 5721 28203 5779 28209
rect 5721 28200 5733 28203
rect 4764 28172 5733 28200
rect 4764 28160 4770 28172
rect 5721 28169 5733 28172
rect 5767 28169 5779 28203
rect 5721 28163 5779 28169
rect 9033 28203 9091 28209
rect 9033 28169 9045 28203
rect 9079 28200 9091 28203
rect 9490 28200 9496 28212
rect 9079 28172 9496 28200
rect 9079 28169 9091 28172
rect 9033 28163 9091 28169
rect 9490 28160 9496 28172
rect 9548 28200 9554 28212
rect 9858 28200 9864 28212
rect 9548 28172 9864 28200
rect 9548 28160 9554 28172
rect 9858 28160 9864 28172
rect 9916 28160 9922 28212
rect 3326 28092 3332 28144
rect 3384 28132 3390 28144
rect 3605 28135 3663 28141
rect 3605 28132 3617 28135
rect 3384 28104 3617 28132
rect 3384 28092 3390 28104
rect 3605 28101 3617 28104
rect 3651 28101 3663 28135
rect 3605 28095 3663 28101
rect 6178 28092 6184 28144
rect 6236 28132 6242 28144
rect 11238 28132 11244 28144
rect 6236 28104 11244 28132
rect 6236 28092 6242 28104
rect 11238 28092 11244 28104
rect 11296 28092 11302 28144
rect 2685 28067 2743 28073
rect 2685 28064 2697 28067
rect 2215 28036 2697 28064
rect 2215 28005 2243 28036
rect 2685 28033 2697 28036
rect 2731 28064 2743 28067
rect 4522 28064 4528 28076
rect 2731 28036 4528 28064
rect 2731 28033 2743 28036
rect 2685 28027 2743 28033
rect 4522 28024 4528 28036
rect 4580 28024 4586 28076
rect 9677 28067 9735 28073
rect 9677 28064 9689 28067
rect 8956 28036 9689 28064
rect 2200 27999 2258 28005
rect 2200 27965 2212 27999
rect 2246 27965 2258 27999
rect 2200 27959 2258 27965
rect 3212 27999 3270 28005
rect 3212 27965 3224 27999
rect 3258 27996 3270 27999
rect 3326 27996 3332 28008
rect 3258 27968 3332 27996
rect 3258 27965 3270 27968
rect 3212 27959 3270 27965
rect 3326 27956 3332 27968
rect 3384 27956 3390 28008
rect 4157 27999 4215 28005
rect 4157 27965 4169 27999
rect 4203 27996 4215 27999
rect 4246 27996 4252 28008
rect 4203 27968 4252 27996
rect 4203 27965 4215 27968
rect 4157 27959 4215 27965
rect 4246 27956 4252 27968
rect 4304 27956 4310 28008
rect 4982 27996 4988 28008
rect 4448 27968 4988 27996
rect 2682 27888 2688 27940
rect 2740 27928 2746 27940
rect 4448 27928 4476 27968
rect 4982 27956 4988 27968
rect 5040 27956 5046 28008
rect 5534 27956 5540 28008
rect 5592 27996 5598 28008
rect 6876 27999 6934 28005
rect 6876 27996 6888 27999
rect 5592 27968 6888 27996
rect 5592 27956 5598 27968
rect 6876 27965 6888 27968
rect 6922 27996 6934 27999
rect 7285 27999 7343 28005
rect 7285 27996 7297 27999
rect 6922 27968 7297 27996
rect 6922 27965 6934 27968
rect 6876 27959 6934 27965
rect 7285 27965 7297 27968
rect 7331 27965 7343 27999
rect 7285 27959 7343 27965
rect 8113 27999 8171 28005
rect 8113 27965 8125 27999
rect 8159 27996 8171 27999
rect 8846 27996 8852 28008
rect 8159 27968 8852 27996
rect 8159 27965 8171 27968
rect 8113 27959 8171 27965
rect 8846 27956 8852 27968
rect 8904 27956 8910 28008
rect 2740 27900 4476 27928
rect 4519 27931 4577 27937
rect 2740 27888 2746 27900
rect 4519 27897 4531 27931
rect 4565 27928 4577 27931
rect 4706 27928 4712 27940
rect 4565 27900 4712 27928
rect 4565 27897 4577 27900
rect 4519 27891 4577 27897
rect 2866 27820 2872 27872
rect 2924 27860 2930 27872
rect 3053 27863 3111 27869
rect 3053 27860 3065 27863
rect 2924 27832 3065 27860
rect 2924 27820 2930 27832
rect 3053 27829 3065 27832
rect 3099 27860 3111 27863
rect 3878 27860 3884 27872
rect 3099 27832 3884 27860
rect 3099 27829 3111 27832
rect 3053 27823 3111 27829
rect 3878 27820 3884 27832
rect 3936 27820 3942 27872
rect 4065 27863 4123 27869
rect 4065 27829 4077 27863
rect 4111 27860 4123 27863
rect 4534 27860 4562 27891
rect 4706 27888 4712 27900
rect 4764 27928 4770 27940
rect 6181 27931 6239 27937
rect 6181 27928 6193 27931
rect 4764 27900 6193 27928
rect 4764 27888 4770 27900
rect 6181 27897 6193 27900
rect 6227 27928 6239 27931
rect 6546 27928 6552 27940
rect 6227 27900 6552 27928
rect 6227 27897 6239 27900
rect 6181 27891 6239 27897
rect 6546 27888 6552 27900
rect 6604 27928 6610 27940
rect 6963 27931 7021 27937
rect 6604 27900 6919 27928
rect 6604 27888 6610 27900
rect 5074 27860 5080 27872
rect 4111 27832 4562 27860
rect 5035 27832 5080 27860
rect 4111 27829 4123 27832
rect 4065 27823 4123 27829
rect 5074 27820 5080 27832
rect 5132 27860 5138 27872
rect 5353 27863 5411 27869
rect 5353 27860 5365 27863
rect 5132 27832 5365 27860
rect 5132 27820 5138 27832
rect 5353 27829 5365 27832
rect 5399 27829 5411 27863
rect 6638 27860 6644 27872
rect 6599 27832 6644 27860
rect 5353 27823 5411 27829
rect 6638 27820 6644 27832
rect 6696 27820 6702 27872
rect 6891 27860 6919 27900
rect 6963 27897 6975 27931
rect 7009 27928 7021 27931
rect 7650 27928 7656 27940
rect 7009 27900 7656 27928
rect 7009 27897 7021 27900
rect 6963 27891 7021 27897
rect 7650 27888 7656 27900
rect 7708 27888 7714 27940
rect 8434 27931 8492 27937
rect 8434 27928 8446 27931
rect 7944 27900 8446 27928
rect 7944 27869 7972 27900
rect 8434 27897 8446 27900
rect 8480 27928 8492 27931
rect 8956 27928 8984 28036
rect 9677 28033 9689 28036
rect 9723 28064 9735 28067
rect 9723 28036 10225 28064
rect 9723 28033 9735 28036
rect 9677 28027 9735 28033
rect 9861 27999 9919 28005
rect 9861 27996 9873 27999
rect 8480 27900 8984 27928
rect 9324 27968 9873 27996
rect 8480 27897 8492 27900
rect 8434 27891 8492 27897
rect 7929 27863 7987 27869
rect 7929 27860 7941 27863
rect 6891 27832 7941 27860
rect 7929 27829 7941 27832
rect 7975 27829 7987 27863
rect 7929 27823 7987 27829
rect 8018 27820 8024 27872
rect 8076 27860 8082 27872
rect 9324 27869 9352 27968
rect 9861 27965 9873 27968
rect 9907 27965 9919 27999
rect 9861 27959 9919 27965
rect 10197 27937 10225 28036
rect 10182 27931 10240 27937
rect 10182 27897 10194 27931
rect 10228 27897 10240 27931
rect 10182 27891 10240 27897
rect 9309 27863 9367 27869
rect 9309 27860 9321 27863
rect 8076 27832 9321 27860
rect 8076 27820 8082 27832
rect 9309 27829 9321 27832
rect 9355 27829 9367 27863
rect 9309 27823 9367 27829
rect 9858 27820 9864 27872
rect 9916 27860 9922 27872
rect 10781 27863 10839 27869
rect 10781 27860 10793 27863
rect 9916 27832 10793 27860
rect 9916 27820 9922 27832
rect 10781 27829 10793 27832
rect 10827 27829 10839 27863
rect 12618 27860 12624 27872
rect 12579 27832 12624 27860
rect 10781 27823 10839 27829
rect 12618 27820 12624 27832
rect 12676 27820 12682 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 4982 27616 4988 27668
rect 5040 27656 5046 27668
rect 7650 27656 7656 27668
rect 5040 27628 7052 27656
rect 7611 27628 7656 27656
rect 5040 27616 5046 27628
rect 4706 27548 4712 27600
rect 4764 27588 4770 27600
rect 6270 27588 6276 27600
rect 4764 27560 4809 27588
rect 5368 27560 6276 27588
rect 4764 27548 4770 27560
rect 2682 27520 2688 27532
rect 2643 27492 2688 27520
rect 2682 27480 2688 27492
rect 2740 27480 2746 27532
rect 2958 27520 2964 27532
rect 2919 27492 2964 27520
rect 2958 27480 2964 27492
rect 3016 27480 3022 27532
rect 3970 27480 3976 27532
rect 4028 27520 4034 27532
rect 5368 27529 5396 27560
rect 6270 27548 6276 27560
rect 6328 27588 6334 27600
rect 6365 27591 6423 27597
rect 6365 27588 6377 27591
rect 6328 27560 6377 27588
rect 6328 27548 6334 27560
rect 6365 27557 6377 27560
rect 6411 27557 6423 27591
rect 6914 27588 6920 27600
rect 6875 27560 6920 27588
rect 6365 27551 6423 27557
rect 6914 27548 6920 27560
rect 6972 27548 6978 27600
rect 5353 27523 5411 27529
rect 5353 27520 5365 27523
rect 4028 27492 5365 27520
rect 4028 27480 4034 27492
rect 5353 27489 5365 27492
rect 5399 27489 5411 27523
rect 7024 27520 7052 27628
rect 7650 27616 7656 27628
rect 7708 27616 7714 27668
rect 9490 27656 9496 27668
rect 9451 27628 9496 27656
rect 9490 27616 9496 27628
rect 9548 27616 9554 27668
rect 8478 27588 8484 27600
rect 8439 27560 8484 27588
rect 8478 27548 8484 27560
rect 8536 27548 8542 27600
rect 9858 27588 9864 27600
rect 9819 27560 9864 27588
rect 9858 27548 9864 27560
rect 9916 27548 9922 27600
rect 7742 27520 7748 27532
rect 7024 27492 7748 27520
rect 5353 27483 5411 27489
rect 7742 27480 7748 27492
rect 7800 27480 7806 27532
rect 7834 27480 7840 27532
rect 7892 27520 7898 27532
rect 8205 27523 8263 27529
rect 8205 27520 8217 27523
rect 7892 27492 8217 27520
rect 7892 27480 7898 27492
rect 8205 27489 8217 27492
rect 8251 27489 8263 27523
rect 8205 27483 8263 27489
rect 3145 27455 3203 27461
rect 3145 27421 3157 27455
rect 3191 27452 3203 27455
rect 4430 27452 4436 27464
rect 3191 27424 4436 27452
rect 3191 27421 3203 27424
rect 3145 27415 3203 27421
rect 4430 27412 4436 27424
rect 4488 27412 4494 27464
rect 5994 27412 6000 27464
rect 6052 27452 6058 27464
rect 6273 27455 6331 27461
rect 6273 27452 6285 27455
rect 6052 27424 6285 27452
rect 6052 27412 6058 27424
rect 6273 27421 6285 27424
rect 6319 27421 6331 27455
rect 6273 27415 6331 27421
rect 9769 27455 9827 27461
rect 9769 27421 9781 27455
rect 9815 27452 9827 27455
rect 10226 27452 10232 27464
rect 9815 27424 10232 27452
rect 9815 27421 9827 27424
rect 9769 27415 9827 27421
rect 10226 27412 10232 27424
rect 10284 27412 10290 27464
rect 3418 27344 3424 27396
rect 3476 27384 3482 27396
rect 6730 27384 6736 27396
rect 3476 27356 6736 27384
rect 3476 27344 3482 27356
rect 6730 27344 6736 27356
rect 6788 27344 6794 27396
rect 10318 27384 10324 27396
rect 10279 27356 10324 27384
rect 10318 27344 10324 27356
rect 10376 27344 10382 27396
rect 3142 27276 3148 27328
rect 3200 27316 3206 27328
rect 3436 27316 3464 27344
rect 4246 27316 4252 27328
rect 3200 27288 3464 27316
rect 4207 27288 4252 27316
rect 3200 27276 3206 27288
rect 4246 27276 4252 27288
rect 4304 27276 4310 27328
rect 8846 27316 8852 27328
rect 8807 27288 8852 27316
rect 8846 27276 8852 27288
rect 8904 27276 8910 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 2682 27112 2688 27124
rect 2643 27084 2688 27112
rect 2682 27072 2688 27084
rect 2740 27072 2746 27124
rect 5718 27112 5724 27124
rect 3804 27084 5724 27112
rect 3804 26976 3832 27084
rect 5718 27072 5724 27084
rect 5776 27072 5782 27124
rect 6270 27112 6276 27124
rect 6231 27084 6276 27112
rect 6270 27072 6276 27084
rect 6328 27072 6334 27124
rect 6730 27072 6736 27124
rect 6788 27112 6794 27124
rect 8665 27115 8723 27121
rect 8665 27112 8677 27115
rect 6788 27084 8677 27112
rect 6788 27072 6794 27084
rect 8665 27081 8677 27084
rect 8711 27081 8723 27115
rect 9858 27112 9864 27124
rect 9819 27084 9864 27112
rect 8665 27075 8723 27081
rect 4062 27004 4068 27056
rect 4120 27044 4126 27056
rect 4120 27016 5120 27044
rect 4120 27004 4126 27016
rect 3436 26948 3832 26976
rect 3881 26979 3939 26985
rect 3436 26917 3464 26948
rect 3881 26945 3893 26979
rect 3927 26976 3939 26979
rect 4246 26976 4252 26988
rect 3927 26948 4252 26976
rect 3927 26945 3939 26948
rect 3881 26939 3939 26945
rect 4246 26936 4252 26948
rect 4304 26936 4310 26988
rect 5092 26985 5120 27016
rect 5994 27004 6000 27056
rect 6052 27044 6058 27056
rect 6549 27047 6607 27053
rect 6549 27044 6561 27047
rect 6052 27016 6561 27044
rect 6052 27004 6058 27016
rect 6549 27013 6561 27016
rect 6595 27013 6607 27047
rect 6549 27007 6607 27013
rect 7742 27004 7748 27056
rect 7800 27044 7806 27056
rect 8297 27047 8355 27053
rect 8297 27044 8309 27047
rect 7800 27016 8309 27044
rect 7800 27004 7806 27016
rect 8297 27013 8309 27016
rect 8343 27013 8355 27047
rect 8297 27007 8355 27013
rect 5077 26979 5135 26985
rect 5077 26945 5089 26979
rect 5123 26945 5135 26979
rect 8018 26976 8024 26988
rect 7979 26948 8024 26976
rect 5077 26939 5135 26945
rect 8018 26936 8024 26948
rect 8076 26936 8082 26988
rect 2133 26911 2191 26917
rect 2133 26908 2145 26911
rect 1964 26880 2145 26908
rect 1854 26732 1860 26784
rect 1912 26772 1918 26784
rect 1964 26781 1992 26880
rect 2133 26877 2145 26880
rect 2179 26877 2191 26911
rect 2133 26871 2191 26877
rect 3053 26911 3111 26917
rect 3053 26877 3065 26911
rect 3099 26908 3111 26911
rect 3421 26911 3479 26917
rect 3421 26908 3433 26911
rect 3099 26880 3433 26908
rect 3099 26877 3111 26880
rect 3053 26871 3111 26877
rect 3421 26877 3433 26880
rect 3467 26877 3479 26911
rect 3421 26871 3479 26877
rect 3605 26911 3663 26917
rect 3605 26877 3617 26911
rect 3651 26877 3663 26911
rect 7285 26911 7343 26917
rect 7285 26908 7297 26911
rect 3605 26871 3663 26877
rect 7116 26880 7297 26908
rect 2958 26800 2964 26852
rect 3016 26840 3022 26852
rect 3510 26840 3516 26852
rect 3016 26812 3516 26840
rect 3016 26800 3022 26812
rect 3510 26800 3516 26812
rect 3568 26840 3574 26852
rect 3620 26840 3648 26871
rect 3568 26812 3648 26840
rect 3568 26800 3574 26812
rect 4614 26800 4620 26852
rect 4672 26840 4678 26852
rect 4801 26843 4859 26849
rect 4801 26840 4813 26843
rect 4672 26812 4813 26840
rect 4672 26800 4678 26812
rect 4801 26809 4813 26812
rect 4847 26809 4859 26843
rect 4801 26803 4859 26809
rect 4893 26843 4951 26849
rect 4893 26809 4905 26843
rect 4939 26840 4951 26843
rect 5074 26840 5080 26852
rect 4939 26812 5080 26840
rect 4939 26809 4951 26812
rect 4893 26803 4951 26809
rect 5074 26800 5080 26812
rect 5132 26840 5138 26852
rect 5721 26843 5779 26849
rect 5721 26840 5733 26843
rect 5132 26812 5733 26840
rect 5132 26800 5138 26812
rect 5721 26809 5733 26812
rect 5767 26809 5779 26843
rect 5721 26803 5779 26809
rect 1949 26775 2007 26781
rect 1949 26772 1961 26775
rect 1912 26744 1961 26772
rect 1912 26732 1918 26744
rect 1949 26741 1961 26744
rect 1995 26741 2007 26775
rect 2314 26772 2320 26784
rect 2275 26744 2320 26772
rect 1949 26735 2007 26741
rect 2314 26732 2320 26744
rect 2372 26732 2378 26784
rect 4525 26775 4583 26781
rect 4525 26741 4537 26775
rect 4571 26772 4583 26775
rect 4706 26772 4712 26784
rect 4571 26744 4712 26772
rect 4571 26741 4583 26744
rect 4525 26735 4583 26741
rect 4706 26732 4712 26744
rect 4764 26732 4770 26784
rect 5810 26732 5816 26784
rect 5868 26772 5874 26784
rect 7116 26781 7144 26880
rect 7285 26877 7297 26880
rect 7331 26877 7343 26911
rect 7742 26908 7748 26920
rect 7703 26880 7748 26908
rect 7285 26871 7343 26877
rect 7742 26868 7748 26880
rect 7800 26868 7806 26920
rect 8294 26868 8300 26920
rect 8352 26908 8358 26920
rect 8680 26908 8708 27075
rect 9858 27072 9864 27084
rect 9916 27072 9922 27124
rect 10226 27112 10232 27124
rect 10187 27084 10232 27112
rect 10226 27072 10232 27084
rect 10284 27112 10290 27124
rect 10551 27115 10609 27121
rect 10551 27112 10563 27115
rect 10284 27084 10563 27112
rect 10284 27072 10290 27084
rect 10551 27081 10563 27084
rect 10597 27081 10609 27115
rect 10551 27075 10609 27081
rect 8849 26911 8907 26917
rect 8849 26908 8861 26911
rect 8352 26880 8477 26908
rect 8680 26880 8861 26908
rect 8352 26868 8358 26880
rect 8449 26840 8477 26880
rect 8849 26877 8861 26880
rect 8895 26877 8907 26911
rect 9306 26908 9312 26920
rect 9267 26880 9312 26908
rect 8849 26871 8907 26877
rect 9306 26868 9312 26880
rect 9364 26868 9370 26920
rect 10448 26911 10506 26917
rect 10448 26908 10460 26911
rect 9876 26880 10460 26908
rect 9876 26840 9904 26880
rect 10448 26877 10460 26880
rect 10494 26908 10506 26911
rect 10873 26911 10931 26917
rect 10873 26908 10885 26911
rect 10494 26880 10885 26908
rect 10494 26877 10506 26880
rect 10448 26871 10506 26877
rect 10873 26877 10885 26880
rect 10919 26877 10931 26911
rect 10873 26871 10931 26877
rect 8449 26812 9904 26840
rect 7101 26775 7159 26781
rect 7101 26772 7113 26775
rect 5868 26744 7113 26772
rect 5868 26732 5874 26744
rect 7101 26741 7113 26744
rect 7147 26741 7159 26775
rect 7101 26735 7159 26741
rect 8846 26732 8852 26784
rect 8904 26772 8910 26784
rect 8941 26775 8999 26781
rect 8941 26772 8953 26775
rect 8904 26744 8953 26772
rect 8904 26732 8910 26744
rect 8941 26741 8953 26744
rect 8987 26741 8999 26775
rect 8941 26735 8999 26741
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 3145 26571 3203 26577
rect 3145 26537 3157 26571
rect 3191 26568 3203 26571
rect 4246 26568 4252 26580
rect 3191 26540 4252 26568
rect 3191 26537 3203 26540
rect 3145 26531 3203 26537
rect 4246 26528 4252 26540
rect 4304 26528 4310 26580
rect 4430 26528 4436 26580
rect 4488 26568 4494 26580
rect 5077 26571 5135 26577
rect 5077 26568 5089 26571
rect 4488 26540 5089 26568
rect 4488 26528 4494 26540
rect 5077 26537 5089 26540
rect 5123 26537 5135 26571
rect 7282 26568 7288 26580
rect 7243 26540 7288 26568
rect 5077 26531 5135 26537
rect 7282 26528 7288 26540
rect 7340 26568 7346 26580
rect 7653 26571 7711 26577
rect 7653 26568 7665 26571
rect 7340 26540 7665 26568
rect 7340 26528 7346 26540
rect 7653 26537 7665 26540
rect 7699 26568 7711 26571
rect 7742 26568 7748 26580
rect 7699 26540 7748 26568
rect 7699 26537 7711 26540
rect 7653 26531 7711 26537
rect 7742 26528 7748 26540
rect 7800 26528 7806 26580
rect 8846 26528 8852 26580
rect 8904 26568 8910 26580
rect 9769 26571 9827 26577
rect 9769 26568 9781 26571
rect 8904 26540 9781 26568
rect 8904 26528 8910 26540
rect 9769 26537 9781 26540
rect 9815 26537 9827 26571
rect 9769 26531 9827 26537
rect 2501 26503 2559 26509
rect 2501 26469 2513 26503
rect 2547 26500 2559 26503
rect 3510 26500 3516 26512
rect 2547 26472 3516 26500
rect 2547 26469 2559 26472
rect 2501 26463 2559 26469
rect 3510 26460 3516 26472
rect 3568 26500 3574 26512
rect 4798 26500 4804 26512
rect 3568 26472 4568 26500
rect 4759 26472 4804 26500
rect 3568 26460 3574 26472
rect 2961 26435 3019 26441
rect 2961 26401 2973 26435
rect 3007 26432 3019 26435
rect 3326 26432 3332 26444
rect 3007 26404 3332 26432
rect 3007 26401 3019 26404
rect 2961 26395 3019 26401
rect 3326 26392 3332 26404
rect 3384 26392 3390 26444
rect 4338 26432 4344 26444
rect 4299 26404 4344 26432
rect 4338 26392 4344 26404
rect 4396 26392 4402 26444
rect 4540 26441 4568 26472
rect 4798 26460 4804 26472
rect 4856 26460 4862 26512
rect 6365 26503 6423 26509
rect 6365 26469 6377 26503
rect 6411 26500 6423 26503
rect 6638 26500 6644 26512
rect 6411 26472 6644 26500
rect 6411 26469 6423 26472
rect 6365 26463 6423 26469
rect 6638 26460 6644 26472
rect 6696 26460 6702 26512
rect 8312 26472 10180 26500
rect 4525 26435 4583 26441
rect 4525 26401 4537 26435
rect 4571 26432 4583 26435
rect 4890 26432 4896 26444
rect 4571 26404 4896 26432
rect 4571 26401 4583 26404
rect 4525 26395 4583 26401
rect 4890 26392 4896 26404
rect 4948 26392 4954 26444
rect 5718 26432 5724 26444
rect 5679 26404 5724 26432
rect 5718 26392 5724 26404
rect 5776 26392 5782 26444
rect 6086 26432 6092 26444
rect 6047 26404 6092 26432
rect 6086 26392 6092 26404
rect 6144 26392 6150 26444
rect 8018 26432 8024 26444
rect 7979 26404 8024 26432
rect 8018 26392 8024 26404
rect 8076 26392 8082 26444
rect 8110 26392 8116 26444
rect 8168 26432 8174 26444
rect 8312 26441 8340 26472
rect 8297 26435 8355 26441
rect 8297 26432 8309 26435
rect 8168 26404 8309 26432
rect 8168 26392 8174 26404
rect 8297 26401 8309 26404
rect 8343 26401 8355 26435
rect 9674 26432 9680 26444
rect 9635 26404 9680 26432
rect 8297 26395 8355 26401
rect 9674 26392 9680 26404
rect 9732 26392 9738 26444
rect 10152 26441 10180 26472
rect 10137 26435 10195 26441
rect 10137 26401 10149 26435
rect 10183 26432 10195 26435
rect 10318 26432 10324 26444
rect 10183 26404 10324 26432
rect 10183 26401 10195 26404
rect 10137 26395 10195 26401
rect 10318 26392 10324 26404
rect 10376 26392 10382 26444
rect 11308 26435 11366 26441
rect 11308 26401 11320 26435
rect 11354 26432 11366 26435
rect 11514 26432 11520 26444
rect 11354 26404 11520 26432
rect 11354 26401 11366 26404
rect 11308 26395 11366 26401
rect 11514 26392 11520 26404
rect 11572 26392 11578 26444
rect 2314 26324 2320 26376
rect 2372 26364 2378 26376
rect 6104 26364 6132 26392
rect 8570 26364 8576 26376
rect 2372 26336 6132 26364
rect 8531 26336 8576 26364
rect 2372 26324 2378 26336
rect 8570 26324 8576 26336
rect 8628 26324 8634 26376
rect 11422 26364 11428 26376
rect 11394 26324 11428 26364
rect 11480 26324 11486 26376
rect 4614 26256 4620 26308
rect 4672 26296 4678 26308
rect 5445 26299 5503 26305
rect 5445 26296 5457 26299
rect 4672 26268 5457 26296
rect 4672 26256 4678 26268
rect 5445 26265 5457 26268
rect 5491 26265 5503 26299
rect 5445 26259 5503 26265
rect 7742 26256 7748 26308
rect 7800 26296 7806 26308
rect 8849 26299 8907 26305
rect 8849 26296 8861 26299
rect 7800 26268 8861 26296
rect 7800 26256 7806 26268
rect 8849 26265 8861 26268
rect 8895 26296 8907 26299
rect 9306 26296 9312 26308
rect 8895 26268 9312 26296
rect 8895 26265 8907 26268
rect 8849 26259 8907 26265
rect 9306 26256 9312 26268
rect 9364 26256 9370 26308
rect 10778 26228 10784 26240
rect 10739 26200 10784 26228
rect 10778 26188 10784 26200
rect 10836 26188 10842 26240
rect 11394 26237 11422 26324
rect 11379 26231 11437 26237
rect 11379 26197 11391 26231
rect 11425 26197 11437 26231
rect 11379 26191 11437 26197
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 4203 26027 4261 26033
rect 4203 25993 4215 26027
rect 4249 26024 4261 26027
rect 4614 26024 4620 26036
rect 4249 25996 4620 26024
rect 4249 25993 4261 25996
rect 4203 25987 4261 25993
rect 4614 25984 4620 25996
rect 4672 25984 4678 26036
rect 4890 26024 4896 26036
rect 4851 25996 4896 26024
rect 4890 25984 4896 25996
rect 4948 25984 4954 26036
rect 6086 26024 6092 26036
rect 6047 25996 6092 26024
rect 6086 25984 6092 25996
rect 6144 25984 6150 26036
rect 8662 25984 8668 26036
rect 8720 26024 8726 26036
rect 9674 26024 9680 26036
rect 8720 25996 9680 26024
rect 8720 25984 8726 25996
rect 9674 25984 9680 25996
rect 9732 26024 9738 26036
rect 9953 26027 10011 26033
rect 9953 26024 9965 26027
rect 9732 25996 9965 26024
rect 9732 25984 9738 25996
rect 9953 25993 9965 25996
rect 9999 25993 10011 26027
rect 10318 26024 10324 26036
rect 10279 25996 10324 26024
rect 9953 25987 10011 25993
rect 10318 25984 10324 25996
rect 10376 25984 10382 26036
rect 5258 25956 5264 25968
rect 5171 25928 5264 25956
rect 5258 25916 5264 25928
rect 5316 25956 5322 25968
rect 6822 25956 6828 25968
rect 5316 25928 6828 25956
rect 5316 25916 5322 25928
rect 6822 25916 6828 25928
rect 6880 25916 6886 25968
rect 4798 25848 4804 25900
rect 4856 25888 4862 25900
rect 8018 25888 8024 25900
rect 4856 25860 8024 25888
rect 4856 25848 4862 25860
rect 8018 25848 8024 25860
rect 8076 25888 8082 25900
rect 8205 25891 8263 25897
rect 8205 25888 8217 25891
rect 8076 25860 8217 25888
rect 8076 25848 8082 25860
rect 8205 25857 8217 25860
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 10597 25891 10655 25897
rect 10597 25857 10609 25891
rect 10643 25888 10655 25891
rect 10778 25888 10784 25900
rect 10643 25860 10784 25888
rect 10643 25857 10655 25860
rect 10597 25851 10655 25857
rect 10778 25848 10784 25860
rect 10836 25888 10842 25900
rect 12437 25891 12495 25897
rect 12437 25888 12449 25891
rect 10836 25860 12449 25888
rect 10836 25848 10842 25860
rect 12437 25857 12449 25860
rect 12483 25857 12495 25891
rect 12437 25851 12495 25857
rect 3418 25780 3424 25832
rect 3476 25820 3482 25832
rect 4100 25823 4158 25829
rect 4100 25820 4112 25823
rect 3476 25792 4112 25820
rect 3476 25780 3482 25792
rect 4100 25789 4112 25792
rect 4146 25820 4158 25823
rect 4525 25823 4583 25829
rect 4525 25820 4537 25823
rect 4146 25792 4537 25820
rect 4146 25789 4158 25792
rect 4100 25783 4158 25789
rect 4525 25789 4537 25792
rect 4571 25789 4583 25823
rect 5074 25820 5080 25832
rect 5035 25792 5080 25820
rect 4525 25783 4583 25789
rect 5074 25780 5080 25792
rect 5132 25780 5138 25832
rect 6822 25780 6828 25832
rect 6880 25820 6886 25832
rect 7190 25820 7196 25832
rect 6880 25792 7196 25820
rect 6880 25780 6886 25792
rect 7190 25780 7196 25792
rect 7248 25780 7254 25832
rect 7653 25823 7711 25829
rect 7653 25789 7665 25823
rect 7699 25789 7711 25823
rect 7653 25783 7711 25789
rect 7929 25823 7987 25829
rect 7929 25789 7941 25823
rect 7975 25820 7987 25823
rect 8754 25820 8760 25832
rect 7975 25792 8760 25820
rect 7975 25789 7987 25792
rect 7929 25783 7987 25789
rect 3973 25755 4031 25761
rect 3973 25721 3985 25755
rect 4019 25752 4031 25755
rect 4338 25752 4344 25764
rect 4019 25724 4344 25752
rect 4019 25721 4031 25724
rect 3973 25715 4031 25721
rect 4338 25712 4344 25724
rect 4396 25752 4402 25764
rect 5092 25752 5120 25780
rect 7668 25752 7696 25783
rect 8754 25780 8760 25792
rect 8812 25780 8818 25832
rect 9677 25823 9735 25829
rect 9677 25789 9689 25823
rect 9723 25820 9735 25823
rect 10410 25820 10416 25832
rect 9723 25792 10416 25820
rect 9723 25789 9735 25792
rect 9677 25783 9735 25789
rect 10410 25780 10416 25792
rect 10468 25780 10474 25832
rect 4396 25724 5120 25752
rect 7116 25724 7696 25752
rect 9078 25755 9136 25761
rect 4396 25712 4402 25724
rect 7116 25696 7144 25724
rect 9078 25721 9090 25755
rect 9124 25721 9136 25755
rect 9078 25715 9136 25721
rect 3053 25687 3111 25693
rect 3053 25653 3065 25687
rect 3099 25684 3111 25687
rect 3326 25684 3332 25696
rect 3099 25656 3332 25684
rect 3099 25653 3111 25656
rect 3053 25647 3111 25653
rect 3326 25644 3332 25656
rect 3384 25644 3390 25696
rect 5718 25684 5724 25696
rect 5679 25656 5724 25684
rect 5718 25644 5724 25656
rect 5776 25644 5782 25696
rect 7098 25684 7104 25696
rect 7059 25656 7104 25684
rect 7098 25644 7104 25656
rect 7156 25644 7162 25696
rect 7926 25644 7932 25696
rect 7984 25684 7990 25696
rect 8573 25687 8631 25693
rect 8573 25684 8585 25687
rect 7984 25656 8585 25684
rect 7984 25644 7990 25656
rect 8573 25653 8585 25656
rect 8619 25684 8631 25687
rect 9093 25684 9121 25715
rect 10686 25712 10692 25764
rect 10744 25752 10750 25764
rect 11241 25755 11299 25761
rect 10744 25724 10789 25752
rect 10744 25712 10750 25724
rect 11241 25721 11253 25755
rect 11287 25721 11299 25755
rect 11241 25715 11299 25721
rect 8619 25656 9121 25684
rect 11256 25684 11284 25715
rect 11514 25684 11520 25696
rect 11256 25656 11520 25684
rect 8619 25653 8631 25656
rect 8573 25647 8631 25653
rect 11514 25644 11520 25656
rect 11572 25644 11578 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 4617 25483 4675 25489
rect 4617 25449 4629 25483
rect 4663 25480 4675 25483
rect 4890 25480 4896 25492
rect 4663 25452 4896 25480
rect 4663 25449 4675 25452
rect 4617 25443 4675 25449
rect 4890 25440 4896 25452
rect 4948 25440 4954 25492
rect 7098 25440 7104 25492
rect 7156 25480 7162 25492
rect 8110 25480 8116 25492
rect 7156 25452 8116 25480
rect 7156 25440 7162 25452
rect 8110 25440 8116 25452
rect 8168 25480 8174 25492
rect 8389 25483 8447 25489
rect 8389 25480 8401 25483
rect 8168 25452 8401 25480
rect 8168 25440 8174 25452
rect 8389 25449 8401 25452
rect 8435 25449 8447 25483
rect 8754 25480 8760 25492
rect 8715 25452 8760 25480
rect 8389 25443 8447 25449
rect 8754 25440 8760 25452
rect 8812 25440 8818 25492
rect 9950 25440 9956 25492
rect 10008 25480 10014 25492
rect 10045 25483 10103 25489
rect 10045 25480 10057 25483
rect 10008 25452 10057 25480
rect 10008 25440 10014 25452
rect 10045 25449 10057 25452
rect 10091 25449 10103 25483
rect 10045 25443 10103 25449
rect 10597 25483 10655 25489
rect 10597 25449 10609 25483
rect 10643 25480 10655 25483
rect 10686 25480 10692 25492
rect 10643 25452 10692 25480
rect 10643 25449 10655 25452
rect 10597 25443 10655 25449
rect 10686 25440 10692 25452
rect 10744 25480 10750 25492
rect 10873 25483 10931 25489
rect 10873 25480 10885 25483
rect 10744 25452 10885 25480
rect 10744 25440 10750 25452
rect 10873 25449 10885 25452
rect 10919 25449 10931 25483
rect 10873 25443 10931 25449
rect 5997 25415 6055 25421
rect 5997 25381 6009 25415
rect 6043 25412 6055 25415
rect 6178 25412 6184 25424
rect 6043 25384 6184 25412
rect 6043 25381 6055 25384
rect 5997 25375 6055 25381
rect 6178 25372 6184 25384
rect 6236 25372 6242 25424
rect 7190 25412 7196 25424
rect 7151 25384 7196 25412
rect 7190 25372 7196 25384
rect 7248 25372 7254 25424
rect 7561 25415 7619 25421
rect 7561 25381 7573 25415
rect 7607 25412 7619 25415
rect 7742 25412 7748 25424
rect 7607 25384 7748 25412
rect 7607 25381 7619 25384
rect 7561 25375 7619 25381
rect 7742 25372 7748 25384
rect 7800 25372 7806 25424
rect 10410 25372 10416 25424
rect 10468 25412 10474 25424
rect 11330 25412 11336 25424
rect 10468 25384 11336 25412
rect 10468 25372 10474 25384
rect 11330 25372 11336 25384
rect 11388 25412 11394 25424
rect 11609 25415 11667 25421
rect 11609 25412 11621 25415
rect 11388 25384 11621 25412
rect 11388 25372 11394 25384
rect 11609 25381 11621 25384
rect 11655 25381 11667 25415
rect 11609 25375 11667 25381
rect 4430 25344 4436 25356
rect 4391 25316 4436 25344
rect 4430 25304 4436 25316
rect 4488 25304 4494 25356
rect 8570 25304 8576 25356
rect 8628 25344 8634 25356
rect 9398 25344 9404 25356
rect 8628 25316 9404 25344
rect 8628 25304 8634 25316
rect 9398 25304 9404 25316
rect 9456 25344 9462 25356
rect 9677 25347 9735 25353
rect 9677 25344 9689 25347
rect 9456 25316 9689 25344
rect 9456 25304 9462 25316
rect 9677 25313 9689 25316
rect 9723 25313 9735 25347
rect 9677 25307 9735 25313
rect 4338 25236 4344 25288
rect 4396 25276 4402 25288
rect 5905 25279 5963 25285
rect 5905 25276 5917 25279
rect 4396 25248 5917 25276
rect 4396 25236 4402 25248
rect 5905 25245 5917 25248
rect 5951 25276 5963 25279
rect 6086 25276 6092 25288
rect 5951 25248 6092 25276
rect 5951 25245 5963 25248
rect 5905 25239 5963 25245
rect 6086 25236 6092 25248
rect 6144 25236 6150 25288
rect 6549 25279 6607 25285
rect 6549 25245 6561 25279
rect 6595 25276 6607 25279
rect 7190 25276 7196 25288
rect 6595 25248 7196 25276
rect 6595 25245 6607 25248
rect 6549 25239 6607 25245
rect 7190 25236 7196 25248
rect 7248 25236 7254 25288
rect 7282 25236 7288 25288
rect 7340 25276 7346 25288
rect 7469 25279 7527 25285
rect 7469 25276 7481 25279
rect 7340 25248 7481 25276
rect 7340 25236 7346 25248
rect 7469 25245 7481 25248
rect 7515 25245 7527 25279
rect 7469 25239 7527 25245
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25276 8171 25279
rect 10042 25276 10048 25288
rect 8159 25248 10048 25276
rect 8159 25245 8171 25248
rect 8113 25239 8171 25245
rect 10042 25236 10048 25248
rect 10100 25236 10106 25288
rect 11517 25279 11575 25285
rect 11517 25245 11529 25279
rect 11563 25245 11575 25279
rect 11790 25276 11796 25288
rect 11751 25248 11796 25276
rect 11517 25239 11575 25245
rect 11422 25168 11428 25220
rect 11480 25208 11486 25220
rect 11532 25208 11560 25239
rect 11790 25236 11796 25248
rect 11848 25236 11854 25288
rect 11480 25180 11560 25208
rect 11480 25168 11486 25180
rect 5074 25140 5080 25152
rect 5035 25112 5080 25140
rect 5074 25100 5080 25112
rect 5132 25100 5138 25152
rect 5442 25140 5448 25152
rect 5403 25112 5448 25140
rect 5442 25100 5448 25112
rect 5500 25100 5506 25152
rect 6914 25140 6920 25152
rect 6875 25112 6920 25140
rect 6914 25100 6920 25112
rect 6972 25100 6978 25152
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 3283 24939 3341 24945
rect 3283 24905 3295 24939
rect 3329 24936 3341 24939
rect 4338 24936 4344 24948
rect 3329 24908 4344 24936
rect 3329 24905 3341 24908
rect 3283 24899 3341 24905
rect 4338 24896 4344 24908
rect 4396 24896 4402 24948
rect 4430 24896 4436 24948
rect 4488 24936 4494 24948
rect 4985 24939 5043 24945
rect 4985 24936 4997 24939
rect 4488 24908 4997 24936
rect 4488 24896 4494 24908
rect 4985 24905 4997 24908
rect 5031 24905 5043 24939
rect 4985 24899 5043 24905
rect 7926 24896 7932 24948
rect 7984 24936 7990 24948
rect 8665 24939 8723 24945
rect 8665 24936 8677 24939
rect 7984 24908 8677 24936
rect 7984 24896 7990 24908
rect 8665 24905 8677 24908
rect 8711 24936 8723 24939
rect 9950 24936 9956 24948
rect 8711 24908 9956 24936
rect 8711 24905 8723 24908
rect 8665 24899 8723 24905
rect 3050 24828 3056 24880
rect 3108 24868 3114 24880
rect 3605 24871 3663 24877
rect 3605 24868 3617 24871
rect 3108 24840 3617 24868
rect 3108 24828 3114 24840
rect 3227 24741 3255 24840
rect 3605 24837 3617 24840
rect 3651 24837 3663 24871
rect 3605 24831 3663 24837
rect 4062 24760 4068 24812
rect 4120 24800 4126 24812
rect 4448 24800 4476 24896
rect 8754 24868 8760 24880
rect 7208 24840 8760 24868
rect 7208 24812 7236 24840
rect 8754 24828 8760 24840
rect 8812 24828 8818 24880
rect 4120 24772 4476 24800
rect 4120 24760 4126 24772
rect 5442 24760 5448 24812
rect 5500 24800 5506 24812
rect 6549 24803 6607 24809
rect 6549 24800 6561 24803
rect 5500 24772 6561 24800
rect 5500 24760 5506 24772
rect 6549 24769 6561 24772
rect 6595 24769 6607 24803
rect 7190 24800 7196 24812
rect 7151 24772 7196 24800
rect 6549 24763 6607 24769
rect 3212 24735 3270 24741
rect 3212 24701 3224 24735
rect 3258 24701 3270 24735
rect 3212 24695 3270 24701
rect 4154 24692 4160 24744
rect 4212 24741 4218 24744
rect 4212 24735 4266 24741
rect 4212 24701 4220 24735
rect 4254 24732 4266 24735
rect 4617 24735 4675 24741
rect 4617 24732 4629 24735
rect 4254 24704 4629 24732
rect 4254 24701 4266 24704
rect 4212 24695 4266 24701
rect 4617 24701 4629 24704
rect 4663 24701 4675 24735
rect 4617 24695 4675 24701
rect 4212 24692 4218 24695
rect 4065 24667 4123 24673
rect 4065 24633 4077 24667
rect 4111 24664 4123 24667
rect 4295 24667 4353 24673
rect 4295 24664 4307 24667
rect 4111 24636 4307 24664
rect 4111 24633 4123 24636
rect 4065 24627 4123 24633
rect 4295 24633 4307 24636
rect 4341 24664 4353 24667
rect 5261 24667 5319 24673
rect 5261 24664 5273 24667
rect 4341 24636 5273 24664
rect 4341 24633 4353 24636
rect 4295 24627 4353 24633
rect 5261 24633 5273 24636
rect 5307 24633 5319 24667
rect 5261 24627 5319 24633
rect 5353 24667 5411 24673
rect 5353 24633 5365 24667
rect 5399 24664 5411 24667
rect 5442 24664 5448 24676
rect 5399 24636 5448 24664
rect 5399 24633 5411 24636
rect 5353 24627 5411 24633
rect 5442 24624 5448 24636
rect 5500 24624 5506 24676
rect 5902 24664 5908 24676
rect 5863 24636 5908 24664
rect 5902 24624 5908 24636
rect 5960 24624 5966 24676
rect 6178 24596 6184 24608
rect 6139 24568 6184 24596
rect 6178 24556 6184 24568
rect 6236 24556 6242 24608
rect 6564 24596 6592 24763
rect 7190 24760 7196 24772
rect 7248 24760 7254 24812
rect 7282 24760 7288 24812
rect 7340 24800 7346 24812
rect 8205 24803 8263 24809
rect 8205 24800 8217 24803
rect 7340 24772 8217 24800
rect 7340 24760 7346 24772
rect 8205 24769 8217 24772
rect 8251 24769 8263 24803
rect 8846 24800 8852 24812
rect 8807 24772 8852 24800
rect 8205 24763 8263 24769
rect 8846 24760 8852 24772
rect 8904 24760 8910 24812
rect 6914 24664 6920 24676
rect 6875 24636 6920 24664
rect 6914 24624 6920 24636
rect 6972 24624 6978 24676
rect 7009 24667 7067 24673
rect 7009 24633 7021 24667
rect 7055 24633 7067 24667
rect 8956 24664 8984 24908
rect 9950 24896 9956 24908
rect 10008 24936 10014 24948
rect 10045 24939 10103 24945
rect 10045 24936 10057 24939
rect 10008 24908 10057 24936
rect 10008 24896 10014 24908
rect 10045 24905 10057 24908
rect 10091 24905 10103 24939
rect 10045 24899 10103 24905
rect 11330 24896 11336 24948
rect 11388 24936 11394 24948
rect 11609 24939 11667 24945
rect 11609 24936 11621 24939
rect 11388 24908 11621 24936
rect 11388 24896 11394 24908
rect 11609 24905 11621 24908
rect 11655 24905 11667 24939
rect 11609 24899 11667 24905
rect 10410 24828 10416 24880
rect 10468 24868 10474 24880
rect 11422 24868 11428 24880
rect 10468 24840 11428 24868
rect 10468 24828 10474 24840
rect 11422 24828 11428 24840
rect 11480 24868 11486 24880
rect 11977 24871 12035 24877
rect 11977 24868 11989 24871
rect 11480 24840 11989 24868
rect 11480 24828 11486 24840
rect 11977 24837 11989 24840
rect 12023 24837 12035 24871
rect 11977 24831 12035 24837
rect 11333 24803 11391 24809
rect 11333 24769 11345 24803
rect 11379 24800 11391 24803
rect 11790 24800 11796 24812
rect 11379 24772 11796 24800
rect 11379 24769 11391 24772
rect 11333 24763 11391 24769
rect 11790 24760 11796 24772
rect 11848 24760 11854 24812
rect 9769 24735 9827 24741
rect 9769 24701 9781 24735
rect 9815 24732 9827 24735
rect 10413 24735 10471 24741
rect 10413 24732 10425 24735
rect 9815 24704 10425 24732
rect 9815 24701 9827 24704
rect 9769 24695 9827 24701
rect 10413 24701 10425 24704
rect 10459 24701 10471 24735
rect 10413 24695 10471 24701
rect 9170 24667 9228 24673
rect 9170 24664 9182 24667
rect 8956 24636 9182 24664
rect 7009 24627 7067 24633
rect 9170 24633 9182 24636
rect 9216 24633 9228 24667
rect 9170 24627 9228 24633
rect 7024 24596 7052 24627
rect 6564 24568 7052 24596
rect 7742 24556 7748 24608
rect 7800 24596 7806 24608
rect 7837 24599 7895 24605
rect 7837 24596 7849 24599
rect 7800 24568 7849 24596
rect 7800 24556 7806 24568
rect 7837 24565 7849 24568
rect 7883 24565 7895 24599
rect 10428 24596 10456 24695
rect 10686 24664 10692 24676
rect 10647 24636 10692 24664
rect 10686 24624 10692 24636
rect 10744 24624 10750 24676
rect 10781 24667 10839 24673
rect 10781 24633 10793 24667
rect 10827 24633 10839 24667
rect 10781 24627 10839 24633
rect 10796 24596 10824 24627
rect 10428 24568 10824 24596
rect 7837 24559 7895 24565
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 3099 24395 3157 24401
rect 3099 24361 3111 24395
rect 3145 24392 3157 24395
rect 6914 24392 6920 24404
rect 3145 24364 6920 24392
rect 3145 24361 3157 24364
rect 3099 24355 3157 24361
rect 6914 24352 6920 24364
rect 6972 24352 6978 24404
rect 8846 24392 8852 24404
rect 8807 24364 8852 24392
rect 8846 24352 8852 24364
rect 8904 24352 8910 24404
rect 9398 24392 9404 24404
rect 9359 24364 9404 24392
rect 9398 24352 9404 24364
rect 9456 24352 9462 24404
rect 11379 24395 11437 24401
rect 11379 24361 11391 24395
rect 11425 24392 11437 24395
rect 14826 24392 14832 24404
rect 11425 24364 14832 24392
rect 11425 24361 11437 24364
rect 11379 24355 11437 24361
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 4430 24284 4436 24336
rect 4488 24324 4494 24336
rect 4706 24324 4712 24336
rect 4488 24296 4712 24324
rect 4488 24284 4494 24296
rect 4706 24284 4712 24296
rect 4764 24324 4770 24336
rect 5214 24327 5272 24333
rect 5214 24324 5226 24327
rect 4764 24296 5226 24324
rect 4764 24284 4770 24296
rect 5214 24293 5226 24296
rect 5260 24293 5272 24327
rect 5214 24287 5272 24293
rect 5810 24284 5816 24336
rect 5868 24324 5874 24336
rect 6825 24327 6883 24333
rect 6825 24324 6837 24327
rect 5868 24296 6837 24324
rect 5868 24284 5874 24296
rect 6825 24293 6837 24296
rect 6871 24293 6883 24327
rect 9858 24324 9864 24336
rect 9819 24296 9864 24324
rect 6825 24287 6883 24293
rect 9858 24284 9864 24296
rect 9916 24284 9922 24336
rect 3028 24259 3086 24265
rect 3028 24225 3040 24259
rect 3074 24256 3086 24259
rect 3234 24256 3240 24268
rect 3074 24228 3240 24256
rect 3074 24225 3086 24228
rect 3028 24219 3086 24225
rect 3234 24216 3240 24228
rect 3292 24216 3298 24268
rect 6086 24256 6092 24268
rect 6047 24228 6092 24256
rect 6086 24216 6092 24228
rect 6144 24216 6150 24268
rect 8018 24216 8024 24268
rect 8076 24256 8082 24268
rect 8240 24259 8298 24265
rect 8240 24256 8252 24259
rect 8076 24228 8252 24256
rect 8076 24216 8082 24228
rect 8240 24225 8252 24228
rect 8286 24225 8298 24259
rect 11238 24256 11244 24268
rect 11199 24228 11244 24256
rect 8240 24219 8298 24225
rect 11238 24216 11244 24228
rect 11296 24216 11302 24268
rect 4893 24191 4951 24197
rect 4893 24188 4905 24191
rect 4724 24160 4905 24188
rect 3510 24052 3516 24064
rect 3471 24024 3516 24052
rect 3510 24012 3516 24024
rect 3568 24012 3574 24064
rect 4338 24012 4344 24064
rect 4396 24052 4402 24064
rect 4724 24061 4752 24160
rect 4893 24157 4905 24160
rect 4939 24157 4951 24191
rect 4893 24151 4951 24157
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24188 6607 24191
rect 6733 24191 6791 24197
rect 6733 24188 6745 24191
rect 6595 24160 6745 24188
rect 6595 24157 6607 24160
rect 6549 24151 6607 24157
rect 6733 24157 6745 24160
rect 6779 24188 6791 24191
rect 7834 24188 7840 24200
rect 6779 24160 7840 24188
rect 6779 24157 6791 24160
rect 6733 24151 6791 24157
rect 7834 24148 7840 24160
rect 7892 24148 7898 24200
rect 8754 24148 8760 24200
rect 8812 24188 8818 24200
rect 9766 24188 9772 24200
rect 8812 24160 9772 24188
rect 8812 24148 8818 24160
rect 9766 24148 9772 24160
rect 9824 24148 9830 24200
rect 10042 24188 10048 24200
rect 10003 24160 10048 24188
rect 10042 24148 10048 24160
rect 10100 24148 10106 24200
rect 5902 24080 5908 24132
rect 5960 24120 5966 24132
rect 7282 24120 7288 24132
rect 5960 24092 7288 24120
rect 5960 24080 5966 24092
rect 7282 24080 7288 24092
rect 7340 24080 7346 24132
rect 4709 24055 4767 24061
rect 4709 24052 4721 24055
rect 4396 24024 4721 24052
rect 4396 24012 4402 24024
rect 4709 24021 4721 24024
rect 4755 24021 4767 24055
rect 5810 24052 5816 24064
rect 5771 24024 5816 24052
rect 4709 24015 4767 24021
rect 5810 24012 5816 24024
rect 5868 24012 5874 24064
rect 6914 24012 6920 24064
rect 6972 24052 6978 24064
rect 7650 24052 7656 24064
rect 6972 24024 7656 24052
rect 6972 24012 6978 24024
rect 7650 24012 7656 24024
rect 7708 24052 7714 24064
rect 8343 24055 8401 24061
rect 8343 24052 8355 24055
rect 7708 24024 8355 24052
rect 7708 24012 7714 24024
rect 8343 24021 8355 24024
rect 8389 24021 8401 24055
rect 8343 24015 8401 24021
rect 9950 24012 9956 24064
rect 10008 24052 10014 24064
rect 10686 24052 10692 24064
rect 10008 24024 10692 24052
rect 10008 24012 10014 24024
rect 10686 24012 10692 24024
rect 10744 24012 10750 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 2317 23851 2375 23857
rect 2317 23817 2329 23851
rect 2363 23848 2375 23851
rect 4154 23848 4160 23860
rect 2363 23820 4160 23848
rect 2363 23817 2375 23820
rect 2317 23811 2375 23817
rect 2459 23653 2487 23820
rect 4154 23808 4160 23820
rect 4212 23848 4218 23860
rect 5534 23848 5540 23860
rect 4212 23820 5540 23848
rect 4212 23808 4218 23820
rect 5534 23808 5540 23820
rect 5592 23808 5598 23860
rect 5810 23808 5816 23860
rect 5868 23848 5874 23860
rect 6181 23851 6239 23857
rect 6181 23848 6193 23851
rect 5868 23820 6193 23848
rect 5868 23808 5874 23820
rect 6181 23817 6193 23820
rect 6227 23848 6239 23851
rect 7837 23851 7895 23857
rect 7837 23848 7849 23851
rect 6227 23820 7849 23848
rect 6227 23817 6239 23820
rect 6181 23811 6239 23817
rect 7837 23817 7849 23820
rect 7883 23848 7895 23851
rect 8570 23848 8576 23860
rect 7883 23820 8576 23848
rect 7883 23817 7895 23820
rect 7837 23811 7895 23817
rect 8570 23808 8576 23820
rect 8628 23808 8634 23860
rect 9398 23808 9404 23860
rect 9456 23848 9462 23860
rect 9493 23851 9551 23857
rect 9493 23848 9505 23851
rect 9456 23820 9505 23848
rect 9456 23808 9462 23820
rect 9493 23817 9505 23820
rect 9539 23848 9551 23851
rect 9858 23848 9864 23860
rect 9539 23820 9864 23848
rect 9539 23817 9551 23820
rect 9493 23811 9551 23817
rect 9858 23808 9864 23820
rect 9916 23808 9922 23860
rect 3053 23783 3111 23789
rect 3053 23749 3065 23783
rect 3099 23780 3111 23783
rect 3234 23780 3240 23792
rect 3099 23752 3240 23780
rect 3099 23749 3111 23752
rect 3053 23743 3111 23749
rect 3234 23740 3240 23752
rect 3292 23740 3298 23792
rect 5442 23740 5448 23792
rect 5500 23780 5506 23792
rect 5905 23783 5963 23789
rect 5905 23780 5917 23783
rect 5500 23752 5917 23780
rect 5500 23740 5506 23752
rect 5905 23749 5917 23752
rect 5951 23749 5963 23783
rect 5905 23743 5963 23749
rect 6748 23752 8524 23780
rect 2547 23715 2605 23721
rect 2547 23681 2559 23715
rect 2593 23712 2605 23715
rect 6748 23712 6776 23752
rect 8496 23724 8524 23752
rect 9766 23740 9772 23792
rect 9824 23780 9830 23792
rect 10965 23783 11023 23789
rect 10965 23780 10977 23783
rect 9824 23752 10977 23780
rect 9824 23740 9830 23752
rect 10965 23749 10977 23752
rect 11011 23749 11023 23783
rect 10965 23743 11023 23749
rect 6914 23712 6920 23724
rect 2593 23684 6776 23712
rect 6875 23684 6920 23712
rect 2593 23681 2605 23684
rect 2547 23675 2605 23681
rect 6914 23672 6920 23684
rect 6972 23672 6978 23724
rect 7282 23712 7288 23724
rect 7243 23684 7288 23712
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 8478 23712 8484 23724
rect 8391 23684 8484 23712
rect 8478 23672 8484 23684
rect 8536 23672 8542 23724
rect 8754 23712 8760 23724
rect 8715 23684 8760 23712
rect 8754 23672 8760 23684
rect 8812 23672 8818 23724
rect 10042 23672 10048 23724
rect 10100 23712 10106 23724
rect 10321 23715 10379 23721
rect 10321 23712 10333 23715
rect 10100 23684 10333 23712
rect 10100 23672 10106 23684
rect 10321 23681 10333 23684
rect 10367 23712 10379 23715
rect 11238 23712 11244 23724
rect 10367 23684 11244 23712
rect 10367 23681 10379 23684
rect 10321 23675 10379 23681
rect 11238 23672 11244 23684
rect 11296 23712 11302 23724
rect 11333 23715 11391 23721
rect 11333 23712 11345 23715
rect 11296 23684 11345 23712
rect 11296 23672 11302 23684
rect 11333 23681 11345 23684
rect 11379 23681 11391 23715
rect 11333 23675 11391 23681
rect 2444 23647 2502 23653
rect 2444 23613 2456 23647
rect 2490 23613 2502 23647
rect 2444 23607 2502 23613
rect 3050 23604 3056 23656
rect 3108 23644 3114 23656
rect 3234 23644 3240 23656
rect 3108 23616 3240 23644
rect 3108 23604 3114 23616
rect 3234 23604 3240 23616
rect 3292 23604 3298 23656
rect 3421 23647 3479 23653
rect 3421 23613 3433 23647
rect 3467 23613 3479 23647
rect 3421 23607 3479 23613
rect 3436 23576 3464 23607
rect 3510 23604 3516 23656
rect 3568 23644 3574 23656
rect 3881 23647 3939 23653
rect 3881 23644 3893 23647
rect 3568 23616 3893 23644
rect 3568 23604 3574 23616
rect 3881 23613 3893 23616
rect 3927 23613 3939 23647
rect 4890 23644 4896 23656
rect 3881 23607 3939 23613
rect 4126 23616 4896 23644
rect 3602 23576 3608 23588
rect 3436 23548 3608 23576
rect 3602 23536 3608 23548
rect 3660 23576 3666 23588
rect 4126 23576 4154 23616
rect 4890 23604 4896 23616
rect 4948 23604 4954 23656
rect 4985 23647 5043 23653
rect 4985 23613 4997 23647
rect 5031 23644 5043 23647
rect 5810 23644 5816 23656
rect 5031 23616 5816 23644
rect 5031 23613 5043 23616
rect 4985 23607 5043 23613
rect 3660 23548 4154 23576
rect 4249 23579 4307 23585
rect 3660 23536 3666 23548
rect 4249 23545 4261 23579
rect 4295 23576 4307 23579
rect 5000 23576 5028 23607
rect 5810 23604 5816 23616
rect 5868 23604 5874 23656
rect 4295 23548 5028 23576
rect 7009 23579 7067 23585
rect 4295 23545 4307 23548
rect 4249 23539 4307 23545
rect 7009 23545 7021 23579
rect 7055 23545 7067 23579
rect 7009 23539 7067 23545
rect 4430 23508 4436 23520
rect 4391 23480 4436 23508
rect 4430 23468 4436 23480
rect 4488 23508 4494 23520
rect 4801 23511 4859 23517
rect 4801 23508 4813 23511
rect 4488 23480 4813 23508
rect 4488 23468 4494 23480
rect 4801 23477 4813 23480
rect 4847 23477 4859 23511
rect 4801 23471 4859 23477
rect 5166 23468 5172 23520
rect 5224 23508 5230 23520
rect 5353 23511 5411 23517
rect 5353 23508 5365 23511
rect 5224 23480 5365 23508
rect 5224 23468 5230 23480
rect 5353 23477 5365 23480
rect 5399 23477 5411 23511
rect 5353 23471 5411 23477
rect 5534 23468 5540 23520
rect 5592 23508 5598 23520
rect 6178 23508 6184 23520
rect 5592 23480 6184 23508
rect 5592 23468 5598 23480
rect 6178 23468 6184 23480
rect 6236 23508 6242 23520
rect 6549 23511 6607 23517
rect 6549 23508 6561 23511
rect 6236 23480 6561 23508
rect 6236 23468 6242 23480
rect 6549 23477 6561 23480
rect 6595 23508 6607 23511
rect 7024 23508 7052 23539
rect 8570 23536 8576 23588
rect 8628 23576 8634 23588
rect 10045 23579 10103 23585
rect 8628 23548 8673 23576
rect 8628 23536 8634 23548
rect 10045 23545 10057 23579
rect 10091 23545 10103 23579
rect 10045 23539 10103 23545
rect 6595 23480 7052 23508
rect 6595 23477 6607 23480
rect 6549 23471 6607 23477
rect 8018 23468 8024 23520
rect 8076 23508 8082 23520
rect 8205 23511 8263 23517
rect 8205 23508 8217 23511
rect 8076 23480 8217 23508
rect 8076 23468 8082 23480
rect 8205 23477 8217 23480
rect 8251 23477 8263 23511
rect 8205 23471 8263 23477
rect 9674 23468 9680 23520
rect 9732 23508 9738 23520
rect 9769 23511 9827 23517
rect 9769 23508 9781 23511
rect 9732 23480 9781 23508
rect 9732 23468 9738 23480
rect 9769 23477 9781 23480
rect 9815 23508 9827 23511
rect 10060 23508 10088 23539
rect 10134 23536 10140 23588
rect 10192 23576 10198 23588
rect 10192 23548 10237 23576
rect 10192 23536 10198 23548
rect 9815 23480 10088 23508
rect 9815 23477 9827 23480
rect 9769 23471 9827 23477
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 3053 23307 3111 23313
rect 3053 23273 3065 23307
rect 3099 23304 3111 23307
rect 5534 23304 5540 23316
rect 3099 23276 5390 23304
rect 5495 23276 5540 23304
rect 3099 23273 3111 23276
rect 3053 23267 3111 23273
rect 3510 23236 3516 23248
rect 3471 23208 3516 23236
rect 3510 23196 3516 23208
rect 3568 23196 3574 23248
rect 4430 23196 4436 23248
rect 4488 23236 4494 23248
rect 4979 23239 5037 23245
rect 4979 23236 4991 23239
rect 4488 23208 4991 23236
rect 4488 23196 4494 23208
rect 4979 23205 4991 23208
rect 5025 23236 5037 23239
rect 5166 23236 5172 23248
rect 5025 23208 5172 23236
rect 5025 23205 5037 23208
rect 4979 23199 5037 23205
rect 5166 23196 5172 23208
rect 5224 23196 5230 23248
rect 5362 23236 5390 23276
rect 5534 23264 5540 23276
rect 5592 23264 5598 23316
rect 5810 23304 5816 23316
rect 5771 23276 5816 23304
rect 5810 23264 5816 23276
rect 5868 23264 5874 23316
rect 7650 23304 7656 23316
rect 7611 23276 7656 23304
rect 7650 23264 7656 23276
rect 7708 23264 7714 23316
rect 7834 23264 7840 23316
rect 7892 23304 7898 23316
rect 8251 23307 8309 23313
rect 8251 23304 8263 23307
rect 7892 23276 8263 23304
rect 7892 23264 7898 23276
rect 8251 23273 8263 23276
rect 8297 23273 8309 23307
rect 8251 23267 8309 23273
rect 8478 23264 8484 23316
rect 8536 23304 8542 23316
rect 8573 23307 8631 23313
rect 8573 23304 8585 23307
rect 8536 23276 8585 23304
rect 8536 23264 8542 23276
rect 8573 23273 8585 23276
rect 8619 23273 8631 23307
rect 9674 23304 9680 23316
rect 9635 23276 9680 23304
rect 8573 23267 8631 23273
rect 9674 23264 9680 23276
rect 9732 23264 9738 23316
rect 5626 23236 5632 23248
rect 5362 23208 5632 23236
rect 5626 23196 5632 23208
rect 5684 23196 5690 23248
rect 6546 23196 6552 23248
rect 6604 23236 6610 23248
rect 6686 23239 6744 23245
rect 6686 23236 6698 23239
rect 6604 23208 6698 23236
rect 6604 23196 6610 23208
rect 6686 23205 6698 23208
rect 6732 23205 6744 23239
rect 8018 23236 8024 23248
rect 6686 23199 6744 23205
rect 7852 23208 8024 23236
rect 106 23128 112 23180
rect 164 23168 170 23180
rect 2866 23168 2872 23180
rect 164 23140 2872 23168
rect 164 23128 170 23140
rect 2866 23128 2872 23140
rect 2924 23128 2930 23180
rect 3050 23128 3056 23180
rect 3108 23168 3114 23180
rect 3326 23168 3332 23180
rect 3108 23140 3332 23168
rect 3108 23128 3114 23140
rect 3326 23128 3332 23140
rect 3384 23128 3390 23180
rect 3418 23128 3424 23180
rect 3476 23168 3482 23180
rect 7852 23168 7880 23208
rect 8018 23196 8024 23208
rect 8076 23196 8082 23248
rect 8110 23168 8116 23180
rect 3476 23140 7880 23168
rect 8023 23140 8116 23168
rect 3476 23128 3482 23140
rect 8110 23128 8116 23140
rect 8168 23128 8174 23180
rect 10686 23168 10692 23180
rect 10647 23140 10692 23168
rect 10686 23128 10692 23140
rect 10744 23128 10750 23180
rect 4617 23103 4675 23109
rect 4617 23069 4629 23103
rect 4663 23069 4675 23103
rect 4617 23063 4675 23069
rect 6365 23103 6423 23109
rect 6365 23069 6377 23103
rect 6411 23069 6423 23103
rect 6365 23063 6423 23069
rect 3418 22924 3424 22976
rect 3476 22964 3482 22976
rect 4062 22964 4068 22976
rect 3476 22936 4068 22964
rect 3476 22924 3482 22936
rect 4062 22924 4068 22936
rect 4120 22924 4126 22976
rect 4522 22964 4528 22976
rect 4483 22936 4528 22964
rect 4522 22924 4528 22936
rect 4580 22964 4586 22976
rect 4632 22964 4660 23063
rect 4580 22936 4660 22964
rect 4580 22924 4586 22936
rect 5902 22924 5908 22976
rect 5960 22964 5966 22976
rect 6181 22967 6239 22973
rect 6181 22964 6193 22967
rect 5960 22936 6193 22964
rect 5960 22924 5966 22936
rect 6181 22933 6193 22936
rect 6227 22964 6239 22967
rect 6380 22964 6408 23063
rect 7926 23060 7932 23112
rect 7984 23100 7990 23112
rect 8128 23100 8156 23128
rect 7984 23072 8156 23100
rect 7984 23060 7990 23072
rect 7285 23035 7343 23041
rect 7285 23001 7297 23035
rect 7331 23032 7343 23035
rect 9398 23032 9404 23044
rect 7331 23004 9404 23032
rect 7331 23001 7343 23004
rect 7285 22995 7343 23001
rect 9398 22992 9404 23004
rect 9456 22992 9462 23044
rect 10134 22964 10140 22976
rect 6227 22936 6408 22964
rect 10095 22936 10140 22964
rect 6227 22933 6239 22936
rect 6181 22927 6239 22933
rect 10134 22924 10140 22936
rect 10192 22924 10198 22976
rect 10226 22924 10232 22976
rect 10284 22964 10290 22976
rect 10827 22967 10885 22973
rect 10827 22964 10839 22967
rect 10284 22936 10839 22964
rect 10284 22924 10290 22936
rect 10827 22933 10839 22936
rect 10873 22933 10885 22967
rect 10827 22927 10885 22933
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 2866 22760 2872 22772
rect 2827 22732 2872 22760
rect 2866 22720 2872 22732
rect 2924 22720 2930 22772
rect 3510 22760 3516 22772
rect 3471 22732 3516 22760
rect 3510 22720 3516 22732
rect 3568 22760 3574 22772
rect 7745 22763 7803 22769
rect 3568 22732 4200 22760
rect 3568 22720 3574 22732
rect 3878 22556 3884 22568
rect 3839 22528 3884 22556
rect 3878 22516 3884 22528
rect 3936 22516 3942 22568
rect 4172 22565 4200 22732
rect 7745 22729 7757 22763
rect 7791 22760 7803 22763
rect 10134 22760 10140 22772
rect 7791 22732 10140 22760
rect 7791 22729 7803 22732
rect 7745 22723 7803 22729
rect 10134 22720 10140 22732
rect 10192 22720 10198 22772
rect 10686 22760 10692 22772
rect 10647 22732 10692 22760
rect 10686 22720 10692 22732
rect 10744 22720 10750 22772
rect 4801 22695 4859 22701
rect 4801 22661 4813 22695
rect 4847 22692 4859 22695
rect 4847 22664 10364 22692
rect 4847 22661 4859 22664
rect 4801 22655 4859 22661
rect 4338 22624 4344 22636
rect 4299 22596 4344 22624
rect 4338 22584 4344 22596
rect 4396 22584 4402 22636
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22624 4767 22627
rect 5166 22624 5172 22636
rect 4755 22596 5172 22624
rect 4755 22593 4767 22596
rect 4709 22587 4767 22593
rect 5166 22584 5172 22596
rect 5224 22624 5230 22636
rect 5902 22624 5908 22636
rect 5224 22596 5764 22624
rect 5863 22596 5908 22624
rect 5224 22584 5230 22596
rect 4157 22559 4215 22565
rect 4157 22525 4169 22559
rect 4203 22556 4215 22559
rect 5258 22556 5264 22568
rect 4203 22528 4936 22556
rect 5219 22528 5264 22556
rect 4203 22525 4215 22528
rect 4157 22519 4215 22525
rect 2866 22448 2872 22500
rect 2924 22488 2930 22500
rect 4801 22491 4859 22497
rect 4801 22488 4813 22491
rect 2924 22460 4813 22488
rect 2924 22448 2930 22460
rect 4801 22457 4813 22460
rect 4847 22457 4859 22491
rect 4908 22488 4936 22528
rect 5258 22516 5264 22528
rect 5316 22516 5322 22568
rect 5629 22559 5687 22565
rect 5629 22525 5641 22559
rect 5675 22525 5687 22559
rect 5629 22519 5687 22525
rect 5644 22488 5672 22519
rect 4908 22460 5672 22488
rect 5736 22488 5764 22596
rect 5902 22584 5908 22596
rect 5960 22584 5966 22636
rect 9398 22624 9404 22636
rect 9311 22596 9404 22624
rect 9398 22584 9404 22596
rect 9456 22624 9462 22636
rect 10226 22624 10232 22636
rect 9456 22596 10232 22624
rect 9456 22584 9462 22596
rect 10226 22584 10232 22596
rect 10284 22584 10290 22636
rect 6822 22556 6828 22568
rect 6783 22528 6828 22556
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 10336 22556 10364 22664
rect 10908 22559 10966 22565
rect 10908 22556 10920 22559
rect 10336 22528 10920 22556
rect 10908 22525 10920 22528
rect 10954 22556 10966 22559
rect 11333 22559 11391 22565
rect 11333 22556 11345 22559
rect 10954 22528 11345 22556
rect 10954 22525 10966 22528
rect 10908 22519 10966 22525
rect 11333 22525 11345 22528
rect 11379 22556 11391 22559
rect 11514 22556 11520 22568
rect 11379 22528 11520 22556
rect 11379 22525 11391 22528
rect 11333 22519 11391 22525
rect 11514 22516 11520 22528
rect 11572 22516 11578 22568
rect 6273 22491 6331 22497
rect 6273 22488 6285 22491
rect 5736 22460 6285 22488
rect 4801 22451 4859 22457
rect 5184 22432 5212 22460
rect 6273 22457 6285 22460
rect 6319 22488 6331 22491
rect 6546 22488 6552 22500
rect 6319 22460 6552 22488
rect 6319 22457 6331 22460
rect 6273 22451 6331 22457
rect 6546 22448 6552 22460
rect 6604 22488 6610 22500
rect 6641 22491 6699 22497
rect 6641 22488 6653 22491
rect 6604 22460 6653 22488
rect 6604 22448 6610 22460
rect 6641 22457 6653 22460
rect 6687 22488 6699 22491
rect 7187 22491 7245 22497
rect 7187 22488 7199 22491
rect 6687 22460 7199 22488
rect 6687 22457 6699 22460
rect 6641 22451 6699 22457
rect 7187 22457 7199 22460
rect 7233 22488 7245 22491
rect 8478 22488 8484 22500
rect 7233 22460 8484 22488
rect 7233 22457 7245 22460
rect 7187 22451 7245 22457
rect 8478 22448 8484 22460
rect 8536 22448 8542 22500
rect 9493 22491 9551 22497
rect 9493 22457 9505 22491
rect 9539 22488 9551 22491
rect 9766 22488 9772 22500
rect 9539 22460 9772 22488
rect 9539 22457 9551 22460
rect 9493 22451 9551 22457
rect 5077 22423 5135 22429
rect 5077 22389 5089 22423
rect 5123 22420 5135 22423
rect 5166 22420 5172 22432
rect 5123 22392 5172 22420
rect 5123 22389 5135 22392
rect 5077 22383 5135 22389
rect 5166 22380 5172 22392
rect 5224 22380 5230 22432
rect 7926 22380 7932 22432
rect 7984 22420 7990 22432
rect 8113 22423 8171 22429
rect 8113 22420 8125 22423
rect 7984 22392 8125 22420
rect 7984 22380 7990 22392
rect 8113 22389 8125 22392
rect 8159 22389 8171 22423
rect 8113 22383 8171 22389
rect 9217 22423 9275 22429
rect 9217 22389 9229 22423
rect 9263 22420 9275 22423
rect 9508 22420 9536 22451
rect 9766 22448 9772 22460
rect 9824 22448 9830 22500
rect 10045 22491 10103 22497
rect 10045 22457 10057 22491
rect 10091 22488 10103 22491
rect 10226 22488 10232 22500
rect 10091 22460 10232 22488
rect 10091 22457 10103 22460
rect 10045 22451 10103 22457
rect 10226 22448 10232 22460
rect 10284 22448 10290 22500
rect 9263 22392 9536 22420
rect 9263 22389 9275 22392
rect 9217 22383 9275 22389
rect 10778 22380 10784 22432
rect 10836 22420 10842 22432
rect 11011 22423 11069 22429
rect 11011 22420 11023 22423
rect 10836 22392 11023 22420
rect 10836 22380 10842 22392
rect 11011 22389 11023 22392
rect 11057 22389 11069 22423
rect 11011 22383 11069 22389
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 2682 22176 2688 22228
rect 2740 22216 2746 22228
rect 4249 22219 4307 22225
rect 4249 22216 4261 22219
rect 2740 22188 4261 22216
rect 2740 22176 2746 22188
rect 4249 22185 4261 22188
rect 4295 22185 4307 22219
rect 4522 22216 4528 22228
rect 4483 22188 4528 22216
rect 4249 22179 4307 22185
rect 4264 22148 4292 22179
rect 4522 22176 4528 22188
rect 4580 22176 4586 22228
rect 5258 22176 5264 22228
rect 5316 22216 5322 22228
rect 5445 22219 5503 22225
rect 5445 22216 5457 22219
rect 5316 22188 5457 22216
rect 5316 22176 5322 22188
rect 5445 22185 5457 22188
rect 5491 22185 5503 22219
rect 9398 22216 9404 22228
rect 9359 22188 9404 22216
rect 5445 22179 5503 22185
rect 9398 22176 9404 22188
rect 9456 22176 9462 22228
rect 8199 22151 8257 22157
rect 4264 22120 6316 22148
rect 4264 22080 4292 22120
rect 6288 22092 6316 22120
rect 8199 22117 8211 22151
rect 8245 22148 8257 22151
rect 8478 22148 8484 22160
rect 8245 22120 8484 22148
rect 8245 22117 8257 22120
rect 8199 22111 8257 22117
rect 8478 22108 8484 22120
rect 8536 22108 8542 22160
rect 9766 22148 9772 22160
rect 8772 22120 9772 22148
rect 4433 22083 4491 22089
rect 4433 22080 4445 22083
rect 4264 22052 4445 22080
rect 4433 22049 4445 22052
rect 4479 22049 4491 22083
rect 4433 22043 4491 22049
rect 4985 22083 5043 22089
rect 4985 22049 4997 22083
rect 5031 22080 5043 22083
rect 5166 22080 5172 22092
rect 5031 22052 5172 22080
rect 5031 22049 5043 22052
rect 4985 22043 5043 22049
rect 5166 22040 5172 22052
rect 5224 22040 5230 22092
rect 6270 22080 6276 22092
rect 6183 22052 6276 22080
rect 6270 22040 6276 22052
rect 6328 22040 6334 22092
rect 6825 22083 6883 22089
rect 6825 22049 6837 22083
rect 6871 22080 6883 22083
rect 7098 22080 7104 22092
rect 6871 22052 7104 22080
rect 6871 22049 6883 22052
rect 6825 22043 6883 22049
rect 7098 22040 7104 22052
rect 7156 22040 7162 22092
rect 8772 22089 8800 22120
rect 9766 22108 9772 22120
rect 9824 22148 9830 22160
rect 9861 22151 9919 22157
rect 9861 22148 9873 22151
rect 9824 22120 9873 22148
rect 9824 22108 9830 22120
rect 9861 22117 9873 22120
rect 9907 22117 9919 22151
rect 9861 22111 9919 22117
rect 9950 22108 9956 22160
rect 10008 22148 10014 22160
rect 10413 22151 10471 22157
rect 10413 22148 10425 22151
rect 10008 22120 10425 22148
rect 10008 22108 10014 22120
rect 10413 22117 10425 22120
rect 10459 22148 10471 22151
rect 10594 22148 10600 22160
rect 10459 22120 10600 22148
rect 10459 22117 10471 22120
rect 10413 22111 10471 22117
rect 10594 22108 10600 22120
rect 10652 22108 10658 22160
rect 8757 22083 8815 22089
rect 8757 22049 8769 22083
rect 8803 22049 8815 22083
rect 11238 22080 11244 22092
rect 11199 22052 11244 22080
rect 8757 22043 8815 22049
rect 11238 22040 11244 22052
rect 11296 22080 11302 22092
rect 12618 22080 12624 22092
rect 11296 22052 12624 22080
rect 11296 22040 11302 22052
rect 12618 22040 12624 22052
rect 12676 22040 12682 22092
rect 7009 22015 7067 22021
rect 7009 21981 7021 22015
rect 7055 22012 7067 22015
rect 7834 22012 7840 22024
rect 7055 21984 7840 22012
rect 7055 21981 7067 21984
rect 7009 21975 7067 21981
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 9490 21972 9496 22024
rect 9548 22012 9554 22024
rect 9769 22015 9827 22021
rect 9769 22012 9781 22015
rect 9548 21984 9781 22012
rect 9548 21972 9554 21984
rect 9769 21981 9781 21984
rect 9815 22012 9827 22015
rect 10778 22012 10784 22024
rect 9815 21984 10784 22012
rect 9815 21981 9827 21984
rect 9769 21975 9827 21981
rect 10778 21972 10784 21984
rect 10836 21972 10842 22024
rect 3697 21947 3755 21953
rect 3697 21913 3709 21947
rect 3743 21944 3755 21947
rect 3878 21944 3884 21956
rect 3743 21916 3884 21944
rect 3743 21913 3755 21916
rect 3697 21907 3755 21913
rect 3878 21904 3884 21916
rect 3936 21944 3942 21956
rect 5718 21944 5724 21956
rect 3936 21916 5724 21944
rect 3936 21904 3942 21916
rect 5718 21904 5724 21916
rect 5776 21944 5782 21956
rect 6638 21944 6644 21956
rect 5776 21916 6644 21944
rect 5776 21904 5782 21916
rect 6638 21904 6644 21916
rect 6696 21904 6702 21956
rect 8386 21904 8392 21956
rect 8444 21944 8450 21956
rect 11054 21944 11060 21956
rect 8444 21916 11060 21944
rect 8444 21904 8450 21916
rect 11054 21904 11060 21916
rect 11112 21904 11118 21956
rect 5902 21836 5908 21888
rect 5960 21876 5966 21888
rect 6822 21876 6828 21888
rect 5960 21848 6828 21876
rect 5960 21836 5966 21848
rect 6822 21836 6828 21848
rect 6880 21876 6886 21888
rect 7285 21879 7343 21885
rect 7285 21876 7297 21879
rect 6880 21848 7297 21876
rect 6880 21836 6886 21848
rect 7285 21845 7297 21848
rect 7331 21845 7343 21879
rect 10778 21876 10784 21888
rect 10739 21848 10784 21876
rect 7285 21839 7343 21845
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 10870 21836 10876 21888
rect 10928 21876 10934 21888
rect 11379 21879 11437 21885
rect 11379 21876 11391 21879
rect 10928 21848 11391 21876
rect 10928 21836 10934 21848
rect 11379 21845 11391 21848
rect 11425 21845 11437 21879
rect 11379 21839 11437 21845
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 6270 21672 6276 21684
rect 6231 21644 6276 21672
rect 6270 21632 6276 21644
rect 6328 21672 6334 21684
rect 6822 21672 6828 21684
rect 6328 21644 6828 21672
rect 6328 21632 6334 21644
rect 6822 21632 6828 21644
rect 6880 21632 6886 21684
rect 7009 21675 7067 21681
rect 7009 21641 7021 21675
rect 7055 21672 7067 21675
rect 7098 21672 7104 21684
rect 7055 21644 7104 21672
rect 7055 21641 7067 21644
rect 7009 21635 7067 21641
rect 7098 21632 7104 21644
rect 7156 21632 7162 21684
rect 9766 21672 9772 21684
rect 9727 21644 9772 21672
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 4614 21564 4620 21616
rect 4672 21604 4678 21616
rect 10410 21604 10416 21616
rect 4672 21576 10416 21604
rect 4672 21564 4678 21576
rect 10410 21564 10416 21576
rect 10468 21564 10474 21616
rect 10594 21604 10600 21616
rect 10555 21576 10600 21604
rect 10594 21564 10600 21576
rect 10652 21564 10658 21616
rect 5902 21536 5908 21548
rect 5863 21508 5908 21536
rect 5902 21496 5908 21508
rect 5960 21496 5966 21548
rect 10045 21539 10103 21545
rect 10045 21505 10057 21539
rect 10091 21536 10103 21539
rect 10778 21536 10784 21548
rect 10091 21508 10784 21536
rect 10091 21505 10103 21508
rect 10045 21499 10103 21505
rect 10778 21496 10784 21508
rect 10836 21496 10842 21548
rect 1486 21428 1492 21480
rect 1544 21468 1550 21480
rect 3548 21471 3606 21477
rect 3548 21468 3560 21471
rect 1544 21440 3560 21468
rect 1544 21428 1550 21440
rect 3548 21437 3560 21440
rect 3594 21468 3606 21471
rect 3973 21471 4031 21477
rect 3973 21468 3985 21471
rect 3594 21440 3985 21468
rect 3594 21437 3606 21440
rect 3548 21431 3606 21437
rect 3973 21437 3985 21440
rect 4019 21468 4031 21471
rect 4154 21468 4160 21480
rect 4019 21440 4160 21468
rect 4019 21437 4031 21440
rect 3973 21431 4031 21437
rect 4154 21428 4160 21440
rect 4212 21428 4218 21480
rect 4890 21428 4896 21480
rect 4948 21468 4954 21480
rect 5077 21471 5135 21477
rect 5077 21468 5089 21471
rect 4948 21440 5089 21468
rect 4948 21428 4954 21440
rect 5077 21437 5089 21440
rect 5123 21468 5135 21471
rect 5445 21471 5503 21477
rect 5445 21468 5457 21471
rect 5123 21440 5457 21468
rect 5123 21437 5135 21440
rect 5077 21431 5135 21437
rect 5445 21437 5457 21440
rect 5491 21468 5503 21471
rect 5534 21468 5540 21480
rect 5491 21440 5540 21468
rect 5491 21437 5503 21440
rect 5445 21431 5503 21437
rect 5534 21428 5540 21440
rect 5592 21428 5598 21480
rect 5629 21471 5687 21477
rect 5629 21437 5641 21471
rect 5675 21437 5687 21471
rect 5629 21431 5687 21437
rect 4525 21403 4583 21409
rect 4525 21369 4537 21403
rect 4571 21400 4583 21403
rect 5644 21400 5672 21431
rect 6730 21428 6736 21480
rect 6788 21468 6794 21480
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 6788 21440 6837 21468
rect 6788 21428 6794 21440
rect 6825 21437 6837 21440
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 4571 21372 5672 21400
rect 6840 21400 6868 21431
rect 7190 21428 7196 21480
rect 7248 21468 7254 21480
rect 8205 21471 8263 21477
rect 8205 21468 8217 21471
rect 7248 21440 8217 21468
rect 7248 21428 7254 21440
rect 8205 21437 8217 21440
rect 8251 21468 8263 21471
rect 9030 21468 9036 21480
rect 8251 21440 9036 21468
rect 8251 21437 8263 21440
rect 8205 21431 8263 21437
rect 9030 21428 9036 21440
rect 9088 21428 9094 21480
rect 7285 21403 7343 21409
rect 7285 21400 7297 21403
rect 6840 21372 7297 21400
rect 4571 21369 4583 21372
rect 4525 21363 4583 21369
rect 5184 21344 5212 21372
rect 7285 21369 7297 21372
rect 7331 21369 7343 21403
rect 7285 21363 7343 21369
rect 7745 21403 7803 21409
rect 7745 21369 7757 21403
rect 7791 21400 7803 21403
rect 8021 21403 8079 21409
rect 8021 21400 8033 21403
rect 7791 21372 8033 21400
rect 7791 21369 7803 21372
rect 7745 21363 7803 21369
rect 8021 21369 8033 21372
rect 8067 21400 8079 21403
rect 8478 21400 8484 21412
rect 8067 21372 8484 21400
rect 8067 21369 8079 21372
rect 8021 21363 8079 21369
rect 8478 21360 8484 21372
rect 8536 21409 8542 21412
rect 8536 21403 8584 21409
rect 8536 21369 8538 21403
rect 8572 21369 8584 21403
rect 10134 21400 10140 21412
rect 10095 21372 10140 21400
rect 8536 21363 8584 21369
rect 8536 21360 8542 21363
rect 10134 21360 10140 21372
rect 10192 21360 10198 21412
rect 3510 21292 3516 21344
rect 3568 21332 3574 21344
rect 3651 21335 3709 21341
rect 3651 21332 3663 21335
rect 3568 21304 3663 21332
rect 3568 21292 3574 21304
rect 3651 21301 3663 21304
rect 3697 21301 3709 21335
rect 3651 21295 3709 21301
rect 5166 21292 5172 21344
rect 5224 21292 5230 21344
rect 8202 21292 8208 21344
rect 8260 21332 8266 21344
rect 9125 21335 9183 21341
rect 9125 21332 9137 21335
rect 8260 21304 9137 21332
rect 8260 21292 8266 21304
rect 9125 21301 9137 21304
rect 9171 21301 9183 21335
rect 11238 21332 11244 21344
rect 11199 21304 11244 21332
rect 9125 21295 9183 21301
rect 11238 21292 11244 21304
rect 11296 21292 11302 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 3510 21088 3516 21140
rect 3568 21128 3574 21140
rect 3605 21131 3663 21137
rect 3605 21128 3617 21131
rect 3568 21100 3617 21128
rect 3568 21088 3574 21100
rect 3605 21097 3617 21100
rect 3651 21097 3663 21131
rect 7834 21128 7840 21140
rect 7795 21100 7840 21128
rect 3605 21091 3663 21097
rect 7834 21088 7840 21100
rect 7892 21088 7898 21140
rect 9030 21128 9036 21140
rect 8991 21100 9036 21128
rect 9030 21088 9036 21100
rect 9088 21088 9094 21140
rect 9490 21128 9496 21140
rect 9451 21100 9496 21128
rect 9490 21088 9496 21100
rect 9548 21088 9554 21140
rect 10134 21088 10140 21140
rect 10192 21128 10198 21140
rect 10318 21128 10324 21140
rect 10192 21100 10324 21128
rect 10192 21088 10198 21100
rect 10318 21088 10324 21100
rect 10376 21128 10382 21140
rect 10689 21131 10747 21137
rect 10689 21128 10701 21131
rect 10376 21100 10701 21128
rect 10376 21088 10382 21100
rect 10689 21097 10701 21100
rect 10735 21097 10747 21131
rect 10689 21091 10747 21097
rect 10778 21088 10784 21140
rect 10836 21128 10842 21140
rect 11379 21131 11437 21137
rect 11379 21128 11391 21131
rect 10836 21100 11391 21128
rect 10836 21088 10842 21100
rect 11379 21097 11391 21100
rect 11425 21097 11437 21131
rect 11379 21091 11437 21097
rect 4246 21060 4252 21072
rect 4207 21032 4252 21060
rect 4246 21020 4252 21032
rect 4304 21020 4310 21072
rect 6365 21063 6423 21069
rect 6365 21029 6377 21063
rect 6411 21060 6423 21063
rect 7190 21060 7196 21072
rect 6411 21032 7052 21060
rect 7151 21032 7196 21060
rect 6411 21029 6423 21032
rect 6365 21023 6423 21029
rect 6638 20992 6644 21004
rect 6599 20964 6644 20992
rect 6638 20952 6644 20964
rect 6696 20952 6702 21004
rect 7024 21001 7052 21032
rect 7190 21020 7196 21032
rect 7248 21020 7254 21072
rect 8202 21060 8208 21072
rect 8163 21032 8208 21060
rect 8202 21020 8208 21032
rect 8260 21020 8266 21072
rect 9858 21060 9864 21072
rect 9819 21032 9864 21060
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 10413 21063 10471 21069
rect 10413 21029 10425 21063
rect 10459 21060 10471 21063
rect 10594 21060 10600 21072
rect 10459 21032 10600 21060
rect 10459 21029 10471 21032
rect 10413 21023 10471 21029
rect 10594 21020 10600 21032
rect 10652 21020 10658 21072
rect 7009 20995 7067 21001
rect 7009 20961 7021 20995
rect 7055 20992 7067 20995
rect 7098 20992 7104 21004
rect 7055 20964 7104 20992
rect 7055 20961 7067 20964
rect 7009 20955 7067 20961
rect 7098 20952 7104 20964
rect 7156 20952 7162 21004
rect 11054 20952 11060 21004
rect 11112 20992 11118 21004
rect 11276 20995 11334 21001
rect 11276 20992 11288 20995
rect 11112 20964 11288 20992
rect 11112 20952 11118 20964
rect 11276 20961 11288 20964
rect 11322 20961 11334 20995
rect 11276 20955 11334 20961
rect 4154 20884 4160 20936
rect 4212 20924 4218 20936
rect 7561 20927 7619 20933
rect 4212 20896 4257 20924
rect 4212 20884 4218 20896
rect 7561 20893 7573 20927
rect 7607 20924 7619 20927
rect 8110 20924 8116 20936
rect 7607 20896 8116 20924
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 8110 20884 8116 20896
rect 8168 20884 8174 20936
rect 8754 20924 8760 20936
rect 8715 20896 8760 20924
rect 8754 20884 8760 20896
rect 8812 20884 8818 20936
rect 9490 20884 9496 20936
rect 9548 20924 9554 20936
rect 9769 20927 9827 20933
rect 9769 20924 9781 20927
rect 9548 20896 9781 20924
rect 9548 20884 9554 20896
rect 9769 20893 9781 20896
rect 9815 20924 9827 20927
rect 10870 20924 10876 20936
rect 9815 20896 10876 20924
rect 9815 20893 9827 20896
rect 9769 20887 9827 20893
rect 10870 20884 10876 20896
rect 10928 20884 10934 20936
rect 4614 20816 4620 20868
rect 4672 20856 4678 20868
rect 4709 20859 4767 20865
rect 4709 20856 4721 20859
rect 4672 20828 4721 20856
rect 4672 20816 4678 20828
rect 4709 20825 4721 20828
rect 4755 20856 4767 20859
rect 4755 20828 5580 20856
rect 4755 20825 4767 20828
rect 4709 20819 4767 20825
rect 5552 20800 5580 20828
rect 5166 20788 5172 20800
rect 5127 20760 5172 20788
rect 5166 20748 5172 20760
rect 5224 20748 5230 20800
rect 5534 20788 5540 20800
rect 5495 20760 5540 20788
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 4982 20544 4988 20596
rect 5040 20584 5046 20596
rect 5718 20584 5724 20596
rect 5040 20556 5724 20584
rect 5040 20544 5046 20556
rect 5718 20544 5724 20556
rect 5776 20584 5782 20596
rect 6549 20587 6607 20593
rect 6549 20584 6561 20587
rect 5776 20556 6561 20584
rect 5776 20544 5782 20556
rect 6549 20553 6561 20556
rect 6595 20553 6607 20587
rect 6549 20547 6607 20553
rect 7929 20587 7987 20593
rect 7929 20553 7941 20587
rect 7975 20584 7987 20587
rect 8202 20584 8208 20596
rect 7975 20556 8208 20584
rect 7975 20553 7987 20556
rect 7929 20547 7987 20553
rect 2731 20519 2789 20525
rect 2731 20485 2743 20519
rect 2777 20516 2789 20519
rect 4154 20516 4160 20528
rect 2777 20488 4160 20516
rect 2777 20485 2789 20488
rect 2731 20479 2789 20485
rect 4154 20476 4160 20488
rect 4212 20476 4218 20528
rect 3510 20408 3516 20460
rect 3568 20448 3574 20460
rect 3697 20451 3755 20457
rect 3697 20448 3709 20451
rect 3568 20420 3709 20448
rect 3568 20408 3574 20420
rect 3697 20417 3709 20420
rect 3743 20417 3755 20451
rect 3697 20411 3755 20417
rect 5261 20451 5319 20457
rect 5261 20417 5273 20451
rect 5307 20448 5319 20451
rect 5534 20448 5540 20460
rect 5307 20420 5540 20448
rect 5307 20417 5319 20420
rect 5261 20411 5319 20417
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 1394 20340 1400 20392
rect 1452 20380 1458 20392
rect 2660 20383 2718 20389
rect 2660 20380 2672 20383
rect 1452 20352 2672 20380
rect 1452 20340 1458 20352
rect 2660 20349 2672 20352
rect 2706 20380 2718 20383
rect 2774 20380 2780 20392
rect 2706 20352 2780 20380
rect 2706 20349 2718 20352
rect 2660 20343 2718 20349
rect 2774 20340 2780 20352
rect 2832 20380 2838 20392
rect 3053 20383 3111 20389
rect 3053 20380 3065 20383
rect 2832 20352 3065 20380
rect 2832 20340 2838 20352
rect 3053 20349 3065 20352
rect 3099 20349 3111 20383
rect 6564 20380 6592 20547
rect 8202 20544 8208 20556
rect 8260 20584 8266 20596
rect 9677 20587 9735 20593
rect 9677 20584 9689 20587
rect 8260 20556 9689 20584
rect 8260 20544 8266 20556
rect 9677 20553 9689 20556
rect 9723 20584 9735 20587
rect 9858 20584 9864 20596
rect 9723 20556 9864 20584
rect 9723 20553 9735 20556
rect 9677 20547 9735 20553
rect 9858 20544 9864 20556
rect 9916 20544 9922 20596
rect 8754 20408 8760 20460
rect 8812 20448 8818 20460
rect 10226 20448 10232 20460
rect 8812 20420 10232 20448
rect 8812 20408 8818 20420
rect 10226 20408 10232 20420
rect 10284 20448 10290 20460
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 10284 20420 10517 20448
rect 10284 20408 10290 20420
rect 10505 20417 10517 20420
rect 10551 20417 10563 20451
rect 10505 20411 10563 20417
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6564 20352 6837 20380
rect 3053 20343 3111 20349
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 7285 20383 7343 20389
rect 7285 20380 7297 20383
rect 7156 20352 7297 20380
rect 7156 20340 7162 20352
rect 7285 20349 7297 20352
rect 7331 20349 7343 20383
rect 7285 20343 7343 20349
rect 7561 20383 7619 20389
rect 7561 20349 7573 20383
rect 7607 20380 7619 20383
rect 8386 20380 8392 20392
rect 7607 20352 8392 20380
rect 7607 20349 7619 20352
rect 7561 20343 7619 20349
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 3513 20315 3571 20321
rect 3513 20281 3525 20315
rect 3559 20312 3571 20315
rect 3789 20315 3847 20321
rect 3789 20312 3801 20315
rect 3559 20284 3801 20312
rect 3559 20281 3571 20284
rect 3513 20275 3571 20281
rect 3789 20281 3801 20284
rect 3835 20312 3847 20315
rect 4341 20315 4399 20321
rect 3835 20284 4154 20312
rect 3835 20281 3847 20284
rect 3789 20275 3847 20281
rect 4126 20244 4154 20284
rect 4341 20281 4353 20315
rect 4387 20312 4399 20315
rect 4890 20312 4896 20324
rect 4387 20284 4896 20312
rect 4387 20281 4399 20284
rect 4341 20275 4399 20281
rect 4890 20272 4896 20284
rect 4948 20272 4954 20324
rect 5350 20272 5356 20324
rect 5408 20312 5414 20324
rect 5905 20315 5963 20321
rect 5408 20284 5453 20312
rect 5408 20272 5414 20284
rect 5905 20281 5917 20315
rect 5951 20312 5963 20315
rect 6086 20312 6092 20324
rect 5951 20284 6092 20312
rect 5951 20281 5963 20284
rect 5905 20275 5963 20281
rect 6086 20272 6092 20284
rect 6144 20272 6150 20324
rect 8478 20312 8484 20324
rect 8220 20284 8484 20312
rect 4246 20244 4252 20256
rect 4126 20216 4252 20244
rect 4246 20204 4252 20216
rect 4304 20244 4310 20256
rect 4706 20244 4712 20256
rect 4304 20216 4712 20244
rect 4304 20204 4310 20216
rect 4706 20204 4712 20216
rect 4764 20204 4770 20256
rect 5077 20247 5135 20253
rect 5077 20213 5089 20247
rect 5123 20244 5135 20247
rect 5368 20244 5396 20272
rect 8220 20256 8248 20284
rect 8478 20272 8484 20284
rect 8536 20312 8542 20324
rect 8710 20315 8768 20321
rect 8710 20312 8722 20315
rect 8536 20284 8722 20312
rect 8536 20272 8542 20284
rect 8710 20281 8722 20284
rect 8756 20281 8768 20315
rect 10226 20312 10232 20324
rect 10187 20284 10232 20312
rect 8710 20275 8768 20281
rect 10226 20272 10232 20284
rect 10284 20272 10290 20324
rect 10318 20272 10324 20324
rect 10376 20312 10382 20324
rect 10376 20284 10421 20312
rect 10376 20272 10382 20284
rect 5123 20216 5396 20244
rect 6273 20247 6331 20253
rect 5123 20213 5135 20216
rect 5077 20207 5135 20213
rect 6273 20213 6285 20247
rect 6319 20244 6331 20247
rect 6638 20244 6644 20256
rect 6319 20216 6644 20244
rect 6319 20213 6331 20216
rect 6273 20207 6331 20213
rect 6638 20204 6644 20216
rect 6696 20244 6702 20256
rect 7006 20244 7012 20256
rect 6696 20216 7012 20244
rect 6696 20204 6702 20216
rect 7006 20204 7012 20216
rect 7064 20204 7070 20256
rect 8202 20244 8208 20256
rect 8163 20216 8208 20244
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 9309 20247 9367 20253
rect 9309 20213 9321 20247
rect 9355 20244 9367 20247
rect 10336 20244 10364 20272
rect 9355 20216 10364 20244
rect 9355 20213 9367 20216
rect 9309 20207 9367 20213
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 11241 20247 11299 20253
rect 11241 20244 11253 20247
rect 11112 20216 11253 20244
rect 11112 20204 11118 20216
rect 11241 20213 11253 20216
rect 11287 20213 11299 20247
rect 11241 20207 11299 20213
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 3881 20043 3939 20049
rect 3881 20009 3893 20043
rect 3927 20040 3939 20043
rect 4154 20040 4160 20052
rect 3927 20012 4160 20040
rect 3927 20009 3939 20012
rect 3881 20003 3939 20009
rect 4154 20000 4160 20012
rect 4212 20000 4218 20052
rect 4433 20043 4491 20049
rect 4433 20009 4445 20043
rect 4479 20009 4491 20043
rect 4433 20003 4491 20009
rect 3418 19932 3424 19984
rect 3476 19972 3482 19984
rect 4448 19972 4476 20003
rect 4706 20000 4712 20052
rect 4764 20040 4770 20052
rect 4985 20043 5043 20049
rect 4985 20040 4997 20043
rect 4764 20012 4997 20040
rect 4764 20000 4770 20012
rect 4985 20009 4997 20012
rect 5031 20009 5043 20043
rect 4985 20003 5043 20009
rect 5258 20000 5264 20052
rect 5316 20040 5322 20052
rect 6917 20043 6975 20049
rect 5316 20012 6729 20040
rect 5316 20000 5322 20012
rect 3476 19944 4476 19972
rect 3476 19932 3482 19944
rect 4890 19932 4896 19984
rect 4948 19972 4954 19984
rect 5902 19972 5908 19984
rect 4948 19944 5908 19972
rect 4948 19932 4954 19944
rect 5902 19932 5908 19944
rect 5960 19932 5966 19984
rect 5997 19975 6055 19981
rect 5997 19941 6009 19975
rect 6043 19972 6055 19975
rect 6178 19972 6184 19984
rect 6043 19944 6184 19972
rect 6043 19941 6055 19944
rect 5997 19935 6055 19941
rect 6178 19932 6184 19944
rect 6236 19932 6242 19984
rect 6701 19972 6729 20012
rect 6917 20009 6929 20043
rect 6963 20040 6975 20043
rect 7098 20040 7104 20052
rect 6963 20012 7104 20040
rect 6963 20009 6975 20012
rect 6917 20003 6975 20009
rect 7098 20000 7104 20012
rect 7156 20040 7162 20052
rect 7193 20043 7251 20049
rect 7193 20040 7205 20043
rect 7156 20012 7205 20040
rect 7156 20000 7162 20012
rect 7193 20009 7205 20012
rect 7239 20009 7251 20043
rect 7466 20040 7472 20052
rect 7427 20012 7472 20040
rect 7193 20003 7251 20009
rect 7466 20000 7472 20012
rect 7524 20000 7530 20052
rect 8386 20000 8392 20052
rect 8444 20040 8450 20052
rect 8941 20043 8999 20049
rect 8941 20040 8953 20043
rect 8444 20012 8953 20040
rect 8444 20000 8450 20012
rect 8941 20009 8953 20012
rect 8987 20009 8999 20043
rect 9490 20040 9496 20052
rect 9451 20012 9496 20040
rect 8941 20003 8999 20009
rect 9490 20000 9496 20012
rect 9548 20000 9554 20052
rect 9815 20043 9873 20049
rect 9815 20009 9827 20043
rect 9861 20040 9873 20043
rect 10042 20040 10048 20052
rect 9861 20012 10048 20040
rect 9861 20009 9873 20012
rect 9815 20003 9873 20009
rect 10042 20000 10048 20012
rect 10100 20000 10106 20052
rect 10226 20000 10232 20052
rect 10284 20040 10290 20052
rect 10505 20043 10563 20049
rect 10505 20040 10517 20043
rect 10284 20012 10517 20040
rect 10284 20000 10290 20012
rect 10505 20009 10517 20012
rect 10551 20040 10563 20043
rect 10827 20043 10885 20049
rect 10827 20040 10839 20043
rect 10551 20012 10839 20040
rect 10551 20009 10563 20012
rect 10505 20003 10563 20009
rect 10827 20009 10839 20012
rect 10873 20009 10885 20043
rect 10827 20003 10885 20009
rect 8570 19972 8576 19984
rect 6701 19944 8576 19972
rect 8570 19932 8576 19944
rect 8628 19932 8634 19984
rect 2682 19904 2688 19916
rect 2643 19876 2688 19904
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 2958 19904 2964 19916
rect 2919 19876 2964 19904
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 3145 19907 3203 19913
rect 3145 19873 3157 19907
rect 3191 19904 3203 19907
rect 4982 19904 4988 19916
rect 3191 19876 4988 19904
rect 3191 19873 3203 19876
rect 3145 19867 3203 19873
rect 4982 19864 4988 19876
rect 5040 19904 5046 19916
rect 5261 19907 5319 19913
rect 5261 19904 5273 19907
rect 5040 19876 5273 19904
rect 5040 19864 5046 19876
rect 5261 19873 5273 19876
rect 5307 19873 5319 19907
rect 5261 19867 5319 19873
rect 6822 19864 6828 19916
rect 6880 19904 6886 19916
rect 7377 19907 7435 19913
rect 7377 19904 7389 19907
rect 6880 19876 7389 19904
rect 6880 19864 6886 19876
rect 7377 19873 7389 19876
rect 7423 19904 7435 19907
rect 7834 19904 7840 19916
rect 7423 19876 7840 19904
rect 7423 19873 7435 19876
rect 7377 19867 7435 19873
rect 7834 19864 7840 19876
rect 7892 19864 7898 19916
rect 7929 19907 7987 19913
rect 7929 19873 7941 19907
rect 7975 19904 7987 19907
rect 8478 19904 8484 19916
rect 7975 19876 8484 19904
rect 7975 19873 7987 19876
rect 7929 19867 7987 19873
rect 8478 19864 8484 19876
rect 8536 19864 8542 19916
rect 9582 19864 9588 19916
rect 9640 19904 9646 19916
rect 9712 19907 9770 19913
rect 9712 19904 9724 19907
rect 9640 19876 9724 19904
rect 9640 19864 9646 19876
rect 9712 19873 9724 19876
rect 9758 19873 9770 19907
rect 9712 19867 9770 19873
rect 10229 19907 10287 19913
rect 10229 19873 10241 19907
rect 10275 19904 10287 19907
rect 10318 19904 10324 19916
rect 10275 19876 10324 19904
rect 10275 19873 10287 19876
rect 10229 19867 10287 19873
rect 10318 19864 10324 19876
rect 10376 19864 10382 19916
rect 10594 19864 10600 19916
rect 10652 19904 10658 19916
rect 10724 19907 10782 19913
rect 10724 19904 10736 19907
rect 10652 19876 10736 19904
rect 10652 19864 10658 19876
rect 10724 19873 10736 19876
rect 10770 19873 10782 19907
rect 10724 19867 10782 19873
rect 2590 19796 2596 19848
rect 2648 19836 2654 19848
rect 4062 19836 4068 19848
rect 2648 19808 4068 19836
rect 2648 19796 2654 19808
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 6086 19796 6092 19848
rect 6144 19836 6150 19848
rect 6181 19839 6239 19845
rect 6181 19836 6193 19839
rect 6144 19808 6193 19836
rect 6144 19796 6150 19808
rect 6181 19805 6193 19808
rect 6227 19805 6239 19839
rect 6181 19799 6239 19805
rect 3510 19700 3516 19712
rect 3471 19672 3516 19700
rect 3510 19660 3516 19672
rect 3568 19660 3574 19712
rect 8662 19660 8668 19712
rect 8720 19700 8726 19712
rect 10318 19700 10324 19712
rect 8720 19672 10324 19700
rect 8720 19660 8726 19672
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 2682 19456 2688 19508
rect 2740 19496 2746 19508
rect 2961 19499 3019 19505
rect 2961 19496 2973 19499
rect 2740 19468 2973 19496
rect 2740 19456 2746 19468
rect 2961 19465 2973 19468
rect 3007 19496 3019 19499
rect 5258 19496 5264 19508
rect 3007 19468 5264 19496
rect 3007 19465 3019 19468
rect 2961 19459 3019 19465
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 5350 19456 5356 19508
rect 5408 19496 5414 19508
rect 5905 19499 5963 19505
rect 5905 19496 5917 19499
rect 5408 19468 5917 19496
rect 5408 19456 5414 19468
rect 5905 19465 5917 19468
rect 5951 19465 5963 19499
rect 7742 19496 7748 19508
rect 7703 19468 7748 19496
rect 5905 19459 5963 19465
rect 7742 19456 7748 19468
rect 7800 19456 7806 19508
rect 7834 19456 7840 19508
rect 7892 19496 7898 19508
rect 8021 19499 8079 19505
rect 8021 19496 8033 19499
rect 7892 19468 8033 19496
rect 7892 19456 7898 19468
rect 8021 19465 8033 19468
rect 8067 19465 8079 19499
rect 8021 19459 8079 19465
rect 8110 19456 8116 19508
rect 8168 19496 8174 19508
rect 10275 19499 10333 19505
rect 10275 19496 10287 19499
rect 8168 19468 10287 19496
rect 8168 19456 8174 19468
rect 10275 19465 10287 19468
rect 10321 19465 10333 19499
rect 10275 19459 10333 19465
rect 3418 19388 3424 19440
rect 3476 19428 3482 19440
rect 4065 19431 4123 19437
rect 3476 19400 3877 19428
rect 3476 19388 3482 19400
rect 2590 19360 2596 19372
rect 2551 19332 2596 19360
rect 2590 19320 2596 19332
rect 2648 19320 2654 19372
rect 3849 19360 3877 19400
rect 4065 19397 4077 19431
rect 4111 19428 4123 19431
rect 4614 19428 4620 19440
rect 4111 19400 4620 19428
rect 4111 19397 4123 19400
rect 4065 19391 4123 19397
rect 4614 19388 4620 19400
rect 4672 19388 4678 19440
rect 4982 19360 4988 19372
rect 3849 19332 4568 19360
rect 4943 19332 4988 19360
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 1857 19295 1915 19301
rect 1857 19292 1869 19295
rect 1811 19264 1869 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 1857 19261 1869 19264
rect 1903 19261 1915 19295
rect 1857 19255 1915 19261
rect 1872 19224 1900 19255
rect 1946 19252 1952 19304
rect 2004 19292 2010 19304
rect 2317 19295 2375 19301
rect 2317 19292 2329 19295
rect 2004 19264 2329 19292
rect 2004 19252 2010 19264
rect 2317 19261 2329 19264
rect 2363 19261 2375 19295
rect 2317 19255 2375 19261
rect 2958 19224 2964 19236
rect 1872 19196 2964 19224
rect 2958 19184 2964 19196
rect 3016 19224 3022 19236
rect 3237 19227 3295 19233
rect 3237 19224 3249 19227
rect 3016 19196 3249 19224
rect 3016 19184 3022 19196
rect 3237 19193 3249 19196
rect 3283 19193 3295 19227
rect 3510 19224 3516 19236
rect 3471 19196 3516 19224
rect 3237 19187 3295 19193
rect 3510 19184 3516 19196
rect 3568 19184 3574 19236
rect 3602 19184 3608 19236
rect 3660 19224 3666 19236
rect 4540 19233 4568 19332
rect 4982 19320 4988 19332
rect 5040 19320 5046 19372
rect 6086 19320 6092 19372
rect 6144 19360 6150 19372
rect 9582 19360 9588 19372
rect 6144 19332 9588 19360
rect 6144 19320 6150 19332
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 6822 19292 6828 19304
rect 6783 19264 6828 19292
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 8570 19292 8576 19304
rect 8531 19264 8576 19292
rect 8570 19252 8576 19264
rect 8628 19252 8634 19304
rect 9033 19295 9091 19301
rect 9033 19261 9045 19295
rect 9079 19261 9091 19295
rect 10172 19295 10230 19301
rect 10172 19292 10184 19295
rect 9033 19255 9091 19261
rect 9968 19264 10184 19292
rect 4525 19227 4583 19233
rect 3660 19196 3705 19224
rect 3660 19184 3666 19196
rect 4525 19193 4537 19227
rect 4571 19224 4583 19227
rect 4893 19227 4951 19233
rect 4893 19224 4905 19227
rect 4571 19196 4905 19224
rect 4571 19193 4583 19196
rect 4525 19187 4583 19193
rect 4893 19193 4905 19196
rect 4939 19224 4951 19227
rect 5258 19224 5264 19236
rect 4939 19196 5264 19224
rect 4939 19193 4951 19196
rect 4893 19187 4951 19193
rect 5258 19184 5264 19196
rect 5316 19233 5322 19236
rect 5316 19227 5364 19233
rect 5316 19193 5318 19227
rect 5352 19193 5364 19227
rect 5316 19187 5364 19193
rect 7146 19227 7204 19233
rect 7146 19193 7158 19227
rect 7192 19193 7204 19227
rect 9048 19224 9076 19255
rect 7146 19187 7204 19193
rect 8496 19196 9076 19224
rect 5316 19184 5322 19187
rect 6178 19156 6184 19168
rect 6139 19128 6184 19156
rect 6178 19116 6184 19128
rect 6236 19116 6242 19168
rect 6641 19159 6699 19165
rect 6641 19125 6653 19159
rect 6687 19156 6699 19159
rect 7161 19156 7189 19187
rect 8496 19168 8524 19196
rect 7742 19156 7748 19168
rect 6687 19128 7748 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 7742 19116 7748 19128
rect 7800 19156 7806 19168
rect 8202 19156 8208 19168
rect 7800 19128 8208 19156
rect 7800 19116 7806 19128
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 8478 19156 8484 19168
rect 8439 19128 8484 19156
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 8662 19156 8668 19168
rect 8623 19128 8668 19156
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 8754 19116 8760 19168
rect 8812 19156 8818 19168
rect 9968 19165 9996 19264
rect 10172 19261 10184 19264
rect 10218 19261 10230 19295
rect 10172 19255 10230 19261
rect 9953 19159 10011 19165
rect 9953 19156 9965 19159
rect 8812 19128 9965 19156
rect 8812 19116 8818 19128
rect 9953 19125 9965 19128
rect 9999 19125 10011 19159
rect 9953 19119 10011 19125
rect 10594 19116 10600 19168
rect 10652 19156 10658 19168
rect 10689 19159 10747 19165
rect 10689 19156 10701 19159
rect 10652 19128 10701 19156
rect 10652 19116 10658 19128
rect 10689 19125 10701 19128
rect 10735 19125 10747 19159
rect 10689 19119 10747 19125
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 106 18912 112 18964
rect 164 18952 170 18964
rect 1486 18952 1492 18964
rect 164 18924 1492 18952
rect 164 18912 170 18924
rect 1486 18912 1492 18924
rect 1544 18912 1550 18964
rect 2498 18912 2504 18964
rect 2556 18952 2562 18964
rect 3418 18952 3424 18964
rect 2556 18924 3424 18952
rect 2556 18912 2562 18924
rect 3418 18912 3424 18924
rect 3476 18912 3482 18964
rect 4062 18912 4068 18964
rect 4120 18952 4126 18964
rect 4249 18955 4307 18961
rect 4249 18952 4261 18955
rect 4120 18924 4261 18952
rect 4120 18912 4126 18924
rect 4249 18921 4261 18924
rect 4295 18921 4307 18955
rect 4249 18915 4307 18921
rect 5721 18955 5779 18961
rect 5721 18921 5733 18955
rect 5767 18952 5779 18955
rect 6178 18952 6184 18964
rect 5767 18924 6184 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 7742 18952 7748 18964
rect 7703 18924 7748 18952
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 2590 18884 2596 18896
rect 2551 18856 2596 18884
rect 2590 18844 2596 18856
rect 2648 18844 2654 18896
rect 5163 18887 5221 18893
rect 5163 18853 5175 18887
rect 5209 18884 5221 18887
rect 5258 18884 5264 18896
rect 5209 18856 5264 18884
rect 5209 18853 5221 18856
rect 5163 18847 5221 18853
rect 5258 18844 5264 18856
rect 5316 18844 5322 18896
rect 5902 18844 5908 18896
rect 5960 18884 5966 18896
rect 5997 18887 6055 18893
rect 5997 18884 6009 18887
rect 5960 18856 6009 18884
rect 5960 18844 5966 18856
rect 5997 18853 6009 18856
rect 6043 18853 6055 18887
rect 5997 18847 6055 18853
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 1432 18819 1490 18825
rect 1432 18816 1444 18819
rect 1360 18788 1444 18816
rect 1360 18776 1366 18788
rect 1432 18785 1444 18788
rect 1478 18785 1490 18819
rect 1432 18779 1490 18785
rect 3145 18819 3203 18825
rect 3145 18785 3157 18819
rect 3191 18816 3203 18819
rect 4614 18816 4620 18828
rect 3191 18788 4620 18816
rect 3191 18785 3203 18788
rect 3145 18779 3203 18785
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 7377 18819 7435 18825
rect 7377 18785 7389 18819
rect 7423 18816 7435 18819
rect 7466 18816 7472 18828
rect 7423 18788 7472 18816
rect 7423 18785 7435 18788
rect 7377 18779 7435 18785
rect 7466 18776 7472 18788
rect 7524 18776 7530 18828
rect 2498 18748 2504 18760
rect 2459 18720 2504 18748
rect 2498 18708 2504 18720
rect 2556 18708 2562 18760
rect 4062 18748 4068 18760
rect 2792 18720 4068 18748
rect 1535 18683 1593 18689
rect 1535 18649 1547 18683
rect 1581 18680 1593 18683
rect 2792 18680 2820 18720
rect 4062 18708 4068 18720
rect 4120 18748 4126 18760
rect 4709 18751 4767 18757
rect 4709 18748 4721 18751
rect 4120 18720 4721 18748
rect 4120 18708 4126 18720
rect 4709 18717 4721 18720
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18748 4859 18751
rect 5350 18748 5356 18760
rect 4847 18720 5356 18748
rect 4847 18717 4859 18720
rect 4801 18711 4859 18717
rect 5350 18708 5356 18720
rect 5408 18708 5414 18760
rect 1581 18652 2820 18680
rect 1581 18649 1593 18652
rect 1535 18643 1593 18649
rect 3602 18640 3608 18692
rect 3660 18640 3666 18692
rect 1946 18612 1952 18624
rect 1907 18584 1952 18612
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 3513 18615 3571 18621
rect 3513 18581 3525 18615
rect 3559 18612 3571 18615
rect 3620 18612 3648 18640
rect 4246 18612 4252 18624
rect 3559 18584 4252 18612
rect 3559 18581 3571 18584
rect 3513 18575 3571 18581
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 6822 18612 6828 18624
rect 6783 18584 6828 18612
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 7190 18612 7196 18624
rect 7151 18584 7196 18612
rect 7190 18572 7196 18584
rect 7248 18572 7254 18624
rect 8110 18572 8116 18624
rect 8168 18612 8174 18624
rect 8297 18615 8355 18621
rect 8297 18612 8309 18615
rect 8168 18584 8309 18612
rect 8168 18572 8174 18584
rect 8297 18581 8309 18584
rect 8343 18581 8355 18615
rect 8570 18612 8576 18624
rect 8531 18584 8576 18612
rect 8297 18575 8355 18581
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 2314 18368 2320 18420
rect 2372 18408 2378 18420
rect 2409 18411 2467 18417
rect 2409 18408 2421 18411
rect 2372 18380 2421 18408
rect 2372 18368 2378 18380
rect 2409 18377 2421 18380
rect 2455 18377 2467 18411
rect 2409 18371 2467 18377
rect 2590 18368 2596 18420
rect 2648 18408 2654 18420
rect 2777 18411 2835 18417
rect 2777 18408 2789 18411
rect 2648 18380 2789 18408
rect 2648 18368 2654 18380
rect 2777 18377 2789 18380
rect 2823 18408 2835 18411
rect 3697 18411 3755 18417
rect 3697 18408 3709 18411
rect 2823 18380 3709 18408
rect 2823 18377 2835 18380
rect 2777 18371 2835 18377
rect 3697 18377 3709 18380
rect 3743 18408 3755 18411
rect 3789 18411 3847 18417
rect 3789 18408 3801 18411
rect 3743 18380 3801 18408
rect 3743 18377 3755 18380
rect 3697 18371 3755 18377
rect 3789 18377 3801 18380
rect 3835 18377 3847 18411
rect 3789 18371 3847 18377
rect 6641 18411 6699 18417
rect 6641 18377 6653 18411
rect 6687 18408 6699 18411
rect 7466 18408 7472 18420
rect 6687 18380 7472 18408
rect 6687 18377 6699 18380
rect 6641 18371 6699 18377
rect 7466 18368 7472 18380
rect 7524 18368 7530 18420
rect 5721 18343 5779 18349
rect 5721 18309 5733 18343
rect 5767 18340 5779 18343
rect 7650 18340 7656 18352
rect 5767 18312 7656 18340
rect 5767 18309 5779 18312
rect 5721 18303 5779 18309
rect 7650 18300 7656 18312
rect 7708 18300 7714 18352
rect 4062 18272 4068 18284
rect 4023 18244 4068 18272
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18272 4767 18275
rect 4890 18272 4896 18284
rect 4755 18244 4896 18272
rect 4755 18241 4767 18244
rect 4709 18235 4767 18241
rect 4890 18232 4896 18244
rect 4948 18232 4954 18284
rect 8294 18272 8300 18284
rect 5362 18244 8300 18272
rect 2016 18207 2074 18213
rect 2016 18173 2028 18207
rect 2062 18204 2074 18207
rect 2314 18204 2320 18216
rect 2062 18176 2320 18204
rect 2062 18173 2074 18176
rect 2016 18167 2074 18173
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 3012 18207 3070 18213
rect 3012 18204 3024 18207
rect 2424 18176 3024 18204
rect 1394 18096 1400 18148
rect 1452 18136 1458 18148
rect 2424 18136 2452 18176
rect 3012 18173 3024 18176
rect 3058 18204 3070 18207
rect 5362 18204 5390 18244
rect 8294 18232 8300 18244
rect 8352 18232 8358 18284
rect 8662 18272 8668 18284
rect 8623 18244 8668 18272
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 3058 18176 3556 18204
rect 3058 18173 3070 18176
rect 3012 18167 3070 18173
rect 1452 18108 2452 18136
rect 1452 18096 1458 18108
rect 2498 18096 2504 18148
rect 2556 18136 2562 18148
rect 3099 18139 3157 18145
rect 3099 18136 3111 18139
rect 2556 18108 3111 18136
rect 2556 18096 2562 18108
rect 3099 18105 3111 18108
rect 3145 18105 3157 18139
rect 3099 18099 3157 18105
rect 1302 18028 1308 18080
rect 1360 18068 1366 18080
rect 1581 18071 1639 18077
rect 1581 18068 1593 18071
rect 1360 18040 1593 18068
rect 1360 18028 1366 18040
rect 1581 18037 1593 18040
rect 1627 18037 1639 18071
rect 1581 18031 1639 18037
rect 2087 18071 2145 18077
rect 2087 18037 2099 18071
rect 2133 18068 2145 18071
rect 2314 18068 2320 18080
rect 2133 18040 2320 18068
rect 2133 18037 2145 18040
rect 2087 18031 2145 18037
rect 2314 18028 2320 18040
rect 2372 18028 2378 18080
rect 3528 18077 3556 18176
rect 4724 18176 5390 18204
rect 3697 18139 3755 18145
rect 3697 18105 3709 18139
rect 3743 18136 3755 18139
rect 4157 18139 4215 18145
rect 4157 18136 4169 18139
rect 3743 18108 4169 18136
rect 3743 18105 3755 18108
rect 3697 18099 3755 18105
rect 4157 18105 4169 18108
rect 4203 18136 4215 18139
rect 4522 18136 4528 18148
rect 4203 18108 4528 18136
rect 4203 18105 4215 18108
rect 4157 18099 4215 18105
rect 4522 18096 4528 18108
rect 4580 18096 4586 18148
rect 3513 18071 3571 18077
rect 3513 18037 3525 18071
rect 3559 18068 3571 18071
rect 4724 18068 4752 18176
rect 5442 18164 5448 18216
rect 5500 18204 5506 18216
rect 5537 18207 5595 18213
rect 5537 18204 5549 18207
rect 5500 18176 5549 18204
rect 5500 18164 5506 18176
rect 5537 18173 5549 18176
rect 5583 18204 5595 18207
rect 5997 18207 6055 18213
rect 5997 18204 6009 18207
rect 5583 18176 6009 18204
rect 5583 18173 5595 18176
rect 5537 18167 5595 18173
rect 5997 18173 6009 18176
rect 6043 18173 6055 18207
rect 10410 18204 10416 18216
rect 10468 18213 10474 18216
rect 10468 18207 10506 18213
rect 10358 18176 10416 18204
rect 5997 18167 6055 18173
rect 10410 18164 10416 18176
rect 10494 18204 10506 18207
rect 10870 18204 10876 18216
rect 10494 18176 10876 18204
rect 10494 18173 10506 18176
rect 10468 18167 10506 18173
rect 10468 18164 10474 18167
rect 10870 18164 10876 18176
rect 10928 18164 10934 18216
rect 5077 18139 5135 18145
rect 5077 18105 5089 18139
rect 5123 18136 5135 18139
rect 5258 18136 5264 18148
rect 5123 18108 5264 18136
rect 5123 18105 5135 18108
rect 5077 18099 5135 18105
rect 5258 18096 5264 18108
rect 5316 18136 5322 18148
rect 5810 18136 5816 18148
rect 5316 18108 5816 18136
rect 5316 18096 5322 18108
rect 5810 18096 5816 18108
rect 5868 18096 5874 18148
rect 7190 18136 7196 18148
rect 7151 18108 7196 18136
rect 7190 18096 7196 18108
rect 7248 18096 7254 18148
rect 7282 18096 7288 18148
rect 7340 18136 7346 18148
rect 7837 18139 7895 18145
rect 7340 18108 7385 18136
rect 7340 18096 7346 18108
rect 7837 18105 7849 18139
rect 7883 18136 7895 18139
rect 8386 18136 8392 18148
rect 7883 18108 8392 18136
rect 7883 18105 7895 18108
rect 7837 18099 7895 18105
rect 8386 18096 8392 18108
rect 8444 18096 8450 18148
rect 8986 18139 9044 18145
rect 8986 18136 8998 18139
rect 8496 18108 8998 18136
rect 5350 18068 5356 18080
rect 3559 18040 4752 18068
rect 5311 18040 5356 18068
rect 3559 18037 3571 18040
rect 3513 18031 3571 18037
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 7650 18028 7656 18080
rect 7708 18068 7714 18080
rect 8496 18077 8524 18108
rect 8986 18105 8998 18108
rect 9032 18105 9044 18139
rect 8986 18099 9044 18105
rect 8113 18071 8171 18077
rect 8113 18068 8125 18071
rect 7708 18040 8125 18068
rect 7708 18028 7714 18040
rect 8113 18037 8125 18040
rect 8159 18068 8171 18071
rect 8481 18071 8539 18077
rect 8481 18068 8493 18071
rect 8159 18040 8493 18068
rect 8159 18037 8171 18040
rect 8113 18031 8171 18037
rect 8481 18037 8493 18040
rect 8527 18037 8539 18071
rect 9582 18068 9588 18080
rect 9543 18040 9588 18068
rect 8481 18031 8539 18037
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10551 18071 10609 18077
rect 10551 18068 10563 18071
rect 9824 18040 10563 18068
rect 9824 18028 9830 18040
rect 10551 18037 10563 18040
rect 10597 18037 10609 18071
rect 10551 18031 10609 18037
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 2498 17864 2504 17876
rect 2459 17836 2504 17864
rect 2498 17824 2504 17836
rect 2556 17824 2562 17876
rect 3099 17867 3157 17873
rect 3099 17833 3111 17867
rect 3145 17864 3157 17867
rect 3510 17864 3516 17876
rect 3145 17836 3516 17864
rect 3145 17833 3157 17836
rect 3099 17827 3157 17833
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 8662 17824 8668 17876
rect 8720 17864 8726 17876
rect 8757 17867 8815 17873
rect 8757 17864 8769 17867
rect 8720 17836 8769 17864
rect 8720 17824 8726 17836
rect 8757 17833 8769 17836
rect 8803 17833 8815 17867
rect 8757 17827 8815 17833
rect 2314 17756 2320 17808
rect 2372 17796 2378 17808
rect 4154 17796 4160 17808
rect 2372 17768 4160 17796
rect 2372 17756 2378 17768
rect 4154 17756 4160 17768
rect 4212 17756 4218 17808
rect 4246 17756 4252 17808
rect 4304 17796 4310 17808
rect 4801 17799 4859 17805
rect 4304 17768 4349 17796
rect 4304 17756 4310 17768
rect 4801 17765 4813 17799
rect 4847 17796 4859 17799
rect 4890 17796 4896 17808
rect 4847 17768 4896 17796
rect 4847 17765 4859 17768
rect 4801 17759 4859 17765
rect 4890 17756 4896 17768
rect 4948 17756 4954 17808
rect 6086 17796 6092 17808
rect 6047 17768 6092 17796
rect 6086 17756 6092 17768
rect 6144 17756 6150 17808
rect 7650 17756 7656 17808
rect 7708 17796 7714 17808
rect 7882 17799 7940 17805
rect 7882 17796 7894 17799
rect 7708 17768 7894 17796
rect 7708 17756 7714 17768
rect 7882 17765 7894 17768
rect 7928 17765 7940 17799
rect 9766 17796 9772 17808
rect 9727 17768 9772 17796
rect 7882 17759 7940 17765
rect 9766 17756 9772 17768
rect 9824 17756 9830 17808
rect 9858 17756 9864 17808
rect 9916 17796 9922 17808
rect 9916 17768 9961 17796
rect 9916 17756 9922 17768
rect 3028 17731 3086 17737
rect 3028 17697 3040 17731
rect 3074 17728 3086 17731
rect 3234 17728 3240 17740
rect 3074 17700 3240 17728
rect 3074 17697 3086 17700
rect 3028 17691 3086 17697
rect 3234 17688 3240 17700
rect 3292 17688 3298 17740
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 5994 17660 6000 17672
rect 4212 17632 4257 17660
rect 5955 17632 6000 17660
rect 4212 17620 4218 17632
rect 5994 17620 6000 17632
rect 6052 17620 6058 17672
rect 6178 17620 6184 17672
rect 6236 17660 6242 17672
rect 6273 17663 6331 17669
rect 6273 17660 6285 17663
rect 6236 17632 6285 17660
rect 6236 17620 6242 17632
rect 6273 17629 6285 17632
rect 6319 17629 6331 17663
rect 7558 17660 7564 17672
rect 7519 17632 7564 17660
rect 6273 17623 6331 17629
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 10042 17660 10048 17672
rect 8628 17632 10048 17660
rect 8628 17620 8634 17632
rect 10042 17620 10048 17632
rect 10100 17620 10106 17672
rect 3510 17484 3516 17536
rect 3568 17524 3574 17536
rect 5261 17527 5319 17533
rect 5261 17524 5273 17527
rect 3568 17496 5273 17524
rect 3568 17484 3574 17496
rect 5261 17493 5273 17496
rect 5307 17524 5319 17527
rect 5534 17524 5540 17536
rect 5307 17496 5540 17524
rect 5307 17493 5319 17496
rect 5261 17487 5319 17493
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 7193 17527 7251 17533
rect 7193 17493 7205 17527
rect 7239 17524 7251 17527
rect 7282 17524 7288 17536
rect 7239 17496 7288 17524
rect 7239 17493 7251 17496
rect 7193 17487 7251 17493
rect 7282 17484 7288 17496
rect 7340 17524 7346 17536
rect 8110 17524 8116 17536
rect 7340 17496 8116 17524
rect 7340 17484 7346 17496
rect 8110 17484 8116 17496
rect 8168 17484 8174 17536
rect 8202 17484 8208 17536
rect 8260 17524 8266 17536
rect 8481 17527 8539 17533
rect 8481 17524 8493 17527
rect 8260 17496 8493 17524
rect 8260 17484 8266 17496
rect 8481 17493 8493 17496
rect 8527 17524 8539 17527
rect 9858 17524 9864 17536
rect 8527 17496 9864 17524
rect 8527 17493 8539 17496
rect 8481 17487 8539 17493
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 3145 17323 3203 17329
rect 3145 17289 3157 17323
rect 3191 17320 3203 17323
rect 3234 17320 3240 17332
rect 3191 17292 3240 17320
rect 3191 17289 3203 17292
rect 3145 17283 3203 17289
rect 3234 17280 3240 17292
rect 3292 17280 3298 17332
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 4617 17323 4675 17329
rect 4617 17320 4629 17323
rect 4304 17292 4629 17320
rect 4304 17280 4310 17292
rect 4617 17289 4629 17292
rect 4663 17289 4675 17323
rect 4617 17283 4675 17289
rect 6086 17280 6092 17332
rect 6144 17320 6150 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 6144 17292 6561 17320
rect 6144 17280 6150 17292
rect 6549 17289 6561 17292
rect 6595 17289 6607 17323
rect 6549 17283 6607 17289
rect 7469 17323 7527 17329
rect 7469 17289 7481 17323
rect 7515 17320 7527 17323
rect 7834 17320 7840 17332
rect 7515 17292 7840 17320
rect 7515 17289 7527 17292
rect 7469 17283 7527 17289
rect 3510 17184 3516 17196
rect 3471 17156 3516 17184
rect 3510 17144 3516 17156
rect 3568 17184 3574 17196
rect 4341 17187 4399 17193
rect 3568 17156 4108 17184
rect 3568 17144 3574 17156
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 3602 17116 3608 17128
rect 2924 17088 3608 17116
rect 2924 17076 2930 17088
rect 3602 17076 3608 17088
rect 3660 17076 3666 17128
rect 4080 17125 4108 17156
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 5350 17184 5356 17196
rect 4387 17156 5356 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5905 17187 5963 17193
rect 5905 17153 5917 17187
rect 5951 17184 5963 17187
rect 6822 17184 6828 17196
rect 5951 17156 6828 17184
rect 5951 17153 5963 17156
rect 5905 17147 5963 17153
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 4065 17119 4123 17125
rect 4065 17085 4077 17119
rect 4111 17085 4123 17119
rect 4065 17079 4123 17085
rect 4893 17119 4951 17125
rect 4893 17085 4905 17119
rect 4939 17116 4951 17119
rect 5166 17116 5172 17128
rect 4939 17088 5172 17116
rect 4939 17085 4951 17088
rect 4893 17079 4951 17085
rect 5166 17076 5172 17088
rect 5224 17076 5230 17128
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 5629 17119 5687 17125
rect 5629 17116 5641 17119
rect 5592 17088 5641 17116
rect 5592 17076 5598 17088
rect 5629 17085 5641 17088
rect 5675 17085 5687 17119
rect 5629 17079 5687 17085
rect 6984 17119 7042 17125
rect 6984 17085 6996 17119
rect 7030 17116 7042 17119
rect 7484 17116 7512 17283
rect 7834 17280 7840 17292
rect 7892 17320 7898 17332
rect 8018 17320 8024 17332
rect 7892 17292 8024 17320
rect 7892 17280 7898 17292
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 9401 17323 9459 17329
rect 9401 17289 9413 17323
rect 9447 17320 9459 17323
rect 9582 17320 9588 17332
rect 9447 17292 9588 17320
rect 9447 17289 9459 17292
rect 9401 17283 9459 17289
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 10505 17323 10563 17329
rect 10505 17320 10517 17323
rect 9916 17292 10517 17320
rect 9916 17280 9922 17292
rect 10505 17289 10517 17292
rect 10551 17289 10563 17323
rect 11514 17320 11520 17332
rect 11475 17292 11520 17320
rect 10505 17283 10563 17289
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 8570 17252 8576 17264
rect 8531 17224 8576 17252
rect 8570 17212 8576 17224
rect 8628 17212 8634 17264
rect 9490 17212 9496 17264
rect 9548 17212 9554 17264
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 9508 17184 9536 17212
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 8444 17156 9597 17184
rect 8444 17144 8450 17156
rect 9585 17153 9597 17156
rect 9631 17184 9643 17187
rect 10873 17187 10931 17193
rect 10873 17184 10885 17187
rect 9631 17156 10885 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 10873 17153 10885 17156
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 7030 17088 7512 17116
rect 7030 17085 7042 17088
rect 6984 17079 7042 17085
rect 10686 17076 10692 17128
rect 10744 17116 10750 17128
rect 11124 17119 11182 17125
rect 11124 17116 11136 17119
rect 10744 17088 11136 17116
rect 10744 17076 10750 17088
rect 11124 17085 11136 17088
rect 11170 17116 11182 17119
rect 11514 17116 11520 17128
rect 11170 17088 11520 17116
rect 11170 17085 11182 17088
rect 11124 17079 11182 17085
rect 11514 17076 11520 17088
rect 11572 17076 11578 17128
rect 2593 17051 2651 17057
rect 2593 17017 2605 17051
rect 2639 17048 2651 17051
rect 5994 17048 6000 17060
rect 2639 17020 6000 17048
rect 2639 17017 2651 17020
rect 2593 17011 2651 17017
rect 5994 17008 6000 17020
rect 6052 17048 6058 17060
rect 6181 17051 6239 17057
rect 6181 17048 6193 17051
rect 6052 17020 6193 17048
rect 6052 17008 6058 17020
rect 6181 17017 6193 17020
rect 6227 17017 6239 17051
rect 8018 17048 8024 17060
rect 7979 17020 8024 17048
rect 6181 17011 6239 17017
rect 8018 17008 8024 17020
rect 8076 17008 8082 17060
rect 8110 17008 8116 17060
rect 8168 17048 8174 17060
rect 8168 17020 8261 17048
rect 8168 17008 8174 17020
rect 9674 17008 9680 17060
rect 9732 17048 9738 17060
rect 10226 17048 10232 17060
rect 9732 17020 9777 17048
rect 10187 17020 10232 17048
rect 9732 17008 9738 17020
rect 10226 17008 10232 17020
rect 10284 17008 10290 17060
rect 4338 16940 4344 16992
rect 4396 16980 4402 16992
rect 4893 16983 4951 16989
rect 4893 16980 4905 16983
rect 4396 16952 4905 16980
rect 4396 16940 4402 16952
rect 4893 16949 4905 16952
rect 4939 16980 4951 16983
rect 4985 16983 5043 16989
rect 4985 16980 4997 16983
rect 4939 16952 4997 16980
rect 4939 16949 4951 16952
rect 4893 16943 4951 16949
rect 4985 16949 4997 16952
rect 5031 16949 5043 16983
rect 4985 16943 5043 16949
rect 7055 16983 7113 16989
rect 7055 16949 7067 16983
rect 7101 16980 7113 16983
rect 7282 16980 7288 16992
rect 7101 16952 7288 16980
rect 7101 16949 7113 16952
rect 7055 16943 7113 16949
rect 7282 16940 7288 16952
rect 7340 16940 7346 16992
rect 7650 16940 7656 16992
rect 7708 16980 7714 16992
rect 7745 16983 7803 16989
rect 7745 16980 7757 16983
rect 7708 16952 7757 16980
rect 7708 16940 7714 16952
rect 7745 16949 7757 16952
rect 7791 16949 7803 16983
rect 8128 16980 8156 17008
rect 8941 16983 8999 16989
rect 8941 16980 8953 16983
rect 8128 16952 8953 16980
rect 7745 16943 7803 16949
rect 8941 16949 8953 16952
rect 8987 16949 8999 16983
rect 8941 16943 8999 16949
rect 10962 16940 10968 16992
rect 11020 16980 11026 16992
rect 11195 16983 11253 16989
rect 11195 16980 11207 16983
rect 11020 16952 11207 16980
rect 11020 16940 11026 16952
rect 11195 16949 11207 16952
rect 11241 16949 11253 16983
rect 11195 16943 11253 16949
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 3602 16776 3608 16788
rect 3563 16748 3608 16776
rect 3602 16736 3608 16748
rect 3660 16736 3666 16788
rect 4154 16736 4160 16788
rect 4212 16776 4218 16788
rect 4617 16779 4675 16785
rect 4617 16776 4629 16779
rect 4212 16748 4629 16776
rect 4212 16736 4218 16748
rect 4617 16745 4629 16748
rect 4663 16745 4675 16779
rect 4617 16739 4675 16745
rect 5537 16779 5595 16785
rect 5537 16745 5549 16779
rect 5583 16776 5595 16779
rect 5810 16776 5816 16788
rect 5583 16748 5816 16776
rect 5583 16745 5595 16748
rect 5537 16739 5595 16745
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 6086 16776 6092 16788
rect 6047 16748 6092 16776
rect 6086 16736 6092 16748
rect 6144 16736 6150 16788
rect 7055 16779 7113 16785
rect 7055 16745 7067 16779
rect 7101 16776 7113 16779
rect 7190 16776 7196 16788
rect 7101 16748 7196 16776
rect 7101 16745 7113 16748
rect 7055 16739 7113 16745
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 7558 16776 7564 16788
rect 7519 16748 7564 16776
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 8018 16736 8024 16788
rect 8076 16776 8082 16788
rect 8076 16748 9168 16776
rect 8076 16736 8082 16748
rect 3142 16668 3148 16720
rect 3200 16708 3206 16720
rect 4890 16708 4896 16720
rect 3200 16680 4896 16708
rect 3200 16668 3206 16680
rect 4890 16668 4896 16680
rect 4948 16668 4954 16720
rect 7282 16668 7288 16720
rect 7340 16708 7346 16720
rect 8110 16708 8116 16720
rect 7340 16680 8116 16708
rect 7340 16668 7346 16680
rect 8110 16668 8116 16680
rect 8168 16668 8174 16720
rect 8202 16668 8208 16720
rect 8260 16708 8266 16720
rect 9140 16717 9168 16748
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 10137 16779 10195 16785
rect 10137 16776 10149 16779
rect 9824 16748 10149 16776
rect 9824 16736 9830 16748
rect 10137 16745 10149 16748
rect 10183 16745 10195 16779
rect 10137 16739 10195 16745
rect 9125 16711 9183 16717
rect 8260 16680 8305 16708
rect 8260 16668 8266 16680
rect 9125 16677 9137 16711
rect 9171 16708 9183 16711
rect 10962 16708 10968 16720
rect 9171 16680 10968 16708
rect 9171 16677 9183 16680
rect 9125 16671 9183 16677
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 2961 16643 3019 16649
rect 2961 16609 2973 16643
rect 3007 16640 3019 16643
rect 3510 16640 3516 16652
rect 3007 16612 3516 16640
rect 3007 16609 3019 16612
rect 2961 16603 3019 16609
rect 3510 16600 3516 16612
rect 3568 16600 3574 16652
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4706 16640 4712 16652
rect 4203 16612 4712 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 6952 16643 7010 16649
rect 6952 16640 6964 16643
rect 6604 16612 6964 16640
rect 6604 16600 6610 16612
rect 6952 16609 6964 16612
rect 6998 16609 7010 16643
rect 9582 16640 9588 16652
rect 9543 16612 9588 16640
rect 6952 16603 7010 16609
rect 9582 16600 9588 16612
rect 9640 16640 9646 16652
rect 10594 16640 10600 16652
rect 9640 16612 10600 16640
rect 9640 16600 9646 16612
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 10744 16612 10789 16640
rect 10744 16600 10750 16612
rect 5166 16572 5172 16584
rect 5127 16544 5172 16572
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 5994 16532 6000 16584
rect 6052 16572 6058 16584
rect 7926 16572 7932 16584
rect 6052 16544 7932 16572
rect 6052 16532 6058 16544
rect 7926 16532 7932 16544
rect 7984 16532 7990 16584
rect 8386 16572 8392 16584
rect 8347 16544 8392 16572
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 3145 16507 3203 16513
rect 3145 16473 3157 16507
rect 3191 16504 3203 16507
rect 4338 16504 4344 16516
rect 3191 16476 3877 16504
rect 4299 16476 4344 16504
rect 3191 16473 3203 16476
rect 3145 16467 3203 16473
rect 3849 16436 3877 16476
rect 4338 16464 4344 16476
rect 4396 16464 4402 16516
rect 7742 16464 7748 16516
rect 7800 16504 7806 16516
rect 10827 16507 10885 16513
rect 10827 16504 10839 16507
rect 7800 16476 10839 16504
rect 7800 16464 7806 16476
rect 10827 16473 10839 16476
rect 10873 16473 10885 16507
rect 10827 16467 10885 16473
rect 4430 16436 4436 16448
rect 3849 16408 4436 16436
rect 4430 16396 4436 16408
rect 4488 16396 4494 16448
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 9815 16439 9873 16445
rect 9815 16436 9827 16439
rect 9456 16408 9827 16436
rect 9456 16396 9462 16408
rect 9815 16405 9827 16408
rect 9861 16405 9873 16439
rect 9815 16399 9873 16405
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 3053 16235 3111 16241
rect 3053 16201 3065 16235
rect 3099 16232 3111 16235
rect 3510 16232 3516 16244
rect 3099 16204 3516 16232
rect 3099 16201 3111 16204
rect 3053 16195 3111 16201
rect 3510 16192 3516 16204
rect 3568 16192 3574 16244
rect 4246 16192 4252 16244
rect 4304 16232 4310 16244
rect 4433 16235 4491 16241
rect 4433 16232 4445 16235
rect 4304 16204 4445 16232
rect 4304 16192 4310 16204
rect 4433 16201 4445 16204
rect 4479 16201 4491 16235
rect 4433 16195 4491 16201
rect 5445 16235 5503 16241
rect 5445 16201 5457 16235
rect 5491 16232 5503 16235
rect 5718 16232 5724 16244
rect 5491 16204 5724 16232
rect 5491 16201 5503 16204
rect 5445 16195 5503 16201
rect 5718 16192 5724 16204
rect 5776 16192 5782 16244
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 8389 16235 8447 16241
rect 8389 16232 8401 16235
rect 8168 16204 8401 16232
rect 8168 16192 8174 16204
rect 8389 16201 8401 16204
rect 8435 16201 8447 16235
rect 8389 16195 8447 16201
rect 10597 16235 10655 16241
rect 10597 16201 10609 16235
rect 10643 16232 10655 16235
rect 10686 16232 10692 16244
rect 10643 16204 10692 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 5629 16167 5687 16173
rect 5629 16164 5641 16167
rect 4126 16136 5641 16164
rect 2222 16056 2228 16108
rect 2280 16096 2286 16108
rect 4126 16096 4154 16136
rect 5629 16133 5641 16136
rect 5675 16133 5687 16167
rect 5736 16164 5764 16192
rect 10778 16164 10784 16176
rect 5736 16136 10784 16164
rect 5629 16127 5687 16133
rect 10778 16124 10784 16136
rect 10836 16124 10842 16176
rect 10873 16167 10931 16173
rect 10873 16133 10885 16167
rect 10919 16164 10931 16167
rect 15470 16164 15476 16176
rect 10919 16136 15476 16164
rect 10919 16133 10931 16136
rect 10873 16127 10931 16133
rect 15470 16124 15476 16136
rect 15528 16124 15534 16176
rect 2280 16068 4154 16096
rect 2280 16056 2286 16068
rect 4890 16056 4896 16108
rect 4948 16096 4954 16108
rect 6546 16096 6552 16108
rect 4948 16068 6552 16096
rect 4948 16056 4954 16068
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 7558 16096 7564 16108
rect 7519 16068 7564 16096
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 8113 16099 8171 16105
rect 8113 16065 8125 16099
rect 8159 16096 8171 16099
rect 8202 16096 8208 16108
rect 8159 16068 8208 16096
rect 8159 16065 8171 16068
rect 8113 16059 8171 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 9217 16099 9275 16105
rect 9217 16065 9229 16099
rect 9263 16096 9275 16099
rect 9398 16096 9404 16108
rect 9263 16068 9404 16096
rect 9263 16065 9275 16068
rect 9217 16059 9275 16065
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 9490 16056 9496 16108
rect 9548 16096 9554 16108
rect 9548 16068 9593 16096
rect 9548 16056 9554 16068
rect 2685 16031 2743 16037
rect 2685 15997 2697 16031
rect 2731 16028 2743 16031
rect 3510 16028 3516 16040
rect 2731 16000 3516 16028
rect 2731 15997 2743 16000
rect 2685 15991 2743 15997
rect 3510 15988 3516 16000
rect 3568 15988 3574 16040
rect 5261 16031 5319 16037
rect 5261 16028 5273 16031
rect 5092 16000 5273 16028
rect 3834 15963 3892 15969
rect 3834 15960 3846 15963
rect 3344 15932 3846 15960
rect 3344 15904 3372 15932
rect 3834 15929 3846 15932
rect 3880 15929 3892 15963
rect 3834 15923 3892 15929
rect 4614 15920 4620 15972
rect 4672 15960 4678 15972
rect 5092 15969 5120 16000
rect 5261 15997 5273 16000
rect 5307 15997 5319 16031
rect 7006 16028 7012 16040
rect 6967 16000 7012 16028
rect 5261 15991 5319 15997
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 7469 16031 7527 16037
rect 7469 15997 7481 16031
rect 7515 16028 7527 16031
rect 8662 16028 8668 16040
rect 7515 16000 8668 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 5077 15963 5135 15969
rect 5077 15960 5089 15963
rect 4672 15932 5089 15960
rect 4672 15920 4678 15932
rect 5077 15929 5089 15932
rect 5123 15929 5135 15963
rect 5077 15923 5135 15929
rect 5629 15963 5687 15969
rect 5629 15929 5641 15963
rect 5675 15960 5687 15963
rect 6273 15963 6331 15969
rect 6273 15960 6285 15963
rect 5675 15932 6285 15960
rect 5675 15929 5687 15932
rect 5629 15923 5687 15929
rect 6273 15929 6285 15932
rect 6319 15960 6331 15963
rect 7484 15960 7512 15991
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 10502 15988 10508 16040
rect 10560 16028 10566 16040
rect 10689 16031 10747 16037
rect 10689 16028 10701 16031
rect 10560 16000 10701 16028
rect 10560 15988 10566 16000
rect 10689 15997 10701 16000
rect 10735 16028 10747 16031
rect 11241 16031 11299 16037
rect 11241 16028 11253 16031
rect 10735 16000 11253 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 11241 15997 11253 16000
rect 11287 15997 11299 16031
rect 11241 15991 11299 15997
rect 6319 15932 7512 15960
rect 9033 15963 9091 15969
rect 6319 15929 6331 15932
rect 6273 15923 6331 15929
rect 9033 15929 9045 15963
rect 9079 15960 9091 15963
rect 9306 15960 9312 15972
rect 9079 15932 9312 15960
rect 9079 15929 9091 15932
rect 9033 15923 9091 15929
rect 9306 15920 9312 15932
rect 9364 15920 9370 15972
rect 3326 15892 3332 15904
rect 3287 15864 3332 15892
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 4706 15892 4712 15904
rect 4667 15864 4712 15892
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 5810 15892 5816 15904
rect 5723 15864 5816 15892
rect 5810 15852 5816 15864
rect 5868 15892 5874 15904
rect 6178 15892 6184 15904
rect 5868 15864 6184 15892
rect 5868 15852 5874 15864
rect 6178 15852 6184 15864
rect 6236 15852 6242 15904
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 9582 15892 9588 15904
rect 8444 15864 9588 15892
rect 8444 15852 8450 15864
rect 9582 15852 9588 15864
rect 9640 15892 9646 15904
rect 10137 15895 10195 15901
rect 10137 15892 10149 15895
rect 9640 15864 10149 15892
rect 9640 15852 9646 15864
rect 10137 15861 10149 15864
rect 10183 15861 10195 15895
rect 10137 15855 10195 15861
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 2866 15688 2872 15700
rect 2608 15660 2872 15688
rect 2498 15512 2504 15564
rect 2556 15552 2562 15564
rect 2608 15561 2636 15660
rect 2866 15648 2872 15660
rect 2924 15688 2930 15700
rect 2924 15660 3096 15688
rect 2924 15648 2930 15660
rect 2593 15555 2651 15561
rect 2593 15552 2605 15555
rect 2556 15524 2605 15552
rect 2556 15512 2562 15524
rect 2593 15521 2605 15524
rect 2639 15521 2651 15555
rect 2593 15515 2651 15521
rect 2682 15512 2688 15564
rect 2740 15552 2746 15564
rect 2869 15555 2927 15561
rect 2869 15552 2881 15555
rect 2740 15524 2881 15552
rect 2740 15512 2746 15524
rect 2869 15521 2881 15524
rect 2915 15521 2927 15555
rect 3068 15552 3096 15660
rect 3510 15648 3516 15700
rect 3568 15688 3574 15700
rect 4157 15691 4215 15697
rect 4157 15688 4169 15691
rect 3568 15660 4169 15688
rect 3568 15648 3574 15660
rect 4157 15657 4169 15660
rect 4203 15657 4215 15691
rect 5166 15688 5172 15700
rect 5127 15660 5172 15688
rect 4157 15651 4215 15657
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 6178 15648 6184 15700
rect 6236 15688 6242 15700
rect 6273 15691 6331 15697
rect 6273 15688 6285 15691
rect 6236 15660 6285 15688
rect 6236 15648 6242 15660
rect 6273 15657 6285 15660
rect 6319 15657 6331 15691
rect 6273 15651 6331 15657
rect 9217 15691 9275 15697
rect 9217 15657 9229 15691
rect 9263 15688 9275 15691
rect 9398 15688 9404 15700
rect 9263 15660 9404 15688
rect 9263 15657 9275 15660
rect 9217 15651 9275 15657
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 9548 15660 11345 15688
rect 9548 15648 9554 15660
rect 11333 15657 11345 15660
rect 11379 15657 11391 15691
rect 11333 15651 11391 15657
rect 3145 15623 3203 15629
rect 3145 15589 3157 15623
rect 3191 15620 3203 15623
rect 5184 15620 5212 15648
rect 7834 15620 7840 15632
rect 3191 15592 5212 15620
rect 6840 15592 7840 15620
rect 3191 15589 3203 15592
rect 3145 15583 3203 15589
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 3068 15524 4077 15552
rect 2869 15515 2927 15521
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4614 15552 4620 15564
rect 4575 15524 4620 15552
rect 4065 15515 4123 15521
rect 2884 15484 2912 15515
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 6840 15561 6868 15592
rect 7834 15580 7840 15592
rect 7892 15580 7898 15632
rect 9306 15580 9312 15632
rect 9364 15620 9370 15632
rect 9861 15623 9919 15629
rect 9861 15620 9873 15623
rect 9364 15592 9873 15620
rect 9364 15580 9370 15592
rect 9861 15589 9873 15592
rect 9907 15589 9919 15623
rect 9861 15583 9919 15589
rect 6825 15555 6883 15561
rect 6825 15521 6837 15555
rect 6871 15521 6883 15555
rect 6825 15515 6883 15521
rect 8754 15512 8760 15564
rect 8812 15552 8818 15564
rect 9398 15552 9404 15564
rect 8812 15524 9404 15552
rect 8812 15512 8818 15524
rect 9398 15512 9404 15524
rect 9456 15512 9462 15564
rect 10778 15512 10784 15564
rect 10836 15552 10842 15564
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 10836 15524 11253 15552
rect 10836 15512 10842 15524
rect 11241 15521 11253 15524
rect 11287 15552 11299 15555
rect 11330 15552 11336 15564
rect 11287 15524 11336 15552
rect 11287 15521 11299 15524
rect 11241 15515 11299 15521
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 11698 15552 11704 15564
rect 11659 15524 11704 15552
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 5442 15484 5448 15496
rect 2884 15456 5448 15484
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 5902 15484 5908 15496
rect 5863 15456 5908 15484
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 7742 15484 7748 15496
rect 7703 15456 7748 15484
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 7926 15444 7932 15496
rect 7984 15484 7990 15496
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 7984 15456 8033 15484
rect 7984 15444 7990 15456
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 9766 15484 9772 15496
rect 9727 15456 9772 15484
rect 8021 15447 8079 15453
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 10042 15484 10048 15496
rect 10003 15456 10048 15484
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 6914 15376 6920 15428
rect 6972 15416 6978 15428
rect 7469 15419 7527 15425
rect 7469 15416 7481 15419
rect 6972 15388 7481 15416
rect 6972 15376 6978 15388
rect 7469 15385 7481 15388
rect 7515 15385 7527 15419
rect 7469 15379 7527 15385
rect 3510 15308 3516 15360
rect 3568 15348 3574 15360
rect 3605 15351 3663 15357
rect 3605 15348 3617 15351
rect 3568 15320 3617 15348
rect 3568 15308 3574 15320
rect 3605 15317 3617 15320
rect 3651 15317 3663 15351
rect 3605 15311 3663 15317
rect 4338 15308 4344 15360
rect 4396 15348 4402 15360
rect 7006 15348 7012 15360
rect 4396 15320 7012 15348
rect 4396 15308 4402 15320
rect 7006 15308 7012 15320
rect 7064 15348 7070 15360
rect 7101 15351 7159 15357
rect 7101 15348 7113 15351
rect 7064 15320 7113 15348
rect 7064 15308 7070 15320
rect 7101 15317 7113 15320
rect 7147 15317 7159 15351
rect 10686 15348 10692 15360
rect 10647 15320 10692 15348
rect 7101 15311 7159 15317
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 2133 15147 2191 15153
rect 2133 15113 2145 15147
rect 2179 15144 2191 15147
rect 2682 15144 2688 15156
rect 2179 15116 2688 15144
rect 2179 15113 2191 15116
rect 2133 15107 2191 15113
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 2777 15147 2835 15153
rect 2777 15113 2789 15147
rect 2823 15144 2835 15147
rect 4338 15144 4344 15156
rect 2823 15116 4344 15144
rect 2823 15113 2835 15116
rect 2777 15107 2835 15113
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 4522 15144 4528 15156
rect 4483 15116 4528 15144
rect 4522 15104 4528 15116
rect 4580 15104 4586 15156
rect 5537 15147 5595 15153
rect 5537 15113 5549 15147
rect 5583 15144 5595 15147
rect 5626 15144 5632 15156
rect 5583 15116 5632 15144
rect 5583 15113 5595 15116
rect 5537 15107 5595 15113
rect 5626 15104 5632 15116
rect 5684 15144 5690 15156
rect 6457 15147 6515 15153
rect 6457 15144 6469 15147
rect 5684 15116 6469 15144
rect 5684 15104 5690 15116
rect 6457 15113 6469 15116
rect 6503 15113 6515 15147
rect 6457 15107 6515 15113
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 7006 15144 7012 15156
rect 6687 15116 7012 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 7006 15104 7012 15116
rect 7064 15144 7070 15156
rect 7834 15144 7840 15156
rect 7064 15116 7840 15144
rect 7064 15104 7070 15116
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 9306 15144 9312 15156
rect 9267 15116 9312 15144
rect 9306 15104 9312 15116
rect 9364 15144 9370 15156
rect 9677 15147 9735 15153
rect 9677 15144 9689 15147
rect 9364 15116 9689 15144
rect 9364 15104 9370 15116
rect 9677 15113 9689 15116
rect 9723 15113 9735 15147
rect 11330 15144 11336 15156
rect 11291 15116 11336 15144
rect 9677 15107 9735 15113
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 11422 15104 11428 15156
rect 11480 15144 11486 15156
rect 11698 15144 11704 15156
rect 11480 15116 11704 15144
rect 11480 15104 11486 15116
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 2498 15076 2504 15088
rect 2459 15048 2504 15076
rect 2498 15036 2504 15048
rect 2556 15036 2562 15088
rect 3050 15036 3056 15088
rect 3108 15076 3114 15088
rect 7650 15076 7656 15088
rect 3108 15048 7656 15076
rect 3108 15036 3114 15048
rect 7650 15036 7656 15048
rect 7708 15036 7714 15088
rect 10778 15036 10784 15088
rect 10836 15036 10842 15088
rect 6178 15008 6184 15020
rect 4172 14980 6184 15008
rect 2593 14943 2651 14949
rect 2593 14909 2605 14943
rect 2639 14940 2651 14943
rect 2682 14940 2688 14952
rect 2639 14912 2688 14940
rect 2639 14909 2651 14912
rect 2593 14903 2651 14909
rect 2682 14900 2688 14912
rect 2740 14940 2746 14952
rect 3053 14943 3111 14949
rect 3053 14940 3065 14943
rect 2740 14912 3065 14940
rect 2740 14900 2746 14912
rect 3053 14909 3065 14912
rect 3099 14909 3111 14943
rect 3053 14903 3111 14909
rect 3510 14900 3516 14952
rect 3568 14940 3574 14952
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3568 14912 3617 14940
rect 3568 14900 3574 14912
rect 3605 14909 3617 14912
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 3326 14832 3332 14884
rect 3384 14872 3390 14884
rect 3421 14875 3479 14881
rect 3421 14872 3433 14875
rect 3384 14844 3433 14872
rect 3384 14832 3390 14844
rect 3421 14841 3433 14844
rect 3467 14872 3479 14875
rect 3967 14875 4025 14881
rect 3967 14872 3979 14875
rect 3467 14844 3979 14872
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 3967 14841 3979 14844
rect 4013 14872 4025 14875
rect 4172 14872 4200 14980
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 6457 15011 6515 15017
rect 6457 14977 6469 15011
rect 6503 15008 6515 15011
rect 8202 15008 8208 15020
rect 6503 14980 8208 15008
rect 6503 14977 6515 14980
rect 6457 14971 6515 14977
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 8389 15011 8447 15017
rect 8389 14977 8401 15011
rect 8435 15008 8447 15011
rect 8478 15008 8484 15020
rect 8435 14980 8484 15008
rect 8435 14977 8447 14980
rect 8389 14971 8447 14977
rect 8478 14968 8484 14980
rect 8536 15008 8542 15020
rect 9490 15008 9496 15020
rect 8536 14980 9496 15008
rect 8536 14968 8542 14980
rect 9490 14968 9496 14980
rect 9548 14968 9554 15020
rect 10226 14968 10232 15020
rect 10284 15008 10290 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 10284 14980 10517 15008
rect 10284 14968 10290 14980
rect 10505 14977 10517 14980
rect 10551 15008 10563 15011
rect 10796 15008 10824 15036
rect 10551 14980 10824 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 5442 14940 5448 14952
rect 5399 14912 5448 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 7561 14943 7619 14949
rect 7561 14909 7573 14943
rect 7607 14940 7619 14943
rect 7834 14940 7840 14952
rect 7607 14912 7840 14940
rect 7607 14909 7619 14912
rect 7561 14903 7619 14909
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 4013 14844 4200 14872
rect 4013 14841 4025 14844
rect 3967 14835 4025 14841
rect 4246 14832 4252 14884
rect 4304 14872 4310 14884
rect 6914 14872 6920 14884
rect 4304 14844 6920 14872
rect 4304 14832 4310 14844
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 7006 14832 7012 14884
rect 7064 14872 7070 14884
rect 8710 14875 8768 14881
rect 8710 14872 8722 14875
rect 7064 14844 7109 14872
rect 8220 14844 8722 14872
rect 7064 14832 7070 14844
rect 4798 14804 4804 14816
rect 4759 14776 4804 14804
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 5261 14807 5319 14813
rect 5261 14773 5273 14807
rect 5307 14804 5319 14807
rect 5442 14804 5448 14816
rect 5307 14776 5448 14804
rect 5307 14773 5319 14776
rect 5261 14767 5319 14773
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 5997 14807 6055 14813
rect 5997 14773 6009 14807
rect 6043 14804 6055 14807
rect 6178 14804 6184 14816
rect 6043 14776 6184 14804
rect 6043 14773 6055 14776
rect 5997 14767 6055 14773
rect 6178 14764 6184 14776
rect 6236 14804 6242 14816
rect 7558 14804 7564 14816
rect 6236 14776 7564 14804
rect 6236 14764 6242 14776
rect 7558 14764 7564 14776
rect 7616 14804 7622 14816
rect 8220 14813 8248 14844
rect 8710 14841 8722 14844
rect 8756 14872 8768 14875
rect 9858 14872 9864 14884
rect 8756 14844 9864 14872
rect 8756 14841 8768 14844
rect 8710 14835 8768 14841
rect 9858 14832 9864 14844
rect 9916 14832 9922 14884
rect 10042 14832 10048 14884
rect 10100 14872 10106 14884
rect 10226 14872 10232 14884
rect 10100 14844 10232 14872
rect 10100 14832 10106 14844
rect 10226 14832 10232 14844
rect 10284 14832 10290 14884
rect 10321 14875 10379 14881
rect 10321 14841 10333 14875
rect 10367 14872 10379 14875
rect 10686 14872 10692 14884
rect 10367 14844 10692 14872
rect 10367 14841 10379 14844
rect 10321 14835 10379 14841
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 7616 14776 8217 14804
rect 7616 14764 7622 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 3099 14603 3157 14609
rect 3099 14569 3111 14603
rect 3145 14600 3157 14603
rect 4246 14600 4252 14612
rect 3145 14572 4252 14600
rect 3145 14569 3157 14572
rect 3099 14563 3157 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 4341 14603 4399 14609
rect 4341 14569 4353 14603
rect 4387 14600 4399 14603
rect 4798 14600 4804 14612
rect 4387 14572 4804 14600
rect 4387 14569 4399 14572
rect 4341 14563 4399 14569
rect 2498 14492 2504 14544
rect 2556 14532 2562 14544
rect 3605 14535 3663 14541
rect 3605 14532 3617 14535
rect 2556 14504 3617 14532
rect 2556 14492 2562 14504
rect 3605 14501 3617 14504
rect 3651 14532 3663 14535
rect 4062 14532 4068 14544
rect 3651 14504 4068 14532
rect 3651 14501 3663 14504
rect 3605 14495 3663 14501
rect 4062 14492 4068 14504
rect 4120 14532 4126 14544
rect 4356 14532 4384 14563
rect 4798 14560 4804 14572
rect 4856 14560 4862 14612
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 7800 14572 7941 14600
rect 7800 14560 7806 14572
rect 7929 14569 7941 14572
rect 7975 14569 7987 14603
rect 8478 14600 8484 14612
rect 8439 14572 8484 14600
rect 7929 14563 7987 14569
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 10686 14600 10692 14612
rect 10643 14572 10692 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 7098 14532 7104 14544
rect 4120 14504 4384 14532
rect 7059 14504 7104 14532
rect 4120 14492 4126 14504
rect 7098 14492 7104 14504
rect 7156 14492 7162 14544
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 9998 14535 10056 14541
rect 9998 14532 10010 14535
rect 9916 14504 10010 14532
rect 9916 14492 9922 14504
rect 9998 14501 10010 14504
rect 10044 14501 10056 14535
rect 9998 14495 10056 14501
rect 10226 14492 10232 14544
rect 10284 14532 10290 14544
rect 10873 14535 10931 14541
rect 10873 14532 10885 14535
rect 10284 14504 10885 14532
rect 10284 14492 10290 14504
rect 10873 14501 10885 14504
rect 10919 14501 10931 14535
rect 10873 14495 10931 14501
rect 2866 14464 2872 14476
rect 2827 14436 2872 14464
rect 2866 14424 2872 14436
rect 2924 14424 2930 14476
rect 3142 14424 3148 14476
rect 3200 14464 3206 14476
rect 4157 14467 4215 14473
rect 4157 14464 4169 14467
rect 3200 14436 4169 14464
rect 3200 14424 3206 14436
rect 4157 14433 4169 14436
rect 4203 14433 4215 14467
rect 4157 14427 4215 14433
rect 4522 14424 4528 14476
rect 4580 14464 4586 14476
rect 4709 14467 4767 14473
rect 4709 14464 4721 14467
rect 4580 14436 4721 14464
rect 4580 14424 4586 14436
rect 4709 14433 4721 14436
rect 4755 14464 4767 14467
rect 5350 14464 5356 14476
rect 4755 14436 5356 14464
rect 4755 14433 4767 14436
rect 4709 14427 4767 14433
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 5626 14464 5632 14476
rect 5587 14436 5632 14464
rect 5626 14424 5632 14436
rect 5684 14424 5690 14476
rect 8640 14467 8698 14473
rect 8640 14433 8652 14467
rect 8686 14464 8698 14467
rect 8754 14464 8760 14476
rect 8686 14436 8760 14464
rect 8686 14433 8698 14436
rect 8640 14427 8698 14433
rect 8754 14424 8760 14436
rect 8812 14464 8818 14476
rect 9033 14467 9091 14473
rect 9033 14464 9045 14467
rect 8812 14436 9045 14464
rect 8812 14424 8818 14436
rect 9033 14433 9045 14436
rect 9079 14433 9091 14467
rect 9033 14427 9091 14433
rect 11425 14467 11483 14473
rect 11425 14433 11437 14467
rect 11471 14464 11483 14467
rect 11514 14464 11520 14476
rect 11471 14436 11520 14464
rect 11471 14433 11483 14436
rect 11425 14427 11483 14433
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 5810 14396 5816 14408
rect 5771 14368 5816 14396
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 6840 14368 7021 14396
rect 4246 14288 4252 14340
rect 4304 14328 4310 14340
rect 6730 14328 6736 14340
rect 4304 14300 6736 14328
rect 4304 14288 4310 14300
rect 6730 14288 6736 14300
rect 6788 14288 6794 14340
rect 6840 14272 6868 14368
rect 7009 14365 7021 14368
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14396 7711 14399
rect 7926 14396 7932 14408
rect 7699 14368 7932 14396
rect 7699 14365 7711 14368
rect 7653 14359 7711 14365
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 10318 14396 10324 14408
rect 9723 14368 10324 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 8711 14331 8769 14337
rect 8711 14297 8723 14331
rect 8757 14328 8769 14331
rect 8846 14328 8852 14340
rect 8757 14300 8852 14328
rect 8757 14297 8769 14300
rect 8711 14291 8769 14297
rect 8846 14288 8852 14300
rect 8904 14288 8910 14340
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14328 9551 14331
rect 9766 14328 9772 14340
rect 9539 14300 9772 14328
rect 9539 14297 9551 14300
rect 9493 14291 9551 14297
rect 9766 14288 9772 14300
rect 9824 14328 9830 14340
rect 11563 14331 11621 14337
rect 11563 14328 11575 14331
rect 9824 14300 11575 14328
rect 9824 14288 9830 14300
rect 11563 14297 11575 14300
rect 11609 14297 11621 14331
rect 11563 14291 11621 14297
rect 4982 14220 4988 14272
rect 5040 14260 5046 14272
rect 5902 14260 5908 14272
rect 5040 14232 5908 14260
rect 5040 14220 5046 14232
rect 5902 14220 5908 14232
rect 5960 14260 5966 14272
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 5960 14232 6193 14260
rect 5960 14220 5966 14232
rect 6181 14229 6193 14232
rect 6227 14229 6239 14263
rect 6822 14260 6828 14272
rect 6783 14232 6828 14260
rect 6181 14223 6239 14229
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 5077 14059 5135 14065
rect 5077 14056 5089 14059
rect 4488 14028 5089 14056
rect 4488 14016 4494 14028
rect 5077 14025 5089 14028
rect 5123 14056 5135 14059
rect 5166 14056 5172 14068
rect 5123 14028 5172 14056
rect 5123 14025 5135 14028
rect 5077 14019 5135 14025
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 5350 14016 5356 14068
rect 5408 14056 5414 14068
rect 6181 14059 6239 14065
rect 6181 14056 6193 14059
rect 5408 14028 6193 14056
rect 5408 14016 5414 14028
rect 6181 14025 6193 14028
rect 6227 14025 6239 14059
rect 6181 14019 6239 14025
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 9858 14056 9864 14068
rect 9815 14028 9864 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 4126 13960 7027 13988
rect 2866 13880 2872 13932
rect 2924 13920 2930 13932
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 2924 13892 3065 13920
rect 2924 13880 2930 13892
rect 3053 13889 3065 13892
rect 3099 13920 3111 13923
rect 4126 13920 4154 13960
rect 3099 13892 4154 13920
rect 5905 13923 5963 13929
rect 3099 13889 3111 13892
rect 3053 13883 3111 13889
rect 5905 13889 5917 13923
rect 5951 13920 5963 13923
rect 6999 13920 7027 13960
rect 7926 13948 7932 14000
rect 7984 13988 7990 14000
rect 9309 13991 9367 13997
rect 9309 13988 9321 13991
rect 7984 13960 9321 13988
rect 7984 13948 7990 13960
rect 9309 13957 9321 13960
rect 9355 13957 9367 13991
rect 9309 13951 9367 13957
rect 8570 13920 8576 13932
rect 5951 13892 6960 13920
rect 6999 13892 8576 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 3881 13855 3939 13861
rect 3881 13821 3893 13855
rect 3927 13852 3939 13855
rect 4062 13852 4068 13864
rect 3927 13824 4068 13852
rect 3927 13821 3939 13824
rect 3881 13815 3939 13821
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4157 13855 4215 13861
rect 4157 13821 4169 13855
rect 4203 13852 4215 13855
rect 4338 13852 4344 13864
rect 4203 13824 4344 13852
rect 4203 13821 4215 13824
rect 4157 13815 4215 13821
rect 2682 13784 2688 13796
rect 2595 13756 2688 13784
rect 2682 13744 2688 13756
rect 2740 13784 2746 13796
rect 4172 13784 4200 13815
rect 4338 13812 4344 13824
rect 4396 13812 4402 13864
rect 5166 13852 5172 13864
rect 5127 13824 5172 13852
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 5258 13812 5264 13864
rect 5316 13852 5322 13864
rect 5626 13852 5632 13864
rect 5316 13824 5632 13852
rect 5316 13812 5322 13824
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 6932 13861 6960 13892
rect 8570 13880 8576 13892
rect 8628 13880 8634 13932
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13920 8815 13923
rect 8846 13920 8852 13932
rect 8803 13892 8852 13920
rect 8803 13889 8815 13892
rect 8757 13883 8815 13889
rect 8846 13880 8852 13892
rect 8904 13920 8910 13932
rect 8904 13892 9536 13920
rect 8904 13880 8910 13892
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13852 6975 13855
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 6963 13824 8125 13852
rect 6963 13821 6975 13824
rect 6917 13815 6975 13821
rect 8113 13821 8125 13824
rect 8159 13821 8171 13855
rect 8113 13815 8171 13821
rect 9508 13796 9536 13892
rect 9600 13892 10180 13920
rect 2740 13756 4200 13784
rect 7238 13787 7296 13793
rect 2740 13744 2746 13756
rect 7238 13753 7250 13787
rect 7284 13784 7296 13787
rect 7558 13784 7564 13796
rect 7284 13756 7564 13784
rect 7284 13753 7296 13756
rect 7238 13747 7296 13753
rect 3142 13676 3148 13728
rect 3200 13716 3206 13728
rect 3421 13719 3479 13725
rect 3421 13716 3433 13719
rect 3200 13688 3433 13716
rect 3200 13676 3206 13688
rect 3421 13685 3433 13688
rect 3467 13685 3479 13719
rect 3421 13679 3479 13685
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 3697 13719 3755 13725
rect 3697 13716 3709 13719
rect 3568 13688 3709 13716
rect 3568 13676 3574 13688
rect 3697 13685 3709 13688
rect 3743 13685 3755 13719
rect 4706 13716 4712 13728
rect 4667 13688 4712 13716
rect 3697 13679 3755 13685
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 6641 13719 6699 13725
rect 6641 13685 6653 13719
rect 6687 13716 6699 13719
rect 6730 13716 6736 13728
rect 6687 13688 6736 13716
rect 6687 13685 6699 13688
rect 6641 13679 6699 13685
rect 6730 13676 6736 13688
rect 6788 13716 6794 13728
rect 7253 13716 7281 13747
rect 7558 13744 7564 13756
rect 7616 13744 7622 13796
rect 8849 13787 8907 13793
rect 8849 13784 8861 13787
rect 8496 13756 8861 13784
rect 8496 13728 8524 13756
rect 8849 13753 8861 13756
rect 8895 13753 8907 13787
rect 8849 13747 8907 13753
rect 9490 13744 9496 13796
rect 9548 13744 9554 13796
rect 6788 13688 7281 13716
rect 7837 13719 7895 13725
rect 6788 13676 6794 13688
rect 7837 13685 7849 13719
rect 7883 13716 7895 13719
rect 8018 13716 8024 13728
rect 7883 13688 8024 13716
rect 7883 13685 7895 13688
rect 7837 13679 7895 13685
rect 8018 13676 8024 13688
rect 8076 13676 8082 13728
rect 8478 13716 8484 13728
rect 8439 13688 8484 13716
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 8662 13676 8668 13728
rect 8720 13716 8726 13728
rect 9600 13716 9628 13892
rect 10152 13796 10180 13892
rect 10502 13852 10508 13864
rect 10463 13824 10508 13852
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 10781 13855 10839 13861
rect 10781 13821 10793 13855
rect 10827 13852 10839 13855
rect 11422 13852 11428 13864
rect 10827 13824 11428 13852
rect 10827 13821 10839 13824
rect 10781 13815 10839 13821
rect 10134 13784 10140 13796
rect 10047 13756 10140 13784
rect 10134 13744 10140 13756
rect 10192 13784 10198 13796
rect 10796 13784 10824 13815
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 10192 13756 10824 13784
rect 10192 13744 10198 13756
rect 10318 13716 10324 13728
rect 8720 13688 9628 13716
rect 10279 13688 10324 13716
rect 8720 13676 8726 13688
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 11514 13716 11520 13728
rect 11427 13688 11520 13716
rect 11514 13676 11520 13688
rect 11572 13716 11578 13728
rect 13446 13716 13452 13728
rect 11572 13688 13452 13716
rect 11572 13676 11578 13688
rect 13446 13676 13452 13688
rect 13504 13676 13510 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 106 13472 112 13524
rect 164 13512 170 13524
rect 1581 13515 1639 13521
rect 1581 13512 1593 13515
rect 164 13484 1593 13512
rect 164 13472 170 13484
rect 1581 13481 1593 13484
rect 1627 13481 1639 13515
rect 1581 13475 1639 13481
rect 6733 13515 6791 13521
rect 6733 13481 6745 13515
rect 6779 13512 6791 13515
rect 7098 13512 7104 13524
rect 6779 13484 7104 13512
rect 6779 13481 6791 13484
rect 6733 13475 6791 13481
rect 7098 13472 7104 13484
rect 7156 13512 7162 13524
rect 8846 13512 8852 13524
rect 7156 13484 8248 13512
rect 8807 13484 8852 13512
rect 7156 13472 7162 13484
rect 4982 13444 4988 13456
rect 4943 13416 4988 13444
rect 4982 13404 4988 13416
rect 5040 13404 5046 13456
rect 6175 13447 6233 13453
rect 6175 13413 6187 13447
rect 6221 13444 6233 13447
rect 6638 13444 6644 13456
rect 6221 13416 6644 13444
rect 6221 13413 6233 13416
rect 6175 13407 6233 13413
rect 6638 13404 6644 13416
rect 6696 13444 6702 13456
rect 7882 13447 7940 13453
rect 7882 13444 7894 13447
rect 6696 13416 7894 13444
rect 6696 13404 6702 13416
rect 7882 13413 7894 13416
rect 7928 13413 7940 13447
rect 8220 13444 8248 13484
rect 8846 13472 8852 13484
rect 8904 13472 8910 13524
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 10318 13512 10324 13524
rect 9539 13484 10324 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 10318 13472 10324 13484
rect 10376 13472 10382 13524
rect 10502 13472 10508 13524
rect 10560 13512 10566 13524
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10560 13484 10701 13512
rect 10560 13472 10566 13484
rect 10689 13481 10701 13484
rect 10735 13481 10747 13515
rect 10689 13475 10747 13481
rect 9861 13447 9919 13453
rect 9861 13444 9873 13447
rect 8220 13416 9873 13444
rect 7882 13407 7940 13413
rect 9861 13413 9873 13416
rect 9907 13444 9919 13447
rect 10226 13444 10232 13456
rect 9907 13416 10232 13444
rect 9907 13413 9919 13416
rect 9861 13407 9919 13413
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1486 13376 1492 13388
rect 1443 13348 1492 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13376 2927 13379
rect 3050 13376 3056 13388
rect 2915 13348 3056 13376
rect 2915 13345 2927 13348
rect 2869 13339 2927 13345
rect 3050 13336 3056 13348
rect 3108 13336 3114 13388
rect 4249 13379 4307 13385
rect 4249 13345 4261 13379
rect 4295 13345 4307 13379
rect 4249 13339 4307 13345
rect 1946 13268 1952 13320
rect 2004 13308 2010 13320
rect 2682 13308 2688 13320
rect 2004 13280 2688 13308
rect 2004 13268 2010 13280
rect 2682 13268 2688 13280
rect 2740 13308 2746 13320
rect 4264 13308 4292 13339
rect 4706 13336 4712 13388
rect 4764 13376 4770 13388
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 4764 13348 4813 13376
rect 4764 13336 4770 13348
rect 4801 13345 4813 13348
rect 4847 13376 4859 13379
rect 5077 13379 5135 13385
rect 5077 13376 5089 13379
rect 4847 13348 5089 13376
rect 4847 13345 4859 13348
rect 4801 13339 4859 13345
rect 5077 13345 5089 13348
rect 5123 13376 5135 13379
rect 5258 13376 5264 13388
rect 5123 13348 5264 13376
rect 5123 13345 5135 13348
rect 5077 13339 5135 13345
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 5810 13376 5816 13388
rect 5723 13348 5816 13376
rect 5810 13336 5816 13348
rect 5868 13376 5874 13388
rect 7377 13379 7435 13385
rect 7377 13376 7389 13379
rect 5868 13348 7389 13376
rect 5868 13336 5874 13348
rect 7377 13345 7389 13348
rect 7423 13345 7435 13379
rect 7377 13339 7435 13345
rect 7558 13308 7564 13320
rect 2740 13280 4292 13308
rect 7519 13280 7564 13308
rect 2740 13268 2746 13280
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 8864 13280 9781 13308
rect 8864 13252 8892 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 10042 13308 10048 13320
rect 10003 13280 10048 13308
rect 9769 13271 9827 13277
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 3099 13243 3157 13249
rect 3099 13209 3111 13243
rect 3145 13240 3157 13243
rect 8846 13240 8852 13252
rect 3145 13212 8852 13240
rect 3145 13209 3157 13212
rect 3099 13203 3157 13209
rect 8846 13200 8852 13212
rect 8904 13200 8910 13252
rect 3697 13175 3755 13181
rect 3697 13141 3709 13175
rect 3743 13172 3755 13175
rect 4062 13172 4068 13184
rect 3743 13144 4068 13172
rect 3743 13141 3755 13144
rect 3697 13135 3755 13141
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 5077 13175 5135 13181
rect 5077 13141 5089 13175
rect 5123 13172 5135 13175
rect 5353 13175 5411 13181
rect 5353 13172 5365 13175
rect 5123 13144 5365 13172
rect 5123 13141 5135 13144
rect 5077 13135 5135 13141
rect 5353 13141 5365 13144
rect 5399 13172 5411 13175
rect 5718 13172 5724 13184
rect 5399 13144 5724 13172
rect 5399 13141 5411 13144
rect 5353 13135 5411 13141
rect 5718 13132 5724 13144
rect 5776 13132 5782 13184
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 8478 13172 8484 13184
rect 7248 13144 8484 13172
rect 7248 13132 7254 13144
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 1486 12928 1492 12980
rect 1544 12968 1550 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 1544 12940 1593 12968
rect 1544 12928 1550 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 3050 12968 3056 12980
rect 3011 12940 3056 12968
rect 1581 12931 1639 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3418 12968 3424 12980
rect 3379 12940 3424 12968
rect 3418 12928 3424 12940
rect 3476 12968 3482 12980
rect 3743 12971 3801 12977
rect 3743 12968 3755 12971
rect 3476 12940 3755 12968
rect 3476 12928 3482 12940
rect 3743 12937 3755 12940
rect 3789 12937 3801 12971
rect 3743 12931 3801 12937
rect 3970 12928 3976 12980
rect 4028 12928 4034 12980
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 6963 12971 7021 12977
rect 6963 12968 6975 12971
rect 6880 12940 6975 12968
rect 6880 12928 6886 12940
rect 6963 12937 6975 12940
rect 7009 12937 7021 12971
rect 6963 12931 7021 12937
rect 8846 12928 8852 12980
rect 8904 12968 8910 12980
rect 9217 12971 9275 12977
rect 9217 12968 9229 12971
rect 8904 12940 9229 12968
rect 8904 12928 8910 12940
rect 9217 12937 9229 12940
rect 9263 12937 9275 12971
rect 9217 12931 9275 12937
rect 9490 12928 9496 12980
rect 9548 12968 9554 12980
rect 10551 12971 10609 12977
rect 10551 12968 10563 12971
rect 9548 12940 10563 12968
rect 9548 12928 9554 12940
rect 10551 12937 10563 12940
rect 10597 12937 10609 12971
rect 10551 12931 10609 12937
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 3326 12900 3332 12912
rect 2832 12872 3332 12900
rect 2832 12860 2838 12872
rect 3326 12860 3332 12872
rect 3384 12860 3390 12912
rect 3878 12900 3884 12912
rect 3839 12872 3884 12900
rect 3878 12860 3884 12872
rect 3936 12860 3942 12912
rect 3988 12900 4016 12928
rect 10226 12900 10232 12912
rect 3988 12872 6868 12900
rect 3973 12835 4031 12841
rect 3973 12801 3985 12835
rect 4019 12832 4031 12835
rect 4062 12832 4068 12844
rect 4019 12804 4068 12832
rect 4019 12801 4031 12804
rect 3973 12795 4031 12801
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4338 12792 4344 12844
rect 4396 12832 4402 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 4396 12804 6561 12832
rect 4396 12792 4402 12804
rect 5184 12776 5212 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12764 3663 12767
rect 4706 12764 4712 12776
rect 3651 12736 4712 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 5166 12764 5172 12776
rect 5079 12736 5172 12764
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5718 12764 5724 12776
rect 5631 12736 5724 12764
rect 5718 12724 5724 12736
rect 5776 12764 5782 12776
rect 6178 12764 6184 12776
rect 5776 12736 6184 12764
rect 5776 12724 5782 12736
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 6840 12773 6868 12872
rect 7300 12872 9674 12900
rect 10187 12872 10232 12900
rect 7300 12773 7328 12872
rect 7926 12832 7932 12844
rect 7887 12804 7932 12832
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 9646 12832 9674 12872
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 11514 12832 11520 12844
rect 9646 12804 11520 12832
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 6840 12767 6918 12773
rect 6840 12736 6872 12767
rect 6860 12733 6872 12736
rect 6906 12764 6918 12767
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 6906 12736 7297 12764
rect 6906 12733 6918 12736
rect 6860 12727 6918 12733
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12764 8631 12767
rect 8846 12764 8852 12776
rect 8619 12736 8852 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 8846 12724 8852 12736
rect 8904 12724 8910 12776
rect 9398 12764 9404 12776
rect 9456 12773 9462 12776
rect 9456 12767 9494 12773
rect 9346 12736 9404 12764
rect 9398 12724 9404 12736
rect 9482 12764 9494 12767
rect 9861 12767 9919 12773
rect 9861 12764 9873 12767
rect 9482 12736 9873 12764
rect 9482 12733 9494 12736
rect 9456 12727 9494 12733
rect 9861 12733 9873 12736
rect 9907 12733 9919 12767
rect 9861 12727 9919 12733
rect 10480 12767 10538 12773
rect 10480 12733 10492 12767
rect 10526 12764 10538 12767
rect 10870 12764 10876 12776
rect 10526 12736 10876 12764
rect 10526 12733 10538 12736
rect 10480 12727 10538 12733
rect 9456 12724 9462 12727
rect 10870 12724 10876 12736
rect 10928 12764 10934 12776
rect 10928 12736 11008 12764
rect 10928 12724 10934 12736
rect 1578 12656 1584 12708
rect 1636 12696 1642 12708
rect 5077 12699 5135 12705
rect 5077 12696 5089 12699
rect 1636 12668 5089 12696
rect 1636 12656 1642 12668
rect 5077 12665 5089 12668
rect 5123 12696 5135 12699
rect 5736 12696 5764 12724
rect 5123 12668 5764 12696
rect 5905 12699 5963 12705
rect 5123 12665 5135 12668
rect 5077 12659 5135 12665
rect 5905 12665 5917 12699
rect 5951 12696 5963 12699
rect 7558 12696 7564 12708
rect 5951 12668 7564 12696
rect 5951 12665 5963 12668
rect 5905 12659 5963 12665
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 8018 12656 8024 12708
rect 8076 12696 8082 12708
rect 8076 12668 8121 12696
rect 8076 12656 8082 12668
rect 8662 12656 8668 12708
rect 8720 12696 8726 12708
rect 9539 12699 9597 12705
rect 9539 12696 9551 12699
rect 8720 12668 9551 12696
rect 8720 12656 8726 12668
rect 9539 12665 9551 12668
rect 9585 12665 9597 12699
rect 9539 12659 9597 12665
rect 2682 12628 2688 12640
rect 2643 12600 2688 12628
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 4249 12631 4307 12637
rect 4249 12628 4261 12631
rect 3568 12600 4261 12628
rect 3568 12588 3574 12600
rect 4249 12597 4261 12600
rect 4295 12597 4307 12631
rect 4706 12628 4712 12640
rect 4667 12600 4712 12628
rect 4249 12591 4307 12597
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 6273 12631 6331 12637
rect 6273 12597 6285 12631
rect 6319 12628 6331 12631
rect 6730 12628 6736 12640
rect 6319 12600 6736 12628
rect 6319 12597 6331 12600
rect 6273 12591 6331 12597
rect 6730 12588 6736 12600
rect 6788 12628 6794 12640
rect 7653 12631 7711 12637
rect 7653 12628 7665 12631
rect 6788 12600 7665 12628
rect 6788 12588 6794 12600
rect 7653 12597 7665 12600
rect 7699 12597 7711 12631
rect 8036 12628 8064 12656
rect 10980 12640 11008 12736
rect 8849 12631 8907 12637
rect 8849 12628 8861 12631
rect 8036 12600 8861 12628
rect 7653 12591 7711 12597
rect 8849 12597 8861 12600
rect 8895 12597 8907 12631
rect 10962 12628 10968 12640
rect 10923 12600 10968 12628
rect 8849 12591 8907 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 4798 12424 4804 12436
rect 4759 12396 4804 12424
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 7558 12424 7564 12436
rect 7519 12396 7564 12424
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 8757 12427 8815 12433
rect 8757 12424 8769 12427
rect 8076 12396 8769 12424
rect 8076 12384 8082 12396
rect 8757 12393 8769 12396
rect 8803 12393 8815 12427
rect 9766 12424 9772 12436
rect 9727 12396 9772 12424
rect 8757 12387 8815 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 13630 12424 13636 12436
rect 13591 12396 13636 12424
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 3142 12356 3148 12368
rect 3103 12328 3148 12356
rect 3142 12316 3148 12328
rect 3200 12316 3206 12368
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 7926 12356 7932 12368
rect 4120 12328 4568 12356
rect 7887 12328 7932 12356
rect 4120 12316 4126 12328
rect 1670 12248 1676 12300
rect 1728 12288 1734 12300
rect 2590 12288 2596 12300
rect 1728 12260 2596 12288
rect 1728 12248 1734 12260
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 4157 12291 4215 12297
rect 4157 12288 4169 12291
rect 2823 12260 4169 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 4157 12257 4169 12260
rect 4203 12288 4215 12291
rect 4338 12288 4344 12300
rect 4203 12260 4344 12288
rect 4203 12257 4215 12260
rect 4157 12251 4215 12257
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12220 2559 12223
rect 2792 12220 2820 12251
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 2547 12192 2820 12220
rect 3697 12223 3755 12229
rect 2547 12189 2559 12192
rect 2501 12183 2559 12189
rect 3697 12189 3709 12223
rect 3743 12220 3755 12223
rect 3878 12220 3884 12232
rect 3743 12192 3884 12220
rect 3743 12189 3755 12192
rect 3697 12183 3755 12189
rect 3878 12180 3884 12192
rect 3936 12220 3942 12232
rect 4062 12220 4068 12232
rect 3936 12192 4068 12220
rect 3936 12180 3942 12192
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4430 12180 4436 12232
rect 4488 12220 4494 12232
rect 4540 12229 4568 12328
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 8260 12328 9720 12356
rect 8260 12316 8266 12328
rect 9692 12300 9720 12328
rect 5074 12248 5080 12300
rect 5132 12288 5138 12300
rect 5718 12288 5724 12300
rect 5132 12260 5724 12288
rect 5132 12248 5138 12260
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 6178 12288 6184 12300
rect 6139 12260 6184 12288
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 9674 12288 9680 12300
rect 9587 12260 9680 12288
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 13446 12288 13452 12300
rect 13407 12260 13452 12288
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 4488 12192 4537 12220
rect 4488 12180 4494 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4706 12180 4712 12232
rect 4764 12220 4770 12232
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 4764 12192 5181 12220
rect 4764 12180 4770 12192
rect 5169 12189 5181 12192
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 6457 12223 6515 12229
rect 6457 12189 6469 12223
rect 6503 12220 6515 12223
rect 6638 12220 6644 12232
rect 6503 12192 6644 12220
rect 6503 12189 6515 12192
rect 6457 12183 6515 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7834 12220 7840 12232
rect 7747 12192 7840 12220
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12220 8539 12223
rect 8846 12220 8852 12232
rect 8527 12192 8852 12220
rect 8527 12189 8539 12192
rect 8481 12183 8539 12189
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 1854 12112 1860 12164
rect 1912 12152 1918 12164
rect 4798 12152 4804 12164
rect 1912 12124 4804 12152
rect 1912 12112 1918 12124
rect 4798 12112 4804 12124
rect 4856 12112 4862 12164
rect 5537 12155 5595 12161
rect 5537 12152 5549 12155
rect 4908 12124 5549 12152
rect 3970 12044 3976 12096
rect 4028 12084 4034 12096
rect 4295 12087 4353 12093
rect 4295 12084 4307 12087
rect 4028 12056 4307 12084
rect 4028 12044 4034 12056
rect 4295 12053 4307 12056
rect 4341 12053 4353 12087
rect 4295 12047 4353 12053
rect 4433 12087 4491 12093
rect 4433 12053 4445 12087
rect 4479 12084 4491 12087
rect 4614 12084 4620 12096
rect 4479 12056 4620 12084
rect 4479 12053 4491 12056
rect 4433 12047 4491 12053
rect 4614 12044 4620 12056
rect 4672 12084 4678 12096
rect 4908 12084 4936 12124
rect 5537 12121 5549 12124
rect 5583 12121 5595 12155
rect 7852 12152 7880 12180
rect 10042 12152 10048 12164
rect 7852 12124 10048 12152
rect 5537 12115 5595 12121
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 4672 12056 4936 12084
rect 7101 12087 7159 12093
rect 4672 12044 4678 12056
rect 7101 12053 7113 12087
rect 7147 12084 7159 12087
rect 7190 12084 7196 12096
rect 7147 12056 7196 12084
rect 7147 12053 7159 12056
rect 7101 12047 7159 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 9398 12084 9404 12096
rect 7524 12056 9404 12084
rect 7524 12044 7530 12056
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 1670 11880 1676 11892
rect 1631 11852 1676 11880
rect 1670 11840 1676 11852
rect 1728 11840 1734 11892
rect 1949 11883 2007 11889
rect 1949 11849 1961 11883
rect 1995 11880 2007 11883
rect 2222 11880 2228 11892
rect 1995 11852 2228 11880
rect 1995 11849 2007 11852
rect 1949 11843 2007 11849
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 3510 11880 3516 11892
rect 2363 11852 3516 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 1765 11679 1823 11685
rect 1765 11645 1777 11679
rect 1811 11676 1823 11679
rect 2332 11676 2360 11843
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 3881 11883 3939 11889
rect 3881 11849 3893 11883
rect 3927 11880 3939 11883
rect 4249 11883 4307 11889
rect 4249 11880 4261 11883
rect 3927 11852 4261 11880
rect 3927 11849 3939 11852
rect 3881 11843 3939 11849
rect 4249 11849 4261 11852
rect 4295 11880 4307 11883
rect 4430 11880 4436 11892
rect 4295 11852 4436 11880
rect 4295 11849 4307 11852
rect 4249 11843 4307 11849
rect 4430 11840 4436 11852
rect 4488 11840 4494 11892
rect 4798 11880 4804 11892
rect 4759 11852 4804 11880
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 5718 11840 5724 11892
rect 5776 11880 5782 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 5776 11852 6469 11880
rect 5776 11840 5782 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 8665 11883 8723 11889
rect 8665 11880 8677 11883
rect 6788 11852 8677 11880
rect 6788 11840 6794 11852
rect 8665 11849 8677 11852
rect 8711 11849 8723 11883
rect 8665 11843 8723 11849
rect 2498 11772 2504 11824
rect 2556 11812 2562 11824
rect 2685 11815 2743 11821
rect 2685 11812 2697 11815
rect 2556 11784 2697 11812
rect 2556 11772 2562 11784
rect 2685 11781 2697 11784
rect 2731 11812 2743 11815
rect 3418 11812 3424 11824
rect 2731 11784 3424 11812
rect 2731 11781 2743 11784
rect 2685 11775 2743 11781
rect 3418 11772 3424 11784
rect 3476 11772 3482 11824
rect 3436 11685 3464 11772
rect 4448 11744 4476 11840
rect 4614 11812 4620 11824
rect 4575 11784 4620 11812
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 7653 11815 7711 11821
rect 7653 11781 7665 11815
rect 7699 11812 7711 11815
rect 7834 11812 7840 11824
rect 7699 11784 7840 11812
rect 7699 11781 7711 11784
rect 7653 11775 7711 11781
rect 7834 11772 7840 11784
rect 7892 11772 7898 11824
rect 8680 11812 8708 11843
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 10045 11883 10103 11889
rect 10045 11880 10057 11883
rect 9732 11852 10057 11880
rect 9732 11840 9738 11852
rect 10045 11849 10057 11852
rect 10091 11849 10103 11883
rect 10045 11843 10103 11849
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 10192 11852 10425 11880
rect 10192 11840 10198 11852
rect 10413 11849 10425 11852
rect 10459 11849 10471 11883
rect 13446 11880 13452 11892
rect 13407 11852 13452 11880
rect 10413 11843 10471 11849
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 8680 11784 8800 11812
rect 4709 11747 4767 11753
rect 4709 11744 4721 11747
rect 4448 11716 4721 11744
rect 4709 11713 4721 11716
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 8662 11744 8668 11756
rect 7147 11716 8668 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 1811 11648 2360 11676
rect 3421 11679 3479 11685
rect 1811 11645 1823 11648
rect 1765 11639 1823 11645
rect 3421 11645 3433 11679
rect 3467 11645 3479 11679
rect 3421 11639 3479 11645
rect 3513 11679 3571 11685
rect 3513 11645 3525 11679
rect 3559 11676 3571 11679
rect 3970 11676 3976 11688
rect 3559 11648 3976 11676
rect 3559 11645 3571 11648
rect 3513 11639 3571 11645
rect 3970 11636 3976 11648
rect 4028 11676 4034 11688
rect 4488 11679 4546 11685
rect 4488 11676 4500 11679
rect 4028 11648 4500 11676
rect 4028 11636 4034 11648
rect 4488 11645 4500 11648
rect 4534 11676 4546 11679
rect 5445 11679 5503 11685
rect 5445 11676 5457 11679
rect 4534 11648 5457 11676
rect 4534 11645 4546 11648
rect 4488 11639 4546 11645
rect 5445 11645 5457 11648
rect 5491 11676 5503 11679
rect 5721 11679 5779 11685
rect 5721 11676 5733 11679
rect 5491 11648 5733 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 5721 11645 5733 11648
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 4341 11611 4399 11617
rect 4341 11577 4353 11611
rect 4387 11608 4399 11611
rect 4706 11608 4712 11620
rect 4387 11580 4712 11608
rect 4387 11577 4399 11580
rect 4341 11571 4399 11577
rect 4706 11568 4712 11580
rect 4764 11568 4770 11620
rect 7190 11608 7196 11620
rect 7151 11580 7196 11608
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 8772 11608 8800 11784
rect 8849 11747 8907 11753
rect 8849 11713 8861 11747
rect 8895 11744 8907 11747
rect 8938 11744 8944 11756
rect 8895 11716 8944 11744
rect 8895 11713 8907 11716
rect 8849 11707 8907 11713
rect 8938 11704 8944 11716
rect 8996 11744 9002 11756
rect 9766 11744 9772 11756
rect 8996 11716 9772 11744
rect 8996 11704 9002 11716
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 9170 11611 9228 11617
rect 9170 11608 9182 11611
rect 8772 11580 9182 11608
rect 9170 11577 9182 11580
rect 9216 11577 9228 11611
rect 9170 11571 9228 11577
rect 6178 11540 6184 11552
rect 6139 11512 6184 11540
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 7926 11540 7932 11552
rect 7616 11512 7932 11540
rect 7616 11500 7622 11512
rect 7926 11500 7932 11512
rect 7984 11540 7990 11552
rect 8021 11543 8079 11549
rect 8021 11540 8033 11543
rect 7984 11512 8033 11540
rect 7984 11500 7990 11512
rect 8021 11509 8033 11512
rect 8067 11509 8079 11543
rect 9766 11540 9772 11552
rect 9727 11512 9772 11540
rect 8021 11503 8079 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10594 11540 10600 11552
rect 10555 11512 10600 11540
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 1728 11308 4537 11336
rect 1728 11296 1734 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 4525 11299 4583 11305
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 4672 11308 5457 11336
rect 4672 11296 4678 11308
rect 5445 11305 5457 11308
rect 5491 11305 5503 11339
rect 7558 11336 7564 11348
rect 7519 11308 7564 11336
rect 5445 11299 5503 11305
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 7929 11339 7987 11345
rect 7929 11305 7941 11339
rect 7975 11336 7987 11339
rect 8662 11336 8668 11348
rect 7975 11308 8668 11336
rect 7975 11305 7987 11308
rect 7929 11299 7987 11305
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 8938 11336 8944 11348
rect 8899 11308 8944 11336
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 1949 11271 2007 11277
rect 1949 11237 1961 11271
rect 1995 11268 2007 11271
rect 4798 11268 4804 11280
rect 1995 11240 4804 11268
rect 1995 11237 2007 11240
rect 1949 11231 2007 11237
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1964 11200 1992 11231
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 6730 11228 6736 11280
rect 6788 11268 6794 11280
rect 6962 11271 7020 11277
rect 6962 11268 6974 11271
rect 6788 11240 6974 11268
rect 6788 11228 6794 11240
rect 6962 11237 6974 11240
rect 7008 11237 7020 11271
rect 6962 11231 7020 11237
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 8205 11271 8263 11277
rect 8205 11268 8217 11271
rect 7892 11240 8217 11268
rect 7892 11228 7898 11240
rect 8205 11237 8217 11240
rect 8251 11237 8263 11271
rect 8205 11231 8263 11237
rect 9766 11228 9772 11280
rect 9824 11268 9830 11280
rect 9861 11271 9919 11277
rect 9861 11268 9873 11271
rect 9824 11240 9873 11268
rect 9824 11228 9830 11240
rect 9861 11237 9873 11240
rect 9907 11237 9919 11271
rect 9861 11231 9919 11237
rect 10413 11271 10471 11277
rect 10413 11237 10425 11271
rect 10459 11268 10471 11271
rect 10778 11268 10784 11280
rect 10459 11240 10784 11268
rect 10459 11237 10471 11240
rect 10413 11231 10471 11237
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 1443 11172 1992 11200
rect 2409 11203 2467 11209
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 2409 11169 2421 11203
rect 2455 11200 2467 11203
rect 2498 11200 2504 11212
rect 2455 11172 2504 11200
rect 2455 11169 2467 11172
rect 2409 11163 2467 11169
rect 2498 11160 2504 11172
rect 2556 11160 2562 11212
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11169 2743 11203
rect 2685 11163 2743 11169
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2700 11132 2728 11163
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 4028 11172 4077 11200
rect 4028 11160 4034 11172
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 4295 11203 4353 11209
rect 4295 11169 4307 11203
rect 4341 11169 4353 11203
rect 5626 11200 5632 11212
rect 5587 11172 5632 11200
rect 4295 11163 4353 11169
rect 2958 11132 2964 11144
rect 2280 11104 2728 11132
rect 2919 11104 2964 11132
rect 2280 11092 2286 11104
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 2317 11067 2375 11073
rect 2317 11033 2329 11067
rect 2363 11064 2375 11067
rect 2501 11067 2559 11073
rect 2501 11064 2513 11067
rect 2363 11036 2513 11064
rect 2363 11033 2375 11036
rect 2317 11027 2375 11033
rect 2501 11033 2513 11036
rect 2547 11064 2559 11067
rect 3050 11064 3056 11076
rect 2547 11036 3056 11064
rect 2547 11033 2559 11036
rect 2501 11027 2559 11033
rect 3050 11024 3056 11036
rect 3108 11024 3114 11076
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4157 11067 4215 11073
rect 4157 11064 4169 11067
rect 4120 11036 4169 11064
rect 4120 11024 4126 11036
rect 4157 11033 4169 11036
rect 4203 11033 4215 11067
rect 4310 11064 4338 11163
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 6638 11200 6644 11212
rect 6599 11172 6644 11200
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 8386 11132 8392 11144
rect 8347 11104 8392 11132
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 10594 11132 10600 11144
rect 9815 11104 10600 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 4430 11064 4436 11076
rect 4310 11036 4436 11064
rect 4157 11027 4215 11033
rect 4430 11024 4436 11036
rect 4488 11064 4494 11076
rect 5074 11064 5080 11076
rect 4488 11036 5080 11064
rect 4488 11024 4494 11036
rect 5074 11024 5080 11036
rect 5132 11064 5138 11076
rect 5813 11067 5871 11073
rect 5813 11064 5825 11067
rect 5132 11036 5825 11064
rect 5132 11024 5138 11036
rect 5813 11033 5825 11036
rect 5859 11033 5871 11067
rect 5813 11027 5871 11033
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 9784 11064 9812 11095
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 9732 11036 9812 11064
rect 9732 11024 9738 11036
rect 3513 10999 3571 11005
rect 3513 10965 3525 10999
rect 3559 10996 3571 10999
rect 3789 10999 3847 11005
rect 3789 10996 3801 10999
rect 3559 10968 3801 10996
rect 3559 10965 3571 10968
rect 3513 10959 3571 10965
rect 3789 10965 3801 10968
rect 3835 10996 3847 10999
rect 4338 10996 4344 11008
rect 3835 10968 4344 10996
rect 3835 10965 3847 10968
rect 3789 10959 3847 10965
rect 4338 10956 4344 10968
rect 4396 10956 4402 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 1670 10792 1676 10804
rect 1631 10764 1676 10792
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 2498 10792 2504 10804
rect 2459 10764 2504 10792
rect 2498 10752 2504 10764
rect 2556 10792 2562 10804
rect 4157 10795 4215 10801
rect 4157 10792 4169 10795
rect 2556 10764 4169 10792
rect 2556 10752 2562 10764
rect 4157 10761 4169 10764
rect 4203 10792 4215 10795
rect 4430 10792 4436 10804
rect 4203 10764 4436 10792
rect 4203 10761 4215 10764
rect 4157 10755 4215 10761
rect 4430 10752 4436 10764
rect 4488 10801 4494 10804
rect 4488 10795 4537 10801
rect 4488 10761 4491 10795
rect 4525 10761 4537 10795
rect 4798 10792 4804 10804
rect 4759 10764 4804 10792
rect 4488 10755 4537 10761
rect 4488 10752 4494 10755
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 8386 10752 8392 10804
rect 8444 10792 8450 10804
rect 8481 10795 8539 10801
rect 8481 10792 8493 10795
rect 8444 10764 8493 10792
rect 8444 10752 8450 10764
rect 8481 10761 8493 10764
rect 8527 10761 8539 10795
rect 9674 10792 9680 10804
rect 9635 10764 9680 10792
rect 8481 10755 8539 10761
rect 4062 10724 4068 10736
rect 3804 10696 4068 10724
rect 3804 10665 3832 10696
rect 4062 10684 4068 10696
rect 4120 10724 4126 10736
rect 4617 10727 4675 10733
rect 4617 10724 4629 10727
rect 4120 10696 4629 10724
rect 4120 10684 4126 10696
rect 4617 10693 4629 10696
rect 4663 10724 4675 10727
rect 4982 10724 4988 10736
rect 4663 10696 4988 10724
rect 4663 10693 4675 10696
rect 4617 10687 4675 10693
rect 4982 10684 4988 10696
rect 5040 10724 5046 10736
rect 5353 10727 5411 10733
rect 5353 10724 5365 10727
rect 5040 10696 5365 10724
rect 5040 10684 5046 10696
rect 5353 10693 5365 10696
rect 5399 10693 5411 10727
rect 5353 10687 5411 10693
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 2884 10628 3801 10656
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1728 10560 1777 10588
rect 1728 10548 1734 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 2884 10597 2912 10628
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10656 4767 10659
rect 5074 10656 5080 10668
rect 4755 10628 5080 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 5074 10616 5080 10628
rect 5132 10656 5138 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5132 10628 5733 10656
rect 5132 10616 5138 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 8496 10656 8524 10755
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 9824 10764 10057 10792
rect 9824 10752 9830 10764
rect 10045 10761 10057 10764
rect 10091 10761 10103 10795
rect 10045 10755 10103 10761
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 8496 10628 8769 10656
rect 5721 10619 5779 10625
rect 8757 10625 8769 10628
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 9033 10659 9091 10665
rect 9033 10656 9045 10659
rect 8904 10628 9045 10656
rect 8904 10616 8910 10628
rect 9033 10625 9045 10628
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 2869 10591 2927 10597
rect 2869 10588 2881 10591
rect 2832 10560 2881 10588
rect 2832 10548 2838 10560
rect 2869 10557 2881 10560
rect 2915 10557 2927 10591
rect 2869 10551 2927 10557
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 3513 10591 3571 10597
rect 3513 10588 3525 10591
rect 3108 10560 3525 10588
rect 3108 10548 3114 10560
rect 3513 10557 3525 10560
rect 3559 10588 3571 10591
rect 4614 10588 4620 10600
rect 3559 10560 4620 10588
rect 3559 10557 3571 10560
rect 3513 10551 3571 10557
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 6914 10588 6920 10600
rect 6875 10560 6920 10588
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 4338 10480 4344 10532
rect 4396 10520 4402 10532
rect 4396 10492 4441 10520
rect 4396 10480 4402 10492
rect 4522 10480 4528 10532
rect 4580 10520 4586 10532
rect 4798 10520 4804 10532
rect 4580 10492 4804 10520
rect 4580 10480 4586 10492
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 7238 10523 7296 10529
rect 7238 10489 7250 10523
rect 7284 10489 7296 10523
rect 7238 10483 7296 10489
rect 8849 10523 8907 10529
rect 8849 10489 8861 10523
rect 8895 10489 8907 10523
rect 8849 10483 8907 10489
rect 1946 10452 1952 10464
rect 1907 10424 1952 10452
rect 1946 10412 1952 10424
rect 2004 10412 2010 10464
rect 6273 10455 6331 10461
rect 6273 10421 6285 10455
rect 6319 10452 6331 10455
rect 6641 10455 6699 10461
rect 6641 10452 6653 10455
rect 6319 10424 6653 10452
rect 6319 10421 6331 10424
rect 6273 10415 6331 10421
rect 6641 10421 6653 10424
rect 6687 10452 6699 10455
rect 6730 10452 6736 10464
rect 6687 10424 6736 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 6730 10412 6736 10424
rect 6788 10452 6794 10464
rect 7253 10452 7281 10483
rect 6788 10424 7281 10452
rect 7837 10455 7895 10461
rect 6788 10412 6794 10424
rect 7837 10421 7849 10455
rect 7883 10452 7895 10455
rect 8662 10452 8668 10464
rect 7883 10424 8668 10452
rect 7883 10421 7895 10424
rect 7837 10415 7895 10421
rect 8662 10412 8668 10424
rect 8720 10452 8726 10464
rect 8864 10452 8892 10483
rect 8720 10424 8892 10452
rect 8720 10412 8726 10424
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 2590 10208 2596 10260
rect 2648 10248 2654 10260
rect 3142 10248 3148 10260
rect 2648 10220 3148 10248
rect 2648 10208 2654 10220
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 3878 10248 3884 10260
rect 3839 10220 3884 10248
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4893 10251 4951 10257
rect 4893 10248 4905 10251
rect 4212 10220 4905 10248
rect 4212 10208 4218 10220
rect 4893 10217 4905 10220
rect 4939 10217 4951 10251
rect 5626 10248 5632 10260
rect 5587 10220 5632 10248
rect 4893 10211 4951 10217
rect 5626 10208 5632 10220
rect 5684 10208 5690 10260
rect 6638 10208 6644 10260
rect 6696 10248 6702 10260
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 6696 10220 6837 10248
rect 6696 10208 6702 10220
rect 6825 10217 6837 10220
rect 6871 10217 6883 10251
rect 7650 10248 7656 10260
rect 7611 10220 7656 10248
rect 6825 10211 6883 10217
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 8662 10248 8668 10260
rect 8623 10220 8668 10248
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 4706 10180 4712 10192
rect 4028 10152 4712 10180
rect 4028 10140 4034 10152
rect 4706 10140 4712 10152
rect 4764 10180 4770 10192
rect 6549 10183 6607 10189
rect 4764 10152 6408 10180
rect 4764 10140 4770 10152
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10112 1458 10124
rect 1670 10112 1676 10124
rect 1452 10084 1676 10112
rect 1452 10072 1458 10084
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 2958 10112 2964 10124
rect 2919 10084 2964 10112
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 3510 10072 3516 10124
rect 3568 10112 3574 10124
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 3568 10084 4261 10112
rect 3568 10072 3574 10084
rect 4249 10081 4261 10084
rect 4295 10081 4307 10115
rect 6086 10112 6092 10124
rect 6047 10084 6092 10112
rect 4249 10075 4307 10081
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 6270 10112 6276 10124
rect 6231 10084 6276 10112
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6380 10112 6408 10152
rect 6549 10149 6561 10183
rect 6595 10180 6607 10183
rect 6914 10180 6920 10192
rect 6595 10152 6920 10180
rect 6595 10149 6607 10152
rect 6549 10143 6607 10149
rect 6914 10140 6920 10152
rect 6972 10180 6978 10192
rect 7193 10183 7251 10189
rect 7193 10180 7205 10183
rect 6972 10152 7205 10180
rect 6972 10140 6978 10152
rect 7193 10149 7205 10152
rect 7239 10149 7251 10183
rect 7193 10143 7251 10149
rect 7374 10112 7380 10124
rect 6380 10084 7380 10112
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 7558 10112 7564 10124
rect 7519 10084 7564 10112
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 9744 10115 9802 10121
rect 9744 10081 9756 10115
rect 9790 10081 9802 10115
rect 9744 10075 9802 10081
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 10778 10112 10784 10124
rect 10735 10084 10784 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4617 10047 4675 10053
rect 4617 10044 4629 10047
rect 4120 10016 4629 10044
rect 4120 10004 4126 10016
rect 4617 10013 4629 10016
rect 4663 10044 4675 10047
rect 5074 10044 5080 10056
rect 4663 10016 5080 10044
rect 4663 10013 4675 10016
rect 4617 10007 4675 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 9759 10044 9787 10075
rect 10778 10072 10784 10084
rect 10836 10072 10842 10124
rect 11054 10044 11060 10056
rect 9759 10016 11060 10044
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 4430 9985 4436 9988
rect 4414 9979 4436 9985
rect 4414 9945 4426 9979
rect 4414 9939 4436 9945
rect 4430 9936 4436 9939
rect 4488 9936 4494 9988
rect 4525 9979 4583 9985
rect 4525 9945 4537 9979
rect 4571 9976 4583 9979
rect 4982 9976 4988 9988
rect 4571 9948 4988 9976
rect 4571 9945 4583 9948
rect 4525 9939 4583 9945
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 1394 9868 1400 9920
rect 1452 9908 1458 9920
rect 2222 9908 2228 9920
rect 1452 9880 2228 9908
rect 1452 9868 1458 9880
rect 2222 9868 2228 9880
rect 2280 9908 2286 9920
rect 2409 9911 2467 9917
rect 2409 9908 2421 9911
rect 2280 9880 2421 9908
rect 2280 9868 2286 9880
rect 2409 9877 2421 9880
rect 2455 9877 2467 9911
rect 2774 9908 2780 9920
rect 2735 9880 2780 9908
rect 2409 9871 2467 9877
rect 2774 9868 2780 9880
rect 2832 9868 2838 9920
rect 5353 9911 5411 9917
rect 5353 9877 5365 9911
rect 5399 9908 5411 9911
rect 5626 9908 5632 9920
rect 5399 9880 5632 9908
rect 5399 9877 5411 9880
rect 5353 9871 5411 9877
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 8386 9908 8392 9920
rect 8343 9880 8392 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9815 9911 9873 9917
rect 9815 9908 9827 9911
rect 9732 9880 9827 9908
rect 9732 9868 9738 9880
rect 9815 9877 9827 9880
rect 9861 9877 9873 9911
rect 9815 9871 9873 9877
rect 10919 9911 10977 9917
rect 10919 9877 10931 9911
rect 10965 9908 10977 9911
rect 12342 9908 12348 9920
rect 10965 9880 12348 9908
rect 10965 9877 10977 9880
rect 10919 9871 10977 9877
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 2958 9704 2964 9716
rect 2919 9676 2964 9704
rect 2958 9664 2964 9676
rect 3016 9664 3022 9716
rect 3697 9707 3755 9713
rect 3697 9673 3709 9707
rect 3743 9704 3755 9707
rect 4062 9704 4068 9716
rect 3743 9676 4068 9704
rect 3743 9673 3755 9676
rect 3697 9667 3755 9673
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 4982 9704 4988 9716
rect 4943 9676 4988 9704
rect 4982 9664 4988 9676
rect 5040 9664 5046 9716
rect 6270 9704 6276 9716
rect 6231 9676 6276 9704
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 7374 9664 7380 9716
rect 7432 9704 7438 9716
rect 7929 9707 7987 9713
rect 7929 9704 7941 9707
rect 7432 9676 7941 9704
rect 7432 9664 7438 9676
rect 7929 9673 7941 9676
rect 7975 9673 7987 9707
rect 7929 9667 7987 9673
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 10134 9704 10140 9716
rect 8076 9676 10140 9704
rect 8076 9664 8082 9676
rect 1946 9596 1952 9648
rect 2004 9636 2010 9648
rect 3237 9639 3295 9645
rect 3237 9636 3249 9639
rect 2004 9608 3249 9636
rect 2004 9596 2010 9608
rect 3237 9605 3249 9608
rect 3283 9605 3295 9639
rect 3237 9599 3295 9605
rect 3252 9500 3280 9599
rect 3326 9596 3332 9648
rect 3384 9636 3390 9648
rect 4614 9636 4620 9648
rect 3384 9608 4531 9636
rect 4575 9608 4620 9636
rect 3384 9596 3390 9608
rect 4246 9568 4252 9580
rect 4207 9540 4252 9568
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 4503 9568 4531 9608
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 7239 9639 7297 9645
rect 7239 9605 7251 9639
rect 7285 9636 7297 9639
rect 9582 9636 9588 9648
rect 7285 9608 9588 9636
rect 7285 9605 7297 9608
rect 7239 9599 7297 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 8018 9568 8024 9580
rect 4503 9540 8024 9568
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9568 8263 9571
rect 8846 9568 8852 9580
rect 8251 9540 8852 9568
rect 8251 9537 8263 9540
rect 8205 9531 8263 9537
rect 8846 9528 8852 9540
rect 8904 9568 8910 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 8904 9540 9137 9568
rect 8904 9528 8910 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 3252 9472 3801 9500
rect 3789 9469 3801 9472
rect 3835 9469 3847 9503
rect 3970 9500 3976 9512
rect 3931 9472 3976 9500
rect 3789 9463 3847 9469
rect 3804 9432 3832 9463
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 5166 9500 5172 9512
rect 5127 9472 5172 9500
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5626 9500 5632 9512
rect 5587 9472 5632 9500
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 7168 9503 7226 9509
rect 7168 9469 7180 9503
rect 7214 9500 7226 9503
rect 7466 9500 7472 9512
rect 7214 9472 7472 9500
rect 7214 9469 7226 9472
rect 7168 9463 7226 9469
rect 7466 9460 7472 9472
rect 7524 9500 7530 9512
rect 9759 9509 9787 9676
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 10873 9707 10931 9713
rect 10873 9704 10885 9707
rect 10836 9676 10885 9704
rect 10836 9664 10842 9676
rect 10873 9673 10885 9676
rect 10919 9673 10931 9707
rect 10873 9667 10931 9673
rect 10597 9639 10655 9645
rect 10597 9605 10609 9639
rect 10643 9636 10655 9639
rect 11054 9636 11060 9648
rect 10643 9608 11060 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 7561 9503 7619 9509
rect 7561 9500 7573 9503
rect 7524 9472 7573 9500
rect 7524 9460 7530 9472
rect 7561 9469 7573 9472
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 9744 9503 9802 9509
rect 9744 9469 9756 9503
rect 9790 9469 9802 9503
rect 9744 9463 9802 9469
rect 4154 9432 4160 9444
rect 3804 9404 4160 9432
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 5902 9432 5908 9444
rect 5863 9404 5908 9432
rect 5902 9392 5908 9404
rect 5960 9392 5966 9444
rect 8297 9435 8355 9441
rect 8297 9401 8309 9435
rect 8343 9432 8355 9435
rect 8386 9432 8392 9444
rect 8343 9404 8392 9432
rect 8343 9401 8355 9404
rect 8297 9395 8355 9401
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 8662 9392 8668 9444
rect 8720 9432 8726 9444
rect 8849 9435 8907 9441
rect 8849 9432 8861 9435
rect 8720 9404 8861 9432
rect 8720 9392 8726 9404
rect 8849 9401 8861 9404
rect 8895 9401 8907 9435
rect 8849 9395 8907 9401
rect 1670 9364 1676 9376
rect 1631 9336 1676 9364
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 6086 9364 6092 9376
rect 3200 9336 6092 9364
rect 3200 9324 3206 9336
rect 6086 9324 6092 9336
rect 6144 9364 6150 9376
rect 6641 9367 6699 9373
rect 6641 9364 6653 9367
rect 6144 9336 6653 9364
rect 6144 9324 6150 9336
rect 6641 9333 6653 9336
rect 6687 9364 6699 9367
rect 6822 9364 6828 9376
rect 6687 9336 6828 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 9815 9367 9873 9373
rect 9815 9364 9827 9367
rect 8076 9336 9827 9364
rect 8076 9324 8082 9336
rect 9815 9333 9827 9336
rect 9861 9333 9873 9367
rect 9815 9327 9873 9333
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 3145 9163 3203 9169
rect 3145 9129 3157 9163
rect 3191 9160 3203 9163
rect 3191 9132 4154 9160
rect 3191 9129 3203 9132
rect 3145 9123 3203 9129
rect 2866 9052 2872 9104
rect 2924 9092 2930 9104
rect 3510 9092 3516 9104
rect 2924 9064 3516 9092
rect 2924 9052 2930 9064
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 3881 9095 3939 9101
rect 3881 9061 3893 9095
rect 3927 9092 3939 9095
rect 3970 9092 3976 9104
rect 3927 9064 3976 9092
rect 3927 9061 3939 9064
rect 3881 9055 3939 9061
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 4126 9092 4154 9132
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 5353 9163 5411 9169
rect 5353 9160 5365 9163
rect 4856 9132 5365 9160
rect 4856 9120 4862 9132
rect 5353 9129 5365 9132
rect 5399 9129 5411 9163
rect 5353 9123 5411 9129
rect 7469 9163 7527 9169
rect 7469 9129 7481 9163
rect 7515 9160 7527 9163
rect 7558 9160 7564 9172
rect 7515 9132 7564 9160
rect 7515 9129 7527 9132
rect 7469 9123 7527 9129
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 9732 9132 9812 9160
rect 9732 9120 9738 9132
rect 5626 9092 5632 9104
rect 4126 9064 5632 9092
rect 2958 9024 2964 9036
rect 2919 8996 2964 9024
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 4908 9033 4936 9064
rect 5626 9052 5632 9064
rect 5684 9092 5690 9104
rect 8110 9092 8116 9104
rect 5684 9064 6132 9092
rect 8071 9064 8116 9092
rect 5684 9052 5690 9064
rect 6104 9036 6132 9064
rect 8110 9052 8116 9064
rect 8168 9052 8174 9104
rect 8662 9092 8668 9104
rect 8623 9064 8668 9092
rect 8662 9052 8668 9064
rect 8720 9052 8726 9104
rect 9784 9101 9812 9132
rect 9769 9095 9827 9101
rect 9769 9061 9781 9095
rect 9815 9061 9827 9095
rect 9769 9055 9827 9061
rect 9858 9052 9864 9104
rect 9916 9092 9922 9104
rect 9916 9064 9961 9092
rect 9916 9052 9922 9064
rect 12342 9052 12348 9104
rect 12400 9092 12406 9104
rect 15562 9092 15568 9104
rect 12400 9064 15568 9092
rect 12400 9052 12406 9064
rect 15562 9052 15568 9064
rect 15620 9052 15626 9104
rect 4341 9027 4399 9033
rect 4341 9024 4353 9027
rect 4126 8996 4353 9024
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 4126 8956 4154 8996
rect 4341 8993 4353 8996
rect 4387 8993 4399 9027
rect 4341 8987 4399 8993
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 8993 4951 9027
rect 5166 9024 5172 9036
rect 4893 8987 4951 8993
rect 5000 8996 5172 9024
rect 2740 8928 4154 8956
rect 2740 8916 2746 8928
rect 3050 8848 3056 8900
rect 3108 8888 3114 8900
rect 5000 8888 5028 8996
rect 5166 8984 5172 8996
rect 5224 9024 5230 9036
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 5224 8996 5733 9024
rect 5224 8984 5230 8996
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 5810 8984 5816 9036
rect 5868 9024 5874 9036
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 5868 8996 5917 9024
rect 5868 8984 5874 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 6086 8984 6092 9036
rect 6144 9024 6150 9036
rect 6365 9027 6423 9033
rect 6365 9024 6377 9027
rect 6144 8996 6377 9024
rect 6144 8984 6150 8996
rect 6365 8993 6377 8996
rect 6411 8993 6423 9027
rect 11238 9024 11244 9036
rect 11199 8996 11244 9024
rect 6365 8987 6423 8993
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 6178 8956 6184 8968
rect 5123 8928 6184 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 6178 8916 6184 8928
rect 6236 8916 6242 8968
rect 6638 8956 6644 8968
rect 6599 8928 6644 8956
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 8018 8956 8024 8968
rect 7979 8928 8024 8956
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 10042 8956 10048 8968
rect 10003 8928 10048 8956
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 3108 8860 5028 8888
rect 3108 8848 3114 8860
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 5166 8820 5172 8832
rect 4028 8792 5172 8820
rect 4028 8780 4034 8792
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8812 8792 8953 8820
rect 8812 8780 8818 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 11379 8823 11437 8829
rect 11379 8820 11391 8823
rect 10836 8792 11391 8820
rect 10836 8780 10842 8792
rect 11379 8789 11391 8792
rect 11425 8789 11437 8823
rect 11379 8783 11437 8789
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 2958 8576 2964 8628
rect 3016 8616 3022 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 3016 8588 3249 8616
rect 3016 8576 3022 8588
rect 3237 8585 3249 8588
rect 3283 8616 3295 8619
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 3283 8588 4077 8616
rect 3283 8585 3295 8588
rect 3237 8579 3295 8585
rect 4065 8585 4077 8588
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 8110 8616 8116 8628
rect 7791 8588 8116 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 8110 8576 8116 8588
rect 8168 8616 8174 8628
rect 9677 8619 9735 8625
rect 9677 8616 9689 8619
rect 8168 8588 9689 8616
rect 8168 8576 8174 8588
rect 9677 8585 9689 8588
rect 9723 8616 9735 8619
rect 9858 8616 9864 8628
rect 9723 8588 9864 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 11238 8616 11244 8628
rect 11199 8588 11244 8616
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 9217 8551 9275 8557
rect 9217 8517 9229 8551
rect 9263 8548 9275 8551
rect 10042 8548 10048 8560
rect 9263 8520 10048 8548
rect 9263 8517 9275 8520
rect 9217 8511 9275 8517
rect 10042 8508 10048 8520
rect 10100 8548 10106 8560
rect 10410 8548 10416 8560
rect 10100 8520 10416 8548
rect 10100 8508 10106 8520
rect 10410 8508 10416 8520
rect 10468 8548 10474 8560
rect 10781 8551 10839 8557
rect 10781 8548 10793 8551
rect 10468 8520 10793 8548
rect 10468 8508 10474 8520
rect 10781 8517 10793 8520
rect 10827 8517 10839 8551
rect 10781 8511 10839 8517
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 4798 8480 4804 8492
rect 1636 8452 4804 8480
rect 1636 8440 1642 8452
rect 4798 8440 4804 8452
rect 4856 8480 4862 8492
rect 5905 8483 5963 8489
rect 4856 8452 5212 8480
rect 4856 8440 4862 8452
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8381 2835 8415
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 2777 8375 2835 8381
rect 3620 8384 3985 8412
rect 2792 8288 2820 8375
rect 2685 8279 2743 8285
rect 2685 8245 2697 8279
rect 2731 8276 2743 8279
rect 2774 8276 2780 8288
rect 2731 8248 2780 8276
rect 2731 8245 2743 8248
rect 2685 8239 2743 8245
rect 2774 8236 2780 8248
rect 2832 8236 2838 8288
rect 2961 8279 3019 8285
rect 2961 8245 2973 8279
rect 3007 8276 3019 8279
rect 3050 8276 3056 8288
rect 3007 8248 3056 8276
rect 3007 8245 3019 8248
rect 2961 8239 3019 8245
rect 3050 8236 3056 8248
rect 3108 8236 3114 8288
rect 3510 8236 3516 8288
rect 3568 8276 3574 8288
rect 3620 8285 3648 8384
rect 3973 8381 3985 8384
rect 4019 8412 4031 8415
rect 4338 8412 4344 8424
rect 4019 8384 4344 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 4338 8372 4344 8384
rect 4396 8372 4402 8424
rect 5184 8421 5212 8452
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 6825 8483 6883 8489
rect 6825 8480 6837 8483
rect 5951 8452 6837 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 6825 8449 6837 8452
rect 6871 8480 6883 8483
rect 6914 8480 6920 8492
rect 6871 8452 6920 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8480 8723 8483
rect 8754 8480 8760 8492
rect 8711 8452 8760 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 8754 8440 8760 8452
rect 8812 8480 8818 8492
rect 9950 8480 9956 8492
rect 8812 8452 9956 8480
rect 8812 8440 8818 8452
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10686 8480 10692 8492
rect 10275 8452 10692 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 3789 8347 3847 8353
rect 3789 8313 3801 8347
rect 3835 8344 3847 8347
rect 4154 8344 4160 8356
rect 3835 8316 4160 8344
rect 3835 8313 3847 8316
rect 3789 8307 3847 8313
rect 4126 8304 4160 8316
rect 4212 8304 4218 8356
rect 3605 8279 3663 8285
rect 3605 8276 3617 8279
rect 3568 8248 3617 8276
rect 3568 8236 3574 8248
rect 3605 8245 3617 8248
rect 3651 8245 3663 8279
rect 4126 8276 4154 8304
rect 4614 8276 4620 8288
rect 4126 8248 4620 8276
rect 3605 8239 3663 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 5077 8279 5135 8285
rect 5077 8245 5089 8279
rect 5123 8276 5135 8279
rect 5534 8276 5540 8288
rect 5123 8248 5540 8276
rect 5123 8245 5135 8248
rect 5077 8239 5135 8245
rect 5534 8236 5540 8248
rect 5592 8276 5598 8288
rect 5644 8276 5672 8375
rect 7187 8347 7245 8353
rect 7187 8313 7199 8347
rect 7233 8313 7245 8347
rect 7187 8307 7245 8313
rect 8757 8347 8815 8353
rect 8757 8313 8769 8347
rect 8803 8313 8815 8347
rect 8757 8307 8815 8313
rect 10321 8347 10379 8353
rect 10321 8313 10333 8347
rect 10367 8313 10379 8347
rect 10321 8307 10379 8313
rect 6086 8276 6092 8288
rect 5592 8248 6092 8276
rect 5592 8236 5598 8248
rect 6086 8236 6092 8248
rect 6144 8276 6150 8288
rect 6181 8279 6239 8285
rect 6181 8276 6193 8279
rect 6144 8248 6193 8276
rect 6144 8236 6150 8248
rect 6181 8245 6193 8248
rect 6227 8245 6239 8279
rect 6181 8239 6239 8245
rect 6641 8279 6699 8285
rect 6641 8245 6653 8279
rect 6687 8276 6699 8279
rect 6730 8276 6736 8288
rect 6687 8248 6736 8276
rect 6687 8245 6699 8248
rect 6641 8239 6699 8245
rect 6730 8236 6736 8248
rect 6788 8276 6794 8288
rect 7202 8276 7230 8307
rect 7282 8276 7288 8288
rect 6788 8248 7288 8276
rect 6788 8236 6794 8248
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 8386 8276 8392 8288
rect 7800 8248 8392 8276
rect 7800 8236 7806 8248
rect 8386 8236 8392 8248
rect 8444 8276 8450 8288
rect 8772 8276 8800 8307
rect 8444 8248 8800 8276
rect 8444 8236 8450 8248
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 9953 8279 10011 8285
rect 9953 8276 9965 8279
rect 9824 8248 9965 8276
rect 9824 8236 9830 8248
rect 9953 8245 9965 8248
rect 9999 8276 10011 8279
rect 10336 8276 10364 8307
rect 9999 8248 10364 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 2682 8072 2688 8084
rect 2179 8044 2688 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2682 8032 2688 8044
rect 2740 8072 2746 8084
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2740 8044 2789 8072
rect 2740 8032 2746 8044
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 3142 8072 3148 8084
rect 3103 8044 3148 8072
rect 2777 8035 2835 8041
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 5813 8075 5871 8081
rect 5813 8072 5825 8075
rect 5408 8044 5825 8072
rect 5408 8032 5414 8044
rect 5813 8041 5825 8044
rect 5859 8041 5871 8075
rect 5813 8035 5871 8041
rect 5902 8032 5908 8084
rect 5960 8072 5966 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 5960 8044 6653 8072
rect 5960 8032 5966 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 8018 8072 8024 8084
rect 7979 8044 8024 8072
rect 6641 8035 6699 8041
rect 2590 7964 2596 8016
rect 2648 8004 2654 8016
rect 2648 7976 5856 8004
rect 2648 7964 2654 7976
rect 5828 7948 5856 7976
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 2038 7936 2044 7948
rect 1995 7908 2044 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 2961 7939 3019 7945
rect 2961 7905 2973 7939
rect 3007 7905 3019 7939
rect 2961 7899 3019 7905
rect 3881 7939 3939 7945
rect 3881 7905 3893 7939
rect 3927 7936 3939 7939
rect 4062 7936 4068 7948
rect 3927 7908 4068 7936
rect 3927 7905 3939 7908
rect 3881 7899 3939 7905
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 2976 7868 3004 7899
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4338 7936 4344 7948
rect 4299 7908 4344 7936
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 5626 7936 5632 7948
rect 5587 7908 5632 7936
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 6089 7939 6147 7945
rect 6089 7936 6101 7939
rect 5868 7908 6101 7936
rect 5868 7896 5874 7908
rect 6089 7905 6101 7908
rect 6135 7905 6147 7939
rect 6656 7936 6684 8035
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9674 8072 9680 8084
rect 9539 8044 9680 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 10778 8072 10784 8084
rect 10739 8044 10784 8072
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 7187 8007 7245 8013
rect 7187 7973 7199 8007
rect 7233 8004 7245 8007
rect 7282 8004 7288 8016
rect 7233 7976 7288 8004
rect 7233 7973 7245 7976
rect 7187 7967 7245 7973
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 8711 8007 8769 8013
rect 8711 7973 8723 8007
rect 8757 8004 8769 8007
rect 8846 8004 8852 8016
rect 8757 7976 8852 8004
rect 8757 7973 8769 7976
rect 8711 7967 8769 7973
rect 8846 7964 8852 7976
rect 8904 7964 8910 8016
rect 9766 8004 9772 8016
rect 9185 7976 9772 8004
rect 6825 7939 6883 7945
rect 6825 7936 6837 7939
rect 6656 7908 6837 7936
rect 6089 7899 6147 7905
rect 6825 7905 6837 7908
rect 6871 7905 6883 7939
rect 8570 7936 8576 7948
rect 8531 7908 8576 7936
rect 6825 7899 6883 7905
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 3970 7868 3976 7880
rect 2547 7840 3976 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4522 7868 4528 7880
rect 4483 7840 4528 7868
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4157 7803 4215 7809
rect 4157 7800 4169 7803
rect 3436 7772 4169 7800
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3436 7741 3464 7772
rect 4157 7769 4169 7772
rect 4203 7769 4215 7803
rect 4157 7763 4215 7769
rect 7745 7803 7803 7809
rect 7745 7769 7757 7803
rect 7791 7800 7803 7803
rect 9185 7800 9213 7976
rect 9766 7964 9772 7976
rect 9824 8004 9830 8016
rect 9861 8007 9919 8013
rect 9861 8004 9873 8007
rect 9824 7976 9873 8004
rect 9824 7964 9830 7976
rect 9861 7973 9873 7976
rect 9907 7973 9919 8007
rect 9861 7967 9919 7973
rect 9950 7964 9956 8016
rect 10008 8004 10014 8016
rect 11379 8007 11437 8013
rect 11379 8004 11391 8007
rect 10008 7976 11391 8004
rect 10008 7964 10014 7976
rect 11379 7973 11391 7976
rect 11425 7973 11437 8007
rect 11379 7967 11437 7973
rect 11238 7936 11244 7948
rect 11199 7908 11244 7936
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 9582 7828 9588 7880
rect 9640 7868 9646 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 9640 7840 9781 7868
rect 9640 7828 9646 7840
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 10060 7800 10088 7831
rect 7791 7772 9213 7800
rect 9692 7772 10088 7800
rect 7791 7769 7803 7772
rect 7745 7763 7803 7769
rect 9692 7744 9720 7772
rect 3421 7735 3479 7741
rect 3421 7732 3433 7735
rect 3108 7704 3433 7732
rect 3108 7692 3114 7704
rect 3421 7701 3433 7704
rect 3467 7701 3479 7735
rect 3421 7695 3479 7701
rect 5261 7735 5319 7741
rect 5261 7701 5273 7735
rect 5307 7732 5319 7735
rect 5534 7732 5540 7744
rect 5307 7704 5540 7732
rect 5307 7701 5319 7704
rect 5261 7695 5319 7701
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 9674 7732 9680 7744
rect 8720 7704 9680 7732
rect 8720 7692 8726 7704
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2590 7528 2596 7540
rect 2551 7500 2596 7528
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 2961 7531 3019 7537
rect 2961 7497 2973 7531
rect 3007 7528 3019 7531
rect 4522 7528 4528 7540
rect 3007 7500 4528 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 2409 7327 2467 7333
rect 1443 7296 1992 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 1964 7200 1992 7296
rect 2409 7293 2421 7327
rect 2455 7324 2467 7327
rect 2976 7324 3004 7491
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 6086 7528 6092 7540
rect 5684 7500 6092 7528
rect 5684 7488 5690 7500
rect 6086 7488 6092 7500
rect 6144 7528 6150 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 6144 7500 6193 7528
rect 6144 7488 6150 7500
rect 6181 7497 6193 7500
rect 6227 7497 6239 7531
rect 7742 7528 7748 7540
rect 7703 7500 7748 7528
rect 6181 7491 6239 7497
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 8481 7531 8539 7537
rect 8481 7497 8493 7531
rect 8527 7528 8539 7531
rect 8570 7528 8576 7540
rect 8527 7500 8576 7528
rect 8527 7497 8539 7500
rect 8481 7491 8539 7497
rect 3326 7420 3332 7472
rect 3384 7460 3390 7472
rect 8496 7460 8524 7491
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 3384 7432 8524 7460
rect 3384 7420 3390 7432
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 10100 7432 10732 7460
rect 10100 7420 10106 7432
rect 3050 7352 3056 7404
rect 3108 7392 3114 7404
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 3108 7364 3525 7392
rect 3108 7352 3114 7364
rect 3513 7361 3525 7364
rect 3559 7392 3571 7395
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 3559 7364 4445 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 8573 7395 8631 7401
rect 8573 7392 8585 7395
rect 5951 7364 8585 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 8573 7361 8585 7364
rect 8619 7392 8631 7395
rect 8938 7392 8944 7404
rect 8619 7364 8944 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 10410 7392 10416 7404
rect 10371 7364 10416 7392
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 10704 7401 10732 7432
rect 10689 7395 10747 7401
rect 10689 7361 10701 7395
rect 10735 7361 10747 7395
rect 10689 7355 10747 7361
rect 2455 7296 3004 7324
rect 3145 7327 3203 7333
rect 2455 7293 2467 7296
rect 2409 7287 2467 7293
rect 3145 7293 3157 7327
rect 3191 7324 3203 7327
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3191 7296 3433 7324
rect 3191 7293 3203 7296
rect 3145 7287 3203 7293
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3694 7324 3700 7336
rect 3655 7296 3700 7324
rect 3421 7287 3479 7293
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7324 5135 7327
rect 5350 7324 5356 7336
rect 5123 7296 5356 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5592 7296 5641 7324
rect 5592 7284 5598 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 6178 7284 6184 7336
rect 6236 7324 6242 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6236 7296 6837 7324
rect 6236 7284 6242 7296
rect 6825 7293 6837 7296
rect 6871 7324 6883 7327
rect 8021 7327 8079 7333
rect 8021 7324 8033 7327
rect 6871 7296 8033 7324
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 8021 7293 8033 7296
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 9493 7327 9551 7333
rect 9493 7293 9505 7327
rect 9539 7324 9551 7327
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 9539 7296 10149 7324
rect 9539 7293 9551 7296
rect 9493 7287 9551 7293
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 2038 7216 2044 7268
rect 2096 7256 2102 7268
rect 2317 7259 2375 7265
rect 2317 7256 2329 7259
rect 2096 7228 2329 7256
rect 2096 7216 2102 7228
rect 2317 7225 2329 7228
rect 2363 7256 2375 7259
rect 6641 7259 6699 7265
rect 2363 7228 3648 7256
rect 2363 7225 2375 7228
rect 2317 7219 2375 7225
rect 1946 7188 1952 7200
rect 1907 7160 1952 7188
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 2498 7148 2504 7200
rect 2556 7188 2562 7200
rect 3145 7191 3203 7197
rect 3145 7188 3157 7191
rect 2556 7160 3157 7188
rect 2556 7148 2562 7160
rect 3145 7157 3157 7160
rect 3191 7188 3203 7191
rect 3237 7191 3295 7197
rect 3237 7188 3249 7191
rect 3191 7160 3249 7188
rect 3191 7157 3203 7160
rect 3145 7151 3203 7157
rect 3237 7157 3249 7160
rect 3283 7157 3295 7191
rect 3620 7188 3648 7228
rect 6641 7225 6653 7259
rect 6687 7256 6699 7259
rect 7187 7259 7245 7265
rect 7187 7256 7199 7259
rect 6687 7228 7199 7256
rect 6687 7225 6699 7228
rect 6641 7219 6699 7225
rect 7187 7225 7199 7228
rect 7233 7256 7245 7259
rect 7282 7256 7288 7268
rect 7233 7228 7288 7256
rect 7233 7225 7245 7228
rect 7187 7219 7245 7225
rect 7282 7216 7288 7228
rect 7340 7216 7346 7268
rect 8570 7216 8576 7268
rect 8628 7256 8634 7268
rect 8894 7259 8952 7265
rect 8894 7256 8906 7259
rect 8628 7228 8906 7256
rect 8628 7216 8634 7228
rect 8894 7225 8906 7228
rect 8940 7225 8952 7259
rect 8894 7219 8952 7225
rect 3881 7191 3939 7197
rect 3881 7188 3893 7191
rect 3620 7160 3893 7188
rect 3237 7151 3295 7157
rect 3881 7157 3893 7160
rect 3927 7157 3939 7191
rect 10152 7188 10180 7287
rect 10505 7259 10563 7265
rect 10505 7225 10517 7259
rect 10551 7225 10563 7259
rect 10505 7219 10563 7225
rect 10520 7188 10548 7219
rect 11330 7188 11336 7200
rect 10152 7160 10548 7188
rect 11291 7160 11336 7188
rect 3881 7151 3939 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 2869 6987 2927 6993
rect 2869 6984 2881 6987
rect 2004 6956 2881 6984
rect 2004 6944 2010 6956
rect 2869 6953 2881 6956
rect 2915 6953 2927 6987
rect 2869 6947 2927 6953
rect 3513 6987 3571 6993
rect 3513 6953 3525 6987
rect 3559 6984 3571 6987
rect 3694 6984 3700 6996
rect 3559 6956 3700 6984
rect 3559 6953 3571 6956
rect 3513 6947 3571 6953
rect 3694 6944 3700 6956
rect 3752 6944 3758 6996
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 4525 6987 4583 6993
rect 4525 6984 4537 6987
rect 4028 6956 4537 6984
rect 4028 6944 4034 6956
rect 4525 6953 4537 6956
rect 4571 6953 4583 6987
rect 6086 6984 6092 6996
rect 6047 6956 6092 6984
rect 4525 6947 4583 6953
rect 6086 6944 6092 6956
rect 6144 6944 6150 6996
rect 8113 6987 8171 6993
rect 8113 6953 8125 6987
rect 8159 6984 8171 6987
rect 9674 6984 9680 6996
rect 8159 6956 9680 6984
rect 8159 6953 8171 6956
rect 8113 6947 8171 6953
rect 9674 6944 9680 6956
rect 9732 6984 9738 6996
rect 9732 6956 9904 6984
rect 9732 6944 9738 6956
rect 3712 6916 3740 6944
rect 6917 6919 6975 6925
rect 3712 6888 5948 6916
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2498 6848 2504 6860
rect 2455 6820 2504 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2682 6848 2688 6860
rect 2643 6820 2688 6848
rect 2682 6808 2688 6820
rect 2740 6848 2746 6860
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 2740 6820 3801 6848
rect 2740 6808 2746 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 4062 6848 4068 6860
rect 4023 6820 4068 6848
rect 3789 6811 3847 6817
rect 2501 6715 2559 6721
rect 2501 6681 2513 6715
rect 2547 6712 2559 6715
rect 2590 6712 2596 6724
rect 2547 6684 2596 6712
rect 2547 6681 2559 6684
rect 2501 6675 2559 6681
rect 2590 6672 2596 6684
rect 2648 6712 2654 6724
rect 3050 6712 3056 6724
rect 2648 6684 3056 6712
rect 2648 6672 2654 6684
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 3804 6644 3832 6811
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4356 6857 4384 6888
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6848 4399 6851
rect 4522 6848 4528 6860
rect 4387 6820 4528 6848
rect 4387 6817 4399 6820
rect 4341 6811 4399 6817
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 5626 6848 5632 6860
rect 5587 6820 5632 6848
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5920 6857 5948 6888
rect 6917 6885 6929 6919
rect 6963 6916 6975 6919
rect 7282 6916 7288 6928
rect 6963 6888 7288 6916
rect 6963 6885 6975 6888
rect 6917 6879 6975 6885
rect 7282 6876 7288 6888
rect 7340 6916 7346 6928
rect 7514 6919 7572 6925
rect 7514 6916 7526 6919
rect 7340 6888 7526 6916
rect 7340 6876 7346 6888
rect 7514 6885 7526 6888
rect 7560 6916 7572 6919
rect 8570 6916 8576 6928
rect 7560 6888 8576 6916
rect 7560 6885 7572 6888
rect 7514 6879 7572 6885
rect 8570 6876 8576 6888
rect 8628 6876 8634 6928
rect 8938 6916 8944 6928
rect 8899 6888 8944 6916
rect 8938 6876 8944 6888
rect 8996 6876 9002 6928
rect 9493 6919 9551 6925
rect 9493 6885 9505 6919
rect 9539 6916 9551 6919
rect 9582 6916 9588 6928
rect 9539 6888 9588 6916
rect 9539 6885 9551 6888
rect 9493 6879 9551 6885
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 9766 6916 9772 6928
rect 9727 6888 9772 6916
rect 9766 6876 9772 6888
rect 9824 6876 9830 6928
rect 9876 6925 9904 6956
rect 10410 6944 10416 6996
rect 10468 6984 10474 6996
rect 10689 6987 10747 6993
rect 10689 6984 10701 6987
rect 10468 6956 10701 6984
rect 10468 6944 10474 6956
rect 10689 6953 10701 6956
rect 10735 6953 10747 6987
rect 10689 6947 10747 6953
rect 9861 6919 9919 6925
rect 9861 6885 9873 6919
rect 9907 6885 9919 6919
rect 9861 6879 9919 6885
rect 5905 6851 5963 6857
rect 5905 6817 5917 6851
rect 5951 6817 5963 6851
rect 5905 6811 5963 6817
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 7193 6851 7251 6857
rect 7193 6848 7205 6851
rect 6696 6820 7205 6848
rect 6696 6808 6702 6820
rect 7193 6817 7205 6820
rect 7239 6848 7251 6851
rect 8754 6848 8760 6860
rect 7239 6820 8760 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6780 5319 6783
rect 5534 6780 5540 6792
rect 5307 6752 5540 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5534 6740 5540 6752
rect 5592 6780 5598 6792
rect 6914 6780 6920 6792
rect 5592 6752 6920 6780
rect 5592 6740 5598 6752
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 10042 6780 10048 6792
rect 10003 6752 10048 6780
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 5718 6712 5724 6724
rect 4212 6684 4257 6712
rect 5679 6684 5724 6712
rect 4212 6672 4218 6684
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 4338 6644 4344 6656
rect 3804 6616 4344 6644
rect 4338 6604 4344 6616
rect 4396 6644 4402 6656
rect 4982 6644 4988 6656
rect 4396 6616 4988 6644
rect 4396 6604 4402 6616
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 2133 6443 2191 6449
rect 2133 6409 2145 6443
rect 2179 6440 2191 6443
rect 2682 6440 2688 6452
rect 2179 6412 2688 6440
rect 2179 6409 2191 6412
rect 2133 6403 2191 6409
rect 2682 6400 2688 6412
rect 2740 6400 2746 6452
rect 9674 6440 9680 6452
rect 9635 6412 9680 6440
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 9824 6412 10425 6440
rect 9824 6400 9830 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 10413 6403 10471 6409
rect 1670 6332 1676 6384
rect 1728 6372 1734 6384
rect 8938 6372 8944 6384
rect 1728 6344 8944 6372
rect 1728 6332 1734 6344
rect 8938 6332 8944 6344
rect 8996 6332 9002 6384
rect 9033 6375 9091 6381
rect 9033 6341 9045 6375
rect 9079 6372 9091 6375
rect 10042 6372 10048 6384
rect 9079 6344 10048 6372
rect 9079 6341 9091 6344
rect 9033 6335 9091 6341
rect 10042 6332 10048 6344
rect 10100 6332 10106 6384
rect 4982 6304 4988 6316
rect 4943 6276 4988 6304
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 8478 6304 8484 6316
rect 8391 6276 8484 6304
rect 8478 6264 8484 6276
rect 8536 6304 8542 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 8536 6276 9965 6304
rect 8536 6264 8542 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 3513 6239 3571 6245
rect 3513 6236 3525 6239
rect 3252 6208 3525 6236
rect 2498 6168 2504 6180
rect 2411 6140 2504 6168
rect 2498 6128 2504 6140
rect 2556 6168 2562 6180
rect 3142 6168 3148 6180
rect 2556 6140 3148 6168
rect 2556 6128 2562 6140
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 2590 6060 2596 6112
rect 2648 6100 2654 6112
rect 3252 6109 3280 6208
rect 3513 6205 3525 6208
rect 3559 6205 3571 6239
rect 5077 6239 5135 6245
rect 5077 6236 5089 6239
rect 3513 6199 3571 6205
rect 4816 6208 5089 6236
rect 4154 6128 4160 6180
rect 4212 6168 4218 6180
rect 4212 6140 4257 6168
rect 4212 6128 4218 6140
rect 2777 6103 2835 6109
rect 2777 6100 2789 6103
rect 2648 6072 2789 6100
rect 2648 6060 2654 6072
rect 2777 6069 2789 6072
rect 2823 6100 2835 6103
rect 3237 6103 3295 6109
rect 3237 6100 3249 6103
rect 2823 6072 3249 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 3237 6069 3249 6072
rect 3283 6069 3295 6103
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 3237 6063 3295 6069
rect 4522 6060 4528 6072
rect 4580 6100 4586 6112
rect 4816 6109 4844 6208
rect 5077 6205 5089 6208
rect 5123 6236 5135 6239
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5123 6208 6377 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6822 6236 6828 6248
rect 6735 6208 6828 6236
rect 6365 6199 6423 6205
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6972 6208 7297 6236
rect 6972 6196 6978 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 6840 6168 6868 6196
rect 8205 6171 8263 6177
rect 8205 6168 8217 6171
rect 6840 6140 8217 6168
rect 8205 6137 8217 6140
rect 8251 6137 8263 6171
rect 8205 6131 8263 6137
rect 8570 6128 8576 6180
rect 8628 6168 8634 6180
rect 8628 6140 8673 6168
rect 8628 6128 8634 6140
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 4580 6072 4813 6100
rect 4580 6060 4586 6072
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 4801 6063 4859 6069
rect 5626 6060 5632 6112
rect 5684 6100 5690 6112
rect 5997 6103 6055 6109
rect 5997 6100 6009 6103
rect 5684 6072 6009 6100
rect 5684 6060 5690 6072
rect 5997 6069 6009 6072
rect 6043 6069 6055 6103
rect 7098 6100 7104 6112
rect 7059 6072 7104 6100
rect 5997 6063 6055 6069
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 7340 6072 7849 6100
rect 7340 6060 7346 6072
rect 7837 6069 7849 6072
rect 7883 6069 7895 6103
rect 7837 6063 7895 6069
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 4154 5896 4160 5908
rect 3559 5868 4160 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 4154 5856 4160 5868
rect 4212 5896 4218 5908
rect 5718 5896 5724 5908
rect 4212 5868 5724 5896
rect 4212 5856 4218 5868
rect 5718 5856 5724 5868
rect 5776 5896 5782 5908
rect 6457 5899 6515 5905
rect 6457 5896 6469 5899
rect 5776 5868 6469 5896
rect 5776 5856 5782 5868
rect 6457 5865 6469 5868
rect 6503 5865 6515 5899
rect 6914 5896 6920 5908
rect 6875 5868 6920 5896
rect 6457 5859 6515 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 8021 5899 8079 5905
rect 8021 5865 8033 5899
rect 8067 5896 8079 5899
rect 8570 5896 8576 5908
rect 8067 5868 8576 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 8570 5856 8576 5868
rect 8628 5896 8634 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8628 5868 9137 5896
rect 8628 5856 8634 5868
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 7282 5788 7288 5840
rect 7340 5828 7346 5840
rect 7422 5831 7480 5837
rect 7422 5828 7434 5831
rect 7340 5800 7434 5828
rect 7340 5788 7346 5800
rect 7422 5797 7434 5800
rect 7468 5797 7480 5831
rect 8478 5828 8484 5840
rect 8439 5800 8484 5828
rect 7422 5791 7480 5797
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 8754 5828 8760 5840
rect 8715 5800 8760 5828
rect 8754 5788 8760 5800
rect 8812 5788 8818 5840
rect 4062 5769 4068 5772
rect 3881 5763 3939 5769
rect 3881 5729 3893 5763
rect 3927 5760 3939 5763
rect 4053 5763 4068 5769
rect 4053 5760 4065 5763
rect 3927 5732 4065 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 4053 5729 4065 5732
rect 4053 5723 4068 5729
rect 4062 5720 4068 5723
rect 4120 5720 4126 5772
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 4430 5760 4436 5772
rect 4387 5732 4436 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 5629 5763 5687 5769
rect 5629 5760 5641 5763
rect 5592 5732 5641 5760
rect 5592 5720 5598 5732
rect 5629 5729 5641 5732
rect 5675 5729 5687 5763
rect 5810 5760 5816 5772
rect 5771 5732 5816 5760
rect 5629 5723 5687 5729
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 7098 5760 7104 5772
rect 7059 5732 7104 5760
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 8938 5720 8944 5772
rect 8996 5760 9002 5772
rect 9582 5760 9588 5772
rect 8996 5732 9588 5760
rect 8996 5720 9002 5732
rect 9582 5720 9588 5732
rect 9640 5760 9646 5772
rect 9712 5763 9770 5769
rect 9712 5760 9724 5763
rect 9640 5732 9724 5760
rect 9640 5720 9646 5732
rect 9712 5729 9724 5732
rect 9758 5760 9770 5763
rect 11330 5760 11336 5772
rect 9758 5732 11336 5760
rect 9758 5729 9770 5732
rect 9712 5723 9770 5729
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 2832 5664 4537 5692
rect 2832 5652 2838 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 5169 5695 5227 5701
rect 5169 5692 5181 5695
rect 5132 5664 5181 5692
rect 5132 5652 5138 5664
rect 5169 5661 5181 5664
rect 5215 5692 5227 5695
rect 5828 5692 5856 5720
rect 5215 5664 5856 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 2590 5584 2596 5636
rect 2648 5624 2654 5636
rect 4154 5624 4160 5636
rect 2648 5596 4160 5624
rect 2648 5584 2654 5596
rect 4154 5584 4160 5596
rect 4212 5624 4218 5636
rect 4212 5596 4257 5624
rect 4212 5584 4218 5596
rect 5534 5556 5540 5568
rect 5495 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 5902 5556 5908 5568
rect 5863 5528 5908 5556
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 9815 5559 9873 5565
rect 9815 5556 9827 5559
rect 9548 5528 9827 5556
rect 9548 5516 9554 5528
rect 9815 5525 9827 5528
rect 9861 5525 9873 5559
rect 9815 5519 9873 5525
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 2685 5355 2743 5361
rect 2685 5321 2697 5355
rect 2731 5352 2743 5355
rect 2866 5352 2872 5364
rect 2731 5324 2872 5352
rect 2731 5321 2743 5324
rect 2685 5315 2743 5321
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 5902 5352 5908 5364
rect 3099 5324 5908 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 3068 5148 3096 5315
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 9582 5352 9588 5364
rect 9543 5324 9588 5352
rect 9582 5312 9588 5324
rect 9640 5352 9646 5364
rect 9950 5352 9956 5364
rect 9640 5324 9956 5352
rect 9640 5312 9646 5324
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 4154 5244 4160 5296
rect 4212 5284 4218 5296
rect 4893 5287 4951 5293
rect 4893 5284 4905 5287
rect 4212 5256 4905 5284
rect 4212 5244 4218 5256
rect 4893 5253 4905 5256
rect 4939 5253 4951 5287
rect 5166 5284 5172 5296
rect 5127 5256 5172 5284
rect 4893 5247 4951 5253
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 9861 5287 9919 5293
rect 9861 5253 9873 5287
rect 9907 5284 9919 5287
rect 10686 5284 10692 5296
rect 9907 5256 10692 5284
rect 9907 5253 9919 5256
rect 9861 5247 9919 5253
rect 10686 5244 10692 5256
rect 10744 5244 10750 5296
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 5316 5188 7389 5216
rect 5316 5176 5322 5188
rect 3418 5148 3424 5160
rect 2547 5120 3096 5148
rect 3331 5120 3424 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 3418 5108 3424 5120
rect 3476 5148 3482 5160
rect 4062 5148 4068 5160
rect 3476 5120 4068 5148
rect 3476 5108 3482 5120
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 5353 5151 5411 5157
rect 5353 5148 5365 5151
rect 4295 5120 5365 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 5353 5117 5365 5120
rect 5399 5117 5411 5151
rect 5810 5148 5816 5160
rect 5723 5120 5816 5148
rect 5353 5111 5411 5117
rect 5368 5080 5396 5111
rect 5810 5108 5816 5120
rect 5868 5148 5874 5160
rect 6178 5148 6184 5160
rect 5868 5120 6184 5148
rect 5868 5108 5874 5120
rect 6178 5108 6184 5120
rect 6236 5108 6242 5160
rect 6840 5157 6868 5188
rect 7377 5185 7389 5188
rect 7423 5216 7435 5219
rect 7466 5216 7472 5228
rect 7423 5188 7472 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 9456 5188 10241 5216
rect 9456 5176 9462 5188
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5148 9091 5151
rect 9582 5148 9588 5160
rect 9079 5120 9588 5148
rect 9079 5117 9091 5120
rect 9033 5111 9091 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 9692 5157 9720 5188
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 9677 5151 9735 5157
rect 9677 5117 9689 5151
rect 9723 5117 9735 5151
rect 9677 5111 9735 5117
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10816 5151 10874 5157
rect 10816 5148 10828 5151
rect 10100 5120 10828 5148
rect 10100 5108 10106 5120
rect 10816 5117 10828 5120
rect 10862 5148 10874 5151
rect 11241 5151 11299 5157
rect 11241 5148 11253 5151
rect 10862 5120 11253 5148
rect 10862 5117 10874 5120
rect 10816 5111 10874 5117
rect 11241 5117 11253 5120
rect 11287 5117 11299 5151
rect 11241 5111 11299 5117
rect 5534 5080 5540 5092
rect 5368 5052 5540 5080
rect 5534 5040 5540 5052
rect 5592 5080 5598 5092
rect 6457 5083 6515 5089
rect 6457 5080 6469 5083
rect 5592 5052 6469 5080
rect 5592 5040 5598 5052
rect 6457 5049 6469 5052
rect 6503 5049 6515 5083
rect 6457 5043 6515 5049
rect 7282 5040 7288 5092
rect 7340 5080 7346 5092
rect 7745 5083 7803 5089
rect 7745 5080 7757 5083
rect 7340 5052 7757 5080
rect 7340 5040 7346 5052
rect 7745 5049 7757 5052
rect 7791 5049 7803 5083
rect 8018 5080 8024 5092
rect 7979 5052 8024 5080
rect 7745 5043 7803 5049
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 8113 5083 8171 5089
rect 8113 5049 8125 5083
rect 8159 5049 8171 5083
rect 8113 5043 8171 5049
rect 8665 5083 8723 5089
rect 8665 5049 8677 5083
rect 8711 5080 8723 5083
rect 9398 5080 9404 5092
rect 8711 5052 9404 5080
rect 8711 5049 8723 5052
rect 8665 5043 8723 5049
rect 3234 4972 3240 5024
rect 3292 5012 3298 5024
rect 4062 5012 4068 5024
rect 3292 4984 4068 5012
rect 3292 4972 3298 4984
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4522 5012 4528 5024
rect 4483 4984 4528 5012
rect 4522 4972 4528 4984
rect 4580 4972 4586 5024
rect 6178 5012 6184 5024
rect 6139 4984 6184 5012
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 7009 5015 7067 5021
rect 7009 4981 7021 5015
rect 7055 5012 7067 5015
rect 7098 5012 7104 5024
rect 7055 4984 7104 5012
rect 7055 4981 7067 4984
rect 7009 4975 7067 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 8128 5012 8156 5043
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 10919 5083 10977 5089
rect 10919 5049 10931 5083
rect 10965 5080 10977 5083
rect 14642 5080 14648 5092
rect 10965 5052 14648 5080
rect 10965 5049 10977 5052
rect 10919 5043 10977 5049
rect 14642 5040 14648 5052
rect 14700 5040 14706 5092
rect 7892 4984 8156 5012
rect 7892 4972 7898 4984
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 3510 4808 3516 4820
rect 2915 4780 3516 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4246 4808 4252 4820
rect 4028 4780 4154 4808
rect 4207 4780 4252 4808
rect 4028 4768 4034 4780
rect 2593 4743 2651 4749
rect 2593 4709 2605 4743
rect 2639 4740 2651 4743
rect 2682 4740 2688 4752
rect 2639 4712 2688 4740
rect 2639 4709 2651 4712
rect 2593 4703 2651 4709
rect 2682 4700 2688 4712
rect 2740 4740 2746 4752
rect 3418 4740 3424 4752
rect 2740 4712 3424 4740
rect 2740 4700 2746 4712
rect 3418 4700 3424 4712
rect 3476 4700 3482 4752
rect 4126 4740 4154 4780
rect 4246 4768 4252 4780
rect 4304 4768 4310 4820
rect 4706 4808 4712 4820
rect 4667 4780 4712 4808
rect 4706 4768 4712 4780
rect 4764 4808 4770 4820
rect 4982 4808 4988 4820
rect 4764 4780 4988 4808
rect 4764 4768 4770 4780
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 6012 4780 7144 4808
rect 6012 4740 6040 4780
rect 7116 4749 7144 4780
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 7248 4780 7389 4808
rect 7248 4768 7254 4780
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 8941 4811 8999 4817
rect 8941 4808 8953 4811
rect 7377 4771 7435 4777
rect 8036 4780 8953 4808
rect 8036 4752 8064 4780
rect 8941 4777 8953 4780
rect 8987 4777 8999 4811
rect 8941 4771 8999 4777
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9364 4780 9413 4808
rect 9364 4768 9370 4780
rect 9401 4777 9413 4780
rect 9447 4808 9459 4811
rect 9490 4808 9496 4820
rect 9447 4780 9496 4808
rect 9447 4777 9459 4780
rect 9401 4771 9459 4777
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 6549 4743 6607 4749
rect 6549 4740 6561 4743
rect 4126 4712 6040 4740
rect 6104 4712 6561 4740
rect 2774 4672 2780 4684
rect 2687 4644 2780 4672
rect 2774 4632 2780 4644
rect 2832 4672 2838 4684
rect 5074 4672 5080 4684
rect 2832 4644 5080 4672
rect 2832 4632 2838 4644
rect 5074 4632 5080 4644
rect 5132 4632 5138 4684
rect 5445 4675 5503 4681
rect 5445 4641 5457 4675
rect 5491 4672 5503 4675
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 5491 4644 5825 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 5813 4641 5825 4644
rect 5859 4672 5871 4675
rect 5902 4672 5908 4684
rect 5859 4644 5908 4672
rect 5859 4641 5871 4644
rect 5813 4635 5871 4641
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 6104 4616 6132 4712
rect 6549 4709 6561 4712
rect 6595 4709 6607 4743
rect 6549 4703 6607 4709
rect 7101 4743 7159 4749
rect 7101 4709 7113 4743
rect 7147 4740 7159 4743
rect 8018 4740 8024 4752
rect 7147 4712 8024 4740
rect 7147 4709 7159 4712
rect 7101 4703 7159 4709
rect 8018 4700 8024 4712
rect 8076 4700 8082 4752
rect 8113 4743 8171 4749
rect 8113 4709 8125 4743
rect 8159 4740 8171 4743
rect 8202 4740 8208 4752
rect 8159 4712 8208 4740
rect 8159 4709 8171 4712
rect 8113 4703 8171 4709
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 9858 4672 9864 4684
rect 9819 4644 9864 4672
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 10134 4632 10140 4684
rect 10192 4672 10198 4684
rect 11238 4672 11244 4684
rect 11296 4681 11302 4684
rect 11296 4675 11334 4681
rect 10192 4644 11244 4672
rect 10192 4632 10198 4644
rect 11238 4632 11244 4644
rect 11322 4641 11334 4675
rect 11296 4635 11334 4641
rect 11296 4632 11302 4635
rect 2498 4564 2504 4616
rect 2556 4604 2562 4616
rect 4522 4604 4528 4616
rect 2556 4576 4528 4604
rect 2556 4564 2562 4576
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4604 5595 4607
rect 6086 4604 6092 4616
rect 5583 4576 6092 4604
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4604 6515 4607
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 6503 4576 7757 4604
rect 6503 4573 6515 4576
rect 6457 4567 6515 4573
rect 7745 4573 7757 4576
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4604 8079 4607
rect 8110 4604 8116 4616
rect 8067 4576 8116 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 5718 4496 5724 4548
rect 5776 4536 5782 4548
rect 6472 4536 6500 4567
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 8846 4604 8852 4616
rect 8711 4576 8852 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 9490 4564 9496 4616
rect 9548 4604 9554 4616
rect 9677 4607 9735 4613
rect 9677 4604 9689 4607
rect 9548 4576 9689 4604
rect 9548 4564 9554 4576
rect 9677 4573 9689 4576
rect 9723 4573 9735 4607
rect 9677 4567 9735 4573
rect 5776 4508 6500 4536
rect 5776 4496 5782 4508
rect 6178 4468 6184 4480
rect 6139 4440 6184 4468
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 10502 4428 10508 4480
rect 10560 4468 10566 4480
rect 11379 4471 11437 4477
rect 11379 4468 11391 4471
rect 10560 4440 11391 4468
rect 10560 4428 10566 4440
rect 11379 4437 11391 4440
rect 11425 4437 11437 4471
rect 11379 4431 11437 4437
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 2774 4264 2780 4276
rect 2735 4236 2780 4264
rect 2774 4224 2780 4236
rect 2832 4224 2838 4276
rect 2866 4224 2872 4276
rect 2924 4264 2930 4276
rect 4249 4267 4307 4273
rect 4249 4264 4261 4267
rect 2924 4236 4261 4264
rect 2924 4224 2930 4236
rect 4249 4233 4261 4236
rect 4295 4264 4307 4267
rect 4706 4264 4712 4276
rect 4295 4236 4712 4264
rect 4295 4233 4307 4236
rect 4249 4227 4307 4233
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 6086 4224 6092 4276
rect 6144 4264 6150 4276
rect 6181 4267 6239 4273
rect 6181 4264 6193 4267
rect 6144 4236 6193 4264
rect 6144 4224 6150 4236
rect 6181 4233 6193 4236
rect 6227 4233 6239 4267
rect 6181 4227 6239 4233
rect 7745 4267 7803 4273
rect 7745 4233 7757 4267
rect 7791 4264 7803 4267
rect 9858 4264 9864 4276
rect 7791 4236 9864 4264
rect 7791 4233 7803 4236
rect 7745 4227 7803 4233
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 11238 4264 11244 4276
rect 11199 4236 11244 4264
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 8846 4156 8852 4208
rect 8904 4196 8910 4208
rect 9217 4199 9275 4205
rect 9217 4196 9229 4199
rect 8904 4168 9229 4196
rect 8904 4156 8910 4168
rect 9217 4165 9229 4168
rect 9263 4165 9275 4199
rect 9217 4159 9275 4165
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4128 4031 4131
rect 4246 4128 4252 4140
rect 4019 4100 4252 4128
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 8665 4131 8723 4137
rect 4764 4100 5304 4128
rect 4764 4088 4770 4100
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 2292 4063 2350 4069
rect 2292 4060 2304 4063
rect 2179 4032 2304 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 2292 4029 2304 4032
rect 2338 4060 2350 4063
rect 3234 4060 3240 4072
rect 2338 4032 3240 4060
rect 2338 4029 2350 4032
rect 2292 4023 2350 4029
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 3329 4063 3387 4069
rect 3329 4029 3341 4063
rect 3375 4029 3387 4063
rect 5074 4060 5080 4072
rect 5035 4032 5080 4060
rect 3329 4023 3387 4029
rect 3142 3992 3148 4004
rect 3055 3964 3148 3992
rect 3142 3952 3148 3964
rect 3200 3992 3206 4004
rect 3344 3992 3372 4023
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 5276 4069 5304 4100
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 9306 4128 9312 4140
rect 8711 4100 9312 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 5261 4063 5319 4069
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 5442 4060 5448 4072
rect 5307 4032 5448 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5626 4060 5632 4072
rect 5587 4032 5632 4060
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 6822 4060 6828 4072
rect 6783 4032 6828 4060
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 9582 4020 9588 4072
rect 9640 4060 9646 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 9640 4032 10057 4060
rect 9640 4020 9646 4032
rect 10045 4029 10057 4032
rect 10091 4060 10103 4063
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 10091 4032 10241 4060
rect 10091 4029 10103 4032
rect 10045 4023 10103 4029
rect 10229 4029 10241 4032
rect 10275 4029 10287 4063
rect 10229 4023 10287 4029
rect 4709 3995 4767 4001
rect 4709 3992 4721 3995
rect 3200 3964 4721 3992
rect 3200 3952 3206 3964
rect 4709 3961 4721 3964
rect 4755 3992 4767 3995
rect 5644 3992 5672 4020
rect 4755 3964 5672 3992
rect 5905 3995 5963 4001
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 5905 3961 5917 3995
rect 5951 3992 5963 3995
rect 6730 3992 6736 4004
rect 5951 3964 6736 3992
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 6730 3952 6736 3964
rect 6788 3952 6794 4004
rect 7190 4001 7196 4004
rect 7146 3995 7196 4001
rect 7146 3992 7158 3995
rect 7024 3964 7158 3992
rect 7024 3936 7052 3964
rect 7146 3961 7158 3964
rect 7192 3961 7196 3995
rect 7146 3955 7196 3961
rect 7190 3952 7196 3955
rect 7248 3952 7254 4004
rect 8481 3995 8539 4001
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 8757 3995 8815 4001
rect 8757 3992 8769 3995
rect 8527 3964 8769 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 8757 3961 8769 3964
rect 8803 3992 8815 3995
rect 9950 3992 9956 4004
rect 8803 3964 9956 3992
rect 8803 3961 8815 3964
rect 8757 3955 8815 3961
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 10134 3992 10140 4004
rect 10095 3964 10140 3992
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 2363 3927 2421 3933
rect 2363 3893 2375 3927
rect 2409 3924 2421 3927
rect 2590 3924 2596 3936
rect 2409 3896 2596 3924
rect 2409 3893 2421 3896
rect 2363 3887 2421 3893
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 6641 3927 6699 3933
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 7006 3924 7012 3936
rect 6687 3896 7012 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8202 3924 8208 3936
rect 8159 3896 8208 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 9858 3924 9864 3936
rect 9723 3896 9864 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 2682 3720 2688 3732
rect 2643 3692 2688 3720
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 3099 3723 3157 3729
rect 3099 3689 3111 3723
rect 3145 3720 3157 3723
rect 5718 3720 5724 3732
rect 3145 3692 5724 3720
rect 3145 3689 3157 3692
rect 3099 3683 3157 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 5997 3723 6055 3729
rect 5997 3689 6009 3723
rect 6043 3720 6055 3723
rect 6178 3720 6184 3732
rect 6043 3692 6184 3720
rect 6043 3689 6055 3692
rect 5997 3683 6055 3689
rect 6178 3680 6184 3692
rect 6236 3720 6242 3732
rect 6822 3720 6828 3732
rect 6236 3692 6828 3720
rect 6236 3680 6242 3692
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 8110 3720 8116 3732
rect 8071 3692 8116 3720
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 8260 3692 11836 3720
rect 8260 3680 8266 3692
rect 5166 3652 5172 3664
rect 4126 3624 5172 3652
rect 3050 3593 3056 3596
rect 3028 3587 3056 3593
rect 3028 3584 3040 3587
rect 2963 3556 3040 3584
rect 3028 3553 3040 3556
rect 3108 3584 3114 3596
rect 4126 3584 4154 3624
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 6641 3655 6699 3661
rect 6641 3652 6653 3655
rect 5276 3624 6653 3652
rect 3108 3556 4154 3584
rect 3028 3547 3056 3553
rect 3050 3544 3056 3547
rect 3108 3544 3114 3556
rect 4246 3544 4252 3596
rect 4304 3584 4310 3596
rect 4341 3587 4399 3593
rect 4341 3584 4353 3587
rect 4304 3556 4353 3584
rect 4304 3544 4310 3556
rect 4341 3553 4353 3556
rect 4387 3553 4399 3587
rect 4706 3584 4712 3596
rect 4667 3556 4712 3584
rect 4341 3547 4399 3553
rect 4356 3516 4384 3547
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 5074 3584 5080 3596
rect 4987 3556 5080 3584
rect 5074 3544 5080 3556
rect 5132 3584 5138 3596
rect 5276 3584 5304 3624
rect 6641 3621 6653 3624
rect 6687 3621 6699 3655
rect 6641 3615 6699 3621
rect 7006 3612 7012 3664
rect 7064 3652 7070 3664
rect 7146 3655 7204 3661
rect 7146 3652 7158 3655
rect 7064 3624 7158 3652
rect 7064 3612 7070 3624
rect 7146 3621 7158 3624
rect 7192 3621 7204 3655
rect 7146 3615 7204 3621
rect 5718 3584 5724 3596
rect 5132 3556 5304 3584
rect 5368 3556 5724 3584
rect 5132 3544 5138 3556
rect 5368 3516 5396 3556
rect 5718 3544 5724 3556
rect 5776 3584 5782 3596
rect 6273 3587 6331 3593
rect 6273 3584 6285 3587
rect 5776 3556 6285 3584
rect 5776 3544 5782 3556
rect 6273 3553 6285 3556
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 7745 3587 7803 3593
rect 7745 3553 7757 3587
rect 7791 3584 7803 3587
rect 8220 3584 8248 3680
rect 9858 3652 9864 3664
rect 9819 3624 9864 3652
rect 9858 3612 9864 3624
rect 9916 3612 9922 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 11241 3655 11299 3661
rect 11241 3652 11253 3655
rect 10008 3624 11253 3652
rect 10008 3612 10014 3624
rect 11241 3621 11253 3624
rect 11287 3621 11299 3655
rect 11241 3615 11299 3621
rect 11808 3596 11836 3692
rect 11790 3584 11796 3596
rect 7791 3556 8248 3584
rect 11751 3556 11796 3584
rect 7791 3553 7803 3556
rect 7745 3547 7803 3553
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 12805 3587 12863 3593
rect 12805 3553 12817 3587
rect 12851 3584 12863 3587
rect 12894 3584 12900 3596
rect 12851 3556 12900 3584
rect 12851 3553 12863 3556
rect 12805 3547 12863 3553
rect 12894 3544 12900 3556
rect 12952 3544 12958 3596
rect 4356 3488 5396 3516
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 5500 3488 5641 3516
rect 5500 3476 5506 3488
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 6822 3516 6828 3528
rect 6783 3488 6828 3516
rect 5629 3479 5687 3485
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 8570 3516 8576 3528
rect 8531 3488 8576 3516
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9769 3519 9827 3525
rect 9769 3516 9781 3519
rect 8904 3488 9781 3516
rect 8904 3476 8910 3488
rect 9769 3485 9781 3488
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 10318 3448 10324 3460
rect 10279 3420 10324 3448
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 9398 3380 9404 3392
rect 9359 3352 9404 3380
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 12943 3383 13001 3389
rect 12943 3380 12955 3383
rect 12860 3352 12955 3380
rect 12860 3340 12866 3352
rect 12943 3349 12955 3352
rect 12989 3349 13001 3383
rect 12943 3343 13001 3349
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 2590 3176 2596 3188
rect 2551 3148 2596 3176
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 3050 3176 3056 3188
rect 3011 3148 3056 3176
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 4614 3176 4620 3188
rect 4575 3148 4620 3176
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 8389 3179 8447 3185
rect 8389 3176 8401 3179
rect 6880 3148 8401 3176
rect 6880 3136 6886 3148
rect 8389 3145 8401 3148
rect 8435 3145 8447 3179
rect 8846 3176 8852 3188
rect 8807 3148 8852 3176
rect 8389 3139 8447 3145
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10321 3179 10379 3185
rect 10321 3176 10333 3179
rect 9916 3148 10333 3176
rect 9916 3136 9922 3148
rect 10321 3145 10333 3148
rect 10367 3145 10379 3179
rect 11790 3176 11796 3188
rect 11751 3148 11796 3176
rect 10321 3139 10379 3145
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 12894 3176 12900 3188
rect 12855 3148 12900 3176
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 2608 3040 2636 3136
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 4706 3108 4712 3120
rect 4387 3080 4712 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 4706 3068 4712 3080
rect 4764 3068 4770 3120
rect 5902 3068 5908 3120
rect 5960 3108 5966 3120
rect 7745 3111 7803 3117
rect 7745 3108 7757 3111
rect 5960 3080 7757 3108
rect 5960 3068 5966 3080
rect 7745 3077 7757 3080
rect 7791 3077 7803 3111
rect 7745 3071 7803 3077
rect 8202 3068 8208 3120
rect 8260 3108 8266 3120
rect 11057 3111 11115 3117
rect 11057 3108 11069 3111
rect 8260 3080 11069 3108
rect 8260 3068 8266 3080
rect 11057 3077 11069 3080
rect 11103 3077 11115 3111
rect 11057 3071 11115 3077
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 2608 3012 3341 3040
rect 3329 3009 3341 3012
rect 3375 3009 3387 3043
rect 3970 3040 3976 3052
rect 3931 3012 3976 3040
rect 3329 3003 3387 3009
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 5920 3040 5948 3068
rect 9398 3040 9404 3052
rect 4126 3012 5948 3040
rect 9359 3012 9404 3040
rect 3418 2864 3424 2916
rect 3476 2904 3482 2916
rect 4126 2904 4154 3012
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3040 10103 3043
rect 10318 3040 10324 3052
rect 10091 3012 10324 3040
rect 10091 3009 10103 3012
rect 10045 3003 10103 3009
rect 10318 3000 10324 3012
rect 10376 3040 10382 3052
rect 10376 3012 12531 3040
rect 10376 3000 10382 3012
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 4801 2975 4859 2981
rect 4801 2972 4813 2975
rect 4672 2944 4813 2972
rect 4672 2932 4678 2944
rect 4801 2941 4813 2944
rect 4847 2941 4859 2975
rect 5442 2972 5448 2984
rect 5403 2944 5448 2972
rect 4801 2935 4859 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 5718 2972 5724 2984
rect 5675 2944 5724 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 6822 2972 6828 2984
rect 6783 2944 6828 2972
rect 6822 2932 6828 2944
rect 6880 2972 6886 2984
rect 12503 2981 12531 3012
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 6880 2944 8033 2972
rect 6880 2932 6886 2944
rect 8021 2941 8033 2944
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 10873 2975 10931 2981
rect 10873 2941 10885 2975
rect 10919 2972 10931 2975
rect 11425 2975 11483 2981
rect 11425 2972 11437 2975
rect 10919 2944 11437 2972
rect 10919 2941 10931 2944
rect 10873 2935 10931 2941
rect 11425 2941 11437 2944
rect 11471 2941 11483 2975
rect 11425 2935 11483 2941
rect 12488 2975 12546 2981
rect 12488 2941 12500 2975
rect 12534 2972 12546 2975
rect 13265 2975 13323 2981
rect 13265 2972 13277 2975
rect 12534 2944 13277 2972
rect 12534 2941 12546 2944
rect 12488 2935 12546 2941
rect 13265 2941 13277 2944
rect 13311 2941 13323 2975
rect 13265 2935 13323 2941
rect 7006 2904 7012 2916
rect 3476 2876 4154 2904
rect 6656 2876 7012 2904
rect 3476 2864 3482 2876
rect 6656 2848 6684 2876
rect 7006 2864 7012 2876
rect 7064 2904 7070 2916
rect 7146 2907 7204 2913
rect 7146 2904 7158 2907
rect 7064 2876 7158 2904
rect 7064 2864 7070 2876
rect 7146 2873 7158 2876
rect 7192 2873 7204 2907
rect 7146 2867 7204 2873
rect 9217 2907 9275 2913
rect 9217 2873 9229 2907
rect 9263 2904 9275 2907
rect 9490 2904 9496 2916
rect 9263 2876 9496 2904
rect 9263 2873 9275 2876
rect 9217 2867 9275 2873
rect 9490 2864 9496 2876
rect 9548 2864 9554 2916
rect 5902 2836 5908 2848
rect 5863 2808 5908 2836
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 6273 2839 6331 2845
rect 6273 2805 6285 2839
rect 6319 2836 6331 2839
rect 6638 2836 6644 2848
rect 6319 2808 6644 2836
rect 6319 2805 6331 2808
rect 6273 2799 6331 2805
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 10888 2836 10916 2935
rect 12575 2907 12633 2913
rect 12575 2873 12587 2907
rect 12621 2904 12633 2907
rect 13722 2904 13728 2916
rect 12621 2876 13728 2904
rect 12621 2873 12633 2876
rect 12575 2867 12633 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 8352 2808 10916 2836
rect 8352 2796 8358 2808
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 3418 2632 3424 2644
rect 3375 2604 3424 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 3881 2635 3939 2641
rect 3881 2601 3893 2635
rect 3927 2632 3939 2635
rect 4614 2632 4620 2644
rect 3927 2604 4620 2632
rect 3927 2601 3939 2604
rect 3881 2595 3939 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 6822 2632 6828 2644
rect 5859 2604 6828 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 7834 2632 7840 2644
rect 7795 2604 7840 2632
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 9398 2632 9404 2644
rect 8711 2604 9404 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 9585 2635 9643 2641
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 9631 2604 9996 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 1302 2524 1308 2576
rect 1360 2564 1366 2576
rect 1949 2567 2007 2573
rect 1949 2564 1961 2567
rect 1360 2536 1961 2564
rect 1360 2524 1366 2536
rect 1949 2533 1961 2536
rect 1995 2533 2007 2567
rect 1949 2527 2007 2533
rect 6638 2524 6644 2576
rect 6696 2564 6702 2576
rect 7238 2567 7296 2573
rect 7238 2564 7250 2567
rect 6696 2536 7250 2564
rect 6696 2524 6702 2536
rect 7238 2533 7250 2536
rect 7284 2533 7296 2567
rect 7238 2527 7296 2533
rect 8570 2524 8576 2576
rect 8628 2564 8634 2576
rect 9968 2573 9996 2604
rect 9125 2567 9183 2573
rect 9125 2564 9137 2567
rect 8628 2536 9137 2564
rect 8628 2524 8634 2536
rect 9125 2533 9137 2536
rect 9171 2564 9183 2567
rect 9861 2567 9919 2573
rect 9861 2564 9873 2567
rect 9171 2536 9873 2564
rect 9171 2533 9183 2536
rect 9125 2527 9183 2533
rect 9861 2533 9873 2536
rect 9907 2533 9919 2567
rect 9861 2527 9919 2533
rect 9953 2567 10011 2573
rect 9953 2533 9965 2567
rect 9999 2564 10011 2567
rect 10134 2564 10140 2576
rect 9999 2536 10140 2564
rect 9999 2533 10011 2536
rect 9953 2527 10011 2533
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 2041 2499 2099 2505
rect 2041 2496 2053 2499
rect 1780 2468 2053 2496
rect 842 2252 848 2304
rect 900 2292 906 2304
rect 1780 2301 1808 2468
rect 2041 2465 2053 2468
rect 2087 2465 2099 2499
rect 2041 2459 2099 2465
rect 4614 2456 4620 2508
rect 4672 2496 4678 2508
rect 4709 2499 4767 2505
rect 4709 2496 4721 2499
rect 4672 2468 4721 2496
rect 4672 2456 4678 2468
rect 4709 2465 4721 2468
rect 4755 2465 4767 2499
rect 5537 2499 5595 2505
rect 5537 2496 5549 2499
rect 4709 2459 4767 2465
rect 4816 2468 5549 2496
rect 4816 2428 4844 2468
rect 5537 2465 5549 2468
rect 5583 2465 5595 2499
rect 5537 2459 5595 2465
rect 5902 2456 5908 2508
rect 5960 2496 5966 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 5960 2468 6929 2496
rect 5960 2456 5966 2468
rect 6917 2465 6929 2468
rect 6963 2496 6975 2499
rect 8113 2499 8171 2505
rect 8113 2496 8125 2499
rect 6963 2468 8125 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 8113 2465 8125 2468
rect 8159 2465 8171 2499
rect 8113 2459 8171 2465
rect 10962 2456 10968 2508
rect 11020 2496 11026 2508
rect 11333 2499 11391 2505
rect 11333 2496 11345 2499
rect 11020 2468 11345 2496
rect 11020 2456 11026 2468
rect 11333 2465 11345 2468
rect 11379 2496 11391 2499
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11379 2468 11897 2496
rect 11379 2465 11391 2468
rect 11333 2459 11391 2465
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 11885 2459 11943 2465
rect 12618 2456 12624 2468
rect 12676 2496 12682 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12676 2468 13185 2496
rect 12676 2456 12682 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 5442 2428 5448 2440
rect 4540 2400 4844 2428
rect 5403 2400 5448 2428
rect 4540 2304 4568 2400
rect 5442 2388 5448 2400
rect 5500 2428 5506 2440
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 5500 2400 6101 2428
rect 5500 2388 5506 2400
rect 6089 2397 6101 2400
rect 6135 2397 6147 2431
rect 6089 2391 6147 2397
rect 9306 2388 9312 2440
rect 9364 2428 9370 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9364 2400 10149 2428
rect 9364 2388 9370 2400
rect 10137 2397 10149 2400
rect 10183 2428 10195 2431
rect 12894 2428 12900 2440
rect 10183 2400 12900 2428
rect 10183 2397 10195 2400
rect 10137 2391 10195 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 1765 2295 1823 2301
rect 1765 2292 1777 2295
rect 900 2264 1777 2292
rect 900 2252 906 2264
rect 1765 2261 1777 2264
rect 1811 2261 1823 2295
rect 4522 2292 4528 2304
rect 4483 2264 4528 2292
rect 1765 2255 1823 2261
rect 4522 2252 4528 2264
rect 4580 2252 4586 2304
rect 6638 2292 6644 2304
rect 6599 2264 6644 2292
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 11514 2292 11520 2304
rect 11475 2264 11520 2292
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 11790 2252 11796 2304
rect 11848 2292 11854 2304
rect 12805 2295 12863 2301
rect 12805 2292 12817 2295
rect 11848 2264 12817 2292
rect 11848 2252 11854 2264
rect 12805 2261 12817 2264
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 1302 2048 1308 2100
rect 1360 2088 1366 2100
rect 6638 2088 6644 2100
rect 1360 2060 6644 2088
rect 1360 2048 1366 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 8938 76 8944 128
rect 8996 116 9002 128
rect 11790 116 11796 128
rect 8996 88 11796 116
rect 8996 76 9002 88
rect 11790 76 11796 88
rect 11848 76 11854 128
<< via1 >>
rect 664 39584 716 39636
rect 2504 39584 2556 39636
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 9772 35980 9824 36032
rect 15476 35980 15528 36032
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 9772 35819 9824 35828
rect 9772 35785 9781 35819
rect 9781 35785 9815 35819
rect 9815 35785 9824 35819
rect 9772 35776 9824 35785
rect 8484 35683 8536 35692
rect 8484 35649 8493 35683
rect 8493 35649 8527 35683
rect 8527 35649 8536 35683
rect 8484 35640 8536 35649
rect 4160 35572 4212 35624
rect 4896 35479 4948 35488
rect 4896 35445 4905 35479
rect 4905 35445 4939 35479
rect 4939 35445 4948 35479
rect 4896 35436 4948 35445
rect 6736 35436 6788 35488
rect 8024 35547 8076 35556
rect 8024 35513 8033 35547
rect 8033 35513 8067 35547
rect 8067 35513 8076 35547
rect 8024 35504 8076 35513
rect 8116 35547 8168 35556
rect 8116 35513 8125 35547
rect 8125 35513 8159 35547
rect 8159 35513 8168 35547
rect 8116 35504 8168 35513
rect 9680 35436 9732 35488
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 112 35232 164 35284
rect 8116 35232 8168 35284
rect 8852 35232 8904 35284
rect 5264 35207 5316 35216
rect 5264 35173 5273 35207
rect 5273 35173 5307 35207
rect 5307 35173 5316 35207
rect 5264 35164 5316 35173
rect 7748 35164 7800 35216
rect 3976 35096 4028 35148
rect 8392 35096 8444 35148
rect 9680 35139 9732 35148
rect 9680 35105 9689 35139
rect 9689 35105 9723 35139
rect 9723 35105 9732 35139
rect 9680 35096 9732 35105
rect 11428 35096 11480 35148
rect 4896 35028 4948 35080
rect 6000 35028 6052 35080
rect 6736 35028 6788 35080
rect 8576 35028 8628 35080
rect 5724 35003 5776 35012
rect 5724 34969 5733 35003
rect 5733 34969 5767 35003
rect 5767 34969 5776 35003
rect 5724 34960 5776 34969
rect 9772 34960 9824 35012
rect 4804 34935 4856 34944
rect 4804 34901 4813 34935
rect 4813 34901 4847 34935
rect 4847 34901 4856 34935
rect 4804 34892 4856 34901
rect 6828 34935 6880 34944
rect 6828 34901 6837 34935
rect 6837 34901 6871 34935
rect 6871 34901 6880 34935
rect 6828 34892 6880 34901
rect 8760 34892 8812 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 3516 34688 3568 34740
rect 5264 34688 5316 34740
rect 5632 34688 5684 34740
rect 6000 34731 6052 34740
rect 6000 34697 6009 34731
rect 6009 34697 6043 34731
rect 6043 34697 6052 34731
rect 6000 34688 6052 34697
rect 8116 34688 8168 34740
rect 9680 34731 9732 34740
rect 9680 34697 9689 34731
rect 9689 34697 9723 34731
rect 9723 34697 9732 34731
rect 9680 34688 9732 34697
rect 13728 34688 13780 34740
rect 3976 34620 4028 34672
rect 7840 34620 7892 34672
rect 8484 34620 8536 34672
rect 4804 34595 4856 34604
rect 4804 34561 4813 34595
rect 4813 34561 4847 34595
rect 4847 34561 4856 34595
rect 4804 34552 4856 34561
rect 8024 34552 8076 34604
rect 6828 34527 6880 34536
rect 6828 34493 6837 34527
rect 6837 34493 6871 34527
rect 6871 34493 6880 34527
rect 6828 34484 6880 34493
rect 4620 34416 4672 34468
rect 7012 34416 7064 34468
rect 3976 34348 4028 34400
rect 7748 34348 7800 34400
rect 8392 34391 8444 34400
rect 8392 34357 8401 34391
rect 8401 34357 8435 34391
rect 8435 34357 8444 34391
rect 8392 34348 8444 34357
rect 10784 34484 10836 34536
rect 8668 34459 8720 34468
rect 8668 34425 8677 34459
rect 8677 34425 8711 34459
rect 8711 34425 8720 34459
rect 8668 34416 8720 34425
rect 8760 34459 8812 34468
rect 8760 34425 8769 34459
rect 8769 34425 8803 34459
rect 8803 34425 8812 34459
rect 8760 34416 8812 34425
rect 8852 34348 8904 34400
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 4804 34144 4856 34196
rect 5632 34187 5684 34196
rect 5632 34153 5641 34187
rect 5641 34153 5675 34187
rect 5675 34153 5684 34187
rect 5632 34144 5684 34153
rect 6736 34144 6788 34196
rect 7012 34187 7064 34196
rect 7012 34153 7021 34187
rect 7021 34153 7055 34187
rect 7055 34153 7064 34187
rect 7012 34144 7064 34153
rect 8760 34144 8812 34196
rect 8852 34144 8904 34196
rect 8668 34076 8720 34128
rect 4712 34051 4764 34060
rect 4712 34017 4721 34051
rect 4721 34017 4755 34051
rect 4755 34017 4764 34051
rect 4712 34008 4764 34017
rect 3516 33940 3568 33992
rect 8484 34008 8536 34060
rect 6644 33983 6696 33992
rect 6644 33949 6653 33983
rect 6653 33949 6687 33983
rect 6687 33949 6696 33983
rect 6644 33940 6696 33949
rect 7656 33872 7708 33924
rect 8852 34008 8904 34060
rect 9956 34051 10008 34060
rect 9956 34017 9965 34051
rect 9965 34017 9999 34051
rect 9999 34017 10008 34051
rect 9956 34008 10008 34017
rect 9404 33940 9456 33992
rect 10968 34008 11020 34060
rect 11244 34051 11296 34060
rect 11244 34017 11253 34051
rect 11253 34017 11287 34051
rect 11287 34017 11296 34051
rect 11244 34008 11296 34017
rect 11428 33940 11480 33992
rect 9588 33872 9640 33924
rect 8760 33804 8812 33856
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 4620 33643 4672 33652
rect 4620 33609 4629 33643
rect 4629 33609 4663 33643
rect 4663 33609 4672 33643
rect 4620 33600 4672 33609
rect 8484 33643 8536 33652
rect 8484 33609 8493 33643
rect 8493 33609 8527 33643
rect 8527 33609 8536 33643
rect 8484 33600 8536 33609
rect 9496 33600 9548 33652
rect 9956 33643 10008 33652
rect 9956 33609 9965 33643
rect 9965 33609 9999 33643
rect 9999 33609 10008 33643
rect 9956 33600 10008 33609
rect 9680 33532 9732 33584
rect 10600 33532 10652 33584
rect 4712 33464 4764 33516
rect 7656 33464 7708 33516
rect 8760 33507 8812 33516
rect 8760 33473 8769 33507
rect 8769 33473 8803 33507
rect 8803 33473 8812 33507
rect 8760 33464 8812 33473
rect 10324 33464 10376 33516
rect 11244 33464 11296 33516
rect 3608 33396 3660 33448
rect 4988 33396 5040 33448
rect 5264 33396 5316 33448
rect 9312 33396 9364 33448
rect 10600 33439 10652 33448
rect 4620 33328 4672 33380
rect 6736 33328 6788 33380
rect 10600 33405 10609 33439
rect 10609 33405 10643 33439
rect 10643 33405 10652 33439
rect 10600 33396 10652 33405
rect 10968 33439 11020 33448
rect 10968 33405 10977 33439
rect 10977 33405 11011 33439
rect 11011 33405 11020 33439
rect 10968 33396 11020 33405
rect 5724 33303 5776 33312
rect 5724 33269 5733 33303
rect 5733 33269 5767 33303
rect 5767 33269 5776 33303
rect 5724 33260 5776 33269
rect 7012 33260 7064 33312
rect 7748 33303 7800 33312
rect 7748 33269 7757 33303
rect 7757 33269 7791 33303
rect 7791 33269 7800 33303
rect 7748 33260 7800 33269
rect 9128 33303 9180 33312
rect 9128 33269 9137 33303
rect 9137 33269 9171 33303
rect 9171 33269 9180 33303
rect 9128 33260 9180 33269
rect 9588 33260 9640 33312
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 4988 33099 5040 33108
rect 4988 33065 4997 33099
rect 4997 33065 5031 33099
rect 5031 33065 5040 33099
rect 4988 33056 5040 33065
rect 6644 33099 6696 33108
rect 6644 33065 6653 33099
rect 6653 33065 6687 33099
rect 6687 33065 6696 33099
rect 6644 33056 6696 33065
rect 9312 33056 9364 33108
rect 5264 32988 5316 33040
rect 5540 32988 5592 33040
rect 5724 32988 5776 33040
rect 6736 32988 6788 33040
rect 10784 33056 10836 33108
rect 11428 33099 11480 33108
rect 11428 33065 11437 33099
rect 11437 33065 11471 33099
rect 11471 33065 11480 33099
rect 11428 33056 11480 33065
rect 9496 32988 9548 33040
rect 10048 32988 10100 33040
rect 12164 32988 12216 33040
rect 2688 32963 2740 32972
rect 2688 32929 2697 32963
rect 2697 32929 2731 32963
rect 2731 32929 2740 32963
rect 2688 32920 2740 32929
rect 2872 32920 2924 32972
rect 8668 32920 8720 32972
rect 9404 32963 9456 32972
rect 9404 32929 9413 32963
rect 9413 32929 9447 32963
rect 9447 32929 9456 32963
rect 9404 32920 9456 32929
rect 10600 32920 10652 32972
rect 11612 32920 11664 32972
rect 5448 32852 5500 32904
rect 5632 32895 5684 32904
rect 5632 32861 5641 32895
rect 5641 32861 5675 32895
rect 5675 32861 5684 32895
rect 5632 32852 5684 32861
rect 5908 32852 5960 32904
rect 7104 32852 7156 32904
rect 10324 32895 10376 32904
rect 3516 32716 3568 32768
rect 9128 32784 9180 32836
rect 10324 32861 10333 32895
rect 10333 32861 10367 32895
rect 10367 32861 10376 32895
rect 10324 32852 10376 32861
rect 11520 32852 11572 32904
rect 9956 32784 10008 32836
rect 7656 32759 7708 32768
rect 7656 32725 7665 32759
rect 7665 32725 7699 32759
rect 7699 32725 7708 32759
rect 7656 32716 7708 32725
rect 8024 32716 8076 32768
rect 9312 32716 9364 32768
rect 11520 32716 11572 32768
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 2872 32555 2924 32564
rect 2872 32521 2881 32555
rect 2881 32521 2915 32555
rect 2915 32521 2924 32555
rect 2872 32512 2924 32521
rect 9956 32555 10008 32564
rect 9956 32521 9965 32555
rect 9965 32521 9999 32555
rect 9999 32521 10008 32555
rect 9956 32512 10008 32521
rect 11612 32555 11664 32564
rect 11612 32521 11621 32555
rect 11621 32521 11655 32555
rect 11655 32521 11664 32555
rect 11612 32512 11664 32521
rect 12164 32555 12216 32564
rect 12164 32521 12173 32555
rect 12173 32521 12207 32555
rect 12207 32521 12216 32555
rect 12164 32512 12216 32521
rect 6644 32444 6696 32496
rect 7840 32419 7892 32428
rect 7840 32385 7849 32419
rect 7849 32385 7883 32419
rect 7883 32385 7892 32419
rect 7840 32376 7892 32385
rect 4804 32308 4856 32360
rect 7196 32283 7248 32292
rect 2688 32172 2740 32224
rect 3240 32172 3292 32224
rect 4712 32215 4764 32224
rect 4712 32181 4721 32215
rect 4721 32181 4755 32215
rect 4755 32181 4764 32215
rect 4712 32172 4764 32181
rect 5264 32215 5316 32224
rect 5264 32181 5273 32215
rect 5273 32181 5307 32215
rect 5307 32181 5316 32215
rect 5264 32172 5316 32181
rect 5908 32215 5960 32224
rect 5908 32181 5917 32215
rect 5917 32181 5951 32215
rect 5951 32181 5960 32215
rect 5908 32172 5960 32181
rect 6644 32215 6696 32224
rect 6644 32181 6653 32215
rect 6653 32181 6687 32215
rect 6687 32181 6696 32215
rect 6644 32172 6696 32181
rect 7196 32249 7205 32283
rect 7205 32249 7239 32283
rect 7239 32249 7248 32283
rect 7196 32240 7248 32249
rect 7656 32240 7708 32292
rect 8760 32444 8812 32496
rect 8944 32376 8996 32428
rect 11428 32376 11480 32428
rect 9864 32308 9916 32360
rect 10416 32351 10468 32360
rect 10416 32317 10425 32351
rect 10425 32317 10459 32351
rect 10459 32317 10468 32351
rect 10416 32308 10468 32317
rect 12164 32308 12216 32360
rect 12900 32351 12952 32360
rect 12900 32317 12909 32351
rect 12909 32317 12943 32351
rect 12943 32317 12952 32351
rect 12900 32308 12952 32317
rect 9312 32240 9364 32292
rect 8668 32172 8720 32224
rect 10508 32172 10560 32224
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 2780 32011 2832 32020
rect 2780 31977 2789 32011
rect 2789 31977 2823 32011
rect 2823 31977 2832 32011
rect 2780 31968 2832 31977
rect 5264 31968 5316 32020
rect 5540 31968 5592 32020
rect 8944 32011 8996 32020
rect 8944 31977 8953 32011
rect 8953 31977 8987 32011
rect 8987 31977 8996 32011
rect 8944 31968 8996 31977
rect 9496 32011 9548 32020
rect 9496 31977 9505 32011
rect 9505 31977 9539 32011
rect 9539 31977 9548 32011
rect 9496 31968 9548 31977
rect 10416 31968 10468 32020
rect 4712 31900 4764 31952
rect 7012 31943 7064 31952
rect 7012 31909 7021 31943
rect 7021 31909 7055 31943
rect 7055 31909 7064 31943
rect 7012 31900 7064 31909
rect 9588 31900 9640 31952
rect 10508 31900 10560 31952
rect 2596 31875 2648 31884
rect 2596 31841 2605 31875
rect 2605 31841 2639 31875
rect 2639 31841 2648 31875
rect 2596 31832 2648 31841
rect 8392 31875 8444 31884
rect 8392 31841 8401 31875
rect 8401 31841 8435 31875
rect 8435 31841 8444 31875
rect 8392 31832 8444 31841
rect 11520 31875 11572 31884
rect 11520 31841 11529 31875
rect 11529 31841 11563 31875
rect 11563 31841 11572 31875
rect 11520 31832 11572 31841
rect 11704 31875 11756 31884
rect 11704 31841 11713 31875
rect 11713 31841 11747 31875
rect 11747 31841 11756 31875
rect 11704 31832 11756 31841
rect 12900 31832 12952 31884
rect 4252 31807 4304 31816
rect 4252 31773 4261 31807
rect 4261 31773 4295 31807
rect 4295 31773 4304 31807
rect 4252 31764 4304 31773
rect 8024 31764 8076 31816
rect 9404 31764 9456 31816
rect 7196 31696 7248 31748
rect 10324 31739 10376 31748
rect 10324 31705 10333 31739
rect 10333 31705 10367 31739
rect 10367 31705 10376 31739
rect 10324 31696 10376 31705
rect 5172 31671 5224 31680
rect 5172 31637 5181 31671
rect 5181 31637 5215 31671
rect 5215 31637 5224 31671
rect 5172 31628 5224 31637
rect 7840 31671 7892 31680
rect 7840 31637 7849 31671
rect 7849 31637 7883 31671
rect 7883 31637 7892 31671
rect 7840 31628 7892 31637
rect 7932 31628 7984 31680
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 2596 31467 2648 31476
rect 2596 31433 2605 31467
rect 2605 31433 2639 31467
rect 2639 31433 2648 31467
rect 2596 31424 2648 31433
rect 4712 31424 4764 31476
rect 7012 31424 7064 31476
rect 8024 31424 8076 31476
rect 8484 31424 8536 31476
rect 9588 31467 9640 31476
rect 9588 31433 9597 31467
rect 9597 31433 9631 31467
rect 9631 31433 9640 31467
rect 9588 31424 9640 31433
rect 5632 31399 5684 31408
rect 5632 31365 5641 31399
rect 5641 31365 5675 31399
rect 5675 31365 5684 31399
rect 5632 31356 5684 31365
rect 6736 31356 6788 31408
rect 11520 31424 11572 31476
rect 10324 31399 10376 31408
rect 10324 31365 10333 31399
rect 10333 31365 10367 31399
rect 10367 31365 10376 31399
rect 10324 31356 10376 31365
rect 4252 31288 4304 31340
rect 5172 31288 5224 31340
rect 3240 31127 3292 31136
rect 3240 31093 3249 31127
rect 3249 31093 3283 31127
rect 3283 31093 3292 31127
rect 3516 31220 3568 31272
rect 3240 31084 3292 31093
rect 4436 31084 4488 31136
rect 5264 31152 5316 31204
rect 7932 31288 7984 31340
rect 8484 31220 8536 31272
rect 5632 31084 5684 31136
rect 9128 31152 9180 31204
rect 9772 31195 9824 31204
rect 9772 31161 9781 31195
rect 9781 31161 9815 31195
rect 9815 31161 9824 31195
rect 9772 31152 9824 31161
rect 9864 31195 9916 31204
rect 9864 31161 9873 31195
rect 9873 31161 9907 31195
rect 9907 31161 9916 31195
rect 9864 31152 9916 31161
rect 8392 31127 8444 31136
rect 8392 31093 8401 31127
rect 8401 31093 8435 31127
rect 8435 31093 8444 31127
rect 8392 31084 8444 31093
rect 8944 31084 8996 31136
rect 9312 31084 9364 31136
rect 11704 31152 11756 31204
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 2964 30880 3016 30932
rect 3516 30923 3568 30932
rect 3516 30889 3525 30923
rect 3525 30889 3559 30923
rect 3559 30889 3568 30923
rect 3516 30880 3568 30889
rect 4068 30880 4120 30932
rect 4436 30923 4488 30932
rect 4436 30889 4445 30923
rect 4445 30889 4479 30923
rect 4479 30889 4488 30923
rect 4436 30880 4488 30889
rect 5908 30880 5960 30932
rect 7932 30880 7984 30932
rect 4344 30812 4396 30864
rect 5172 30812 5224 30864
rect 8208 30855 8260 30864
rect 8208 30821 8217 30855
rect 8217 30821 8251 30855
rect 8251 30821 8260 30855
rect 8208 30812 8260 30821
rect 8944 30812 8996 30864
rect 9496 30812 9548 30864
rect 10508 30812 10560 30864
rect 6736 30787 6788 30796
rect 6736 30753 6745 30787
rect 6745 30753 6779 30787
rect 6779 30753 6788 30787
rect 6736 30744 6788 30753
rect 7104 30744 7156 30796
rect 9128 30787 9180 30796
rect 9128 30753 9137 30787
rect 9137 30753 9171 30787
rect 9171 30753 9180 30787
rect 9128 30744 9180 30753
rect 10968 30744 11020 30796
rect 3148 30608 3200 30660
rect 5540 30651 5592 30660
rect 5540 30617 5549 30651
rect 5549 30617 5583 30651
rect 5583 30617 5592 30651
rect 5540 30608 5592 30617
rect 9772 30676 9824 30728
rect 10416 30676 10468 30728
rect 9404 30583 9456 30592
rect 9404 30549 9413 30583
rect 9413 30549 9447 30583
rect 9447 30549 9456 30583
rect 9404 30540 9456 30549
rect 9588 30540 9640 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 4344 30379 4396 30388
rect 4344 30345 4353 30379
rect 4353 30345 4387 30379
rect 4387 30345 4396 30379
rect 4344 30336 4396 30345
rect 6092 30200 6144 30252
rect 7104 30336 7156 30388
rect 9496 30379 9548 30388
rect 9496 30345 9505 30379
rect 9505 30345 9539 30379
rect 9539 30345 9548 30379
rect 9496 30336 9548 30345
rect 10508 30379 10560 30388
rect 10508 30345 10517 30379
rect 10517 30345 10551 30379
rect 10551 30345 10560 30379
rect 10508 30336 10560 30345
rect 10968 30336 11020 30388
rect 9588 30268 9640 30320
rect 7380 30200 7432 30252
rect 8668 30200 8720 30252
rect 6184 30132 6236 30184
rect 8484 30132 8536 30184
rect 5908 30107 5960 30116
rect 5908 30073 5917 30107
rect 5917 30073 5951 30107
rect 5951 30073 5960 30107
rect 5908 30064 5960 30073
rect 3332 29996 3384 30048
rect 3976 29996 4028 30048
rect 4988 30039 5040 30048
rect 4988 30005 4997 30039
rect 4997 30005 5031 30039
rect 5031 30005 5040 30039
rect 4988 29996 5040 30005
rect 7196 29996 7248 30048
rect 7656 29996 7708 30048
rect 8852 30039 8904 30048
rect 8852 30005 8861 30039
rect 8861 30005 8895 30039
rect 8895 30005 8904 30039
rect 8852 29996 8904 30005
rect 10048 29996 10100 30048
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 1584 29835 1636 29844
rect 1584 29801 1593 29835
rect 1593 29801 1627 29835
rect 1627 29801 1636 29835
rect 1584 29792 1636 29801
rect 5908 29792 5960 29844
rect 6828 29835 6880 29844
rect 6828 29801 6837 29835
rect 6837 29801 6871 29835
rect 6871 29801 6880 29835
rect 6828 29792 6880 29801
rect 8208 29792 8260 29844
rect 8852 29792 8904 29844
rect 12440 29792 12492 29844
rect 3976 29724 4028 29776
rect 5632 29767 5684 29776
rect 5632 29733 5641 29767
rect 5641 29733 5675 29767
rect 5675 29733 5684 29767
rect 5632 29724 5684 29733
rect 6736 29724 6788 29776
rect 7104 29724 7156 29776
rect 8760 29724 8812 29776
rect 9864 29767 9916 29776
rect 9864 29733 9873 29767
rect 9873 29733 9907 29767
rect 9907 29733 9916 29767
rect 9864 29724 9916 29733
rect 1400 29699 1452 29708
rect 1400 29665 1409 29699
rect 1409 29665 1443 29699
rect 1443 29665 1452 29699
rect 1400 29656 1452 29665
rect 8208 29656 8260 29708
rect 8392 29656 8444 29708
rect 12072 29699 12124 29708
rect 12072 29665 12081 29699
rect 12081 29665 12115 29699
rect 12115 29665 12124 29699
rect 12072 29656 12124 29665
rect 3424 29452 3476 29504
rect 7472 29588 7524 29640
rect 11152 29588 11204 29640
rect 9404 29520 9456 29572
rect 10324 29563 10376 29572
rect 10324 29529 10333 29563
rect 10333 29529 10367 29563
rect 10367 29529 10376 29563
rect 10324 29520 10376 29529
rect 8484 29495 8536 29504
rect 8484 29461 8493 29495
rect 8493 29461 8527 29495
rect 8527 29461 8536 29495
rect 8484 29452 8536 29461
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 4160 29248 4212 29300
rect 9864 29248 9916 29300
rect 11152 29291 11204 29300
rect 11152 29257 11161 29291
rect 11161 29257 11195 29291
rect 11195 29257 11204 29291
rect 11152 29248 11204 29257
rect 7840 29180 7892 29232
rect 8300 29180 8352 29232
rect 8760 29180 8812 29232
rect 2596 29112 2648 29164
rect 3056 29112 3108 29164
rect 3884 29112 3936 29164
rect 4068 29112 4120 29164
rect 6828 29155 6880 29164
rect 6828 29121 6837 29155
rect 6837 29121 6871 29155
rect 6871 29121 6880 29155
rect 6828 29112 6880 29121
rect 7196 29112 7248 29164
rect 8944 29112 8996 29164
rect 10048 29112 10100 29164
rect 10416 29112 10468 29164
rect 5264 29019 5316 29028
rect 5264 28985 5273 29019
rect 5273 28985 5307 29019
rect 5307 28985 5316 29019
rect 5264 28976 5316 28985
rect 1400 28908 1452 28960
rect 3516 28908 3568 28960
rect 3976 28951 4028 28960
rect 3976 28917 3985 28951
rect 3985 28917 4019 28951
rect 4019 28917 4028 28951
rect 3976 28908 4028 28917
rect 7012 28976 7064 29028
rect 6644 28951 6696 28960
rect 6644 28917 6653 28951
rect 6653 28917 6687 28951
rect 6687 28917 6696 28951
rect 7656 28976 7708 29028
rect 6644 28908 6696 28917
rect 8208 28908 8260 28960
rect 9956 28951 10008 28960
rect 9956 28917 9965 28951
rect 9965 28917 9999 28951
rect 9999 28917 10008 28951
rect 9956 28908 10008 28917
rect 12072 28908 12124 28960
rect 12624 28908 12676 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 3148 28747 3200 28756
rect 3148 28713 3157 28747
rect 3157 28713 3191 28747
rect 3191 28713 3200 28747
rect 3148 28704 3200 28713
rect 5264 28704 5316 28756
rect 6644 28704 6696 28756
rect 7012 28704 7064 28756
rect 7472 28747 7524 28756
rect 5080 28636 5132 28688
rect 7472 28713 7481 28747
rect 7481 28713 7515 28747
rect 7515 28713 7524 28747
rect 7472 28704 7524 28713
rect 8944 28747 8996 28756
rect 8944 28713 8953 28747
rect 8953 28713 8987 28747
rect 8987 28713 8996 28747
rect 8944 28704 8996 28713
rect 10048 28704 10100 28756
rect 11152 28704 11204 28756
rect 9864 28679 9916 28688
rect 9864 28645 9873 28679
rect 9873 28645 9907 28679
rect 9907 28645 9916 28679
rect 9864 28636 9916 28645
rect 10416 28679 10468 28688
rect 10416 28645 10425 28679
rect 10425 28645 10459 28679
rect 10459 28645 10468 28679
rect 10416 28636 10468 28645
rect 112 28568 164 28620
rect 2872 28611 2924 28620
rect 2872 28577 2881 28611
rect 2881 28577 2915 28611
rect 2915 28577 2924 28611
rect 2872 28568 2924 28577
rect 11244 28611 11296 28620
rect 11244 28577 11253 28611
rect 11253 28577 11287 28611
rect 11287 28577 11296 28611
rect 11244 28568 11296 28577
rect 12624 28568 12676 28620
rect 2412 28500 2464 28552
rect 4712 28543 4764 28552
rect 4712 28509 4721 28543
rect 4721 28509 4755 28543
rect 4755 28509 4764 28543
rect 4712 28500 4764 28509
rect 6644 28500 6696 28552
rect 7656 28500 7708 28552
rect 8300 28543 8352 28552
rect 8300 28509 8309 28543
rect 8309 28509 8343 28543
rect 8343 28509 8352 28543
rect 8300 28500 8352 28509
rect 3884 28432 3936 28484
rect 4068 28432 4120 28484
rect 5540 28432 5592 28484
rect 6920 28432 6972 28484
rect 3516 28364 3568 28416
rect 6000 28364 6052 28416
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 2412 28203 2464 28212
rect 2412 28169 2421 28203
rect 2421 28169 2455 28203
rect 2455 28169 2464 28203
rect 2412 28160 2464 28169
rect 3424 28203 3476 28212
rect 3424 28169 3433 28203
rect 3433 28169 3467 28203
rect 3467 28169 3476 28203
rect 3424 28160 3476 28169
rect 4712 28160 4764 28212
rect 9496 28160 9548 28212
rect 9864 28160 9916 28212
rect 3332 28092 3384 28144
rect 6184 28092 6236 28144
rect 11244 28135 11296 28144
rect 11244 28101 11253 28135
rect 11253 28101 11287 28135
rect 11287 28101 11296 28135
rect 11244 28092 11296 28101
rect 4528 28024 4580 28076
rect 3332 27956 3384 28008
rect 4252 27956 4304 28008
rect 2688 27888 2740 27940
rect 4988 27956 5040 28008
rect 5540 27956 5592 28008
rect 8852 27956 8904 28008
rect 2872 27820 2924 27872
rect 3884 27820 3936 27872
rect 4712 27888 4764 27940
rect 6552 27888 6604 27940
rect 5080 27863 5132 27872
rect 5080 27829 5089 27863
rect 5089 27829 5123 27863
rect 5123 27829 5132 27863
rect 5080 27820 5132 27829
rect 6644 27863 6696 27872
rect 6644 27829 6653 27863
rect 6653 27829 6687 27863
rect 6687 27829 6696 27863
rect 6644 27820 6696 27829
rect 7656 27888 7708 27940
rect 8024 27820 8076 27872
rect 9864 27820 9916 27872
rect 12624 27863 12676 27872
rect 12624 27829 12633 27863
rect 12633 27829 12667 27863
rect 12667 27829 12676 27863
rect 12624 27820 12676 27829
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 4988 27616 5040 27668
rect 7656 27659 7708 27668
rect 4712 27591 4764 27600
rect 4712 27557 4721 27591
rect 4721 27557 4755 27591
rect 4755 27557 4764 27591
rect 4712 27548 4764 27557
rect 2688 27523 2740 27532
rect 2688 27489 2697 27523
rect 2697 27489 2731 27523
rect 2731 27489 2740 27523
rect 2688 27480 2740 27489
rect 2964 27523 3016 27532
rect 2964 27489 2973 27523
rect 2973 27489 3007 27523
rect 3007 27489 3016 27523
rect 2964 27480 3016 27489
rect 3976 27480 4028 27532
rect 6276 27548 6328 27600
rect 6920 27591 6972 27600
rect 6920 27557 6929 27591
rect 6929 27557 6963 27591
rect 6963 27557 6972 27591
rect 6920 27548 6972 27557
rect 7656 27625 7665 27659
rect 7665 27625 7699 27659
rect 7699 27625 7708 27659
rect 7656 27616 7708 27625
rect 9496 27659 9548 27668
rect 9496 27625 9505 27659
rect 9505 27625 9539 27659
rect 9539 27625 9548 27659
rect 9496 27616 9548 27625
rect 8484 27591 8536 27600
rect 8484 27557 8493 27591
rect 8493 27557 8527 27591
rect 8527 27557 8536 27591
rect 8484 27548 8536 27557
rect 9864 27591 9916 27600
rect 9864 27557 9873 27591
rect 9873 27557 9907 27591
rect 9907 27557 9916 27591
rect 9864 27548 9916 27557
rect 7748 27523 7800 27532
rect 7748 27489 7757 27523
rect 7757 27489 7791 27523
rect 7791 27489 7800 27523
rect 7748 27480 7800 27489
rect 7840 27480 7892 27532
rect 4436 27455 4488 27464
rect 4436 27421 4445 27455
rect 4445 27421 4479 27455
rect 4479 27421 4488 27455
rect 4436 27412 4488 27421
rect 6000 27412 6052 27464
rect 10232 27412 10284 27464
rect 3424 27344 3476 27396
rect 6736 27344 6788 27396
rect 10324 27387 10376 27396
rect 10324 27353 10333 27387
rect 10333 27353 10367 27387
rect 10367 27353 10376 27387
rect 10324 27344 10376 27353
rect 3148 27276 3200 27328
rect 4252 27319 4304 27328
rect 4252 27285 4261 27319
rect 4261 27285 4295 27319
rect 4295 27285 4304 27319
rect 4252 27276 4304 27285
rect 8852 27319 8904 27328
rect 8852 27285 8861 27319
rect 8861 27285 8895 27319
rect 8895 27285 8904 27319
rect 8852 27276 8904 27285
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 2688 27115 2740 27124
rect 2688 27081 2697 27115
rect 2697 27081 2731 27115
rect 2731 27081 2740 27115
rect 2688 27072 2740 27081
rect 5724 27072 5776 27124
rect 6276 27115 6328 27124
rect 6276 27081 6285 27115
rect 6285 27081 6319 27115
rect 6319 27081 6328 27115
rect 6276 27072 6328 27081
rect 6736 27072 6788 27124
rect 9864 27115 9916 27124
rect 4068 27004 4120 27056
rect 4252 26936 4304 26988
rect 6000 27004 6052 27056
rect 7748 27004 7800 27056
rect 8024 26979 8076 26988
rect 8024 26945 8033 26979
rect 8033 26945 8067 26979
rect 8067 26945 8076 26979
rect 8024 26936 8076 26945
rect 1860 26732 1912 26784
rect 2964 26800 3016 26852
rect 3516 26800 3568 26852
rect 4620 26800 4672 26852
rect 5080 26800 5132 26852
rect 2320 26775 2372 26784
rect 2320 26741 2329 26775
rect 2329 26741 2363 26775
rect 2363 26741 2372 26775
rect 2320 26732 2372 26741
rect 4712 26732 4764 26784
rect 5816 26732 5868 26784
rect 7748 26911 7800 26920
rect 7748 26877 7757 26911
rect 7757 26877 7791 26911
rect 7791 26877 7800 26911
rect 7748 26868 7800 26877
rect 8300 26868 8352 26920
rect 9864 27081 9873 27115
rect 9873 27081 9907 27115
rect 9907 27081 9916 27115
rect 9864 27072 9916 27081
rect 10232 27115 10284 27124
rect 10232 27081 10241 27115
rect 10241 27081 10275 27115
rect 10275 27081 10284 27115
rect 10232 27072 10284 27081
rect 9312 26911 9364 26920
rect 9312 26877 9321 26911
rect 9321 26877 9355 26911
rect 9355 26877 9364 26911
rect 9312 26868 9364 26877
rect 8852 26732 8904 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 4252 26528 4304 26580
rect 4436 26528 4488 26580
rect 7288 26571 7340 26580
rect 7288 26537 7297 26571
rect 7297 26537 7331 26571
rect 7331 26537 7340 26571
rect 7288 26528 7340 26537
rect 7748 26528 7800 26580
rect 8852 26528 8904 26580
rect 3516 26503 3568 26512
rect 3516 26469 3525 26503
rect 3525 26469 3559 26503
rect 3559 26469 3568 26503
rect 4804 26503 4856 26512
rect 3516 26460 3568 26469
rect 3332 26392 3384 26444
rect 4344 26435 4396 26444
rect 4344 26401 4353 26435
rect 4353 26401 4387 26435
rect 4387 26401 4396 26435
rect 4344 26392 4396 26401
rect 4804 26469 4813 26503
rect 4813 26469 4847 26503
rect 4847 26469 4856 26503
rect 4804 26460 4856 26469
rect 6644 26460 6696 26512
rect 4896 26392 4948 26444
rect 5724 26435 5776 26444
rect 5724 26401 5733 26435
rect 5733 26401 5767 26435
rect 5767 26401 5776 26435
rect 5724 26392 5776 26401
rect 6092 26435 6144 26444
rect 6092 26401 6101 26435
rect 6101 26401 6135 26435
rect 6135 26401 6144 26435
rect 6092 26392 6144 26401
rect 8024 26435 8076 26444
rect 8024 26401 8033 26435
rect 8033 26401 8067 26435
rect 8067 26401 8076 26435
rect 8024 26392 8076 26401
rect 8116 26392 8168 26444
rect 9680 26435 9732 26444
rect 9680 26401 9689 26435
rect 9689 26401 9723 26435
rect 9723 26401 9732 26435
rect 9680 26392 9732 26401
rect 10324 26392 10376 26444
rect 11520 26392 11572 26444
rect 2320 26324 2372 26376
rect 8576 26367 8628 26376
rect 8576 26333 8585 26367
rect 8585 26333 8619 26367
rect 8619 26333 8628 26367
rect 8576 26324 8628 26333
rect 11428 26324 11480 26376
rect 4620 26256 4672 26308
rect 7748 26256 7800 26308
rect 9312 26256 9364 26308
rect 10784 26231 10836 26240
rect 10784 26197 10793 26231
rect 10793 26197 10827 26231
rect 10827 26197 10836 26231
rect 10784 26188 10836 26197
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 4620 25984 4672 26036
rect 4896 26027 4948 26036
rect 4896 25993 4905 26027
rect 4905 25993 4939 26027
rect 4939 25993 4948 26027
rect 4896 25984 4948 25993
rect 6092 26027 6144 26036
rect 6092 25993 6101 26027
rect 6101 25993 6135 26027
rect 6135 25993 6144 26027
rect 6092 25984 6144 25993
rect 8668 25984 8720 26036
rect 9680 25984 9732 26036
rect 10324 26027 10376 26036
rect 10324 25993 10333 26027
rect 10333 25993 10367 26027
rect 10367 25993 10376 26027
rect 10324 25984 10376 25993
rect 5264 25959 5316 25968
rect 5264 25925 5273 25959
rect 5273 25925 5307 25959
rect 5307 25925 5316 25959
rect 5264 25916 5316 25925
rect 6828 25916 6880 25968
rect 4804 25848 4856 25900
rect 8024 25848 8076 25900
rect 10784 25848 10836 25900
rect 3424 25780 3476 25832
rect 5080 25823 5132 25832
rect 5080 25789 5089 25823
rect 5089 25789 5123 25823
rect 5123 25789 5132 25823
rect 5080 25780 5132 25789
rect 6828 25780 6880 25832
rect 7196 25823 7248 25832
rect 7196 25789 7205 25823
rect 7205 25789 7239 25823
rect 7239 25789 7248 25823
rect 7196 25780 7248 25789
rect 8760 25823 8812 25832
rect 4344 25712 4396 25764
rect 8760 25789 8769 25823
rect 8769 25789 8803 25823
rect 8803 25789 8812 25823
rect 8760 25780 8812 25789
rect 10416 25780 10468 25832
rect 3332 25644 3384 25696
rect 5724 25687 5776 25696
rect 5724 25653 5733 25687
rect 5733 25653 5767 25687
rect 5767 25653 5776 25687
rect 5724 25644 5776 25653
rect 7104 25687 7156 25696
rect 7104 25653 7113 25687
rect 7113 25653 7147 25687
rect 7147 25653 7156 25687
rect 7104 25644 7156 25653
rect 7932 25644 7984 25696
rect 10692 25755 10744 25764
rect 10692 25721 10701 25755
rect 10701 25721 10735 25755
rect 10735 25721 10744 25755
rect 10692 25712 10744 25721
rect 11520 25687 11572 25696
rect 11520 25653 11529 25687
rect 11529 25653 11563 25687
rect 11563 25653 11572 25687
rect 11520 25644 11572 25653
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 4896 25440 4948 25492
rect 7104 25440 7156 25492
rect 8116 25440 8168 25492
rect 8760 25483 8812 25492
rect 8760 25449 8769 25483
rect 8769 25449 8803 25483
rect 8803 25449 8812 25483
rect 8760 25440 8812 25449
rect 9956 25440 10008 25492
rect 10692 25440 10744 25492
rect 6184 25372 6236 25424
rect 7196 25415 7248 25424
rect 7196 25381 7205 25415
rect 7205 25381 7239 25415
rect 7239 25381 7248 25415
rect 7196 25372 7248 25381
rect 7748 25372 7800 25424
rect 10416 25372 10468 25424
rect 11336 25372 11388 25424
rect 4436 25347 4488 25356
rect 4436 25313 4445 25347
rect 4445 25313 4479 25347
rect 4479 25313 4488 25347
rect 4436 25304 4488 25313
rect 8576 25304 8628 25356
rect 9404 25304 9456 25356
rect 4344 25236 4396 25288
rect 6092 25236 6144 25288
rect 7196 25236 7248 25288
rect 7288 25236 7340 25288
rect 10048 25236 10100 25288
rect 11796 25279 11848 25288
rect 11428 25168 11480 25220
rect 11796 25245 11805 25279
rect 11805 25245 11839 25279
rect 11839 25245 11848 25279
rect 11796 25236 11848 25245
rect 5080 25143 5132 25152
rect 5080 25109 5089 25143
rect 5089 25109 5123 25143
rect 5123 25109 5132 25143
rect 5080 25100 5132 25109
rect 5448 25143 5500 25152
rect 5448 25109 5457 25143
rect 5457 25109 5491 25143
rect 5491 25109 5500 25143
rect 5448 25100 5500 25109
rect 6920 25143 6972 25152
rect 6920 25109 6929 25143
rect 6929 25109 6963 25143
rect 6963 25109 6972 25143
rect 6920 25100 6972 25109
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 4344 24896 4396 24948
rect 4436 24896 4488 24948
rect 7932 24896 7984 24948
rect 3056 24828 3108 24880
rect 4068 24760 4120 24812
rect 8760 24828 8812 24880
rect 5448 24760 5500 24812
rect 7196 24803 7248 24812
rect 4160 24692 4212 24744
rect 5448 24624 5500 24676
rect 5908 24667 5960 24676
rect 5908 24633 5917 24667
rect 5917 24633 5951 24667
rect 5951 24633 5960 24667
rect 5908 24624 5960 24633
rect 6184 24599 6236 24608
rect 6184 24565 6193 24599
rect 6193 24565 6227 24599
rect 6227 24565 6236 24599
rect 6184 24556 6236 24565
rect 7196 24769 7205 24803
rect 7205 24769 7239 24803
rect 7239 24769 7248 24803
rect 7196 24760 7248 24769
rect 7288 24760 7340 24812
rect 8852 24803 8904 24812
rect 8852 24769 8861 24803
rect 8861 24769 8895 24803
rect 8895 24769 8904 24803
rect 8852 24760 8904 24769
rect 6920 24667 6972 24676
rect 6920 24633 6929 24667
rect 6929 24633 6963 24667
rect 6963 24633 6972 24667
rect 6920 24624 6972 24633
rect 9956 24896 10008 24948
rect 11336 24896 11388 24948
rect 10416 24828 10468 24880
rect 11428 24828 11480 24880
rect 11796 24760 11848 24812
rect 7748 24556 7800 24608
rect 10692 24667 10744 24676
rect 10692 24633 10701 24667
rect 10701 24633 10735 24667
rect 10735 24633 10744 24667
rect 10692 24624 10744 24633
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 6920 24352 6972 24404
rect 8852 24395 8904 24404
rect 8852 24361 8861 24395
rect 8861 24361 8895 24395
rect 8895 24361 8904 24395
rect 8852 24352 8904 24361
rect 9404 24395 9456 24404
rect 9404 24361 9413 24395
rect 9413 24361 9447 24395
rect 9447 24361 9456 24395
rect 9404 24352 9456 24361
rect 14832 24352 14884 24404
rect 4436 24284 4488 24336
rect 4712 24284 4764 24336
rect 5816 24284 5868 24336
rect 9864 24327 9916 24336
rect 9864 24293 9873 24327
rect 9873 24293 9907 24327
rect 9907 24293 9916 24327
rect 9864 24284 9916 24293
rect 3240 24216 3292 24268
rect 6092 24259 6144 24268
rect 6092 24225 6101 24259
rect 6101 24225 6135 24259
rect 6135 24225 6144 24259
rect 6092 24216 6144 24225
rect 8024 24216 8076 24268
rect 11244 24259 11296 24268
rect 11244 24225 11253 24259
rect 11253 24225 11287 24259
rect 11287 24225 11296 24259
rect 11244 24216 11296 24225
rect 3516 24055 3568 24064
rect 3516 24021 3525 24055
rect 3525 24021 3559 24055
rect 3559 24021 3568 24055
rect 3516 24012 3568 24021
rect 4344 24012 4396 24064
rect 7840 24148 7892 24200
rect 8760 24148 8812 24200
rect 9772 24191 9824 24200
rect 9772 24157 9781 24191
rect 9781 24157 9815 24191
rect 9815 24157 9824 24191
rect 9772 24148 9824 24157
rect 10048 24191 10100 24200
rect 10048 24157 10057 24191
rect 10057 24157 10091 24191
rect 10091 24157 10100 24191
rect 10048 24148 10100 24157
rect 5908 24080 5960 24132
rect 7288 24123 7340 24132
rect 7288 24089 7297 24123
rect 7297 24089 7331 24123
rect 7331 24089 7340 24123
rect 7288 24080 7340 24089
rect 5816 24055 5868 24064
rect 5816 24021 5825 24055
rect 5825 24021 5859 24055
rect 5859 24021 5868 24055
rect 5816 24012 5868 24021
rect 6920 24012 6972 24064
rect 7656 24012 7708 24064
rect 9956 24012 10008 24064
rect 10692 24055 10744 24064
rect 10692 24021 10701 24055
rect 10701 24021 10735 24055
rect 10735 24021 10744 24055
rect 10692 24012 10744 24021
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 4160 23808 4212 23860
rect 5540 23808 5592 23860
rect 5816 23808 5868 23860
rect 8576 23808 8628 23860
rect 9404 23808 9456 23860
rect 9864 23808 9916 23860
rect 3240 23740 3292 23792
rect 5448 23740 5500 23792
rect 9772 23740 9824 23792
rect 6920 23715 6972 23724
rect 6920 23681 6929 23715
rect 6929 23681 6963 23715
rect 6963 23681 6972 23715
rect 6920 23672 6972 23681
rect 7288 23715 7340 23724
rect 7288 23681 7297 23715
rect 7297 23681 7331 23715
rect 7331 23681 7340 23715
rect 7288 23672 7340 23681
rect 8484 23715 8536 23724
rect 8484 23681 8493 23715
rect 8493 23681 8527 23715
rect 8527 23681 8536 23715
rect 8484 23672 8536 23681
rect 8760 23715 8812 23724
rect 8760 23681 8769 23715
rect 8769 23681 8803 23715
rect 8803 23681 8812 23715
rect 8760 23672 8812 23681
rect 10048 23672 10100 23724
rect 11244 23672 11296 23724
rect 3056 23604 3108 23656
rect 3240 23604 3292 23656
rect 3516 23604 3568 23656
rect 3608 23536 3660 23588
rect 4896 23604 4948 23656
rect 5816 23604 5868 23656
rect 4436 23511 4488 23520
rect 4436 23477 4445 23511
rect 4445 23477 4479 23511
rect 4479 23477 4488 23511
rect 4436 23468 4488 23477
rect 5172 23468 5224 23520
rect 5540 23468 5592 23520
rect 6184 23468 6236 23520
rect 8576 23579 8628 23588
rect 8576 23545 8585 23579
rect 8585 23545 8619 23579
rect 8619 23545 8628 23579
rect 8576 23536 8628 23545
rect 8024 23468 8076 23520
rect 9680 23468 9732 23520
rect 10140 23579 10192 23588
rect 10140 23545 10149 23579
rect 10149 23545 10183 23579
rect 10183 23545 10192 23579
rect 10140 23536 10192 23545
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 5540 23307 5592 23316
rect 3516 23239 3568 23248
rect 3516 23205 3525 23239
rect 3525 23205 3559 23239
rect 3559 23205 3568 23239
rect 3516 23196 3568 23205
rect 4436 23196 4488 23248
rect 5172 23196 5224 23248
rect 5540 23273 5549 23307
rect 5549 23273 5583 23307
rect 5583 23273 5592 23307
rect 5540 23264 5592 23273
rect 5816 23307 5868 23316
rect 5816 23273 5825 23307
rect 5825 23273 5859 23307
rect 5859 23273 5868 23307
rect 5816 23264 5868 23273
rect 7656 23307 7708 23316
rect 7656 23273 7665 23307
rect 7665 23273 7699 23307
rect 7699 23273 7708 23307
rect 7656 23264 7708 23273
rect 7840 23264 7892 23316
rect 8484 23264 8536 23316
rect 9680 23307 9732 23316
rect 9680 23273 9689 23307
rect 9689 23273 9723 23307
rect 9723 23273 9732 23307
rect 9680 23264 9732 23273
rect 5632 23196 5684 23248
rect 6552 23196 6604 23248
rect 112 23128 164 23180
rect 2872 23171 2924 23180
rect 2872 23137 2881 23171
rect 2881 23137 2915 23171
rect 2915 23137 2924 23171
rect 2872 23128 2924 23137
rect 3056 23128 3108 23180
rect 3332 23128 3384 23180
rect 3424 23128 3476 23180
rect 8024 23196 8076 23248
rect 8116 23171 8168 23180
rect 8116 23137 8125 23171
rect 8125 23137 8159 23171
rect 8159 23137 8168 23171
rect 8116 23128 8168 23137
rect 10692 23171 10744 23180
rect 10692 23137 10701 23171
rect 10701 23137 10735 23171
rect 10735 23137 10744 23171
rect 10692 23128 10744 23137
rect 3424 22924 3476 22976
rect 4068 22924 4120 22976
rect 4528 22967 4580 22976
rect 4528 22933 4537 22967
rect 4537 22933 4571 22967
rect 4571 22933 4580 22967
rect 4528 22924 4580 22933
rect 5908 22924 5960 22976
rect 7932 23060 7984 23112
rect 9404 22992 9456 23044
rect 10140 22967 10192 22976
rect 10140 22933 10149 22967
rect 10149 22933 10183 22967
rect 10183 22933 10192 22967
rect 10140 22924 10192 22933
rect 10232 22924 10284 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 2872 22763 2924 22772
rect 2872 22729 2881 22763
rect 2881 22729 2915 22763
rect 2915 22729 2924 22763
rect 2872 22720 2924 22729
rect 3516 22763 3568 22772
rect 3516 22729 3525 22763
rect 3525 22729 3559 22763
rect 3559 22729 3568 22763
rect 3516 22720 3568 22729
rect 3884 22559 3936 22568
rect 3884 22525 3893 22559
rect 3893 22525 3927 22559
rect 3927 22525 3936 22559
rect 3884 22516 3936 22525
rect 10140 22720 10192 22772
rect 10692 22763 10744 22772
rect 10692 22729 10701 22763
rect 10701 22729 10735 22763
rect 10735 22729 10744 22763
rect 10692 22720 10744 22729
rect 4344 22627 4396 22636
rect 4344 22593 4353 22627
rect 4353 22593 4387 22627
rect 4387 22593 4396 22627
rect 4344 22584 4396 22593
rect 5172 22584 5224 22636
rect 5908 22627 5960 22636
rect 5264 22559 5316 22568
rect 2872 22448 2924 22500
rect 5264 22525 5273 22559
rect 5273 22525 5307 22559
rect 5307 22525 5316 22559
rect 5264 22516 5316 22525
rect 5908 22593 5917 22627
rect 5917 22593 5951 22627
rect 5951 22593 5960 22627
rect 5908 22584 5960 22593
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 10232 22584 10284 22636
rect 6828 22559 6880 22568
rect 6828 22525 6837 22559
rect 6837 22525 6871 22559
rect 6871 22525 6880 22559
rect 6828 22516 6880 22525
rect 11520 22516 11572 22568
rect 6552 22448 6604 22500
rect 8484 22448 8536 22500
rect 5172 22380 5224 22432
rect 7932 22380 7984 22432
rect 9772 22448 9824 22500
rect 10232 22448 10284 22500
rect 10784 22380 10836 22432
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 2688 22176 2740 22228
rect 4528 22219 4580 22228
rect 4528 22185 4537 22219
rect 4537 22185 4571 22219
rect 4571 22185 4580 22219
rect 4528 22176 4580 22185
rect 5264 22176 5316 22228
rect 9404 22219 9456 22228
rect 9404 22185 9413 22219
rect 9413 22185 9447 22219
rect 9447 22185 9456 22219
rect 9404 22176 9456 22185
rect 8484 22108 8536 22160
rect 5172 22040 5224 22092
rect 6276 22083 6328 22092
rect 6276 22049 6285 22083
rect 6285 22049 6319 22083
rect 6319 22049 6328 22083
rect 6276 22040 6328 22049
rect 7104 22040 7156 22092
rect 9772 22108 9824 22160
rect 9956 22108 10008 22160
rect 10600 22108 10652 22160
rect 11244 22083 11296 22092
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 12624 22040 12676 22092
rect 7840 22015 7892 22024
rect 7840 21981 7849 22015
rect 7849 21981 7883 22015
rect 7883 21981 7892 22015
rect 7840 21972 7892 21981
rect 9496 21972 9548 22024
rect 10784 21972 10836 22024
rect 3884 21904 3936 21956
rect 5724 21904 5776 21956
rect 6644 21904 6696 21956
rect 8392 21904 8444 21956
rect 11060 21904 11112 21956
rect 5908 21836 5960 21888
rect 6828 21836 6880 21888
rect 10784 21879 10836 21888
rect 10784 21845 10793 21879
rect 10793 21845 10827 21879
rect 10827 21845 10836 21879
rect 10784 21836 10836 21845
rect 10876 21836 10928 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 6276 21675 6328 21684
rect 6276 21641 6285 21675
rect 6285 21641 6319 21675
rect 6319 21641 6328 21675
rect 6276 21632 6328 21641
rect 6828 21632 6880 21684
rect 7104 21632 7156 21684
rect 9772 21675 9824 21684
rect 9772 21641 9781 21675
rect 9781 21641 9815 21675
rect 9815 21641 9824 21675
rect 9772 21632 9824 21641
rect 4620 21564 4672 21616
rect 10416 21564 10468 21616
rect 10600 21607 10652 21616
rect 10600 21573 10609 21607
rect 10609 21573 10643 21607
rect 10643 21573 10652 21607
rect 10600 21564 10652 21573
rect 5908 21539 5960 21548
rect 5908 21505 5917 21539
rect 5917 21505 5951 21539
rect 5951 21505 5960 21539
rect 5908 21496 5960 21505
rect 10784 21496 10836 21548
rect 1492 21428 1544 21480
rect 4160 21428 4212 21480
rect 4896 21428 4948 21480
rect 5540 21428 5592 21480
rect 6736 21428 6788 21480
rect 7196 21428 7248 21480
rect 9036 21428 9088 21480
rect 8484 21360 8536 21412
rect 10140 21403 10192 21412
rect 10140 21369 10149 21403
rect 10149 21369 10183 21403
rect 10183 21369 10192 21403
rect 10140 21360 10192 21369
rect 3516 21292 3568 21344
rect 5172 21292 5224 21344
rect 8208 21292 8260 21344
rect 11244 21335 11296 21344
rect 11244 21301 11253 21335
rect 11253 21301 11287 21335
rect 11287 21301 11296 21335
rect 11244 21292 11296 21301
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 3516 21088 3568 21140
rect 7840 21131 7892 21140
rect 7840 21097 7849 21131
rect 7849 21097 7883 21131
rect 7883 21097 7892 21131
rect 7840 21088 7892 21097
rect 9036 21131 9088 21140
rect 9036 21097 9045 21131
rect 9045 21097 9079 21131
rect 9079 21097 9088 21131
rect 9036 21088 9088 21097
rect 9496 21131 9548 21140
rect 9496 21097 9505 21131
rect 9505 21097 9539 21131
rect 9539 21097 9548 21131
rect 9496 21088 9548 21097
rect 10140 21088 10192 21140
rect 10324 21088 10376 21140
rect 10784 21088 10836 21140
rect 4252 21063 4304 21072
rect 4252 21029 4261 21063
rect 4261 21029 4295 21063
rect 4295 21029 4304 21063
rect 4252 21020 4304 21029
rect 7196 21063 7248 21072
rect 6644 20995 6696 21004
rect 6644 20961 6653 20995
rect 6653 20961 6687 20995
rect 6687 20961 6696 20995
rect 6644 20952 6696 20961
rect 7196 21029 7205 21063
rect 7205 21029 7239 21063
rect 7239 21029 7248 21063
rect 7196 21020 7248 21029
rect 8208 21063 8260 21072
rect 8208 21029 8217 21063
rect 8217 21029 8251 21063
rect 8251 21029 8260 21063
rect 8208 21020 8260 21029
rect 9864 21063 9916 21072
rect 9864 21029 9873 21063
rect 9873 21029 9907 21063
rect 9907 21029 9916 21063
rect 9864 21020 9916 21029
rect 10600 21020 10652 21072
rect 7104 20952 7156 21004
rect 11060 20952 11112 21004
rect 4160 20927 4212 20936
rect 4160 20893 4169 20927
rect 4169 20893 4203 20927
rect 4203 20893 4212 20927
rect 4160 20884 4212 20893
rect 8116 20927 8168 20936
rect 8116 20893 8125 20927
rect 8125 20893 8159 20927
rect 8159 20893 8168 20927
rect 8116 20884 8168 20893
rect 8760 20927 8812 20936
rect 8760 20893 8769 20927
rect 8769 20893 8803 20927
rect 8803 20893 8812 20927
rect 8760 20884 8812 20893
rect 9496 20884 9548 20936
rect 10876 20884 10928 20936
rect 4620 20816 4672 20868
rect 5172 20791 5224 20800
rect 5172 20757 5181 20791
rect 5181 20757 5215 20791
rect 5215 20757 5224 20791
rect 5172 20748 5224 20757
rect 5540 20791 5592 20800
rect 5540 20757 5549 20791
rect 5549 20757 5583 20791
rect 5583 20757 5592 20791
rect 5540 20748 5592 20757
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 4988 20544 5040 20596
rect 5724 20544 5776 20596
rect 4160 20476 4212 20528
rect 3516 20408 3568 20460
rect 5540 20408 5592 20460
rect 1400 20340 1452 20392
rect 2780 20340 2832 20392
rect 8208 20544 8260 20596
rect 9864 20544 9916 20596
rect 8760 20408 8812 20460
rect 10232 20408 10284 20460
rect 7104 20340 7156 20392
rect 8392 20383 8444 20392
rect 8392 20349 8401 20383
rect 8401 20349 8435 20383
rect 8435 20349 8444 20383
rect 8392 20340 8444 20349
rect 4896 20272 4948 20324
rect 5356 20315 5408 20324
rect 5356 20281 5365 20315
rect 5365 20281 5399 20315
rect 5399 20281 5408 20315
rect 5356 20272 5408 20281
rect 6092 20272 6144 20324
rect 4252 20204 4304 20256
rect 4712 20247 4764 20256
rect 4712 20213 4721 20247
rect 4721 20213 4755 20247
rect 4755 20213 4764 20247
rect 4712 20204 4764 20213
rect 8484 20272 8536 20324
rect 10232 20315 10284 20324
rect 10232 20281 10241 20315
rect 10241 20281 10275 20315
rect 10275 20281 10284 20315
rect 10232 20272 10284 20281
rect 10324 20315 10376 20324
rect 10324 20281 10333 20315
rect 10333 20281 10367 20315
rect 10367 20281 10376 20315
rect 10324 20272 10376 20281
rect 6644 20204 6696 20256
rect 7012 20204 7064 20256
rect 8208 20247 8260 20256
rect 8208 20213 8217 20247
rect 8217 20213 8251 20247
rect 8251 20213 8260 20247
rect 8208 20204 8260 20213
rect 11060 20204 11112 20256
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 4160 20000 4212 20052
rect 3424 19932 3476 19984
rect 4712 20000 4764 20052
rect 5264 20000 5316 20052
rect 4896 19932 4948 19984
rect 5908 19975 5960 19984
rect 5908 19941 5917 19975
rect 5917 19941 5951 19975
rect 5951 19941 5960 19975
rect 5908 19932 5960 19941
rect 6184 19932 6236 19984
rect 7104 20000 7156 20052
rect 7472 20043 7524 20052
rect 7472 20009 7481 20043
rect 7481 20009 7515 20043
rect 7515 20009 7524 20043
rect 7472 20000 7524 20009
rect 8392 20000 8444 20052
rect 9496 20043 9548 20052
rect 9496 20009 9505 20043
rect 9505 20009 9539 20043
rect 9539 20009 9548 20043
rect 9496 20000 9548 20009
rect 10048 20000 10100 20052
rect 10232 20000 10284 20052
rect 8576 19975 8628 19984
rect 8576 19941 8585 19975
rect 8585 19941 8619 19975
rect 8619 19941 8628 19975
rect 8576 19932 8628 19941
rect 2688 19907 2740 19916
rect 2688 19873 2697 19907
rect 2697 19873 2731 19907
rect 2731 19873 2740 19907
rect 2688 19864 2740 19873
rect 2964 19907 3016 19916
rect 2964 19873 2973 19907
rect 2973 19873 3007 19907
rect 3007 19873 3016 19907
rect 2964 19864 3016 19873
rect 4988 19864 5040 19916
rect 6828 19864 6880 19916
rect 7840 19864 7892 19916
rect 8484 19864 8536 19916
rect 9588 19864 9640 19916
rect 10324 19864 10376 19916
rect 10600 19864 10652 19916
rect 2596 19796 2648 19848
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 6092 19796 6144 19848
rect 3516 19703 3568 19712
rect 3516 19669 3525 19703
rect 3525 19669 3559 19703
rect 3559 19669 3568 19703
rect 3516 19660 3568 19669
rect 8668 19660 8720 19712
rect 10324 19660 10376 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 2688 19456 2740 19508
rect 5264 19456 5316 19508
rect 5356 19456 5408 19508
rect 7748 19499 7800 19508
rect 7748 19465 7757 19499
rect 7757 19465 7791 19499
rect 7791 19465 7800 19499
rect 7748 19456 7800 19465
rect 7840 19456 7892 19508
rect 8116 19456 8168 19508
rect 3424 19388 3476 19440
rect 2596 19363 2648 19372
rect 2596 19329 2605 19363
rect 2605 19329 2639 19363
rect 2639 19329 2648 19363
rect 2596 19320 2648 19329
rect 4620 19388 4672 19440
rect 4988 19363 5040 19372
rect 1952 19252 2004 19304
rect 2964 19184 3016 19236
rect 3516 19227 3568 19236
rect 3516 19193 3525 19227
rect 3525 19193 3559 19227
rect 3559 19193 3568 19227
rect 3516 19184 3568 19193
rect 3608 19227 3660 19236
rect 3608 19193 3617 19227
rect 3617 19193 3651 19227
rect 3651 19193 3660 19227
rect 4988 19329 4997 19363
rect 4997 19329 5031 19363
rect 5031 19329 5040 19363
rect 4988 19320 5040 19329
rect 6092 19320 6144 19372
rect 9588 19363 9640 19372
rect 9588 19329 9597 19363
rect 9597 19329 9631 19363
rect 9631 19329 9640 19363
rect 9588 19320 9640 19329
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 8576 19295 8628 19304
rect 8576 19261 8585 19295
rect 8585 19261 8619 19295
rect 8619 19261 8628 19295
rect 8576 19252 8628 19261
rect 3608 19184 3660 19193
rect 5264 19184 5316 19236
rect 6184 19159 6236 19168
rect 6184 19125 6193 19159
rect 6193 19125 6227 19159
rect 6227 19125 6236 19159
rect 6184 19116 6236 19125
rect 7748 19116 7800 19168
rect 8208 19116 8260 19168
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 8668 19159 8720 19168
rect 8668 19125 8677 19159
rect 8677 19125 8711 19159
rect 8711 19125 8720 19159
rect 8668 19116 8720 19125
rect 8760 19116 8812 19168
rect 10600 19116 10652 19168
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 112 18912 164 18964
rect 1492 18912 1544 18964
rect 2504 18912 2556 18964
rect 3424 18912 3476 18964
rect 4068 18912 4120 18964
rect 6184 18912 6236 18964
rect 7748 18955 7800 18964
rect 7748 18921 7757 18955
rect 7757 18921 7791 18955
rect 7791 18921 7800 18955
rect 7748 18912 7800 18921
rect 2596 18887 2648 18896
rect 2596 18853 2605 18887
rect 2605 18853 2639 18887
rect 2639 18853 2648 18887
rect 2596 18844 2648 18853
rect 5264 18844 5316 18896
rect 5908 18844 5960 18896
rect 1308 18776 1360 18828
rect 4620 18776 4672 18828
rect 7472 18776 7524 18828
rect 2504 18751 2556 18760
rect 2504 18717 2513 18751
rect 2513 18717 2547 18751
rect 2547 18717 2556 18751
rect 2504 18708 2556 18717
rect 4068 18708 4120 18760
rect 5356 18708 5408 18760
rect 3608 18640 3660 18692
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 4252 18572 4304 18624
rect 6828 18615 6880 18624
rect 6828 18581 6837 18615
rect 6837 18581 6871 18615
rect 6871 18581 6880 18615
rect 6828 18572 6880 18581
rect 7196 18615 7248 18624
rect 7196 18581 7205 18615
rect 7205 18581 7239 18615
rect 7239 18581 7248 18615
rect 7196 18572 7248 18581
rect 8116 18572 8168 18624
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 8576 18572 8628 18581
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 2320 18368 2372 18420
rect 2596 18368 2648 18420
rect 7472 18368 7524 18420
rect 7656 18300 7708 18352
rect 4068 18275 4120 18284
rect 4068 18241 4077 18275
rect 4077 18241 4111 18275
rect 4111 18241 4120 18275
rect 4068 18232 4120 18241
rect 4896 18232 4948 18284
rect 2320 18164 2372 18216
rect 1400 18096 1452 18148
rect 8300 18232 8352 18284
rect 8668 18275 8720 18284
rect 8668 18241 8677 18275
rect 8677 18241 8711 18275
rect 8711 18241 8720 18275
rect 8668 18232 8720 18241
rect 2504 18096 2556 18148
rect 1308 18028 1360 18080
rect 2320 18028 2372 18080
rect 4528 18096 4580 18148
rect 5448 18164 5500 18216
rect 10416 18207 10468 18216
rect 10416 18173 10460 18207
rect 10460 18173 10468 18207
rect 10876 18207 10928 18216
rect 10416 18164 10468 18173
rect 10876 18173 10885 18207
rect 10885 18173 10919 18207
rect 10919 18173 10928 18207
rect 10876 18164 10928 18173
rect 5264 18096 5316 18148
rect 5816 18096 5868 18148
rect 7196 18139 7248 18148
rect 7196 18105 7205 18139
rect 7205 18105 7239 18139
rect 7239 18105 7248 18139
rect 7196 18096 7248 18105
rect 7288 18139 7340 18148
rect 7288 18105 7297 18139
rect 7297 18105 7331 18139
rect 7331 18105 7340 18139
rect 7288 18096 7340 18105
rect 8392 18096 8444 18148
rect 5356 18071 5408 18080
rect 5356 18037 5365 18071
rect 5365 18037 5399 18071
rect 5399 18037 5408 18071
rect 5356 18028 5408 18037
rect 7656 18028 7708 18080
rect 9588 18071 9640 18080
rect 9588 18037 9597 18071
rect 9597 18037 9631 18071
rect 9631 18037 9640 18071
rect 9588 18028 9640 18037
rect 9772 18028 9824 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 2504 17867 2556 17876
rect 2504 17833 2513 17867
rect 2513 17833 2547 17867
rect 2547 17833 2556 17867
rect 2504 17824 2556 17833
rect 3516 17824 3568 17876
rect 8668 17824 8720 17876
rect 2320 17756 2372 17808
rect 4160 17756 4212 17808
rect 4252 17799 4304 17808
rect 4252 17765 4261 17799
rect 4261 17765 4295 17799
rect 4295 17765 4304 17799
rect 4252 17756 4304 17765
rect 4896 17756 4948 17808
rect 6092 17799 6144 17808
rect 6092 17765 6101 17799
rect 6101 17765 6135 17799
rect 6135 17765 6144 17799
rect 6092 17756 6144 17765
rect 7656 17756 7708 17808
rect 9772 17799 9824 17808
rect 9772 17765 9781 17799
rect 9781 17765 9815 17799
rect 9815 17765 9824 17799
rect 9772 17756 9824 17765
rect 9864 17799 9916 17808
rect 9864 17765 9873 17799
rect 9873 17765 9907 17799
rect 9907 17765 9916 17799
rect 9864 17756 9916 17765
rect 3240 17688 3292 17740
rect 4160 17663 4212 17672
rect 4160 17629 4169 17663
rect 4169 17629 4203 17663
rect 4203 17629 4212 17663
rect 6000 17663 6052 17672
rect 4160 17620 4212 17629
rect 6000 17629 6009 17663
rect 6009 17629 6043 17663
rect 6043 17629 6052 17663
rect 6000 17620 6052 17629
rect 6184 17620 6236 17672
rect 7564 17663 7616 17672
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 8576 17620 8628 17672
rect 10048 17663 10100 17672
rect 10048 17629 10057 17663
rect 10057 17629 10091 17663
rect 10091 17629 10100 17663
rect 10048 17620 10100 17629
rect 3516 17484 3568 17536
rect 5540 17484 5592 17536
rect 7288 17484 7340 17536
rect 8116 17484 8168 17536
rect 8208 17484 8260 17536
rect 9864 17484 9916 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 3240 17280 3292 17332
rect 4252 17280 4304 17332
rect 6092 17280 6144 17332
rect 3516 17187 3568 17196
rect 3516 17153 3525 17187
rect 3525 17153 3559 17187
rect 3559 17153 3568 17187
rect 3516 17144 3568 17153
rect 2872 17076 2924 17128
rect 3608 17119 3660 17128
rect 3608 17085 3617 17119
rect 3617 17085 3651 17119
rect 3651 17085 3660 17119
rect 3608 17076 3660 17085
rect 5356 17144 5408 17196
rect 6828 17144 6880 17196
rect 5172 17119 5224 17128
rect 5172 17085 5181 17119
rect 5181 17085 5215 17119
rect 5215 17085 5224 17119
rect 5172 17076 5224 17085
rect 5540 17076 5592 17128
rect 7840 17280 7892 17332
rect 8024 17280 8076 17332
rect 9588 17280 9640 17332
rect 9864 17280 9916 17332
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 8576 17255 8628 17264
rect 8576 17221 8585 17255
rect 8585 17221 8619 17255
rect 8619 17221 8628 17255
rect 8576 17212 8628 17221
rect 9496 17212 9548 17264
rect 8392 17144 8444 17196
rect 10692 17076 10744 17128
rect 11520 17076 11572 17128
rect 6000 17008 6052 17060
rect 8024 17051 8076 17060
rect 8024 17017 8033 17051
rect 8033 17017 8067 17051
rect 8067 17017 8076 17051
rect 8024 17008 8076 17017
rect 8116 17051 8168 17060
rect 8116 17017 8125 17051
rect 8125 17017 8159 17051
rect 8159 17017 8168 17051
rect 8116 17008 8168 17017
rect 9680 17051 9732 17060
rect 9680 17017 9689 17051
rect 9689 17017 9723 17051
rect 9723 17017 9732 17051
rect 10232 17051 10284 17060
rect 9680 17008 9732 17017
rect 10232 17017 10241 17051
rect 10241 17017 10275 17051
rect 10275 17017 10284 17051
rect 10232 17008 10284 17017
rect 4344 16940 4396 16992
rect 7288 16940 7340 16992
rect 7656 16940 7708 16992
rect 10968 16940 11020 16992
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 3608 16779 3660 16788
rect 3608 16745 3617 16779
rect 3617 16745 3651 16779
rect 3651 16745 3660 16779
rect 3608 16736 3660 16745
rect 4160 16736 4212 16788
rect 5816 16736 5868 16788
rect 6092 16779 6144 16788
rect 6092 16745 6101 16779
rect 6101 16745 6135 16779
rect 6135 16745 6144 16779
rect 6092 16736 6144 16745
rect 7196 16736 7248 16788
rect 7564 16779 7616 16788
rect 7564 16745 7573 16779
rect 7573 16745 7607 16779
rect 7607 16745 7616 16779
rect 7564 16736 7616 16745
rect 8024 16736 8076 16788
rect 3148 16668 3200 16720
rect 4896 16668 4948 16720
rect 7288 16668 7340 16720
rect 8116 16711 8168 16720
rect 8116 16677 8125 16711
rect 8125 16677 8159 16711
rect 8159 16677 8168 16711
rect 8116 16668 8168 16677
rect 8208 16711 8260 16720
rect 8208 16677 8217 16711
rect 8217 16677 8251 16711
rect 8251 16677 8260 16711
rect 9772 16736 9824 16788
rect 8208 16668 8260 16677
rect 10968 16668 11020 16720
rect 3516 16600 3568 16652
rect 4712 16600 4764 16652
rect 6552 16600 6604 16652
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 10600 16600 10652 16652
rect 10692 16643 10744 16652
rect 10692 16609 10701 16643
rect 10701 16609 10735 16643
rect 10735 16609 10744 16643
rect 10692 16600 10744 16609
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 5172 16532 5224 16541
rect 6000 16532 6052 16584
rect 7932 16532 7984 16584
rect 8392 16575 8444 16584
rect 8392 16541 8401 16575
rect 8401 16541 8435 16575
rect 8435 16541 8444 16575
rect 8392 16532 8444 16541
rect 4344 16507 4396 16516
rect 4344 16473 4353 16507
rect 4353 16473 4387 16507
rect 4387 16473 4396 16507
rect 4344 16464 4396 16473
rect 7748 16464 7800 16516
rect 4436 16396 4488 16448
rect 9404 16396 9456 16448
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 3516 16192 3568 16244
rect 4252 16192 4304 16244
rect 5724 16192 5776 16244
rect 8116 16192 8168 16244
rect 10692 16192 10744 16244
rect 2228 16056 2280 16108
rect 10784 16124 10836 16176
rect 15476 16124 15528 16176
rect 4896 16056 4948 16108
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 8208 16056 8260 16108
rect 9404 16056 9456 16108
rect 9496 16099 9548 16108
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 3516 16031 3568 16040
rect 3516 15997 3525 16031
rect 3525 15997 3559 16031
rect 3559 15997 3568 16031
rect 3516 15988 3568 15997
rect 4620 15920 4672 15972
rect 7012 16031 7064 16040
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 8668 15988 8720 16040
rect 10508 15988 10560 16040
rect 9312 15963 9364 15972
rect 9312 15929 9321 15963
rect 9321 15929 9355 15963
rect 9355 15929 9364 15963
rect 9312 15920 9364 15929
rect 3332 15895 3384 15904
rect 3332 15861 3341 15895
rect 3341 15861 3375 15895
rect 3375 15861 3384 15895
rect 3332 15852 3384 15861
rect 4712 15895 4764 15904
rect 4712 15861 4721 15895
rect 4721 15861 4755 15895
rect 4755 15861 4764 15895
rect 4712 15852 4764 15861
rect 5816 15895 5868 15904
rect 5816 15861 5825 15895
rect 5825 15861 5859 15895
rect 5859 15861 5868 15895
rect 5816 15852 5868 15861
rect 6184 15852 6236 15904
rect 8392 15852 8444 15904
rect 9588 15852 9640 15904
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 2504 15512 2556 15564
rect 2872 15648 2924 15700
rect 2688 15512 2740 15564
rect 3516 15648 3568 15700
rect 5172 15691 5224 15700
rect 5172 15657 5181 15691
rect 5181 15657 5215 15691
rect 5215 15657 5224 15691
rect 5172 15648 5224 15657
rect 6184 15648 6236 15700
rect 9404 15648 9456 15700
rect 9496 15648 9548 15700
rect 7840 15623 7892 15632
rect 4620 15555 4672 15564
rect 4620 15521 4629 15555
rect 4629 15521 4663 15555
rect 4663 15521 4672 15555
rect 4620 15512 4672 15521
rect 7840 15589 7849 15623
rect 7849 15589 7883 15623
rect 7883 15589 7892 15623
rect 7840 15580 7892 15589
rect 9312 15580 9364 15632
rect 8760 15512 8812 15564
rect 9404 15512 9456 15564
rect 10784 15512 10836 15564
rect 11336 15512 11388 15564
rect 11704 15555 11756 15564
rect 11704 15521 11713 15555
rect 11713 15521 11747 15555
rect 11747 15521 11756 15555
rect 11704 15512 11756 15521
rect 5448 15444 5500 15496
rect 5908 15487 5960 15496
rect 5908 15453 5917 15487
rect 5917 15453 5951 15487
rect 5951 15453 5960 15487
rect 5908 15444 5960 15453
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 7932 15444 7984 15496
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 6920 15376 6972 15428
rect 3516 15308 3568 15360
rect 4344 15308 4396 15360
rect 7012 15308 7064 15360
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 2688 15104 2740 15156
rect 4344 15104 4396 15156
rect 4528 15147 4580 15156
rect 4528 15113 4537 15147
rect 4537 15113 4571 15147
rect 4571 15113 4580 15147
rect 4528 15104 4580 15113
rect 5632 15104 5684 15156
rect 7012 15104 7064 15156
rect 7840 15147 7892 15156
rect 7840 15113 7849 15147
rect 7849 15113 7883 15147
rect 7883 15113 7892 15147
rect 7840 15104 7892 15113
rect 9312 15147 9364 15156
rect 9312 15113 9321 15147
rect 9321 15113 9355 15147
rect 9355 15113 9364 15147
rect 9312 15104 9364 15113
rect 11336 15147 11388 15156
rect 11336 15113 11345 15147
rect 11345 15113 11379 15147
rect 11379 15113 11388 15147
rect 11336 15104 11388 15113
rect 11428 15104 11480 15156
rect 11704 15147 11756 15156
rect 11704 15113 11713 15147
rect 11713 15113 11747 15147
rect 11747 15113 11756 15147
rect 11704 15104 11756 15113
rect 2504 15079 2556 15088
rect 2504 15045 2513 15079
rect 2513 15045 2547 15079
rect 2547 15045 2556 15079
rect 2504 15036 2556 15045
rect 3056 15036 3108 15088
rect 7656 15036 7708 15088
rect 10784 15036 10836 15088
rect 2688 14900 2740 14952
rect 3516 14900 3568 14952
rect 3332 14832 3384 14884
rect 6184 14968 6236 15020
rect 8208 14968 8260 15020
rect 8484 14968 8536 15020
rect 9496 14968 9548 15020
rect 10232 14968 10284 15020
rect 5448 14900 5500 14952
rect 7840 14900 7892 14952
rect 4252 14832 4304 14884
rect 6920 14875 6972 14884
rect 6920 14841 6929 14875
rect 6929 14841 6963 14875
rect 6963 14841 6972 14875
rect 6920 14832 6972 14841
rect 7012 14875 7064 14884
rect 7012 14841 7021 14875
rect 7021 14841 7055 14875
rect 7055 14841 7064 14875
rect 7012 14832 7064 14841
rect 4804 14807 4856 14816
rect 4804 14773 4813 14807
rect 4813 14773 4847 14807
rect 4847 14773 4856 14807
rect 4804 14764 4856 14773
rect 5448 14764 5500 14816
rect 6184 14764 6236 14816
rect 7564 14764 7616 14816
rect 9864 14832 9916 14884
rect 10048 14832 10100 14884
rect 10232 14875 10284 14884
rect 10232 14841 10241 14875
rect 10241 14841 10275 14875
rect 10275 14841 10284 14875
rect 10232 14832 10284 14841
rect 10692 14832 10744 14884
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 4252 14560 4304 14612
rect 2504 14492 2556 14544
rect 4068 14492 4120 14544
rect 4804 14560 4856 14612
rect 7748 14560 7800 14612
rect 8484 14603 8536 14612
rect 8484 14569 8493 14603
rect 8493 14569 8527 14603
rect 8527 14569 8536 14603
rect 8484 14560 8536 14569
rect 10692 14560 10744 14612
rect 7104 14535 7156 14544
rect 7104 14501 7113 14535
rect 7113 14501 7147 14535
rect 7147 14501 7156 14535
rect 7104 14492 7156 14501
rect 9864 14492 9916 14544
rect 10232 14492 10284 14544
rect 2872 14467 2924 14476
rect 2872 14433 2881 14467
rect 2881 14433 2915 14467
rect 2915 14433 2924 14467
rect 2872 14424 2924 14433
rect 3148 14424 3200 14476
rect 4528 14424 4580 14476
rect 5356 14467 5408 14476
rect 5356 14433 5365 14467
rect 5365 14433 5399 14467
rect 5399 14433 5408 14467
rect 5356 14424 5408 14433
rect 5632 14467 5684 14476
rect 5632 14433 5641 14467
rect 5641 14433 5675 14467
rect 5675 14433 5684 14467
rect 5632 14424 5684 14433
rect 8760 14424 8812 14476
rect 11520 14424 11572 14476
rect 5816 14399 5868 14408
rect 5816 14365 5825 14399
rect 5825 14365 5859 14399
rect 5859 14365 5868 14399
rect 5816 14356 5868 14365
rect 4252 14288 4304 14340
rect 6736 14288 6788 14340
rect 7932 14356 7984 14408
rect 10324 14356 10376 14408
rect 8852 14288 8904 14340
rect 9772 14288 9824 14340
rect 4988 14220 5040 14272
rect 5908 14220 5960 14272
rect 6828 14263 6880 14272
rect 6828 14229 6837 14263
rect 6837 14229 6871 14263
rect 6871 14229 6880 14263
rect 6828 14220 6880 14229
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 4436 14016 4488 14068
rect 5172 14016 5224 14068
rect 5356 14016 5408 14068
rect 9864 14016 9916 14068
rect 2872 13880 2924 13932
rect 7932 13948 7984 14000
rect 4068 13812 4120 13864
rect 2688 13787 2740 13796
rect 2688 13753 2697 13787
rect 2697 13753 2731 13787
rect 2731 13753 2740 13787
rect 4344 13812 4396 13864
rect 5172 13855 5224 13864
rect 5172 13821 5181 13855
rect 5181 13821 5215 13855
rect 5215 13821 5224 13855
rect 5172 13812 5224 13821
rect 5264 13812 5316 13864
rect 5632 13855 5684 13864
rect 5632 13821 5641 13855
rect 5641 13821 5675 13855
rect 5675 13821 5684 13855
rect 5632 13812 5684 13821
rect 8576 13880 8628 13932
rect 8852 13880 8904 13932
rect 2688 13744 2740 13753
rect 3148 13676 3200 13728
rect 3516 13676 3568 13728
rect 4712 13719 4764 13728
rect 4712 13685 4721 13719
rect 4721 13685 4755 13719
rect 4755 13685 4764 13719
rect 4712 13676 4764 13685
rect 6736 13676 6788 13728
rect 7564 13744 7616 13796
rect 9496 13744 9548 13796
rect 8024 13676 8076 13728
rect 8484 13719 8536 13728
rect 8484 13685 8493 13719
rect 8493 13685 8527 13719
rect 8527 13685 8536 13719
rect 8484 13676 8536 13685
rect 8668 13676 8720 13728
rect 10508 13855 10560 13864
rect 10508 13821 10517 13855
rect 10517 13821 10551 13855
rect 10551 13821 10560 13855
rect 10508 13812 10560 13821
rect 10140 13787 10192 13796
rect 10140 13753 10149 13787
rect 10149 13753 10183 13787
rect 10183 13753 10192 13787
rect 11428 13812 11480 13864
rect 10140 13744 10192 13753
rect 10324 13719 10376 13728
rect 10324 13685 10333 13719
rect 10333 13685 10367 13719
rect 10367 13685 10376 13719
rect 10324 13676 10376 13685
rect 11520 13719 11572 13728
rect 11520 13685 11529 13719
rect 11529 13685 11563 13719
rect 11563 13685 11572 13719
rect 11520 13676 11572 13685
rect 13452 13676 13504 13728
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 112 13472 164 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 8852 13515 8904 13524
rect 7104 13472 7156 13481
rect 4988 13447 5040 13456
rect 4988 13413 4997 13447
rect 4997 13413 5031 13447
rect 5031 13413 5040 13447
rect 4988 13404 5040 13413
rect 6644 13404 6696 13456
rect 8852 13481 8861 13515
rect 8861 13481 8895 13515
rect 8895 13481 8904 13515
rect 8852 13472 8904 13481
rect 10324 13472 10376 13524
rect 10508 13472 10560 13524
rect 10232 13404 10284 13456
rect 1492 13336 1544 13388
rect 3056 13336 3108 13388
rect 1952 13268 2004 13320
rect 2688 13268 2740 13320
rect 4712 13336 4764 13388
rect 5264 13336 5316 13388
rect 5816 13379 5868 13388
rect 5816 13345 5825 13379
rect 5825 13345 5859 13379
rect 5859 13345 5868 13379
rect 5816 13336 5868 13345
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 10048 13311 10100 13320
rect 10048 13277 10057 13311
rect 10057 13277 10091 13311
rect 10091 13277 10100 13311
rect 10048 13268 10100 13277
rect 8852 13200 8904 13252
rect 4068 13132 4120 13184
rect 5724 13175 5776 13184
rect 5724 13141 5733 13175
rect 5733 13141 5767 13175
rect 5767 13141 5776 13175
rect 5724 13132 5776 13141
rect 7196 13132 7248 13184
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 1492 12928 1544 12980
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 3424 12971 3476 12980
rect 3424 12937 3433 12971
rect 3433 12937 3467 12971
rect 3467 12937 3476 12971
rect 3424 12928 3476 12937
rect 3976 12928 4028 12980
rect 6828 12928 6880 12980
rect 8852 12928 8904 12980
rect 9496 12928 9548 12980
rect 2780 12860 2832 12912
rect 3332 12860 3384 12912
rect 3884 12903 3936 12912
rect 3884 12869 3893 12903
rect 3893 12869 3927 12903
rect 3927 12869 3936 12903
rect 3884 12860 3936 12869
rect 10232 12903 10284 12912
rect 4068 12792 4120 12844
rect 4344 12792 4396 12844
rect 4712 12724 4764 12776
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 5724 12767 5776 12776
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 5724 12724 5776 12733
rect 6184 12724 6236 12776
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 10232 12869 10241 12903
rect 10241 12869 10275 12903
rect 10275 12869 10284 12903
rect 10232 12860 10284 12869
rect 11520 12792 11572 12844
rect 8852 12724 8904 12776
rect 9404 12767 9456 12776
rect 9404 12733 9448 12767
rect 9448 12733 9456 12767
rect 9404 12724 9456 12733
rect 10876 12724 10928 12776
rect 1584 12656 1636 12708
rect 7564 12656 7616 12708
rect 8024 12699 8076 12708
rect 8024 12665 8033 12699
rect 8033 12665 8067 12699
rect 8067 12665 8076 12699
rect 8024 12656 8076 12665
rect 8668 12656 8720 12708
rect 2688 12631 2740 12640
rect 2688 12597 2697 12631
rect 2697 12597 2731 12631
rect 2731 12597 2740 12631
rect 2688 12588 2740 12597
rect 3516 12588 3568 12640
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 6736 12588 6788 12640
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 4804 12427 4856 12436
rect 4804 12393 4813 12427
rect 4813 12393 4847 12427
rect 4847 12393 4856 12427
rect 4804 12384 4856 12393
rect 7564 12427 7616 12436
rect 7564 12393 7573 12427
rect 7573 12393 7607 12427
rect 7607 12393 7616 12427
rect 7564 12384 7616 12393
rect 8024 12384 8076 12436
rect 9772 12427 9824 12436
rect 9772 12393 9781 12427
rect 9781 12393 9815 12427
rect 9815 12393 9824 12427
rect 9772 12384 9824 12393
rect 13636 12427 13688 12436
rect 13636 12393 13645 12427
rect 13645 12393 13679 12427
rect 13679 12393 13688 12427
rect 13636 12384 13688 12393
rect 3148 12359 3200 12368
rect 3148 12325 3157 12359
rect 3157 12325 3191 12359
rect 3191 12325 3200 12359
rect 3148 12316 3200 12325
rect 4068 12316 4120 12368
rect 7932 12359 7984 12368
rect 1676 12248 1728 12300
rect 2596 12291 2648 12300
rect 2596 12257 2605 12291
rect 2605 12257 2639 12291
rect 2639 12257 2648 12291
rect 2596 12248 2648 12257
rect 4344 12248 4396 12300
rect 3884 12180 3936 12232
rect 4068 12180 4120 12232
rect 4436 12180 4488 12232
rect 7932 12325 7941 12359
rect 7941 12325 7975 12359
rect 7975 12325 7984 12359
rect 7932 12316 7984 12325
rect 8208 12316 8260 12368
rect 5080 12248 5132 12300
rect 5724 12291 5776 12300
rect 5724 12257 5733 12291
rect 5733 12257 5767 12291
rect 5767 12257 5776 12291
rect 5724 12248 5776 12257
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 6184 12248 6236 12257
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 13452 12291 13504 12300
rect 13452 12257 13461 12291
rect 13461 12257 13495 12291
rect 13495 12257 13504 12291
rect 13452 12248 13504 12257
rect 4712 12180 4764 12232
rect 6644 12180 6696 12232
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 8852 12180 8904 12232
rect 1860 12112 1912 12164
rect 4804 12112 4856 12164
rect 3976 12044 4028 12096
rect 4620 12044 4672 12096
rect 10048 12112 10100 12164
rect 7196 12044 7248 12096
rect 7472 12044 7524 12096
rect 9404 12044 9456 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 1676 11883 1728 11892
rect 1676 11849 1685 11883
rect 1685 11849 1719 11883
rect 1719 11849 1728 11883
rect 1676 11840 1728 11849
rect 2228 11840 2280 11892
rect 3516 11840 3568 11892
rect 4436 11840 4488 11892
rect 4804 11883 4856 11892
rect 4804 11849 4813 11883
rect 4813 11849 4847 11883
rect 4847 11849 4856 11883
rect 4804 11840 4856 11849
rect 5724 11840 5776 11892
rect 6736 11840 6788 11892
rect 2504 11772 2556 11824
rect 3424 11772 3476 11824
rect 4620 11815 4672 11824
rect 4620 11781 4629 11815
rect 4629 11781 4663 11815
rect 4663 11781 4672 11815
rect 4620 11772 4672 11781
rect 7840 11772 7892 11824
rect 9680 11840 9732 11892
rect 10140 11840 10192 11892
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 8668 11704 8720 11756
rect 3976 11636 4028 11688
rect 4712 11568 4764 11620
rect 7196 11611 7248 11620
rect 7196 11577 7205 11611
rect 7205 11577 7239 11611
rect 7239 11577 7248 11611
rect 7196 11568 7248 11577
rect 8944 11704 8996 11756
rect 9772 11704 9824 11756
rect 6184 11543 6236 11552
rect 6184 11509 6193 11543
rect 6193 11509 6227 11543
rect 6227 11509 6236 11543
rect 6184 11500 6236 11509
rect 7564 11500 7616 11552
rect 7932 11500 7984 11552
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 1676 11296 1728 11348
rect 4620 11296 4672 11348
rect 7564 11339 7616 11348
rect 7564 11305 7573 11339
rect 7573 11305 7607 11339
rect 7607 11305 7616 11339
rect 7564 11296 7616 11305
rect 8668 11296 8720 11348
rect 8944 11339 8996 11348
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 4804 11228 4856 11280
rect 6736 11228 6788 11280
rect 7840 11228 7892 11280
rect 9772 11228 9824 11280
rect 10784 11228 10836 11280
rect 2504 11160 2556 11212
rect 2228 11092 2280 11144
rect 3976 11160 4028 11212
rect 5632 11203 5684 11212
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 3056 11024 3108 11076
rect 4068 11024 4120 11076
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 6644 11203 6696 11212
rect 6644 11169 6653 11203
rect 6653 11169 6687 11203
rect 6687 11169 6696 11203
rect 6644 11160 6696 11169
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 4436 11024 4488 11076
rect 5080 11067 5132 11076
rect 5080 11033 5089 11067
rect 5089 11033 5123 11067
rect 5123 11033 5132 11067
rect 5080 11024 5132 11033
rect 9680 11024 9732 11076
rect 10600 11092 10652 11144
rect 4344 10956 4396 11008
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 4436 10752 4488 10804
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 8392 10752 8444 10804
rect 9680 10795 9732 10804
rect 4068 10684 4120 10736
rect 4988 10684 5040 10736
rect 1676 10548 1728 10600
rect 2780 10548 2832 10600
rect 5080 10616 5132 10668
rect 9680 10761 9689 10795
rect 9689 10761 9723 10795
rect 9723 10761 9732 10795
rect 9680 10752 9732 10761
rect 9772 10752 9824 10804
rect 8852 10616 8904 10668
rect 3056 10548 3108 10600
rect 4620 10548 4672 10600
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 4344 10523 4396 10532
rect 4344 10489 4353 10523
rect 4353 10489 4387 10523
rect 4387 10489 4396 10523
rect 4344 10480 4396 10489
rect 4528 10480 4580 10532
rect 4804 10480 4856 10532
rect 1952 10455 2004 10464
rect 1952 10421 1961 10455
rect 1961 10421 1995 10455
rect 1995 10421 2004 10455
rect 1952 10412 2004 10421
rect 6736 10412 6788 10464
rect 8668 10412 8720 10464
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 2596 10208 2648 10260
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 3884 10251 3936 10260
rect 3884 10217 3893 10251
rect 3893 10217 3927 10251
rect 3927 10217 3936 10251
rect 3884 10208 3936 10217
rect 4160 10208 4212 10260
rect 5632 10251 5684 10260
rect 5632 10217 5641 10251
rect 5641 10217 5675 10251
rect 5675 10217 5684 10251
rect 5632 10208 5684 10217
rect 6644 10208 6696 10260
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 8668 10251 8720 10260
rect 8668 10217 8677 10251
rect 8677 10217 8711 10251
rect 8711 10217 8720 10251
rect 8668 10208 8720 10217
rect 3976 10140 4028 10192
rect 4712 10140 4764 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 1676 10072 1728 10124
rect 2964 10115 3016 10124
rect 2964 10081 2973 10115
rect 2973 10081 3007 10115
rect 3007 10081 3016 10115
rect 2964 10072 3016 10081
rect 3516 10072 3568 10124
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 6276 10115 6328 10124
rect 6276 10081 6285 10115
rect 6285 10081 6319 10115
rect 6319 10081 6328 10115
rect 6276 10072 6328 10081
rect 6920 10140 6972 10192
rect 7380 10115 7432 10124
rect 7380 10081 7389 10115
rect 7389 10081 7423 10115
rect 7423 10081 7432 10115
rect 7380 10072 7432 10081
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 4068 10004 4120 10056
rect 5080 10004 5132 10056
rect 10784 10072 10836 10124
rect 11060 10004 11112 10056
rect 4436 9979 4488 9988
rect 4436 9945 4460 9979
rect 4460 9945 4488 9979
rect 4436 9936 4488 9945
rect 4988 9936 5040 9988
rect 1400 9868 1452 9920
rect 2228 9868 2280 9920
rect 2780 9911 2832 9920
rect 2780 9877 2789 9911
rect 2789 9877 2823 9911
rect 2823 9877 2832 9911
rect 2780 9868 2832 9877
rect 5632 9868 5684 9920
rect 8392 9868 8444 9920
rect 9680 9868 9732 9920
rect 12348 9868 12400 9920
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 2964 9707 3016 9716
rect 2964 9673 2973 9707
rect 2973 9673 3007 9707
rect 3007 9673 3016 9707
rect 2964 9664 3016 9673
rect 4068 9664 4120 9716
rect 4988 9707 5040 9716
rect 4988 9673 4997 9707
rect 4997 9673 5031 9707
rect 5031 9673 5040 9707
rect 4988 9664 5040 9673
rect 6276 9707 6328 9716
rect 6276 9673 6285 9707
rect 6285 9673 6319 9707
rect 6319 9673 6328 9707
rect 6276 9664 6328 9673
rect 7380 9664 7432 9716
rect 8024 9664 8076 9716
rect 10140 9707 10192 9716
rect 1952 9596 2004 9648
rect 3332 9596 3384 9648
rect 4620 9639 4672 9648
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 4620 9605 4629 9639
rect 4629 9605 4663 9639
rect 4663 9605 4672 9639
rect 4620 9596 4672 9605
rect 9588 9596 9640 9648
rect 8024 9528 8076 9580
rect 8852 9528 8904 9580
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 5172 9503 5224 9512
rect 5172 9469 5181 9503
rect 5181 9469 5215 9503
rect 5215 9469 5224 9503
rect 5172 9460 5224 9469
rect 5632 9503 5684 9512
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 7472 9460 7524 9512
rect 10140 9673 10149 9707
rect 10149 9673 10183 9707
rect 10183 9673 10192 9707
rect 10140 9664 10192 9673
rect 10784 9664 10836 9716
rect 11060 9596 11112 9648
rect 4160 9392 4212 9444
rect 5908 9435 5960 9444
rect 5908 9401 5917 9435
rect 5917 9401 5951 9435
rect 5951 9401 5960 9435
rect 5908 9392 5960 9401
rect 8392 9392 8444 9444
rect 8668 9392 8720 9444
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 3148 9324 3200 9376
rect 6092 9324 6144 9376
rect 6828 9324 6880 9376
rect 8024 9324 8076 9376
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 2872 9052 2924 9104
rect 3516 9095 3568 9104
rect 3516 9061 3525 9095
rect 3525 9061 3559 9095
rect 3559 9061 3568 9095
rect 3516 9052 3568 9061
rect 3976 9052 4028 9104
rect 4804 9120 4856 9172
rect 7564 9120 7616 9172
rect 9680 9120 9732 9172
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 5632 9052 5684 9104
rect 8116 9095 8168 9104
rect 8116 9061 8125 9095
rect 8125 9061 8159 9095
rect 8159 9061 8168 9095
rect 8116 9052 8168 9061
rect 8668 9095 8720 9104
rect 8668 9061 8677 9095
rect 8677 9061 8711 9095
rect 8711 9061 8720 9095
rect 8668 9052 8720 9061
rect 9864 9095 9916 9104
rect 9864 9061 9873 9095
rect 9873 9061 9907 9095
rect 9907 9061 9916 9095
rect 9864 9052 9916 9061
rect 12348 9052 12400 9104
rect 15568 9052 15620 9104
rect 2688 8916 2740 8968
rect 3056 8848 3108 8900
rect 5172 8984 5224 9036
rect 5816 8984 5868 9036
rect 6092 8984 6144 9036
rect 11244 9027 11296 9036
rect 11244 8993 11253 9027
rect 11253 8993 11287 9027
rect 11287 8993 11296 9027
rect 11244 8984 11296 8993
rect 6184 8916 6236 8968
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 8024 8959 8076 8968
rect 8024 8925 8033 8959
rect 8033 8925 8067 8959
rect 8067 8925 8076 8959
rect 8024 8916 8076 8925
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 3976 8780 4028 8832
rect 5172 8780 5224 8832
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 8760 8780 8812 8832
rect 10784 8780 10836 8832
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 2964 8576 3016 8628
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 9864 8576 9916 8628
rect 11244 8619 11296 8628
rect 11244 8585 11253 8619
rect 11253 8585 11287 8619
rect 11287 8585 11296 8619
rect 11244 8576 11296 8585
rect 10048 8508 10100 8560
rect 10416 8508 10468 8560
rect 1584 8440 1636 8492
rect 4804 8440 4856 8492
rect 2780 8236 2832 8288
rect 3056 8236 3108 8288
rect 3516 8236 3568 8288
rect 4344 8372 4396 8424
rect 6920 8440 6972 8492
rect 8760 8440 8812 8492
rect 9956 8440 10008 8492
rect 10692 8440 10744 8492
rect 4160 8304 4212 8356
rect 4620 8279 4672 8288
rect 4620 8245 4629 8279
rect 4629 8245 4663 8279
rect 4663 8245 4672 8279
rect 4620 8236 4672 8245
rect 5540 8236 5592 8288
rect 6092 8236 6144 8288
rect 6736 8236 6788 8288
rect 7288 8236 7340 8288
rect 7748 8236 7800 8288
rect 8392 8279 8444 8288
rect 8392 8245 8401 8279
rect 8401 8245 8435 8279
rect 8435 8245 8444 8279
rect 8392 8236 8444 8245
rect 9772 8236 9824 8288
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 2688 8032 2740 8084
rect 3148 8075 3200 8084
rect 3148 8041 3157 8075
rect 3157 8041 3191 8075
rect 3191 8041 3200 8075
rect 3148 8032 3200 8041
rect 5356 8032 5408 8084
rect 5908 8032 5960 8084
rect 8024 8075 8076 8084
rect 2596 7964 2648 8016
rect 2044 7896 2096 7948
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 5632 7939 5684 7948
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 5816 7896 5868 7948
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 9680 8032 9732 8084
rect 10784 8075 10836 8084
rect 10784 8041 10793 8075
rect 10793 8041 10827 8075
rect 10827 8041 10836 8075
rect 10784 8032 10836 8041
rect 7288 7964 7340 8016
rect 8852 7964 8904 8016
rect 8576 7939 8628 7948
rect 8576 7905 8585 7939
rect 8585 7905 8619 7939
rect 8619 7905 8628 7939
rect 8576 7896 8628 7905
rect 3976 7828 4028 7880
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 3056 7692 3108 7744
rect 9772 7964 9824 8016
rect 9956 7964 10008 8016
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 9588 7828 9640 7880
rect 5540 7692 5592 7744
rect 8668 7692 8720 7744
rect 9680 7692 9732 7744
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 2596 7531 2648 7540
rect 2596 7497 2605 7531
rect 2605 7497 2639 7531
rect 2639 7497 2648 7531
rect 2596 7488 2648 7497
rect 4528 7488 4580 7540
rect 5632 7488 5684 7540
rect 6092 7488 6144 7540
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 3332 7420 3384 7472
rect 8576 7488 8628 7540
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 10048 7420 10100 7472
rect 3056 7352 3108 7404
rect 8944 7352 8996 7404
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 5356 7327 5408 7336
rect 5356 7293 5365 7327
rect 5365 7293 5399 7327
rect 5399 7293 5408 7327
rect 5356 7284 5408 7293
rect 5540 7284 5592 7336
rect 6184 7284 6236 7336
rect 2044 7216 2096 7268
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 2504 7148 2556 7200
rect 7288 7216 7340 7268
rect 8576 7216 8628 7268
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 1952 6944 2004 6996
rect 3700 6944 3752 6996
rect 3976 6944 4028 6996
rect 6092 6987 6144 6996
rect 6092 6953 6101 6987
rect 6101 6953 6135 6987
rect 6135 6953 6144 6987
rect 6092 6944 6144 6953
rect 9680 6944 9732 6996
rect 2504 6808 2556 6860
rect 2688 6851 2740 6860
rect 2688 6817 2697 6851
rect 2697 6817 2731 6851
rect 2731 6817 2740 6851
rect 2688 6808 2740 6817
rect 4068 6851 4120 6860
rect 2596 6672 2648 6724
rect 3056 6672 3108 6724
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 4528 6808 4580 6860
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 7288 6876 7340 6928
rect 8576 6919 8628 6928
rect 8576 6885 8585 6919
rect 8585 6885 8619 6919
rect 8619 6885 8628 6919
rect 8576 6876 8628 6885
rect 8944 6919 8996 6928
rect 8944 6885 8953 6919
rect 8953 6885 8987 6919
rect 8987 6885 8996 6919
rect 8944 6876 8996 6885
rect 9588 6876 9640 6928
rect 9772 6919 9824 6928
rect 9772 6885 9781 6919
rect 9781 6885 9815 6919
rect 9815 6885 9824 6919
rect 9772 6876 9824 6885
rect 10416 6944 10468 6996
rect 6644 6808 6696 6860
rect 8760 6808 8812 6860
rect 5540 6740 5592 6792
rect 6920 6740 6972 6792
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 4160 6715 4212 6724
rect 4160 6681 4169 6715
rect 4169 6681 4203 6715
rect 4203 6681 4212 6715
rect 5724 6715 5776 6724
rect 4160 6672 4212 6681
rect 5724 6681 5733 6715
rect 5733 6681 5767 6715
rect 5767 6681 5776 6715
rect 5724 6672 5776 6681
rect 4344 6604 4396 6656
rect 4988 6604 5040 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 2688 6400 2740 6452
rect 9680 6443 9732 6452
rect 9680 6409 9689 6443
rect 9689 6409 9723 6443
rect 9723 6409 9732 6443
rect 9680 6400 9732 6409
rect 9772 6400 9824 6452
rect 1676 6332 1728 6384
rect 8944 6332 8996 6384
rect 10048 6332 10100 6384
rect 4988 6307 5040 6316
rect 4988 6273 4997 6307
rect 4997 6273 5031 6307
rect 5031 6273 5040 6307
rect 4988 6264 5040 6273
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 2504 6171 2556 6180
rect 2504 6137 2513 6171
rect 2513 6137 2547 6171
rect 2547 6137 2556 6171
rect 2504 6128 2556 6137
rect 3148 6128 3200 6180
rect 2596 6060 2648 6112
rect 4160 6171 4212 6180
rect 4160 6137 4169 6171
rect 4169 6137 4203 6171
rect 4203 6137 4212 6171
rect 4160 6128 4212 6137
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 6920 6196 6972 6248
rect 8576 6171 8628 6180
rect 8576 6137 8585 6171
rect 8585 6137 8619 6171
rect 8619 6137 8628 6171
rect 8576 6128 8628 6137
rect 4528 6060 4580 6069
rect 5632 6060 5684 6112
rect 7104 6103 7156 6112
rect 7104 6069 7113 6103
rect 7113 6069 7147 6103
rect 7147 6069 7156 6103
rect 7104 6060 7156 6069
rect 7288 6060 7340 6112
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 4160 5856 4212 5908
rect 5724 5856 5776 5908
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 8576 5856 8628 5908
rect 7288 5788 7340 5840
rect 8484 5831 8536 5840
rect 8484 5797 8493 5831
rect 8493 5797 8527 5831
rect 8527 5797 8536 5831
rect 8484 5788 8536 5797
rect 8760 5831 8812 5840
rect 8760 5797 8769 5831
rect 8769 5797 8803 5831
rect 8803 5797 8812 5831
rect 8760 5788 8812 5797
rect 4068 5763 4120 5772
rect 4068 5729 4099 5763
rect 4099 5729 4120 5763
rect 4068 5720 4120 5729
rect 4436 5720 4488 5772
rect 5540 5720 5592 5772
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 7104 5763 7156 5772
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 8944 5720 8996 5772
rect 9588 5720 9640 5772
rect 11336 5720 11388 5772
rect 2780 5652 2832 5704
rect 5080 5652 5132 5704
rect 2596 5584 2648 5636
rect 4160 5627 4212 5636
rect 4160 5593 4169 5627
rect 4169 5593 4203 5627
rect 4203 5593 4212 5627
rect 4160 5584 4212 5593
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 5908 5559 5960 5568
rect 5908 5525 5917 5559
rect 5917 5525 5951 5559
rect 5951 5525 5960 5559
rect 5908 5516 5960 5525
rect 9496 5516 9548 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 2872 5312 2924 5364
rect 5908 5312 5960 5364
rect 9588 5355 9640 5364
rect 9588 5321 9597 5355
rect 9597 5321 9631 5355
rect 9631 5321 9640 5355
rect 9588 5312 9640 5321
rect 9956 5312 10008 5364
rect 4160 5244 4212 5296
rect 5172 5287 5224 5296
rect 5172 5253 5181 5287
rect 5181 5253 5215 5287
rect 5215 5253 5224 5287
rect 5172 5244 5224 5253
rect 10692 5244 10744 5296
rect 5264 5176 5316 5228
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 4068 5151 4120 5160
rect 3424 5108 3476 5117
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 4068 5108 4120 5117
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 6184 5108 6236 5160
rect 7472 5176 7524 5228
rect 9404 5176 9456 5228
rect 9588 5108 9640 5160
rect 10048 5108 10100 5160
rect 5540 5040 5592 5092
rect 7288 5040 7340 5092
rect 8024 5083 8076 5092
rect 8024 5049 8033 5083
rect 8033 5049 8067 5083
rect 8067 5049 8076 5083
rect 8024 5040 8076 5049
rect 3240 4972 3292 5024
rect 4068 4972 4120 5024
rect 4528 5015 4580 5024
rect 4528 4981 4537 5015
rect 4537 4981 4571 5015
rect 4571 4981 4580 5015
rect 4528 4972 4580 4981
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 7104 4972 7156 5024
rect 7840 4972 7892 5024
rect 9404 5040 9456 5092
rect 14648 5040 14700 5092
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 3516 4768 3568 4820
rect 3976 4768 4028 4820
rect 4252 4811 4304 4820
rect 2688 4700 2740 4752
rect 3424 4700 3476 4752
rect 4252 4777 4261 4811
rect 4261 4777 4295 4811
rect 4295 4777 4304 4811
rect 4252 4768 4304 4777
rect 4712 4811 4764 4820
rect 4712 4777 4721 4811
rect 4721 4777 4755 4811
rect 4755 4777 4764 4811
rect 4712 4768 4764 4777
rect 4988 4768 5040 4820
rect 7196 4768 7248 4820
rect 9312 4768 9364 4820
rect 9496 4768 9548 4820
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 5080 4632 5132 4684
rect 5908 4632 5960 4684
rect 8024 4700 8076 4752
rect 8208 4700 8260 4752
rect 9864 4675 9916 4684
rect 9864 4641 9873 4675
rect 9873 4641 9907 4675
rect 9907 4641 9916 4675
rect 9864 4632 9916 4641
rect 10140 4632 10192 4684
rect 11244 4675 11296 4684
rect 11244 4641 11288 4675
rect 11288 4641 11296 4675
rect 11244 4632 11296 4641
rect 2504 4564 2556 4616
rect 4528 4564 4580 4616
rect 6092 4564 6144 4616
rect 5724 4496 5776 4548
rect 8116 4564 8168 4616
rect 8852 4564 8904 4616
rect 9496 4564 9548 4616
rect 6184 4471 6236 4480
rect 6184 4437 6193 4471
rect 6193 4437 6227 4471
rect 6227 4437 6236 4471
rect 6184 4428 6236 4437
rect 10508 4428 10560 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 2780 4267 2832 4276
rect 2780 4233 2789 4267
rect 2789 4233 2823 4267
rect 2823 4233 2832 4267
rect 2780 4224 2832 4233
rect 2872 4224 2924 4276
rect 4712 4224 4764 4276
rect 6092 4224 6144 4276
rect 9864 4224 9916 4276
rect 11244 4267 11296 4276
rect 11244 4233 11253 4267
rect 11253 4233 11287 4267
rect 11287 4233 11296 4267
rect 11244 4224 11296 4233
rect 8852 4156 8904 4208
rect 4252 4088 4304 4140
rect 4712 4088 4764 4140
rect 3240 4020 3292 4072
rect 5080 4063 5132 4072
rect 3148 3995 3200 4004
rect 3148 3961 3157 3995
rect 3157 3961 3191 3995
rect 3191 3961 3200 3995
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 9312 4088 9364 4140
rect 5448 4020 5500 4072
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 9588 4020 9640 4072
rect 3148 3952 3200 3961
rect 6736 3952 6788 4004
rect 7196 3952 7248 4004
rect 9956 3952 10008 4004
rect 10140 3995 10192 4004
rect 10140 3961 10149 3995
rect 10149 3961 10183 3995
rect 10183 3961 10192 3995
rect 10140 3952 10192 3961
rect 2596 3884 2648 3936
rect 7012 3884 7064 3936
rect 8208 3884 8260 3936
rect 9864 3884 9916 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 2688 3723 2740 3732
rect 2688 3689 2697 3723
rect 2697 3689 2731 3723
rect 2731 3689 2740 3723
rect 2688 3680 2740 3689
rect 5724 3680 5776 3732
rect 6184 3680 6236 3732
rect 6828 3680 6880 3732
rect 8116 3723 8168 3732
rect 8116 3689 8125 3723
rect 8125 3689 8159 3723
rect 8159 3689 8168 3723
rect 8116 3680 8168 3689
rect 8208 3680 8260 3732
rect 3056 3587 3108 3596
rect 3056 3553 3074 3587
rect 3074 3553 3108 3587
rect 5172 3612 5224 3664
rect 3056 3544 3108 3553
rect 4252 3544 4304 3596
rect 4712 3587 4764 3596
rect 4712 3553 4721 3587
rect 4721 3553 4755 3587
rect 4755 3553 4764 3587
rect 4712 3544 4764 3553
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 7012 3612 7064 3664
rect 5724 3587 5776 3596
rect 5080 3544 5132 3553
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 9864 3655 9916 3664
rect 9864 3621 9873 3655
rect 9873 3621 9907 3655
rect 9907 3621 9916 3655
rect 9864 3612 9916 3621
rect 9956 3612 10008 3664
rect 11796 3587 11848 3596
rect 11796 3553 11805 3587
rect 11805 3553 11839 3587
rect 11839 3553 11848 3587
rect 11796 3544 11848 3553
rect 12900 3544 12952 3596
rect 5448 3476 5500 3528
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 8852 3476 8904 3528
rect 10324 3451 10376 3460
rect 10324 3417 10333 3451
rect 10333 3417 10367 3451
rect 10367 3417 10376 3451
rect 10324 3408 10376 3417
rect 9404 3383 9456 3392
rect 9404 3349 9413 3383
rect 9413 3349 9447 3383
rect 9447 3349 9456 3383
rect 9404 3340 9456 3349
rect 12808 3340 12860 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 2596 3179 2648 3188
rect 2596 3145 2605 3179
rect 2605 3145 2639 3179
rect 2639 3145 2648 3179
rect 2596 3136 2648 3145
rect 3056 3179 3108 3188
rect 3056 3145 3065 3179
rect 3065 3145 3099 3179
rect 3099 3145 3108 3179
rect 3056 3136 3108 3145
rect 4620 3179 4672 3188
rect 4620 3145 4629 3179
rect 4629 3145 4663 3179
rect 4663 3145 4672 3179
rect 4620 3136 4672 3145
rect 6828 3136 6880 3188
rect 8852 3179 8904 3188
rect 8852 3145 8861 3179
rect 8861 3145 8895 3179
rect 8895 3145 8904 3179
rect 8852 3136 8904 3145
rect 9864 3136 9916 3188
rect 11796 3179 11848 3188
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 12900 3179 12952 3188
rect 12900 3145 12909 3179
rect 12909 3145 12943 3179
rect 12943 3145 12952 3179
rect 12900 3136 12952 3145
rect 4712 3068 4764 3120
rect 5908 3068 5960 3120
rect 8208 3068 8260 3120
rect 3976 3043 4028 3052
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 9404 3043 9456 3052
rect 3424 2907 3476 2916
rect 3424 2873 3433 2907
rect 3433 2873 3467 2907
rect 3467 2873 3476 2907
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 10324 3000 10376 3052
rect 4620 2932 4672 2984
rect 5448 2975 5500 2984
rect 5448 2941 5457 2975
rect 5457 2941 5491 2975
rect 5491 2941 5500 2975
rect 5448 2932 5500 2941
rect 5724 2932 5776 2984
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 3424 2864 3476 2873
rect 7012 2864 7064 2916
rect 9496 2907 9548 2916
rect 9496 2873 9505 2907
rect 9505 2873 9539 2907
rect 9539 2873 9548 2907
rect 9496 2864 9548 2873
rect 5908 2839 5960 2848
rect 5908 2805 5917 2839
rect 5917 2805 5951 2839
rect 5951 2805 5960 2839
rect 5908 2796 5960 2805
rect 6644 2839 6696 2848
rect 6644 2805 6653 2839
rect 6653 2805 6687 2839
rect 6687 2805 6696 2839
rect 6644 2796 6696 2805
rect 8300 2796 8352 2848
rect 13728 2864 13780 2916
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 3424 2592 3476 2644
rect 4620 2592 4672 2644
rect 6828 2592 6880 2644
rect 7840 2635 7892 2644
rect 7840 2601 7849 2635
rect 7849 2601 7883 2635
rect 7883 2601 7892 2635
rect 7840 2592 7892 2601
rect 9404 2592 9456 2644
rect 1308 2524 1360 2576
rect 6644 2524 6696 2576
rect 8576 2524 8628 2576
rect 10140 2524 10192 2576
rect 848 2252 900 2304
rect 4620 2456 4672 2508
rect 5908 2456 5960 2508
rect 10968 2456 11020 2508
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 9312 2388 9364 2440
rect 12900 2388 12952 2440
rect 4528 2295 4580 2304
rect 4528 2261 4537 2295
rect 4537 2261 4571 2295
rect 4571 2261 4580 2295
rect 4528 2252 4580 2261
rect 6644 2295 6696 2304
rect 6644 2261 6653 2295
rect 6653 2261 6687 2295
rect 6687 2261 6696 2295
rect 6644 2252 6696 2261
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 11796 2252 11848 2304
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 1308 2048 1360 2100
rect 6644 2048 6696 2100
rect 8944 76 8996 128
rect 11796 76 11848 128
<< metal2 >>
rect 662 39636 718 40000
rect 1950 39658 2006 40000
rect 3330 39658 3386 40000
rect 4618 39658 4674 40000
rect 5998 39658 6054 40000
rect 662 39584 664 39636
rect 716 39584 718 39636
rect 662 39520 718 39584
rect 1596 39630 2006 39658
rect 110 38720 166 38729
rect 110 38655 166 38664
rect 124 35290 152 38655
rect 112 35284 164 35290
rect 112 35226 164 35232
rect 1596 33134 1624 39630
rect 1950 39520 2006 39630
rect 2504 39636 2556 39642
rect 2504 39578 2556 39584
rect 2976 39630 3386 39658
rect 1504 33106 1624 33134
rect 1398 31376 1454 31385
rect 1398 31311 1454 31320
rect 1412 29714 1440 31311
rect 1400 29708 1452 29714
rect 1400 29650 1452 29656
rect 1412 28966 1440 29650
rect 1400 28960 1452 28966
rect 1400 28902 1452 28908
rect 110 28792 166 28801
rect 110 28727 166 28736
rect 124 28626 152 28727
rect 112 28620 164 28626
rect 112 28562 164 28568
rect 110 23760 166 23769
rect 110 23695 166 23704
rect 124 23186 152 23695
rect 112 23180 164 23186
rect 112 23122 164 23128
rect 1412 20398 1440 28902
rect 1504 23089 1532 33106
rect 1582 30696 1638 30705
rect 1582 30631 1638 30640
rect 1596 29850 1624 30631
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 2412 28552 2464 28558
rect 2412 28494 2464 28500
rect 2424 28218 2452 28494
rect 2412 28212 2464 28218
rect 2412 28154 2464 28160
rect 1860 26784 1912 26790
rect 1860 26726 1912 26732
rect 2320 26784 2372 26790
rect 2320 26726 2372 26732
rect 1490 23080 1546 23089
rect 1490 23015 1546 23024
rect 1492 21480 1544 21486
rect 1492 21422 1544 21428
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1504 18970 1532 21422
rect 112 18964 164 18970
rect 112 18906 164 18912
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 124 18737 152 18906
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18737 1348 18770
rect 110 18728 166 18737
rect 110 18663 166 18672
rect 1306 18728 1362 18737
rect 1306 18663 1362 18672
rect 1320 18086 1348 18663
rect 1400 18148 1452 18154
rect 1400 18090 1452 18096
rect 1308 18080 1360 18086
rect 1308 18022 1360 18028
rect 110 13696 166 13705
rect 110 13631 166 13640
rect 124 13530 152 13631
rect 112 13524 164 13530
rect 112 13466 164 13472
rect 1320 9353 1348 18022
rect 1412 10130 1440 18090
rect 1504 13394 1532 18906
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 1504 12986 1532 13330
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1584 12708 1636 12714
rect 1584 12650 1636 12656
rect 1596 11354 1624 12650
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1688 11898 1716 12242
rect 1872 12170 1900 26726
rect 2332 26382 2360 26726
rect 2320 26376 2372 26382
rect 2320 26318 2372 26324
rect 2318 25936 2374 25945
rect 2318 25871 2374 25880
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18630 1992 19246
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1964 18329 1992 18566
rect 2332 18426 2360 25871
rect 2516 18970 2544 39578
rect 2778 33144 2834 33153
rect 2778 33079 2834 33088
rect 2688 32972 2740 32978
rect 2688 32914 2740 32920
rect 2700 32230 2728 32914
rect 2688 32224 2740 32230
rect 2688 32166 2740 32172
rect 2792 32026 2820 33079
rect 2872 32972 2924 32978
rect 2872 32914 2924 32920
rect 2884 32570 2912 32914
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 2780 32020 2832 32026
rect 2780 31962 2832 31968
rect 2596 31884 2648 31890
rect 2596 31826 2648 31832
rect 2608 31482 2636 31826
rect 2596 31476 2648 31482
rect 2596 31418 2648 31424
rect 2608 29170 2636 31418
rect 2976 31385 3004 39630
rect 3330 39520 3386 39630
rect 4540 39630 4674 39658
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3514 35728 3570 35737
rect 3514 35663 3570 35672
rect 3528 34746 3556 35663
rect 4160 35624 4212 35630
rect 4160 35566 4212 35572
rect 3976 35148 4028 35154
rect 3976 35090 4028 35096
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 3516 34740 3568 34746
rect 3516 34682 3568 34688
rect 3988 34678 4016 35090
rect 3976 34672 4028 34678
rect 3976 34614 4028 34620
rect 3976 34400 4028 34406
rect 3976 34342 4028 34348
rect 3516 33992 3568 33998
rect 3516 33934 3568 33940
rect 3528 33436 3556 33934
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3608 33448 3660 33454
rect 3528 33408 3608 33436
rect 3528 32774 3556 33408
rect 3608 33390 3660 33396
rect 3516 32768 3568 32774
rect 3516 32710 3568 32716
rect 3240 32224 3292 32230
rect 3240 32166 3292 32172
rect 2962 31376 3018 31385
rect 2962 31311 3018 31320
rect 3252 31142 3280 32166
rect 3528 31278 3556 32710
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3516 31272 3568 31278
rect 3516 31214 3568 31220
rect 3240 31136 3292 31142
rect 3240 31078 3292 31084
rect 2964 30932 3016 30938
rect 2964 30874 3016 30880
rect 2596 29164 2648 29170
rect 2596 29106 2648 29112
rect 2872 28620 2924 28626
rect 2872 28562 2924 28568
rect 2688 27940 2740 27946
rect 2688 27882 2740 27888
rect 2700 27538 2728 27882
rect 2884 27878 2912 28562
rect 2872 27872 2924 27878
rect 2872 27814 2924 27820
rect 2976 27538 3004 30874
rect 3148 30660 3200 30666
rect 3148 30602 3200 30608
rect 3056 29164 3108 29170
rect 3056 29106 3108 29112
rect 2688 27532 2740 27538
rect 2688 27474 2740 27480
rect 2964 27532 3016 27538
rect 2964 27474 3016 27480
rect 2700 27130 2728 27474
rect 2688 27124 2740 27130
rect 2688 27066 2740 27072
rect 2700 22234 2728 27066
rect 2976 26858 3004 27474
rect 2964 26852 3016 26858
rect 2964 26794 3016 26800
rect 3068 24886 3096 29106
rect 3160 28762 3188 30602
rect 3148 28756 3200 28762
rect 3148 28698 3200 28704
rect 3252 28234 3280 31078
rect 3528 30938 3556 31214
rect 3516 30932 3568 30938
rect 3516 30874 3568 30880
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3988 30054 4016 34342
rect 4068 30932 4120 30938
rect 4068 30874 4120 30880
rect 3332 30048 3384 30054
rect 3332 29990 3384 29996
rect 3976 30048 4028 30054
rect 3976 29990 4028 29996
rect 3160 28206 3280 28234
rect 3160 27334 3188 28206
rect 3344 28150 3372 29990
rect 3976 29776 4028 29782
rect 3976 29718 4028 29724
rect 3424 29504 3476 29510
rect 3424 29446 3476 29452
rect 3436 28218 3464 29446
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3884 29164 3936 29170
rect 3884 29106 3936 29112
rect 3516 28960 3568 28966
rect 3516 28902 3568 28908
rect 3528 28422 3556 28902
rect 3896 28490 3924 29106
rect 3988 28966 4016 29718
rect 4080 29170 4108 30874
rect 4172 29306 4200 35566
rect 4252 31816 4304 31822
rect 4252 31758 4304 31764
rect 4264 31346 4292 31758
rect 4252 31340 4304 31346
rect 4252 31282 4304 31288
rect 4436 31136 4488 31142
rect 4436 31078 4488 31084
rect 4448 30938 4476 31078
rect 4436 30932 4488 30938
rect 4436 30874 4488 30880
rect 4344 30864 4396 30870
rect 4344 30806 4396 30812
rect 4356 30394 4384 30806
rect 4344 30388 4396 30394
rect 4344 30330 4396 30336
rect 4160 29300 4212 29306
rect 4160 29242 4212 29248
rect 4068 29164 4120 29170
rect 4068 29106 4120 29112
rect 3976 28960 4028 28966
rect 3976 28902 4028 28908
rect 3884 28484 3936 28490
rect 3884 28426 3936 28432
rect 3516 28416 3568 28422
rect 3516 28358 3568 28364
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3424 28212 3476 28218
rect 3424 28154 3476 28160
rect 3332 28144 3384 28150
rect 3332 28086 3384 28092
rect 3344 28014 3372 28086
rect 3332 28008 3384 28014
rect 3252 27968 3332 27996
rect 3148 27328 3200 27334
rect 3148 27270 3200 27276
rect 3056 24880 3108 24886
rect 3056 24822 3108 24828
rect 3068 23662 3096 24822
rect 3252 24274 3280 27968
rect 3332 27950 3384 27956
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3896 27418 3924 27814
rect 3988 27538 4016 28902
rect 4068 28484 4120 28490
rect 4068 28426 4120 28432
rect 3976 27532 4028 27538
rect 3976 27474 4028 27480
rect 3424 27396 3476 27402
rect 3896 27390 4016 27418
rect 3424 27338 3476 27344
rect 3332 26444 3384 26450
rect 3332 26386 3384 26392
rect 3344 25702 3372 26386
rect 3436 26058 3464 27338
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3516 26852 3568 26858
rect 3516 26794 3568 26800
rect 3528 26518 3556 26794
rect 3516 26512 3568 26518
rect 3516 26454 3568 26460
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3436 26030 3556 26058
rect 3424 25832 3476 25838
rect 3424 25774 3476 25780
rect 3332 25696 3384 25702
rect 3332 25638 3384 25644
rect 3240 24268 3292 24274
rect 3240 24210 3292 24216
rect 3252 23798 3280 24210
rect 3240 23792 3292 23798
rect 3160 23740 3240 23746
rect 3160 23734 3292 23740
rect 3160 23718 3280 23734
rect 3056 23656 3108 23662
rect 3056 23598 3108 23604
rect 2872 23180 2924 23186
rect 2872 23122 2924 23128
rect 3056 23180 3108 23186
rect 3056 23122 3108 23128
rect 2884 22778 2912 23122
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 2884 22506 2912 22714
rect 2872 22500 2924 22506
rect 2872 22442 2924 22448
rect 2688 22228 2740 22234
rect 2688 22170 2740 22176
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2608 19378 2636 19790
rect 2700 19514 2728 19858
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 2596 19372 2648 19378
rect 2596 19314 2648 19320
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2596 18896 2648 18902
rect 2596 18838 2648 18844
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 1950 18320 2006 18329
rect 1950 18255 2006 18264
rect 1964 13326 1992 18255
rect 2332 18222 2360 18362
rect 2320 18216 2372 18222
rect 2372 18176 2452 18204
rect 2320 18158 2372 18164
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2332 17814 2360 18022
rect 2320 17808 2372 17814
rect 2320 17750 2372 17756
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1860 12164 1912 12170
rect 1860 12106 1912 12112
rect 2240 11898 2268 16050
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1688 10810 1716 11290
rect 2228 11144 2280 11150
rect 2226 11112 2228 11121
rect 2280 11112 2282 11121
rect 2226 11047 2282 11056
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1582 10704 1638 10713
rect 1582 10639 1638 10648
rect 1596 10266 1624 10639
rect 1688 10606 1716 10746
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 1412 4154 1440 9862
rect 1688 9382 1716 10066
rect 1964 9654 1992 10406
rect 2240 9926 2268 11047
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 7546 1624 8434
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1688 6390 1716 9318
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2056 7274 2084 7890
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1964 7002 1992 7142
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 2424 4154 2452 18176
rect 2516 18154 2544 18702
rect 2608 18426 2636 18838
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2516 17882 2544 18090
rect 2504 17876 2556 17882
rect 2504 17818 2556 17824
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2516 15094 2544 15506
rect 2700 15162 2728 15506
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2516 14550 2544 15030
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2504 14544 2556 14550
rect 2504 14486 2556 14492
rect 2700 13802 2728 14894
rect 2688 13796 2740 13802
rect 2688 13738 2740 13744
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2700 12646 2728 13262
rect 2792 12918 2820 20334
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 2976 19242 3004 19858
rect 2964 19236 3016 19242
rect 2884 19196 2964 19224
rect 2884 17134 2912 19196
rect 2964 19178 3016 19184
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2884 15706 2912 17070
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 3068 15094 3096 23122
rect 3160 16726 3188 23718
rect 3240 23656 3292 23662
rect 3240 23598 3292 23604
rect 3252 17746 3280 23598
rect 3344 23186 3372 25638
rect 3436 23186 3464 25774
rect 3528 24070 3556 26030
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3516 24064 3568 24070
rect 3516 24006 3568 24012
rect 3528 23848 3556 24006
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3528 23820 3648 23848
rect 3516 23656 3568 23662
rect 3516 23598 3568 23604
rect 3528 23254 3556 23598
rect 3620 23594 3648 23820
rect 3608 23588 3660 23594
rect 3608 23530 3660 23536
rect 3516 23248 3568 23254
rect 3516 23190 3568 23196
rect 3332 23180 3384 23186
rect 3332 23122 3384 23128
rect 3424 23180 3476 23186
rect 3424 23122 3476 23128
rect 3436 23066 3464 23122
rect 3344 23038 3464 23066
rect 3344 21865 3372 23038
rect 3424 22976 3476 22982
rect 3424 22918 3476 22924
rect 3330 21856 3386 21865
rect 3330 21791 3386 21800
rect 3436 20369 3464 22918
rect 3528 22778 3556 23190
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3884 22568 3936 22574
rect 3884 22510 3936 22516
rect 3896 21962 3924 22510
rect 3884 21956 3936 21962
rect 3884 21898 3936 21904
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3516 21344 3568 21350
rect 3516 21286 3568 21292
rect 3528 21146 3556 21286
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3528 20466 3556 21082
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3422 20360 3478 20369
rect 3422 20295 3478 20304
rect 3424 19984 3476 19990
rect 3424 19926 3476 19932
rect 3436 19446 3464 19926
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 3528 19242 3556 19654
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3516 19236 3568 19242
rect 3516 19178 3568 19184
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 3252 17338 3280 17682
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3056 15088 3108 15094
rect 3056 15030 3108 15036
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 2884 13938 2912 14418
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 3160 13734 3188 14418
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3068 12986 3096 13330
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2780 12912 2832 12918
rect 3068 12889 3096 12922
rect 2780 12854 2832 12860
rect 3054 12880 3110 12889
rect 3054 12815 3110 12824
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 2516 11218 2544 11766
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2516 10810 2544 11154
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2608 10266 2636 12242
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2700 8974 2728 12582
rect 3160 12374 3188 13670
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 9926 2820 10542
rect 2976 10130 3004 11086
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 3068 10606 3096 11018
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2700 8090 2728 8910
rect 2792 8537 2820 9862
rect 2976 9722 3004 10066
rect 3160 10033 3188 10202
rect 3146 10024 3202 10033
rect 3146 9959 3202 9968
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2778 8528 2834 8537
rect 2778 8463 2834 8472
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2608 7546 2636 7958
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2516 6866 2544 7142
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2516 6186 2544 6802
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2608 6118 2636 6666
rect 2700 6458 2728 6802
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2608 5642 2636 6054
rect 2792 5710 2820 8230
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2596 5636 2648 5642
rect 2596 5578 2648 5584
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 1320 4126 1440 4154
rect 2332 4126 2452 4154
rect 1320 2582 1348 4126
rect 1308 2576 1360 2582
rect 1308 2518 1360 2524
rect 848 2304 900 2310
rect 848 2246 900 2252
rect 478 82 534 480
rect 860 82 888 2246
rect 1308 2100 1360 2106
rect 1308 2042 1360 2048
rect 478 54 888 82
rect 1320 82 1348 2042
rect 2332 2009 2360 4126
rect 2318 2000 2374 2009
rect 2318 1935 2374 1944
rect 1398 82 1454 480
rect 1320 54 1454 82
rect 478 0 534 54
rect 1398 0 1454 54
rect 2318 82 2374 480
rect 2516 82 2544 4558
rect 2608 4185 2636 5578
rect 2884 5370 2912 9046
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2976 8634 3004 8978
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2962 8528 3018 8537
rect 2962 8463 3018 8472
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2594 4176 2650 4185
rect 2594 4111 2650 4120
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2608 3194 2636 3878
rect 2700 3738 2728 4694
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2792 4282 2820 4626
rect 2884 4282 2912 5306
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2976 4154 3004 8463
rect 3068 8294 3096 8842
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 3160 8090 3188 9318
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 7410 3096 7686
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3068 6730 3096 7346
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 2884 4126 3004 4154
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2318 54 2544 82
rect 2884 82 2912 4126
rect 3160 4010 3188 6122
rect 3252 5030 3280 17274
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3344 14890 3372 15846
rect 3332 14884 3384 14890
rect 3332 14826 3384 14832
rect 3436 12986 3464 18906
rect 3528 17882 3556 19178
rect 3620 18698 3648 19178
rect 3608 18692 3660 18698
rect 3608 18634 3660 18640
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3528 17202 3556 17478
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3528 16658 3556 17138
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3620 16794 3648 17070
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 3528 16250 3556 16594
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3528 15706 3556 15982
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 14958 3556 15302
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3528 13734 3556 14894
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3988 12986 4016 27390
rect 4080 27062 4108 28426
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 4080 22982 4108 24754
rect 4172 24750 4200 29242
rect 4540 28082 4568 39630
rect 4618 39520 4674 39630
rect 5828 39630 6054 39658
rect 4896 35488 4948 35494
rect 4896 35430 4948 35436
rect 4908 35086 4936 35430
rect 5264 35216 5316 35222
rect 5264 35158 5316 35164
rect 4896 35080 4948 35086
rect 4896 35022 4948 35028
rect 4804 34944 4856 34950
rect 4804 34886 4856 34892
rect 4816 34610 4844 34886
rect 5276 34746 5304 35158
rect 5724 35012 5776 35018
rect 5724 34954 5776 34960
rect 5264 34740 5316 34746
rect 5264 34682 5316 34688
rect 5632 34740 5684 34746
rect 5632 34682 5684 34688
rect 4804 34604 4856 34610
rect 4804 34546 4856 34552
rect 4620 34468 4672 34474
rect 4620 34410 4672 34416
rect 4632 33658 4660 34410
rect 4816 34202 4844 34546
rect 5644 34202 5672 34682
rect 4804 34196 4856 34202
rect 4804 34138 4856 34144
rect 5632 34196 5684 34202
rect 5632 34138 5684 34144
rect 5736 34082 5764 34954
rect 4712 34060 4764 34066
rect 4712 34002 4764 34008
rect 5644 34054 5764 34082
rect 4620 33652 4672 33658
rect 4620 33594 4672 33600
rect 4632 33386 4660 33594
rect 4724 33522 4752 34002
rect 4712 33516 4764 33522
rect 4712 33458 4764 33464
rect 4988 33448 5040 33454
rect 4988 33390 5040 33396
rect 5264 33448 5316 33454
rect 5264 33390 5316 33396
rect 4620 33380 4672 33386
rect 4620 33322 4672 33328
rect 4632 33134 4660 33322
rect 4632 33106 4752 33134
rect 5000 33114 5028 33390
rect 4724 32230 4752 33106
rect 4988 33108 5040 33114
rect 4988 33050 5040 33056
rect 5276 33046 5304 33390
rect 5264 33040 5316 33046
rect 5264 32982 5316 32988
rect 5540 33040 5592 33046
rect 5540 32982 5592 32988
rect 5448 32904 5500 32910
rect 5448 32846 5500 32852
rect 4804 32360 4856 32366
rect 4804 32302 4856 32308
rect 4712 32224 4764 32230
rect 4712 32166 4764 32172
rect 4724 31958 4752 32166
rect 4712 31952 4764 31958
rect 4712 31894 4764 31900
rect 4724 31482 4752 31894
rect 4712 31476 4764 31482
rect 4712 31418 4764 31424
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 4724 28218 4752 28494
rect 4712 28212 4764 28218
rect 4712 28154 4764 28160
rect 4528 28076 4580 28082
rect 4528 28018 4580 28024
rect 4252 28008 4304 28014
rect 4252 27950 4304 27956
rect 4264 27334 4292 27950
rect 4436 27464 4488 27470
rect 4436 27406 4488 27412
rect 4252 27328 4304 27334
rect 4252 27270 4304 27276
rect 4264 26994 4292 27270
rect 4252 26988 4304 26994
rect 4252 26930 4304 26936
rect 4448 26586 4476 27406
rect 4252 26580 4304 26586
rect 4252 26522 4304 26528
rect 4436 26580 4488 26586
rect 4436 26522 4488 26528
rect 4264 26489 4292 26522
rect 4250 26480 4306 26489
rect 4250 26415 4306 26424
rect 4344 26444 4396 26450
rect 4344 26386 4396 26392
rect 4356 25770 4384 26386
rect 4344 25764 4396 25770
rect 4344 25706 4396 25712
rect 4436 25356 4488 25362
rect 4436 25298 4488 25304
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4356 24954 4384 25230
rect 4448 24954 4476 25298
rect 4344 24948 4396 24954
rect 4344 24890 4396 24896
rect 4436 24948 4488 24954
rect 4436 24890 4488 24896
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 4436 24336 4488 24342
rect 4436 24278 4488 24284
rect 4344 24064 4396 24070
rect 4344 24006 4396 24012
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 4172 21486 4200 23802
rect 4356 22642 4384 24006
rect 4448 23633 4476 24278
rect 4434 23624 4490 23633
rect 4434 23559 4490 23568
rect 4448 23526 4476 23559
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 4540 23474 4568 28018
rect 4712 27940 4764 27946
rect 4712 27882 4764 27888
rect 4724 27606 4752 27882
rect 4712 27600 4764 27606
rect 4712 27542 4764 27548
rect 4620 26852 4672 26858
rect 4620 26794 4672 26800
rect 4632 26314 4660 26794
rect 4724 26790 4752 27542
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4620 26308 4672 26314
rect 4620 26250 4672 26256
rect 4632 26042 4660 26250
rect 4620 26036 4672 26042
rect 4620 25978 4672 25984
rect 4724 24342 4752 26726
rect 4816 26518 4844 32302
rect 5264 32224 5316 32230
rect 5264 32166 5316 32172
rect 5276 32026 5304 32166
rect 5264 32020 5316 32026
rect 5264 31962 5316 31968
rect 5172 31680 5224 31686
rect 5172 31622 5224 31628
rect 5184 31346 5212 31622
rect 5172 31340 5224 31346
rect 5172 31282 5224 31288
rect 5184 30870 5212 31282
rect 5276 31210 5304 31962
rect 5460 31634 5488 32846
rect 5552 32026 5580 32982
rect 5644 32910 5672 34054
rect 5724 33312 5776 33318
rect 5724 33254 5776 33260
rect 5736 33046 5764 33254
rect 5724 33040 5776 33046
rect 5724 32982 5776 32988
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5540 32020 5592 32026
rect 5540 31962 5592 31968
rect 5460 31606 5580 31634
rect 5264 31204 5316 31210
rect 5264 31146 5316 31152
rect 5172 30864 5224 30870
rect 5172 30806 5224 30812
rect 5552 30666 5580 31606
rect 5644 31414 5672 32846
rect 5632 31408 5684 31414
rect 5632 31350 5684 31356
rect 5632 31136 5684 31142
rect 5632 31078 5684 31084
rect 5540 30660 5592 30666
rect 5540 30602 5592 30608
rect 4988 30048 5040 30054
rect 4988 29990 5040 29996
rect 5000 28014 5028 29990
rect 5264 29028 5316 29034
rect 5264 28970 5316 28976
rect 5276 28762 5304 28970
rect 5264 28756 5316 28762
rect 5264 28698 5316 28704
rect 5080 28688 5132 28694
rect 5080 28630 5132 28636
rect 4988 28008 5040 28014
rect 4988 27950 5040 27956
rect 5000 27674 5028 27950
rect 5092 27878 5120 28630
rect 5552 28490 5580 30602
rect 5644 29782 5672 31078
rect 5632 29776 5684 29782
rect 5632 29718 5684 29724
rect 5540 28484 5592 28490
rect 5540 28426 5592 28432
rect 5828 28370 5856 39630
rect 5998 39520 6054 39630
rect 7286 39658 7342 40000
rect 8666 39658 8722 40000
rect 9954 39658 10010 40000
rect 7286 39630 7696 39658
rect 7286 39520 7342 39630
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6736 35488 6788 35494
rect 6736 35430 6788 35436
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6748 35086 6776 35430
rect 6000 35080 6052 35086
rect 6000 35022 6052 35028
rect 6736 35080 6788 35086
rect 6736 35022 6788 35028
rect 6012 34746 6040 35022
rect 6000 34740 6052 34746
rect 6000 34682 6052 34688
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6748 34202 6776 35022
rect 6828 34944 6880 34950
rect 6828 34886 6880 34892
rect 6840 34542 6868 34886
rect 6828 34536 6880 34542
rect 6828 34478 6880 34484
rect 7012 34468 7064 34474
rect 7012 34410 7064 34416
rect 7024 34202 7052 34410
rect 6736 34196 6788 34202
rect 6736 34138 6788 34144
rect 7012 34196 7064 34202
rect 7012 34138 7064 34144
rect 6644 33992 6696 33998
rect 6644 33934 6696 33940
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6656 33114 6684 33934
rect 7668 33930 7696 39630
rect 8666 39630 8892 39658
rect 8666 39520 8722 39630
rect 8484 35692 8536 35698
rect 8484 35634 8536 35640
rect 8024 35556 8076 35562
rect 8024 35498 8076 35504
rect 8116 35556 8168 35562
rect 8116 35498 8168 35504
rect 7748 35216 7800 35222
rect 7748 35158 7800 35164
rect 7760 34406 7788 35158
rect 7840 34672 7892 34678
rect 7840 34614 7892 34620
rect 7748 34400 7800 34406
rect 7748 34342 7800 34348
rect 7656 33924 7708 33930
rect 7656 33866 7708 33872
rect 7656 33516 7708 33522
rect 7656 33458 7708 33464
rect 6736 33380 6788 33386
rect 6736 33322 6788 33328
rect 6644 33108 6696 33114
rect 6644 33050 6696 33056
rect 6748 33046 6776 33322
rect 7012 33312 7064 33318
rect 7012 33254 7064 33260
rect 6736 33040 6788 33046
rect 6736 32982 6788 32988
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 5920 32230 5948 32846
rect 6644 32496 6696 32502
rect 6748 32484 6776 32982
rect 6696 32456 6776 32484
rect 6644 32438 6696 32444
rect 6656 32230 6684 32438
rect 5908 32224 5960 32230
rect 5908 32166 5960 32172
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 5920 30938 5948 32166
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 5908 30932 5960 30938
rect 5908 30874 5960 30880
rect 6092 30252 6144 30258
rect 6092 30194 6144 30200
rect 5908 30116 5960 30122
rect 5908 30058 5960 30064
rect 5920 29850 5948 30058
rect 5908 29844 5960 29850
rect 5908 29786 5960 29792
rect 5644 28342 5856 28370
rect 6000 28416 6052 28422
rect 6000 28358 6052 28364
rect 5540 28008 5592 28014
rect 5540 27950 5592 27956
rect 5080 27872 5132 27878
rect 5080 27814 5132 27820
rect 4988 27668 5040 27674
rect 4988 27610 5040 27616
rect 5092 26858 5120 27814
rect 5080 26852 5132 26858
rect 5080 26794 5132 26800
rect 4804 26512 4856 26518
rect 4804 26454 4856 26460
rect 4896 26444 4948 26450
rect 4896 26386 4948 26392
rect 4908 26042 4936 26386
rect 4896 26036 4948 26042
rect 4896 25978 4948 25984
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4712 24336 4764 24342
rect 4712 24278 4764 24284
rect 4816 23474 4844 25842
rect 4908 25498 4936 25978
rect 5264 25968 5316 25974
rect 5264 25910 5316 25916
rect 5080 25832 5132 25838
rect 5080 25774 5132 25780
rect 4896 25492 4948 25498
rect 4896 25434 4948 25440
rect 5092 25158 5120 25774
rect 5080 25152 5132 25158
rect 5080 25094 5132 25100
rect 4896 23656 4948 23662
rect 4948 23616 5028 23644
rect 4896 23598 4948 23604
rect 4448 23254 4476 23462
rect 4540 23446 4660 23474
rect 4816 23446 4936 23474
rect 4436 23248 4488 23254
rect 4436 23190 4488 23196
rect 4528 22976 4580 22982
rect 4528 22918 4580 22924
rect 4344 22636 4396 22642
rect 4344 22578 4396 22584
rect 4540 22234 4568 22918
rect 4528 22228 4580 22234
rect 4528 22170 4580 22176
rect 4632 21622 4660 23446
rect 4620 21616 4672 21622
rect 4620 21558 4672 21564
rect 4908 21486 4936 23446
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4896 21480 4948 21486
rect 4896 21422 4948 21428
rect 4252 21072 4304 21078
rect 4252 21014 4304 21020
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 4172 20534 4200 20878
rect 4160 20528 4212 20534
rect 4160 20470 4212 20476
rect 4066 20360 4122 20369
rect 4066 20295 4122 20304
rect 4080 19938 4108 20295
rect 4172 20058 4200 20470
rect 4264 20262 4292 21014
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4080 19910 4200 19938
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 4080 18970 4108 19790
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 4080 18290 4108 18702
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4172 17898 4200 19910
rect 4632 19446 4660 20810
rect 5000 20602 5028 23616
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4724 20058 4752 20198
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4908 19990 4936 20266
rect 4896 19984 4948 19990
rect 4896 19926 4948 19932
rect 4620 19440 4672 19446
rect 4620 19382 4672 19388
rect 4632 18834 4660 19382
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4080 17870 4200 17898
rect 4080 16402 4108 17870
rect 4264 17814 4292 18566
rect 4908 18290 4936 19926
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 5000 19378 5028 19858
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 4528 18148 4580 18154
rect 4528 18090 4580 18096
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4252 17808 4304 17814
rect 4252 17750 4304 17756
rect 4172 17678 4200 17750
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4172 16794 4200 17614
rect 4264 17338 4292 17750
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4080 16374 4200 16402
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 4080 13870 4108 14486
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3332 12912 3384 12918
rect 3332 12854 3384 12860
rect 3344 9654 3372 12854
rect 3436 11830 3464 12922
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3528 11898 3556 12582
rect 3896 12238 3924 12854
rect 4080 12850 4108 13126
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4080 12374 4108 12786
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3988 11694 4016 12038
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3988 11218 4016 11630
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3988 10452 4016 11154
rect 4080 11082 4108 12174
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4080 10742 4108 11018
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3896 10424 4016 10452
rect 3896 10266 3924 10424
rect 4172 10266 4200 16374
rect 4264 16250 4292 17274
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4356 16522 4384 16934
rect 4344 16516 4396 16522
rect 4344 16458 4396 16464
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4356 15162 4384 15302
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4252 14884 4304 14890
rect 4252 14826 4304 14832
rect 4264 14618 4292 14826
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3528 9110 3556 10066
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3988 9518 4016 10134
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9722 4108 9998
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4264 9586 4292 14282
rect 4448 14074 4476 16390
rect 4540 15162 4568 18090
rect 4908 17814 4936 18226
rect 4896 17808 4948 17814
rect 4896 17750 4948 17756
rect 4896 16720 4948 16726
rect 4896 16662 4948 16668
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4632 15570 4660 15914
rect 4724 15910 4752 16594
rect 4908 16114 4936 16662
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4528 14476 4580 14482
rect 4632 14464 4660 15506
rect 4580 14436 4660 14464
rect 4528 14418 4580 14424
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4356 12850 4384 13806
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4356 11014 4384 12242
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4448 11898 4476 12174
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4448 11082 4476 11834
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4356 10538 4384 10950
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 9110 4016 9454
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3988 8838 4016 9046
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 4172 8362 4200 9386
rect 4356 8430 4384 10474
rect 4448 9994 4476 10746
rect 4540 10538 4568 14418
rect 4724 13814 4752 15846
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4816 14618 4844 14758
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4724 13786 4844 13814
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 13394 4752 13670
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4724 12646 4752 12718
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 12238 4752 12582
rect 4816 12442 4844 13786
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4632 11830 4660 12038
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4632 11354 4660 11766
rect 4724 11626 4752 12174
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4816 11898 4844 12106
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4632 10606 4660 11290
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4724 10198 4752 11562
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4816 10810 4844 11222
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4710 10024 4766 10033
rect 4436 9988 4488 9994
rect 4710 9959 4766 9968
rect 4436 9930 4488 9936
rect 4448 9674 4476 9930
rect 4448 9654 4660 9674
rect 4448 9648 4672 9654
rect 4448 9646 4620 9648
rect 4620 9590 4672 9596
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3240 4072 3292 4078
rect 3344 4060 3372 7414
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3436 4758 3464 5102
rect 3528 4826 3556 8230
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3712 7002 3740 7278
rect 3988 7002 4016 7822
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 4080 6866 4108 7890
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 4080 5778 4108 6802
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4172 6186 4200 6666
rect 4356 6662 4384 7890
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4540 7546 4568 7822
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4172 5914 4200 6122
rect 4540 6118 4568 6802
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4068 5772 4120 5778
rect 4436 5772 4488 5778
rect 4120 5732 4292 5760
rect 4068 5714 4120 5720
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 4172 5302 4200 5578
rect 4160 5296 4212 5302
rect 4066 5264 4122 5273
rect 4160 5238 4212 5244
rect 4066 5199 4122 5208
rect 4080 5166 4108 5199
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3292 4032 3372 4060
rect 3240 4014 3292 4020
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3068 3194 3096 3538
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3160 1873 3188 3946
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3988 3058 4016 4762
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3436 2650 3464 2858
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3146 1864 3202 1873
rect 3146 1799 3202 1808
rect 3238 82 3294 480
rect 2884 54 3294 82
rect 4080 82 4108 4966
rect 4264 4826 4292 5732
rect 4540 5760 4568 6054
rect 4488 5732 4568 5760
rect 4436 5714 4488 5720
rect 4540 5030 4568 5732
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4264 4146 4292 4762
rect 4540 4622 4568 4966
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4264 3602 4292 4082
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4632 3194 4660 8230
rect 4724 4826 4752 9959
rect 4816 9178 4844 10474
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4816 8498 4844 9114
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4724 4146 4752 4218
rect 4908 4154 4936 16050
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 5000 13462 5028 14214
rect 4988 13456 5040 13462
rect 4988 13398 5040 13404
rect 5092 12306 5120 25094
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5184 23254 5212 23462
rect 5172 23248 5224 23254
rect 5172 23190 5224 23196
rect 5184 22642 5212 23190
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5276 22574 5304 25910
rect 5448 25152 5500 25158
rect 5448 25094 5500 25100
rect 5460 24818 5488 25094
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5460 24682 5488 24754
rect 5448 24676 5500 24682
rect 5448 24618 5500 24624
rect 5460 23798 5488 24618
rect 5552 23866 5580 27950
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5448 23792 5500 23798
rect 5448 23734 5500 23740
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 5552 23322 5580 23462
rect 5540 23316 5592 23322
rect 5540 23258 5592 23264
rect 5644 23254 5672 28342
rect 6012 27470 6040 28358
rect 6000 27464 6052 27470
rect 6000 27406 6052 27412
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 5736 26772 5764 27066
rect 6012 27062 6040 27406
rect 6000 27056 6052 27062
rect 6000 26998 6052 27004
rect 5816 26784 5868 26790
rect 5736 26744 5816 26772
rect 5736 26450 5764 26744
rect 5816 26726 5868 26732
rect 6104 26450 6132 30194
rect 6184 30184 6236 30190
rect 6184 30126 6236 30132
rect 6196 28150 6224 30126
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6656 28966 6684 32166
rect 7024 31958 7052 33254
rect 7668 33134 7696 33458
rect 7760 33318 7788 34342
rect 7748 33312 7800 33318
rect 7748 33254 7800 33260
rect 7746 33144 7802 33153
rect 7668 33106 7746 33134
rect 7746 33079 7802 33088
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 7012 31952 7064 31958
rect 7012 31894 7064 31900
rect 7024 31482 7052 31894
rect 7012 31476 7064 31482
rect 7012 31418 7064 31424
rect 6736 31408 6788 31414
rect 6736 31350 6788 31356
rect 6748 30802 6776 31350
rect 7116 30802 7144 32846
rect 7656 32768 7708 32774
rect 7656 32710 7708 32716
rect 7668 32298 7696 32710
rect 7196 32292 7248 32298
rect 7196 32234 7248 32240
rect 7656 32292 7708 32298
rect 7656 32234 7708 32240
rect 7208 31754 7236 32234
rect 7196 31748 7248 31754
rect 7196 31690 7248 31696
rect 6736 30796 6788 30802
rect 6736 30738 6788 30744
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 6748 29782 6776 30738
rect 7116 30394 7144 30738
rect 7104 30388 7156 30394
rect 7104 30330 7156 30336
rect 7380 30252 7432 30258
rect 7380 30194 7432 30200
rect 7196 30048 7248 30054
rect 7196 29990 7248 29996
rect 6828 29844 6880 29850
rect 6828 29786 6880 29792
rect 6736 29776 6788 29782
rect 6736 29718 6788 29724
rect 6748 28994 6776 29718
rect 6840 29170 6868 29786
rect 7104 29776 7156 29782
rect 7024 29736 7104 29764
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 7024 29034 7052 29736
rect 7104 29718 7156 29724
rect 7208 29170 7236 29990
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 7012 29028 7064 29034
rect 6748 28966 6868 28994
rect 7012 28970 7064 28976
rect 6644 28960 6696 28966
rect 6644 28902 6696 28908
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6656 28762 6684 28902
rect 6644 28756 6696 28762
rect 6564 28716 6644 28744
rect 6184 28144 6236 28150
rect 6184 28086 6236 28092
rect 5724 26444 5776 26450
rect 5724 26386 5776 26392
rect 6092 26444 6144 26450
rect 6092 26386 6144 26392
rect 5736 25702 5764 26386
rect 6104 26042 6132 26386
rect 6092 26036 6144 26042
rect 6092 25978 6144 25984
rect 6196 25945 6224 28086
rect 6564 27946 6592 28716
rect 6644 28698 6696 28704
rect 6656 28633 6684 28698
rect 6644 28552 6696 28558
rect 6644 28494 6696 28500
rect 6552 27940 6604 27946
rect 6552 27882 6604 27888
rect 6656 27878 6684 28494
rect 6644 27872 6696 27878
rect 6644 27814 6696 27820
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6276 27600 6328 27606
rect 6276 27542 6328 27548
rect 6288 27130 6316 27542
rect 6276 27124 6328 27130
rect 6276 27066 6328 27072
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6656 26518 6684 27814
rect 6736 27396 6788 27402
rect 6736 27338 6788 27344
rect 6748 27130 6776 27338
rect 6736 27124 6788 27130
rect 6736 27066 6788 27072
rect 6644 26512 6696 26518
rect 6644 26454 6696 26460
rect 6840 25974 6868 28966
rect 7024 28762 7052 28970
rect 7012 28756 7064 28762
rect 7012 28698 7064 28704
rect 6920 28484 6972 28490
rect 6920 28426 6972 28432
rect 6932 27606 6960 28426
rect 6920 27600 6972 27606
rect 6920 27542 6972 27548
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 7300 26489 7328 26522
rect 7286 26480 7342 26489
rect 7286 26415 7342 26424
rect 6828 25968 6880 25974
rect 6182 25936 6238 25945
rect 6828 25910 6880 25916
rect 6182 25871 6238 25880
rect 6840 25838 6868 25910
rect 6828 25832 6880 25838
rect 6828 25774 6880 25780
rect 7196 25832 7248 25838
rect 7196 25774 7248 25780
rect 5724 25696 5776 25702
rect 5724 25638 5776 25644
rect 7104 25696 7156 25702
rect 7104 25638 7156 25644
rect 5632 23248 5684 23254
rect 5632 23190 5684 23196
rect 5264 22568 5316 22574
rect 5264 22510 5316 22516
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5184 22098 5212 22374
rect 5276 22234 5304 22510
rect 5264 22228 5316 22234
rect 5264 22170 5316 22176
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 5184 21350 5212 22034
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 5184 20806 5212 21286
rect 5172 20800 5224 20806
rect 5172 20742 5224 20748
rect 5184 17134 5212 20742
rect 5276 20058 5304 22170
rect 5736 21962 5764 25638
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 7116 25498 7144 25638
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 6184 25424 6236 25430
rect 6184 25366 6236 25372
rect 6092 25288 6144 25294
rect 6092 25230 6144 25236
rect 5908 24676 5960 24682
rect 5908 24618 5960 24624
rect 5816 24336 5868 24342
rect 5816 24278 5868 24284
rect 5828 24070 5856 24278
rect 5920 24138 5948 24618
rect 6104 24274 6132 25230
rect 6196 24614 6224 25366
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 6932 24682 6960 25094
rect 6920 24676 6972 24682
rect 6920 24618 6972 24624
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 6092 24268 6144 24274
rect 6092 24210 6144 24216
rect 5908 24132 5960 24138
rect 5908 24074 5960 24080
rect 5816 24064 5868 24070
rect 5816 24006 5868 24012
rect 5828 23866 5856 24006
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 5816 23656 5868 23662
rect 5816 23598 5868 23604
rect 5828 23322 5856 23598
rect 6196 23526 6224 24550
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6932 24410 6960 24618
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6932 23730 6960 24006
rect 6920 23724 6972 23730
rect 6920 23666 6972 23672
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 5816 23316 5868 23322
rect 5816 23258 5868 23264
rect 6552 23248 6604 23254
rect 6552 23190 6604 23196
rect 5908 22976 5960 22982
rect 5908 22918 5960 22924
rect 5920 22642 5948 22918
rect 5908 22636 5960 22642
rect 5908 22578 5960 22584
rect 6564 22506 6592 23190
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6552 22500 6604 22506
rect 6552 22442 6604 22448
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6276 22092 6328 22098
rect 6276 22034 6328 22040
rect 5724 21956 5776 21962
rect 5724 21898 5776 21904
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 5920 21554 5948 21830
rect 6288 21690 6316 22034
rect 6644 21956 6696 21962
rect 6644 21898 6696 21904
rect 6276 21684 6328 21690
rect 6276 21626 6328 21632
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 5540 21480 5592 21486
rect 5592 21440 5672 21468
rect 5540 21422 5592 21428
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5552 20466 5580 20742
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5276 19514 5304 19994
rect 5368 19514 5396 20266
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5276 18902 5304 19178
rect 5264 18896 5316 18902
rect 5264 18838 5316 18844
rect 5276 18154 5304 18838
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 5368 18086 5396 18702
rect 5446 18320 5502 18329
rect 5446 18255 5502 18264
rect 5460 18222 5488 18255
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5368 17202 5396 18022
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5552 17134 5580 17478
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5184 15706 5212 16526
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 14958 5488 15438
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5460 14822 5488 14894
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5368 14074 5396 14418
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5184 13977 5212 14010
rect 5170 13968 5226 13977
rect 5170 13903 5226 13912
rect 5184 13870 5212 13903
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5276 13394 5304 13806
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 5000 9994 5028 10678
rect 5092 10674 5120 11018
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 10062 5120 10610
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 5000 9722 5028 9930
rect 4988 9716 5040 9722
rect 4988 9658 5040 9664
rect 5184 9518 5212 12718
rect 5460 10169 5488 14758
rect 5446 10160 5502 10169
rect 5446 10095 5502 10104
rect 5552 9674 5580 17070
rect 5644 15162 5672 21440
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6656 21010 6684 21898
rect 6840 21894 6868 22510
rect 7116 22098 7144 25434
rect 7208 25430 7236 25774
rect 7196 25424 7248 25430
rect 7196 25366 7248 25372
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7288 25288 7340 25294
rect 7288 25230 7340 25236
rect 7208 24818 7236 25230
rect 7300 24818 7328 25230
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7288 24812 7340 24818
rect 7288 24754 7340 24760
rect 7300 24138 7328 24754
rect 7288 24132 7340 24138
rect 7288 24074 7340 24080
rect 7300 23730 7328 24074
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 7116 21690 7144 22034
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 5736 16250 5764 20538
rect 6092 20324 6144 20330
rect 6092 20266 6144 20272
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5920 18902 5948 19926
rect 6104 19854 6132 20266
rect 6656 20262 6684 20946
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6184 19984 6236 19990
rect 6184 19926 6236 19932
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6104 19378 6132 19790
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5828 16794 5856 18090
rect 6104 17898 6132 19314
rect 6196 19174 6224 19926
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6196 18970 6224 19110
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6104 17870 6224 17898
rect 6092 17808 6144 17814
rect 6092 17750 6144 17756
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 6012 17066 6040 17614
rect 6104 17338 6132 17750
rect 6196 17678 6224 17870
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 6104 16794 6132 17274
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5828 15910 5856 16730
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 5644 13870 5672 14418
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5828 13394 5856 14350
rect 5920 14278 5948 15438
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5736 12782 5764 13126
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5736 11898 5764 12242
rect 5724 11892 5776 11898
rect 5776 11852 5856 11880
rect 5724 11834 5776 11840
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5644 11121 5672 11154
rect 5630 11112 5686 11121
rect 5630 11047 5686 11056
rect 5644 10266 5672 11047
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5368 9646 5580 9674
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5184 9042 5212 9454
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5000 6322 5028 6598
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4816 4126 4936 4154
rect 5000 4154 5028 4762
rect 5092 4690 5120 5646
rect 5184 5302 5212 8774
rect 5368 8090 5396 9646
rect 5644 9518 5672 9862
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5644 9110 5672 9454
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5828 9042 5856 11852
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5368 7342 5396 8026
rect 5552 7750 5580 8230
rect 5828 7954 5856 8978
rect 5920 8090 5948 9386
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5552 7342 5580 7686
rect 5644 7546 5672 7890
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5552 6798 5580 7278
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5644 6118 5672 6802
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5552 5574 5580 5714
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5276 4154 5304 5170
rect 5552 5098 5580 5510
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5000 4126 5120 4154
rect 4724 3602 4752 4082
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4632 2990 4660 3130
rect 4724 3126 4752 3538
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4632 2650 4660 2926
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4632 2514 4660 2586
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4540 1873 4568 2246
rect 4526 1864 4582 1873
rect 4526 1799 4582 1808
rect 4158 82 4214 480
rect 4080 54 4214 82
rect 4816 82 4844 4126
rect 5092 4078 5120 4126
rect 5184 4126 5304 4154
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5092 3602 5120 4014
rect 5184 3670 5212 4126
rect 5644 4078 5672 6054
rect 5736 5914 5764 6666
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5828 5166 5856 5714
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5920 5370 5948 5510
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5460 3534 5488 4014
rect 5736 3738 5764 4490
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5460 2990 5488 3470
rect 5736 2990 5764 3538
rect 5920 3126 5948 4626
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5460 2446 5488 2926
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5920 2514 5948 2790
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5170 82 5226 480
rect 4816 54 5226 82
rect 6012 82 6040 16526
rect 6564 16114 6592 16594
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 15706 6224 15846
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6196 15026 6224 15642
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6196 14822 6224 14962
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6748 14346 6776 21422
rect 6840 19922 6868 21626
rect 7116 21010 7144 21626
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7208 21078 7236 21422
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 7116 20398 7144 20946
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6840 18630 6868 19246
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6840 17202 6868 18566
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 7024 16046 7052 20198
rect 7116 20058 7144 20334
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7392 18737 7420 30194
rect 7656 30048 7708 30054
rect 7656 29990 7708 29996
rect 7472 29640 7524 29646
rect 7472 29582 7524 29588
rect 7484 28762 7512 29582
rect 7668 29034 7696 29990
rect 7760 29050 7788 33079
rect 7852 32434 7880 34614
rect 8036 34610 8064 35498
rect 8128 35290 8156 35498
rect 8116 35284 8168 35290
rect 8116 35226 8168 35232
rect 8128 34746 8156 35226
rect 8392 35148 8444 35154
rect 8392 35090 8444 35096
rect 8116 34740 8168 34746
rect 8116 34682 8168 34688
rect 8024 34604 8076 34610
rect 8024 34546 8076 34552
rect 8404 34406 8432 35090
rect 8496 34678 8524 35634
rect 8864 35290 8892 39630
rect 9600 39630 10010 39658
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 8852 35284 8904 35290
rect 8852 35226 8904 35232
rect 8576 35080 8628 35086
rect 8628 35040 8708 35068
rect 8576 35022 8628 35028
rect 8484 34672 8536 34678
rect 8484 34614 8536 34620
rect 8680 34474 8708 35040
rect 8760 34944 8812 34950
rect 8760 34886 8812 34892
rect 8772 34474 8800 34886
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8668 34468 8720 34474
rect 8668 34410 8720 34416
rect 8760 34468 8812 34474
rect 8760 34410 8812 34416
rect 8392 34400 8444 34406
rect 8392 34342 8444 34348
rect 8024 32768 8076 32774
rect 8024 32710 8076 32716
rect 7840 32428 7892 32434
rect 7840 32370 7892 32376
rect 8036 31822 8064 32710
rect 8404 31890 8432 34342
rect 8680 34134 8708 34410
rect 8772 34202 8800 34410
rect 8852 34400 8904 34406
rect 8852 34342 8904 34348
rect 8864 34202 8892 34342
rect 8760 34196 8812 34202
rect 8760 34138 8812 34144
rect 8852 34196 8904 34202
rect 8852 34138 8904 34144
rect 8668 34128 8720 34134
rect 8668 34070 8720 34076
rect 8484 34060 8536 34066
rect 8484 34002 8536 34008
rect 8852 34060 8904 34066
rect 8852 34002 8904 34008
rect 8496 33658 8524 34002
rect 8760 33856 8812 33862
rect 8760 33798 8812 33804
rect 8484 33652 8536 33658
rect 8484 33594 8536 33600
rect 8392 31884 8444 31890
rect 8392 31826 8444 31832
rect 8024 31816 8076 31822
rect 8024 31758 8076 31764
rect 7840 31680 7892 31686
rect 7840 31622 7892 31628
rect 7932 31680 7984 31686
rect 7932 31622 7984 31628
rect 7852 29238 7880 31622
rect 7944 31346 7972 31622
rect 8036 31482 8064 31758
rect 8024 31476 8076 31482
rect 8024 31418 8076 31424
rect 7932 31340 7984 31346
rect 7932 31282 7984 31288
rect 7944 30938 7972 31282
rect 8404 31142 8432 31826
rect 8496 31482 8524 33594
rect 8772 33522 8800 33798
rect 8760 33516 8812 33522
rect 8760 33458 8812 33464
rect 8668 32972 8720 32978
rect 8668 32914 8720 32920
rect 8680 32230 8708 32914
rect 8772 32502 8800 33458
rect 8760 32496 8812 32502
rect 8760 32438 8812 32444
rect 8668 32224 8720 32230
rect 8668 32166 8720 32172
rect 8484 31476 8536 31482
rect 8484 31418 8536 31424
rect 8496 31278 8524 31418
rect 8484 31272 8536 31278
rect 8536 31232 8616 31260
rect 8484 31214 8536 31220
rect 8392 31136 8444 31142
rect 8392 31078 8444 31084
rect 7932 30932 7984 30938
rect 7932 30874 7984 30880
rect 8208 30864 8260 30870
rect 8208 30806 8260 30812
rect 8220 29850 8248 30806
rect 8208 29844 8260 29850
rect 8208 29786 8260 29792
rect 8404 29714 8432 31078
rect 8484 30184 8536 30190
rect 8484 30126 8536 30132
rect 8208 29708 8260 29714
rect 8208 29650 8260 29656
rect 8392 29708 8444 29714
rect 8392 29650 8444 29656
rect 7840 29232 7892 29238
rect 7840 29174 7892 29180
rect 7656 29028 7708 29034
rect 7760 29022 7972 29050
rect 7656 28970 7708 28976
rect 7472 28756 7524 28762
rect 7472 28698 7524 28704
rect 7656 28552 7708 28558
rect 7656 28494 7708 28500
rect 7668 27946 7696 28494
rect 7656 27940 7708 27946
rect 7656 27882 7708 27888
rect 7668 27674 7696 27882
rect 7656 27668 7708 27674
rect 7656 27610 7708 27616
rect 7748 27532 7800 27538
rect 7748 27474 7800 27480
rect 7840 27532 7892 27538
rect 7840 27474 7892 27480
rect 7760 27062 7788 27474
rect 7748 27056 7800 27062
rect 7748 26998 7800 27004
rect 7748 26920 7800 26926
rect 7852 26908 7880 27474
rect 7800 26880 7880 26908
rect 7748 26862 7800 26868
rect 7760 26586 7788 26862
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7760 26314 7788 26522
rect 7944 26432 7972 29022
rect 8220 28966 8248 29650
rect 8496 29510 8524 30126
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8300 29232 8352 29238
rect 8300 29174 8352 29180
rect 8208 28960 8260 28966
rect 8208 28902 8260 28908
rect 8024 27872 8076 27878
rect 8024 27814 8076 27820
rect 8036 26994 8064 27814
rect 8024 26988 8076 26994
rect 8024 26930 8076 26936
rect 8024 26444 8076 26450
rect 7944 26404 8024 26432
rect 8024 26386 8076 26392
rect 8116 26444 8168 26450
rect 8116 26386 8168 26392
rect 7748 26308 7800 26314
rect 7748 26250 7800 26256
rect 8036 25906 8064 26386
rect 8024 25900 8076 25906
rect 8024 25842 8076 25848
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 7748 25424 7800 25430
rect 7748 25366 7800 25372
rect 7760 24614 7788 25366
rect 7944 24954 7972 25638
rect 8128 25498 8156 26386
rect 8116 25492 8168 25498
rect 8116 25434 8168 25440
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7668 23322 7696 24006
rect 7656 23316 7708 23322
rect 7656 23258 7708 23264
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7484 18834 7512 19994
rect 7760 19514 7788 24550
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7852 23322 7880 24142
rect 7944 23633 7972 24890
rect 8024 24268 8076 24274
rect 8024 24210 8076 24216
rect 7930 23624 7986 23633
rect 7930 23559 7986 23568
rect 8036 23526 8064 24210
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 7840 23316 7892 23322
rect 7840 23258 7892 23264
rect 8036 23254 8064 23462
rect 8024 23248 8076 23254
rect 8024 23190 8076 23196
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 7944 22438 7972 23054
rect 7932 22432 7984 22438
rect 7932 22374 7984 22380
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7852 21146 7880 21966
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7852 19514 7880 19858
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7852 19334 7880 19450
rect 7668 19306 7880 19334
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7378 18728 7434 18737
rect 7378 18663 7434 18672
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 18154 7236 18566
rect 7484 18426 7512 18770
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7668 18358 7696 19306
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 18970 7788 19110
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7196 18148 7248 18154
rect 7196 18090 7248 18096
rect 7288 18148 7340 18154
rect 7288 18090 7340 18096
rect 7208 16794 7236 18090
rect 7300 17542 7328 18090
rect 7656 18080 7708 18086
rect 7760 18068 7788 18906
rect 7708 18040 7788 18068
rect 7656 18022 7708 18028
rect 7668 17814 7696 18022
rect 7656 17808 7708 17814
rect 7656 17750 7708 17756
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7300 16726 7328 16934
rect 7576 16794 7604 17614
rect 7668 16998 7696 17750
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7288 16720 7340 16726
rect 7288 16662 7340 16668
rect 7576 16114 7604 16730
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7012 16040 7064 16046
rect 7668 15994 7696 16934
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7012 15982 7064 15988
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6932 14890 6960 15370
rect 7024 15366 7052 15982
rect 7576 15966 7696 15994
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7024 14890 7052 15098
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 7576 14822 7604 15966
rect 7760 15502 7788 16458
rect 7852 15994 7880 17274
rect 7944 16590 7972 22374
rect 8036 17338 8064 23190
rect 8116 23180 8168 23186
rect 8220 23168 8248 28902
rect 8312 28558 8340 29174
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 8496 27606 8524 29446
rect 8484 27600 8536 27606
rect 8484 27542 8536 27548
rect 8588 27452 8616 31232
rect 8680 30258 8708 32166
rect 8668 30252 8720 30258
rect 8668 30194 8720 30200
rect 8864 30138 8892 34002
rect 9404 33992 9456 33998
rect 9404 33934 9456 33940
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 9312 33448 9364 33454
rect 9312 33390 9364 33396
rect 9128 33312 9180 33318
rect 9128 33254 9180 33260
rect 9140 32842 9168 33254
rect 9324 33114 9352 33390
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9416 32978 9444 33934
rect 9600 33930 9628 39630
rect 9954 39520 10010 39630
rect 11334 39658 11390 40000
rect 12622 39658 12678 40000
rect 14002 39658 14058 40000
rect 11334 39630 11468 39658
rect 11334 39520 11390 39630
rect 9772 36032 9824 36038
rect 9772 35974 9824 35980
rect 9784 35834 9812 35974
rect 9772 35828 9824 35834
rect 9772 35770 9824 35776
rect 9680 35488 9732 35494
rect 9680 35430 9732 35436
rect 9692 35154 9720 35430
rect 11440 35154 11468 39630
rect 12452 39630 12678 39658
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 9680 35148 9732 35154
rect 9680 35090 9732 35096
rect 11428 35148 11480 35154
rect 11428 35090 11480 35096
rect 9692 34746 9720 35090
rect 9862 35048 9918 35057
rect 9772 35012 9824 35018
rect 9824 34992 9862 35000
rect 9824 34983 9918 34992
rect 9824 34972 9904 34983
rect 9772 34954 9824 34960
rect 9680 34740 9732 34746
rect 9680 34682 9732 34688
rect 10784 34536 10836 34542
rect 10784 34478 10836 34484
rect 11426 34504 11482 34513
rect 9956 34060 10008 34066
rect 9956 34002 10008 34008
rect 9588 33924 9640 33930
rect 9588 33866 9640 33872
rect 9968 33658 9996 34002
rect 9496 33652 9548 33658
rect 9496 33594 9548 33600
rect 9956 33652 10008 33658
rect 9956 33594 10008 33600
rect 9508 33153 9536 33594
rect 9680 33584 9732 33590
rect 9680 33526 9732 33532
rect 10600 33584 10652 33590
rect 10600 33526 10652 33532
rect 9588 33312 9640 33318
rect 9588 33254 9640 33260
rect 9494 33144 9550 33153
rect 9494 33079 9550 33088
rect 9496 33040 9548 33046
rect 9600 33028 9628 33254
rect 9548 33000 9628 33028
rect 9496 32982 9548 32988
rect 9404 32972 9456 32978
rect 9404 32914 9456 32920
rect 9128 32836 9180 32842
rect 9128 32778 9180 32784
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8944 32428 8996 32434
rect 8944 32370 8996 32376
rect 8956 32026 8984 32370
rect 9324 32298 9352 32710
rect 9312 32292 9364 32298
rect 9312 32234 9364 32240
rect 9508 32026 9536 32982
rect 8944 32020 8996 32026
rect 8944 31962 8996 31968
rect 9496 32020 9548 32026
rect 9496 31962 9548 31968
rect 9588 31952 9640 31958
rect 9588 31894 9640 31900
rect 9404 31816 9456 31822
rect 9404 31758 9456 31764
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9128 31204 9180 31210
rect 9128 31146 9180 31152
rect 8944 31136 8996 31142
rect 8944 31078 8996 31084
rect 8956 30870 8984 31078
rect 8944 30864 8996 30870
rect 8944 30806 8996 30812
rect 9140 30802 9168 31146
rect 9312 31136 9364 31142
rect 9312 31078 9364 31084
rect 9128 30796 9180 30802
rect 9128 30738 9180 30744
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8772 30110 8892 30138
rect 8772 29782 8800 30110
rect 8852 30048 8904 30054
rect 8852 29990 8904 29996
rect 8864 29850 8892 29990
rect 8852 29844 8904 29850
rect 8852 29786 8904 29792
rect 8760 29776 8812 29782
rect 8760 29718 8812 29724
rect 8772 29238 8800 29718
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8760 29232 8812 29238
rect 8760 29174 8812 29180
rect 8944 29164 8996 29170
rect 8944 29106 8996 29112
rect 8956 28762 8984 29106
rect 8944 28756 8996 28762
rect 8944 28698 8996 28704
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8852 28008 8904 28014
rect 8852 27950 8904 27956
rect 8404 27424 8616 27452
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 8168 23140 8248 23168
rect 8116 23122 8168 23128
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 8220 21078 8248 21286
rect 8208 21072 8260 21078
rect 8208 21014 8260 21020
rect 8116 20936 8168 20942
rect 8116 20878 8168 20884
rect 8128 19514 8156 20878
rect 8220 20602 8248 21014
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8220 19174 8248 20198
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 8128 17542 8156 18566
rect 8312 18290 8340 26862
rect 8404 21962 8432 27424
rect 8864 27334 8892 27950
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 8864 26790 8892 27270
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9324 26926 9352 31078
rect 9416 30598 9444 31758
rect 9600 31482 9628 31894
rect 9588 31476 9640 31482
rect 9588 31418 9640 31424
rect 9496 30864 9548 30870
rect 9496 30806 9548 30812
rect 9404 30592 9456 30598
rect 9404 30534 9456 30540
rect 9416 29578 9444 30534
rect 9508 30394 9536 30806
rect 9588 30592 9640 30598
rect 9588 30534 9640 30540
rect 9496 30388 9548 30394
rect 9496 30330 9548 30336
rect 9600 30326 9628 30534
rect 9588 30320 9640 30326
rect 9588 30262 9640 30268
rect 9404 29572 9456 29578
rect 9404 29514 9456 29520
rect 9496 28212 9548 28218
rect 9496 28154 9548 28160
rect 9508 27674 9536 28154
rect 9496 27668 9548 27674
rect 9496 27610 9548 27616
rect 9312 26920 9364 26926
rect 9312 26862 9364 26868
rect 8852 26784 8904 26790
rect 8852 26726 8904 26732
rect 8852 26580 8904 26586
rect 8852 26522 8904 26528
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 8588 25362 8616 26318
rect 8668 26036 8720 26042
rect 8668 25978 8720 25984
rect 8576 25356 8628 25362
rect 8576 25298 8628 25304
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8496 23322 8524 23666
rect 8588 23594 8616 23802
rect 8576 23588 8628 23594
rect 8576 23530 8628 23536
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8484 22500 8536 22506
rect 8484 22442 8536 22448
rect 8496 22166 8524 22442
rect 8484 22160 8536 22166
rect 8484 22102 8536 22108
rect 8392 21956 8444 21962
rect 8392 21898 8444 21904
rect 8496 21418 8524 22102
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8404 20058 8432 20334
rect 8496 20330 8524 21354
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8576 19984 8628 19990
rect 8576 19926 8628 19932
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8496 19174 8524 19858
rect 8588 19310 8616 19926
rect 8680 19718 8708 25978
rect 8760 25832 8812 25838
rect 8760 25774 8812 25780
rect 8772 25498 8800 25774
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8760 24880 8812 24886
rect 8760 24822 8812 24828
rect 8772 24206 8800 24822
rect 8864 24818 8892 26522
rect 9324 26314 9352 26862
rect 9692 26450 9720 33526
rect 10324 33516 10376 33522
rect 10324 33458 10376 33464
rect 10046 33144 10102 33153
rect 10046 33079 10102 33088
rect 10060 33046 10088 33079
rect 10048 33040 10100 33046
rect 10048 32982 10100 32988
rect 10336 32910 10364 33458
rect 10612 33454 10640 33526
rect 10600 33448 10652 33454
rect 10600 33390 10652 33396
rect 10612 32978 10640 33390
rect 10796 33114 10824 34478
rect 11426 34439 11482 34448
rect 10968 34060 11020 34066
rect 10968 34002 11020 34008
rect 11244 34060 11296 34066
rect 11244 34002 11296 34008
rect 10980 33454 11008 34002
rect 11256 33522 11284 34002
rect 11440 33998 11468 34439
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11428 33992 11480 33998
rect 11428 33934 11480 33940
rect 11244 33516 11296 33522
rect 11244 33458 11296 33464
rect 10968 33448 11020 33454
rect 10968 33390 11020 33396
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 10784 33108 10836 33114
rect 10784 33050 10836 33056
rect 11428 33108 11480 33114
rect 11428 33050 11480 33056
rect 10600 32972 10652 32978
rect 10600 32914 10652 32920
rect 10324 32904 10376 32910
rect 10324 32846 10376 32852
rect 9956 32836 10008 32842
rect 9956 32778 10008 32784
rect 9968 32570 9996 32778
rect 9956 32564 10008 32570
rect 9956 32506 10008 32512
rect 9864 32360 9916 32366
rect 9864 32302 9916 32308
rect 9876 31210 9904 32302
rect 10336 31754 10364 32846
rect 11440 32434 11468 33050
rect 12164 33040 12216 33046
rect 12164 32982 12216 32988
rect 11612 32972 11664 32978
rect 11612 32914 11664 32920
rect 11520 32904 11572 32910
rect 11520 32846 11572 32852
rect 11532 32774 11560 32846
rect 11520 32768 11572 32774
rect 11520 32710 11572 32716
rect 11428 32428 11480 32434
rect 11428 32370 11480 32376
rect 10416 32360 10468 32366
rect 10416 32302 10468 32308
rect 10428 32026 10456 32302
rect 10508 32224 10560 32230
rect 10508 32166 10560 32172
rect 10416 32020 10468 32026
rect 10416 31962 10468 31968
rect 10520 31958 10548 32166
rect 11532 32008 11560 32710
rect 11624 32570 11652 32914
rect 12176 32570 12204 32982
rect 11612 32564 11664 32570
rect 11612 32506 11664 32512
rect 12164 32564 12216 32570
rect 12164 32506 12216 32512
rect 12176 32366 12204 32506
rect 12164 32360 12216 32366
rect 12164 32302 12216 32308
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11532 31980 11744 32008
rect 10508 31952 10560 31958
rect 10508 31894 10560 31900
rect 11716 31890 11744 31980
rect 11520 31884 11572 31890
rect 11520 31826 11572 31832
rect 11704 31884 11756 31890
rect 11704 31826 11756 31832
rect 10324 31748 10376 31754
rect 10324 31690 10376 31696
rect 10336 31414 10364 31690
rect 11532 31482 11560 31826
rect 11520 31476 11572 31482
rect 11520 31418 11572 31424
rect 10324 31408 10376 31414
rect 10324 31350 10376 31356
rect 10966 31376 11022 31385
rect 10966 31311 11022 31320
rect 9772 31204 9824 31210
rect 9772 31146 9824 31152
rect 9864 31204 9916 31210
rect 9864 31146 9916 31152
rect 9784 30734 9812 31146
rect 10508 30864 10560 30870
rect 10508 30806 10560 30812
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 10416 30728 10468 30734
rect 10416 30670 10468 30676
rect 10048 30048 10100 30054
rect 10048 29990 10100 29996
rect 9864 29776 9916 29782
rect 9864 29718 9916 29724
rect 9876 29306 9904 29718
rect 9864 29300 9916 29306
rect 9864 29242 9916 29248
rect 9876 28694 9904 29242
rect 10060 29170 10088 29990
rect 10324 29572 10376 29578
rect 10324 29514 10376 29520
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 9956 28960 10008 28966
rect 9956 28902 10008 28908
rect 9864 28688 9916 28694
rect 9864 28630 9916 28636
rect 9876 28218 9904 28630
rect 9864 28212 9916 28218
rect 9864 28154 9916 28160
rect 9864 27872 9916 27878
rect 9968 27860 9996 28902
rect 10060 28762 10088 29106
rect 10048 28756 10100 28762
rect 10048 28698 10100 28704
rect 9916 27832 9996 27860
rect 9864 27814 9916 27820
rect 9876 27606 9904 27814
rect 9864 27600 9916 27606
rect 9864 27542 9916 27548
rect 9876 27130 9904 27542
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 10244 27130 10272 27406
rect 10336 27402 10364 29514
rect 10428 29170 10456 30670
rect 10520 30394 10548 30806
rect 10980 30802 11008 31311
rect 11716 31210 11744 31826
rect 11704 31204 11756 31210
rect 11704 31146 11756 31152
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11426 30832 11482 30841
rect 10968 30796 11020 30802
rect 11426 30767 11482 30776
rect 10968 30738 11020 30744
rect 10980 30394 11008 30738
rect 10508 30388 10560 30394
rect 10508 30330 10560 30336
rect 10968 30388 11020 30394
rect 10968 30330 11020 30336
rect 11152 29640 11204 29646
rect 11152 29582 11204 29588
rect 11164 29306 11192 29582
rect 11152 29300 11204 29306
rect 11152 29242 11204 29248
rect 10416 29164 10468 29170
rect 10416 29106 10468 29112
rect 10428 28694 10456 29106
rect 11164 28762 11192 29242
rect 11152 28756 11204 28762
rect 11152 28698 11204 28704
rect 10416 28688 10468 28694
rect 10416 28630 10468 28636
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 11256 28150 11284 28562
rect 11244 28144 11296 28150
rect 11244 28086 11296 28092
rect 10324 27396 10376 27402
rect 10324 27338 10376 27344
rect 9864 27124 9916 27130
rect 9864 27066 9916 27072
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 9680 26444 9732 26450
rect 9680 26386 9732 26392
rect 10324 26444 10376 26450
rect 10324 26386 10376 26392
rect 9312 26308 9364 26314
rect 9312 26250 9364 26256
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 9692 26042 9720 26386
rect 10336 26042 10364 26386
rect 11440 26382 11468 30767
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 12452 29850 12480 39630
rect 12622 39520 12678 39630
rect 13740 39630 14058 39658
rect 13740 34746 13768 39630
rect 14002 39520 14058 39630
rect 15290 39658 15346 40000
rect 15290 39630 15424 39658
rect 15290 39520 15346 39630
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 15396 35057 15424 39630
rect 15474 38176 15530 38185
rect 15474 38111 15530 38120
rect 15488 36038 15516 38111
rect 15476 36032 15528 36038
rect 15476 35974 15528 35980
rect 15382 35048 15438 35057
rect 15382 34983 15438 34992
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 13728 34740 13780 34746
rect 13728 34682 13780 34688
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 12900 32360 12952 32366
rect 12900 32302 12952 32308
rect 12912 31890 12940 32302
rect 12900 31884 12952 31890
rect 12900 31826 12952 31832
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 12440 29844 12492 29850
rect 12440 29786 12492 29792
rect 12072 29708 12124 29714
rect 12072 29650 12124 29656
rect 12084 28966 12112 29650
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 12072 28960 12124 28966
rect 12072 28902 12124 28908
rect 12624 28960 12676 28966
rect 12624 28902 12676 28908
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 12636 28626 12664 28902
rect 12624 28620 12676 28626
rect 12624 28562 12676 28568
rect 12636 27878 12664 28562
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 12624 27872 12676 27878
rect 12624 27814 12676 27820
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11520 26444 11572 26450
rect 11520 26386 11572 26392
rect 11428 26376 11480 26382
rect 11428 26318 11480 26324
rect 10784 26240 10836 26246
rect 10784 26182 10836 26188
rect 9680 26036 9732 26042
rect 9680 25978 9732 25984
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10796 25906 10824 26182
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10416 25832 10468 25838
rect 10416 25774 10468 25780
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 9404 25356 9456 25362
rect 9404 25298 9456 25304
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 8864 24410 8892 24754
rect 9416 24410 9444 25298
rect 9968 24954 9996 25434
rect 10428 25430 10456 25774
rect 10692 25764 10744 25770
rect 10692 25706 10744 25712
rect 10704 25498 10732 25706
rect 11532 25702 11560 26386
rect 11520 25696 11572 25702
rect 11520 25638 11572 25644
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10416 25424 10468 25430
rect 10416 25366 10468 25372
rect 11336 25424 11388 25430
rect 11336 25366 11388 25372
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 9956 24948 10008 24954
rect 9956 24890 10008 24896
rect 8852 24404 8904 24410
rect 8852 24346 8904 24352
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 9864 24336 9916 24342
rect 9864 24278 9916 24284
rect 8760 24200 8812 24206
rect 8760 24142 8812 24148
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 8772 23730 8800 24142
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 9416 23050 9444 23802
rect 9784 23798 9812 24142
rect 9876 23866 9904 24278
rect 10060 24206 10088 25230
rect 11348 24954 11376 25366
rect 11532 25276 11560 25638
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11796 25288 11848 25294
rect 11532 25248 11796 25276
rect 11796 25230 11848 25236
rect 11428 25220 11480 25226
rect 11428 25162 11480 25168
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 11440 24886 11468 25162
rect 10416 24880 10468 24886
rect 10416 24822 10468 24828
rect 11428 24880 11480 24886
rect 11428 24822 11480 24828
rect 10048 24200 10100 24206
rect 10048 24142 10100 24148
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9772 23792 9824 23798
rect 9772 23734 9824 23740
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9692 23322 9720 23462
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9404 23044 9456 23050
rect 9404 22986 9456 22992
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9416 22234 9444 22578
rect 9772 22500 9824 22506
rect 9772 22442 9824 22448
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9784 22166 9812 22442
rect 9968 22166 9996 24006
rect 10060 23730 10088 24142
rect 10048 23724 10100 23730
rect 10048 23666 10100 23672
rect 10046 23624 10102 23633
rect 10046 23559 10102 23568
rect 10140 23588 10192 23594
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 9956 22160 10008 22166
rect 9956 22102 10008 22108
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 9048 21146 9076 21422
rect 9508 21146 9536 21966
rect 9784 21690 9812 22102
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 8760 20936 8812 20942
rect 8760 20878 8812 20884
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 8772 20466 8800 20878
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 9508 20058 9536 20878
rect 9876 20602 9904 21014
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 10060 20058 10088 23559
rect 10140 23530 10192 23536
rect 10152 22982 10180 23530
rect 10140 22976 10192 22982
rect 10140 22918 10192 22924
rect 10232 22976 10284 22982
rect 10232 22918 10284 22924
rect 10152 22778 10180 22918
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 10244 22642 10272 22918
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 10232 22500 10284 22506
rect 10428 22488 10456 24822
rect 11808 24818 11836 25230
rect 11796 24812 11848 24818
rect 11796 24754 11848 24760
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10704 24070 10732 24618
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 11256 23730 11284 24210
rect 11244 23724 11296 23730
rect 11244 23666 11296 23672
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 10692 23180 10744 23186
rect 10692 23122 10744 23128
rect 10704 23089 10732 23122
rect 10690 23080 10746 23089
rect 10690 23015 10746 23024
rect 10704 22778 10732 23015
rect 10692 22772 10744 22778
rect 10284 22460 10456 22488
rect 10520 22732 10692 22760
rect 10232 22442 10284 22448
rect 10140 21412 10192 21418
rect 10140 21354 10192 21360
rect 10152 21146 10180 21354
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 10244 20466 10272 22442
rect 10416 21616 10468 21622
rect 10416 21558 10468 21564
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10336 20330 10364 21082
rect 10232 20324 10284 20330
rect 10232 20266 10284 20272
rect 10324 20324 10376 20330
rect 10324 20266 10376 20272
rect 10244 20058 10272 20266
rect 9496 20052 9548 20058
rect 9496 19994 9548 20000
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 8850 19952 8906 19961
rect 10336 19922 10364 20266
rect 8850 19887 8906 19896
rect 9588 19916 9640 19922
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8484 19168 8536 19174
rect 8668 19168 8720 19174
rect 8536 19128 8616 19156
rect 8484 19110 8536 19116
rect 8588 18630 8616 19128
rect 8668 19110 8720 19116
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8128 17066 8156 17478
rect 8024 17060 8076 17066
rect 8024 17002 8076 17008
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 8036 16794 8064 17002
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8220 16726 8248 17478
rect 8404 17202 8432 18090
rect 8588 17762 8616 18566
rect 8680 18290 8708 19110
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8680 17882 8708 18226
rect 8668 17876 8720 17882
rect 8668 17818 8720 17824
rect 8588 17734 8708 17762
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8588 17270 8616 17614
rect 8576 17264 8628 17270
rect 8576 17206 8628 17212
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 8128 16250 8156 16662
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8220 16114 8248 16662
rect 8404 16590 8432 17138
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8680 16046 8708 17734
rect 8772 16697 8800 19110
rect 8758 16688 8814 16697
rect 8758 16623 8814 16632
rect 8668 16040 8720 16046
rect 7852 15966 8156 15994
rect 8668 15982 8720 15988
rect 7840 15632 7892 15638
rect 7840 15574 7892 15580
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6644 13456 6696 13462
rect 6748 13444 6776 13670
rect 6696 13416 6776 13444
rect 6644 13398 6696 13404
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6196 12306 6224 12718
rect 6748 12646 6776 13416
rect 6840 12986 6868 14214
rect 7116 13530 7144 14486
rect 7576 13802 7604 14758
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 11558 6224 12242
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6090 10160 6146 10169
rect 6090 10095 6092 10104
rect 6144 10095 6146 10104
rect 6196 10112 6224 11494
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6656 11218 6684 12174
rect 6748 11898 6776 12582
rect 7208 12102 7236 13126
rect 7576 12714 7604 13262
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7576 12442 7604 12650
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6748 11286 6776 11834
rect 7208 11626 7236 12038
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6656 10266 6684 11154
rect 6748 10470 6776 11222
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6276 10124 6328 10130
rect 6196 10084 6276 10112
rect 6092 10066 6144 10072
rect 6276 10066 6328 10072
rect 6104 9382 6132 10066
rect 6288 9722 6316 10066
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6104 8294 6132 8978
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6104 7002 6132 7482
rect 6196 7342 6224 8910
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6656 6866 6684 8910
rect 6748 8294 6776 10406
rect 6932 10198 6960 10542
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7392 9722 7420 10066
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7484 9518 7512 12038
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7576 11354 7604 11494
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7668 10266 7696 15030
rect 7760 14618 7788 15438
rect 7852 15162 7880 15574
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7852 12238 7880 14894
rect 7944 14414 7972 15438
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7944 14006 7972 14350
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 7944 12850 7972 13942
rect 8024 13728 8076 13734
rect 8024 13670 8076 13676
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7944 12458 7972 12786
rect 8036 12714 8064 13670
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 7944 12442 8064 12458
rect 7944 12436 8076 12442
rect 7944 12430 8024 12436
rect 8024 12378 8076 12384
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7852 11830 7880 12174
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7852 11286 7880 11766
rect 7944 11558 7972 12310
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 10033 7604 10066
rect 7562 10024 7618 10033
rect 7562 9959 7618 9968
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6840 6254 6868 9318
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8498 6960 8774
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 8022 7328 8230
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7300 7274 7328 7958
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7300 6934 7328 7210
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6932 6254 6960 6734
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6932 5914 6960 6190
rect 7300 6118 7328 6870
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7116 5778 7144 6054
rect 7300 5846 7328 6054
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7104 5772 7156 5778
rect 7156 5732 7236 5760
rect 7104 5714 7156 5720
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6196 5030 6224 5102
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6196 4729 6224 4966
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6182 4720 6238 4729
rect 6182 4655 6238 4664
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6104 4282 6132 4558
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6196 3738 6224 4422
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6748 3516 6776 3946
rect 6840 3738 6868 4014
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 7024 3670 7052 3878
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 6828 3528 6880 3534
rect 6748 3488 6828 3516
rect 6828 3470 6880 3476
rect 6840 3194 6868 3470
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6656 2582 6684 2790
rect 6840 2650 6868 2926
rect 7024 2922 7052 3606
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6656 2310 6684 2518
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6656 2106 6684 2246
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6090 82 6146 480
rect 6012 54 6146 82
rect 2318 0 2374 54
rect 3238 0 3294 54
rect 4158 0 4214 54
rect 5170 0 5226 54
rect 6090 0 6146 54
rect 7010 82 7066 480
rect 7116 82 7144 4966
rect 7208 4826 7236 5732
rect 7300 5098 7328 5782
rect 7484 5234 7512 9454
rect 7576 9178 7604 9959
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 8036 9586 8064 9658
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 8036 8974 8064 9318
rect 8128 9194 8156 15966
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8220 12374 8248 14962
rect 8404 12889 8432 15846
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8496 14618 8524 14962
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8484 13728 8536 13734
rect 8588 13705 8616 13874
rect 8680 13734 8708 15982
rect 8772 15570 8800 16623
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8668 13728 8720 13734
rect 8484 13670 8536 13676
rect 8574 13696 8630 13705
rect 8496 13190 8524 13670
rect 8668 13670 8720 13676
rect 8574 13631 8630 13640
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8390 12880 8446 12889
rect 8390 12815 8446 12824
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8404 10810 8432 11086
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8404 9450 8432 9862
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8128 9166 8340 9194
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 7546 7788 8230
rect 8036 8090 8064 8910
rect 8128 8634 8156 9046
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7300 4154 7328 5034
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7852 4185 7880 4966
rect 8036 4758 8064 5034
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7208 4126 7328 4154
rect 7838 4176 7894 4185
rect 7208 4010 7236 4126
rect 7838 4111 7894 4120
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7852 2650 7880 4111
rect 8128 4049 8156 4558
rect 8114 4040 8170 4049
rect 8114 3975 8170 3984
rect 8128 3738 8156 3975
rect 8220 3942 8248 4694
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8220 3738 8248 3878
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7010 54 7144 82
rect 7930 82 7986 480
rect 8220 82 8248 3062
rect 8312 2854 8340 9166
rect 8404 8294 8432 9386
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8588 7954 8616 13631
rect 8772 12764 8800 14418
rect 8864 14346 8892 19887
rect 9588 19858 9640 19864
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 9600 19378 9628 19858
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9600 17338 9628 18022
rect 9784 17814 9812 18022
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 9416 16114 9444 16390
rect 9508 16114 9536 17206
rect 9600 17048 9628 17274
rect 9680 17060 9732 17066
rect 9600 17020 9680 17048
rect 9680 17002 9732 17008
rect 9784 16794 9812 17750
rect 9876 17542 9904 17750
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9876 17338 9904 17478
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9312 15972 9364 15978
rect 9312 15914 9364 15920
rect 9324 15638 9352 15914
rect 9416 15706 9444 16050
rect 9600 15910 9628 16594
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9312 15632 9364 15638
rect 9312 15574 9364 15580
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 9324 15162 9352 15574
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8864 13530 8892 13874
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8864 12986 8892 13194
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 9416 12782 9444 15506
rect 9508 15026 9536 15642
rect 10060 15502 10088 17614
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9784 14346 9812 15438
rect 10060 14890 10088 15438
rect 10244 15026 10272 17002
rect 10336 15892 10364 19654
rect 10428 18222 10456 21558
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10520 16046 10548 22732
rect 10692 22714 10744 22720
rect 11520 22568 11572 22574
rect 11520 22510 11572 22516
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10600 22160 10652 22166
rect 10600 22102 10652 22108
rect 10612 21622 10640 22102
rect 10796 22030 10824 22374
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10600 21616 10652 21622
rect 10600 21558 10652 21564
rect 10612 21078 10640 21558
rect 10796 21554 10824 21830
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10796 21146 10824 21490
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10600 21072 10652 21078
rect 10600 21014 10652 21020
rect 10888 20942 10916 21830
rect 11072 21010 11100 21898
rect 11256 21350 11284 22034
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 11072 20262 11100 20946
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10612 19174 10640 19858
rect 10600 19168 10652 19174
rect 10600 19110 10652 19116
rect 10612 16658 10640 19110
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10704 16658 10732 17070
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10704 16250 10732 16594
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10508 16040 10560 16046
rect 10560 16000 10640 16028
rect 10508 15982 10560 15988
rect 10336 15864 10548 15892
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 9876 14550 9904 14826
rect 10244 14550 10272 14826
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9876 14074 9904 14486
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 9508 12986 9536 13738
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 8852 12776 8904 12782
rect 8772 12736 8852 12764
rect 8852 12718 8904 12724
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8680 11762 8708 12650
rect 8864 12238 8892 12718
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8680 11354 8708 11698
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8864 10674 8892 12174
rect 9416 12102 9444 12718
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 9692 11898 9720 12242
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9784 11762 9812 12378
rect 10060 12170 10088 13262
rect 10152 12306 10180 13738
rect 10336 13734 10364 14350
rect 10520 13977 10548 15864
rect 10506 13968 10562 13977
rect 10506 13903 10562 13912
rect 10520 13870 10548 13903
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10336 13530 10364 13670
rect 10520 13530 10548 13806
rect 10612 13705 10640 16000
rect 10796 15570 10824 16118
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 14890 10732 15302
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10704 14618 10732 14826
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10598 13696 10654 13705
rect 10598 13631 10654 13640
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 10244 12918 10272 13398
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 10152 11898 10180 12242
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 8956 11354 8984 11698
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 9784 11286 9812 11494
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 9692 10810 9720 11018
rect 9784 10810 9812 11222
rect 10612 11150 10640 11494
rect 10796 11286 10824 15030
rect 10888 12782 10916 18158
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10980 16726 11008 16934
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8680 10266 8708 10406
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 10796 10130 10824 11222
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8680 9110 8708 9386
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8588 7546 8616 7890
rect 8680 7750 8708 9046
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8498 8800 8774
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8864 8022 8892 9522
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 9600 7886 9628 9590
rect 9692 9178 9720 9862
rect 10796 9722 10824 10066
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9692 8090 9720 9114
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9876 8634 9904 9046
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 10060 8566 10088 8910
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9784 8022 9812 8230
rect 9968 8022 9996 8434
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8588 6934 8616 7210
rect 8956 6934 8984 7346
rect 9600 6934 9628 7822
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9692 7188 9720 7686
rect 9784 7546 9812 7958
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 9692 7160 9812 7188
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8496 5846 8524 6258
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8588 5914 8616 6122
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8772 5846 8800 6802
rect 9402 6760 9458 6769
rect 9402 6695 9458 6704
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8956 5778 8984 6326
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9416 5234 9444 6695
rect 9692 6458 9720 6938
rect 9784 6934 9812 7160
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9784 6458 9812 6870
rect 10060 6798 10088 7414
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 10060 6390 10088 6734
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8864 4214 8892 4558
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8864 3534 8892 4150
rect 9324 4146 9352 4762
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8852 3528 8904 3534
rect 9416 3482 9444 5034
rect 9508 4826 9536 5510
rect 9600 5370 9628 5714
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 8852 3470 8904 3476
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8588 2582 8616 3470
rect 8864 3194 8892 3470
rect 9324 3454 9444 3482
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 9324 2446 9352 3454
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 3058 9444 3334
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9416 2650 9444 2994
rect 9508 2922 9536 4558
rect 9600 4185 9628 5102
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9876 4282 9904 4626
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9586 4176 9642 4185
rect 9586 4111 9642 4120
rect 9600 4078 9628 4111
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9876 3942 9904 4218
rect 9968 4154 9996 5306
rect 10060 5166 10088 6326
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10152 4690 10180 9658
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10428 7410 10456 8502
rect 10692 8492 10744 8498
rect 10796 8480 10824 8774
rect 10744 8452 10824 8480
rect 10692 8434 10744 8440
rect 10796 8090 10824 8452
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10428 7002 10456 7346
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 9968 4126 10088 4154
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9876 3670 9904 3878
rect 9968 3670 9996 3946
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9876 3194 9904 3606
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 7930 54 8248 82
rect 8942 128 8998 480
rect 8942 76 8944 128
rect 8996 76 8998 128
rect 7010 0 7066 54
rect 7930 0 7986 54
rect 8942 0 8998 76
rect 9862 82 9918 480
rect 10060 82 10088 4126
rect 10520 4049 10548 4422
rect 10506 4040 10562 4049
rect 10140 4004 10192 4010
rect 10506 3975 10562 3984
rect 10140 3946 10192 3952
rect 10152 2582 10180 3946
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10336 3058 10364 3402
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 9862 54 10088 82
rect 10704 82 10732 5238
rect 10980 2514 11008 12582
rect 11072 10062 11100 20198
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11072 9654 11100 9998
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11256 9081 11284 21286
rect 11532 17338 11560 22510
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 12636 22098 12664 27814
rect 14830 27296 14886 27305
rect 14289 27228 14585 27248
rect 14830 27231 14886 27240
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14844 24410 14872 27231
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11532 17134 11560 17274
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 15474 16280 15530 16289
rect 15474 16215 15530 16224
rect 15488 16182 15516 16215
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11348 15162 11376 15506
rect 11716 15162 11744 15506
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11440 13870 11468 15098
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11532 13734 11560 14418
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 11532 12850 11560 13670
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 13464 12306 13492 13670
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 13634 12744 13690 12753
rect 13634 12679 13690 12688
rect 13648 12442 13676 12679
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13464 11898 13492 12242
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 12360 9110 12388 9862
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 12348 9104 12400 9110
rect 11242 9072 11298 9081
rect 12348 9046 12400 9052
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 11242 9007 11244 9016
rect 11296 9007 11298 9016
rect 11244 8978 11296 8984
rect 11256 8634 11284 8978
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11256 7188 11284 7890
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 11336 7200 11388 7206
rect 11256 7160 11336 7188
rect 11336 7142 11388 7148
rect 11348 5778 11376 7142
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11256 4282 11284 4626
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 11808 3194 11836 3538
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 10782 82 10838 480
rect 10704 54 10838 82
rect 11532 82 11560 2246
rect 11702 82 11758 480
rect 11808 134 11836 2246
rect 12636 2009 12664 2450
rect 12622 2000 12678 2009
rect 12622 1935 12678 1944
rect 11532 54 11758 82
rect 11796 128 11848 134
rect 11796 70 11848 76
rect 12714 82 12770 480
rect 12820 82 12848 3334
rect 12912 3194 12940 3538
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 12912 2446 12940 3130
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 9862 0 9918 54
rect 10782 0 10838 54
rect 11702 0 11758 54
rect 12714 54 12848 82
rect 13634 82 13690 480
rect 13740 82 13768 2858
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 13634 54 13768 82
rect 14554 82 14610 480
rect 14660 82 14688 5034
rect 14554 54 14688 82
rect 15474 82 15530 480
rect 15580 82 15608 9046
rect 15474 54 15608 82
rect 12714 0 12770 54
rect 13634 0 13690 54
rect 14554 0 14610 54
rect 15474 0 15530 54
<< via2 >>
rect 110 38664 166 38720
rect 1398 31320 1454 31376
rect 110 28736 166 28792
rect 110 23704 166 23760
rect 1582 30640 1638 30696
rect 1490 23024 1546 23080
rect 110 18672 166 18728
rect 1306 18672 1362 18728
rect 110 13640 166 13696
rect 2318 25880 2374 25936
rect 2778 33088 2834 33144
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3514 35672 3570 35728
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 2962 31320 3018 31376
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 1950 18264 2006 18320
rect 2226 11092 2228 11112
rect 2228 11092 2280 11112
rect 2280 11092 2282 11112
rect 2226 11056 2282 11092
rect 1582 10648 1638 10704
rect 1306 9288 1362 9344
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3330 21800 3386 21856
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3422 20304 3478 20360
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3054 12824 3110 12880
rect 3146 9968 3202 10024
rect 2778 8472 2834 8528
rect 2318 1944 2374 2000
rect 2962 8472 3018 8528
rect 2594 4120 2650 4176
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 4250 26424 4306 26480
rect 4434 23568 4490 23624
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 4066 20304 4122 20360
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 4710 9968 4766 10024
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 4066 5208 4122 5264
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 3146 1808 3202 1864
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 7746 33088 7802 33144
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 7286 26424 7342 26480
rect 6182 25880 6238 25936
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 5446 18264 5502 18320
rect 5170 13912 5226 13968
rect 5446 10104 5502 10160
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 5630 11056 5686 11112
rect 4526 1808 4582 1864
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 7930 23568 7986 23624
rect 7378 18672 7434 18728
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 9862 34992 9918 35048
rect 9494 33088 9550 33144
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 10046 33088 10102 33144
rect 11426 34448 11482 34504
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 10966 31320 11022 31376
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11426 30776 11482 30832
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 15474 38120 15530 38176
rect 15382 34992 15438 35048
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 10046 23568 10102 23624
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 10690 23024 10746 23080
rect 8850 19896 8906 19952
rect 8758 16632 8814 16688
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6090 10124 6146 10160
rect 6090 10104 6092 10124
rect 6092 10104 6144 10124
rect 6144 10104 6146 10124
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 7562 9968 7618 10024
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6182 4664 6238 4720
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 8574 13640 8630 13696
rect 8390 12824 8446 12880
rect 7838 4120 7894 4176
rect 8114 3984 8170 4040
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 10506 13912 10562 13968
rect 10598 13640 10654 13696
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 9402 6704 9458 6760
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 9586 4120 9642 4176
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 10506 3984 10562 4040
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 14830 27240 14886 27296
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 15474 16224 15530 16280
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 13634 12688 13690 12744
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 11242 9036 11298 9072
rect 11242 9016 11244 9036
rect 11244 9016 11296 9036
rect 11296 9016 11298 9036
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12622 1944 12678 2000
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
<< metal3 >>
rect 0 38720 480 38752
rect 0 38664 110 38720
rect 166 38664 480 38720
rect 0 38632 480 38664
rect 15520 38181 16000 38208
rect 15469 38178 16000 38181
rect 15388 38176 16000 38178
rect 15388 38120 15474 38176
rect 15530 38120 16000 38176
rect 15388 38118 16000 38120
rect 15469 38115 16000 38118
rect 15520 38088 16000 38115
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 0 36184 480 36304
rect 62 35730 122 36184
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 3509 35730 3575 35733
rect 62 35728 3575 35730
rect 62 35672 3514 35728
rect 3570 35672 3575 35728
rect 62 35670 3575 35672
rect 3509 35667 3575 35670
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 9857 35050 9923 35053
rect 15377 35050 15443 35053
rect 9857 35048 15443 35050
rect 9857 34992 9862 35048
rect 9918 34992 15382 35048
rect 15438 34992 15443 35048
rect 9857 34990 15443 34992
rect 9857 34987 9923 34990
rect 15377 34987 15443 34990
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 11421 34506 11487 34509
rect 15520 34506 16000 34536
rect 11421 34504 16000 34506
rect 11421 34448 11426 34504
rect 11482 34448 16000 34504
rect 11421 34446 16000 34448
rect 11421 34443 11487 34446
rect 15520 34416 16000 34446
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 3610 33760 3930 33761
rect 0 33600 480 33720
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 62 33146 122 33600
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 2773 33146 2839 33149
rect 62 33144 2839 33146
rect 62 33088 2778 33144
rect 2834 33088 2839 33144
rect 62 33086 2839 33088
rect 2773 33083 2839 33086
rect 7741 33146 7807 33149
rect 9489 33146 9555 33149
rect 10041 33146 10107 33149
rect 7741 33144 10107 33146
rect 7741 33088 7746 33144
rect 7802 33088 9494 33144
rect 9550 33088 10046 33144
rect 10102 33088 10107 33144
rect 7741 33086 10107 33088
rect 7741 33083 7807 33086
rect 9489 33083 9555 33086
rect 10041 33083 10107 33086
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 1393 31378 1459 31381
rect 2957 31378 3023 31381
rect 10961 31378 11027 31381
rect 1393 31376 11027 31378
rect 1393 31320 1398 31376
rect 1454 31320 2962 31376
rect 3018 31320 10966 31376
rect 11022 31320 11027 31376
rect 1393 31318 11027 31320
rect 1393 31315 1459 31318
rect 2957 31315 3023 31318
rect 10961 31315 11027 31318
rect 0 31152 480 31272
rect 62 30698 122 31152
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 11421 30834 11487 30837
rect 15520 30834 16000 30864
rect 11421 30832 16000 30834
rect 11421 30776 11426 30832
rect 11482 30776 16000 30832
rect 11421 30774 16000 30776
rect 11421 30771 11487 30774
rect 15520 30744 16000 30774
rect 1577 30698 1643 30701
rect 62 30696 1643 30698
rect 62 30640 1582 30696
rect 1638 30640 1643 30696
rect 62 30638 1643 30640
rect 1577 30635 1643 30638
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 6277 28864 6597 28865
rect 0 28792 480 28824
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 0 28736 110 28792
rect 166 28736 480 28792
rect 0 28704 480 28736
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 14825 27298 14891 27301
rect 15520 27298 16000 27328
rect 14825 27296 16000 27298
rect 14825 27240 14830 27296
rect 14886 27240 16000 27296
rect 14825 27238 16000 27240
rect 14825 27235 14891 27238
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 15520 27208 16000 27238
rect 14277 27167 14597 27168
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 4245 26482 4311 26485
rect 7281 26482 7347 26485
rect 4245 26480 7347 26482
rect 4245 26424 4250 26480
rect 4306 26424 7286 26480
rect 7342 26424 7347 26480
rect 4245 26422 7347 26424
rect 4245 26419 4311 26422
rect 7281 26419 7347 26422
rect 0 26212 480 26240
rect 0 26148 60 26212
rect 124 26148 480 26212
rect 0 26120 480 26148
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 54 25876 60 25940
rect 124 25938 130 25940
rect 2313 25938 2379 25941
rect 6177 25938 6243 25941
rect 124 25936 6243 25938
rect 124 25880 2318 25936
rect 2374 25880 6182 25936
rect 6238 25880 6243 25936
rect 124 25878 6243 25880
rect 124 25876 130 25878
rect 2313 25875 2379 25878
rect 6177 25875 6243 25878
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 0 23760 480 23792
rect 0 23704 110 23760
rect 166 23704 480 23760
rect 0 23672 480 23704
rect 4429 23626 4495 23629
rect 7925 23626 7991 23629
rect 4429 23624 7991 23626
rect 4429 23568 4434 23624
rect 4490 23568 7930 23624
rect 7986 23568 7991 23624
rect 4429 23566 7991 23568
rect 4429 23563 4495 23566
rect 7925 23563 7991 23566
rect 10041 23626 10107 23629
rect 15520 23626 16000 23656
rect 10041 23624 16000 23626
rect 10041 23568 10046 23624
rect 10102 23568 16000 23624
rect 10041 23566 16000 23568
rect 10041 23563 10107 23566
rect 15520 23536 16000 23566
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 1485 23082 1551 23085
rect 10685 23082 10751 23085
rect 1485 23080 10751 23082
rect 1485 23024 1490 23080
rect 1546 23024 10690 23080
rect 10746 23024 10751 23080
rect 1485 23022 10751 23024
rect 1485 23019 1551 23022
rect 10685 23019 10751 23022
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 3325 21858 3391 21861
rect 62 21856 3391 21858
rect 62 21800 3330 21856
rect 3386 21800 3391 21856
rect 62 21798 3391 21800
rect 62 21344 122 21798
rect 3325 21795 3391 21798
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 0 21224 480 21344
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 3417 20362 3483 20365
rect 4061 20362 4127 20365
rect 3417 20360 4127 20362
rect 3417 20304 3422 20360
rect 3478 20304 4066 20360
rect 4122 20304 4127 20360
rect 3417 20302 4127 20304
rect 3417 20299 3483 20302
rect 4061 20299 4127 20302
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 8845 19954 8911 19957
rect 15520 19954 16000 19984
rect 8845 19952 16000 19954
rect 8845 19896 8850 19952
rect 8906 19896 16000 19952
rect 8845 19894 16000 19896
rect 8845 19891 8911 19894
rect 15520 19864 16000 19894
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 0 18728 480 18760
rect 0 18672 110 18728
rect 166 18672 480 18728
rect 0 18640 480 18672
rect 1301 18730 1367 18733
rect 7373 18730 7439 18733
rect 1301 18728 7439 18730
rect 1301 18672 1306 18728
rect 1362 18672 7378 18728
rect 7434 18672 7439 18728
rect 1301 18670 7439 18672
rect 1301 18667 1367 18670
rect 7373 18667 7439 18670
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 1945 18322 2011 18325
rect 5441 18322 5507 18325
rect 1945 18320 5507 18322
rect 1945 18264 1950 18320
rect 2006 18264 5446 18320
rect 5502 18264 5507 18320
rect 1945 18262 5507 18264
rect 1945 18259 2011 18262
rect 5441 18259 5507 18262
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 8753 16690 8819 16693
rect 62 16688 8819 16690
rect 62 16632 8758 16688
rect 8814 16632 8819 16688
rect 62 16630 8819 16632
rect 62 16312 122 16630
rect 8753 16627 8819 16630
rect 3610 16352 3930 16353
rect 0 16192 480 16312
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 15520 16285 16000 16312
rect 15469 16282 16000 16285
rect 15388 16280 16000 16282
rect 15388 16224 15474 16280
rect 15530 16224 16000 16280
rect 15388 16222 16000 16224
rect 15469 16219 16000 16222
rect 15520 16192 16000 16219
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 5165 13970 5231 13973
rect 10501 13970 10567 13973
rect 5165 13968 10567 13970
rect 5165 13912 5170 13968
rect 5226 13912 10506 13968
rect 10562 13912 10567 13968
rect 5165 13910 10567 13912
rect 5165 13907 5231 13910
rect 10501 13907 10567 13910
rect 0 13696 480 13728
rect 0 13640 110 13696
rect 166 13640 480 13696
rect 0 13608 480 13640
rect 8569 13698 8635 13701
rect 10593 13698 10659 13701
rect 8569 13696 10659 13698
rect 8569 13640 8574 13696
rect 8630 13640 10598 13696
rect 10654 13640 10659 13696
rect 8569 13638 10659 13640
rect 8569 13635 8635 13638
rect 10593 13635 10659 13638
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 3049 12882 3115 12885
rect 4102 12882 4108 12884
rect 3049 12880 4108 12882
rect 3049 12824 3054 12880
rect 3110 12824 4108 12880
rect 3049 12822 4108 12824
rect 3049 12819 3115 12822
rect 4102 12820 4108 12822
rect 4172 12882 4178 12884
rect 8385 12882 8451 12885
rect 4172 12880 8451 12882
rect 4172 12824 8390 12880
rect 8446 12824 8451 12880
rect 4172 12822 8451 12824
rect 4172 12820 4178 12822
rect 8385 12819 8451 12822
rect 13629 12746 13695 12749
rect 15520 12746 16000 12776
rect 13629 12744 16000 12746
rect 13629 12688 13634 12744
rect 13690 12688 16000 12744
rect 13629 12686 16000 12688
rect 13629 12683 13695 12686
rect 15520 12656 16000 12686
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 0 11160 480 11280
rect 62 10706 122 11160
rect 2221 11114 2287 11117
rect 5625 11114 5691 11117
rect 2221 11112 5691 11114
rect 2221 11056 2226 11112
rect 2282 11056 5630 11112
rect 5686 11056 5691 11112
rect 2221 11054 5691 11056
rect 2221 11051 2287 11054
rect 5625 11051 5691 11054
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 1577 10706 1643 10709
rect 62 10704 1643 10706
rect 62 10648 1582 10704
rect 1638 10648 1643 10704
rect 62 10646 1643 10648
rect 1577 10643 1643 10646
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 5441 10162 5507 10165
rect 6085 10162 6151 10165
rect 5314 10160 6151 10162
rect 5314 10104 5446 10160
rect 5502 10104 6090 10160
rect 6146 10104 6151 10160
rect 5314 10102 6151 10104
rect 5441 10099 5507 10102
rect 6085 10099 6151 10102
rect 3141 10026 3207 10029
rect 4705 10026 4771 10029
rect 7557 10026 7623 10029
rect 3141 10024 7623 10026
rect 3141 9968 3146 10024
rect 3202 9968 4710 10024
rect 4766 9968 7562 10024
rect 7618 9968 7623 10024
rect 3141 9966 7623 9968
rect 3141 9963 3207 9966
rect 4705 9963 4771 9966
rect 7557 9963 7623 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 1301 9346 1367 9349
rect 62 9344 1367 9346
rect 62 9288 1306 9344
rect 1362 9288 1367 9344
rect 62 9286 1367 9288
rect 62 8832 122 9286
rect 1301 9283 1367 9286
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 11237 9074 11303 9077
rect 15520 9074 16000 9104
rect 11237 9072 16000 9074
rect 11237 9016 11242 9072
rect 11298 9016 16000 9072
rect 11237 9014 16000 9016
rect 11237 9011 11303 9014
rect 15520 8984 16000 9014
rect 0 8712 480 8832
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 2773 8530 2839 8533
rect 2957 8530 3023 8533
rect 2773 8528 3023 8530
rect 2773 8472 2778 8528
rect 2834 8472 2962 8528
rect 3018 8472 3023 8528
rect 2773 8470 3023 8472
rect 2773 8467 2839 8470
rect 2957 8467 3023 8470
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 4102 6762 4108 6764
rect 62 6702 4108 6762
rect 62 6248 122 6702
rect 4102 6700 4108 6702
rect 4172 6762 4178 6764
rect 9397 6762 9463 6765
rect 4172 6760 9463 6762
rect 4172 6704 9402 6760
rect 9458 6704 9463 6760
rect 4172 6702 9463 6704
rect 4172 6700 4178 6702
rect 9397 6699 9463 6702
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 0 6128 480 6248
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 15520 5402 16000 5432
rect 14782 5342 16000 5402
rect 4061 5266 4127 5269
rect 14782 5266 14842 5342
rect 15520 5312 16000 5342
rect 4061 5264 14842 5266
rect 4061 5208 4066 5264
rect 4122 5208 14842 5264
rect 4061 5206 14842 5208
rect 4061 5203 4127 5206
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 6177 4722 6243 4725
rect 9438 4722 9444 4724
rect 6177 4720 9444 4722
rect 6177 4664 6182 4720
rect 6238 4664 9444 4720
rect 6177 4662 9444 4664
rect 6177 4659 6243 4662
rect 9438 4660 9444 4662
rect 9508 4660 9514 4724
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 2589 4178 2655 4181
rect 62 4176 2655 4178
rect 62 4120 2594 4176
rect 2650 4120 2655 4176
rect 62 4118 2655 4120
rect 62 3800 122 4118
rect 2589 4115 2655 4118
rect 7833 4178 7899 4181
rect 9581 4178 9647 4181
rect 7833 4176 9647 4178
rect 7833 4120 7838 4176
rect 7894 4120 9586 4176
rect 9642 4120 9647 4176
rect 7833 4118 9647 4120
rect 7833 4115 7899 4118
rect 9581 4115 9647 4118
rect 8109 4042 8175 4045
rect 10501 4042 10567 4045
rect 8109 4040 10567 4042
rect 8109 3984 8114 4040
rect 8170 3984 10506 4040
rect 10562 3984 10567 4040
rect 8109 3982 10567 3984
rect 8109 3979 8175 3982
rect 10501 3979 10567 3982
rect 6277 3840 6597 3841
rect 0 3680 480 3800
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 2313 2002 2379 2005
rect 12617 2002 12683 2005
rect 2313 2000 12683 2002
rect 2313 1944 2318 2000
rect 2374 1944 12622 2000
rect 12678 1944 12683 2000
rect 2313 1942 12683 1944
rect 2313 1939 2379 1942
rect 12617 1939 12683 1942
rect 3141 1866 3207 1869
rect 4521 1866 4587 1869
rect 62 1864 4587 1866
rect 62 1808 3146 1864
rect 3202 1808 4526 1864
rect 4582 1808 4587 1864
rect 62 1806 4587 1808
rect 62 1352 122 1806
rect 3141 1803 3207 1806
rect 4521 1803 4587 1806
rect 9438 1804 9444 1868
rect 9508 1866 9514 1868
rect 15520 1866 16000 1896
rect 9508 1806 16000 1866
rect 9508 1804 9514 1806
rect 15520 1776 16000 1806
rect 0 1232 480 1352
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 60 26148 124 26212
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 60 25876 124 25940
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 4108 12820 4172 12884
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 4108 6700 4172 6764
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 9444 4660 9508 4724
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
rect 9444 1804 9508 1868
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 59 26212 125 26213
rect 59 26148 60 26212
rect 124 26148 125 26212
rect 59 26147 125 26148
rect 62 25941 122 26147
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 59 25940 125 25941
rect 59 25876 60 25940
rect 124 25876 125 25940
rect 59 25875 125 25876
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 4107 12884 4173 12885
rect 4107 12820 4108 12884
rect 4172 12820 4173 12884
rect 4107 12819 4173 12820
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 4110 6765 4170 12819
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 4107 6764 4173 6765
rect 4107 6700 4108 6764
rect 4172 6700 4173 6764
rect 4107 6699 4173 6700
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 9443 4724 9509 4725
rect 9443 4660 9444 4724
rect 9508 4660 9509 4724
rect 9443 4659 9509 4660
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 9446 1869 9506 4659
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
rect 9443 1868 9509 1869
rect 9443 1804 9444 1868
rect 9508 1804 9509 1868
rect 9443 1803 9509 1804
use scs8hd_inv_8  _073_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__073__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_18 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_18
timestamp 1586364061
transform 1 0 2760 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_22
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_25
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_22
timestamp 1586364061
transform 1 0 3128 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_32
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_36
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__C
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_nor3_4  _156_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 1234 592
use scs8hd_nor3_4  _155_
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_52
timestamp 1586364061
transform 1 0 5888 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_56
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_73
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_81
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _191_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_85
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _197_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_103 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_102
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_115
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_119
timestamp 1586364061
transform 1 0 12052 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_123
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_126
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_130
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_134
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use scs8hd_nor3_4  _157_
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 4324 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_37
timestamp 1586364061
transform 1 0 4508 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_54
timestamp 1586364061
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_58
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 222 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_73
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_77
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _162_
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_119
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_9
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 130 592
use scs8hd_inv_8  _068_
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_nor3_4  _158_
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__158__C
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_32
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _159_
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_or2_4  _072_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 -1 4896
box -38 -48 682 592
use scs8hd_fill_1  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_8  _160_
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_49
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_53
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_66
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_70
timestamp 1586364061
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _161_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_87
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_137
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_inv_8  _108_
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 866 592
use scs8hd_buf_1  _146_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_18
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_22
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_35
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_nand2_4  _109_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_52
timestamp 1586364061
transform 1 0 5888 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_56
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_97
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_108
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_120
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_9
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_12
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_20
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__C
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 774 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _083_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _067_
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use scs8hd_or2_4  _145_
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__098__C
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_60
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _173_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_76
timestamp 1586364061
transform 1 0 8096 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_81
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_89
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_85
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_96
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_108
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_103
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_115
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_11
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 314 592
use scs8hd_or3_4  _080_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_or3_4  _090_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use scs8hd_or3_4  _098_
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_77
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_118
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_130
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_142
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_1  _081_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _070_
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 314 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_21
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _174_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_96
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_12
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_or3_4  _069_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__C
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  _099_
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_52
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_77
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_113
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_or2_4  _171_
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _176_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_94
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_107
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_1  _172_
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__D
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_19
timestamp 1586364061
transform 1 0 2852 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _178_
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _175_
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_48
timestamp 1586364061
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_65
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_70
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_113
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_13
timestamp 1586364061
transform 1 0 2300 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_16
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_1  _076_
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_25
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_21
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_or2_4  _121_
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 682 592
use scs8hd_or4_4  _147_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__C
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__C
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_47
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_60
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_68
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 314 592
use scs8hd_or2_4  _129_
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 682 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_72
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_75
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_85
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_104
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_108
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_1  _120_
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_10
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 406 592
use scs8hd_inv_8  _074_
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_44
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_48
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_52
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6900 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use scs8hd_buf_1  _164_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__D
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_or3_4  _119_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _093_
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_52
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 1050 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_75
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_114
timestamp 1586364061
transform 1 0 11592 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_126
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_10
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_14
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _137_
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_44
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_73
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_131
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_144
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 314 592
use scs8hd_or2_4  _077_
timestamp 1586364061
transform 1 0 2576 0 -1 12512
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 406 592
use scs8hd_or4_4  _095_
timestamp 1586364061
transform 1 0 4140 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__D
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_42
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_59
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_63
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_66
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_81
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_114
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_18
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_43
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_47
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_65
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_69
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_82
timestamp 1586364061
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_81
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_85
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_104
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_108
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_120
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_130
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_142
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6900 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_78
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _078_
timestamp 1586364061
transform 1 0 4140 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_29
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_53
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_57
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_72
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_76
timestamp 1586364061
transform 1 0 8096 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_115
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_127
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_139
timestamp 1586364061
transform 1 0 13892 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_9
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_12
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_19
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_38
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_42
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_49
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_54
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_58
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_90
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_107
timestamp 1586364061
transform 1 0 10948 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_11
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_29
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_63
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_6  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_86
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_143
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_37
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_41
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 5244 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 6900 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_72
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_81
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_108
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_120
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 314 592
use scs8hd_buf_1  _113_
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_23
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_29
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_36
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 4140 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_40
timestamp 1586364061
transform 1 0 4784 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_55
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_66
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_70
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_83
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_87
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_96
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_100
timestamp 1586364061
transform 1 0 10304 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_100
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_104
timestamp 1586364061
transform 1 0 10672 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_121
timestamp 1586364061
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_143
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_143
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_16
timestamp 1586364061
transform 1 0 2576 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_46
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_61
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  FILLER_28_67
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_81
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_85
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_114
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_126
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_138
timestamp 1586364061
transform 1 0 13800 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_44
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_78
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_104
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_108
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_120
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_10
timestamp 1586364061
transform 1 0 2024 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_51
timestamp 1586364061
transform 1 0 5796 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_55
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_61
timestamp 1586364061
transform 1 0 6716 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_79
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_83
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_17
timestamp 1586364061
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_21
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_34
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_38
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_73
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_77
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_90
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_106
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_11
timestamp 1586364061
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_43
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_47
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 406 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_60
timestamp 1586364061
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_77
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_83
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_87
timestamp 1586364061
transform 1 0 9108 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_96
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_100
timestamp 1586364061
transform 1 0 10304 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_107
timestamp 1586364061
transform 1 0 10948 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_119
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_19
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_40
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_29
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_41
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_46
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_50
timestamp 1586364061
transform 1 0 5704 0 -1 21216
box -38 -48 590 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_67
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_71
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_75
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_71
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_90
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_107
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_106
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_120
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_113
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_137
timestamp 1586364061
transform 1 0 13708 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_35_23
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_29
timestamp 1586364061
transform 1 0 3772 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_33
timestamp 1586364061
transform 1 0 4140 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_38
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 406 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 314 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 7268 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_58
timestamp 1586364061
transform 1 0 6440 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_65
timestamp 1586364061
transform 1 0 7084 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_69
timestamp 1586364061
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_73
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_105
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_112
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_120
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_29
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 5428 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_45
timestamp 1586364061
transform 1 0 5244 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_49
timestamp 1586364061
transform 1 0 5612 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_55
timestamp 1586364061
transform 1 0 6164 0 -1 22304
box -38 -48 130 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_65
timestamp 1586364061
transform 1 0 7084 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_69
timestamp 1586364061
transform 1 0 7452 0 -1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_91
timestamp 1586364061
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_113
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 3404 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_37_21
timestamp 1586364061
transform 1 0 3036 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_36
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_40
timestamp 1586364061
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_73
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_78
timestamp 1586364061
transform 1 0 8280 0 1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_143
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4600 0 -1 23392
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_49
timestamp 1586364061
transform 1 0 5612 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_53
timestamp 1586364061
transform 1 0 5980 0 -1 23392
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 23392
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_72
timestamp 1586364061
transform 1 0 7728 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_79
timestamp 1586364061
transform 1 0 8372 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_83
timestamp 1586364061
transform 1 0 8740 0 -1 23392
box -38 -48 774 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_91
timestamp 1586364061
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_96
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_100
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_107
timestamp 1586364061
transform 1 0 10948 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_119
timestamp 1586364061
transform 1 0 12052 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_131
timestamp 1586364061
transform 1 0 13156 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_143
timestamp 1586364061
transform 1 0 14260 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_17
timestamp 1586364061
transform 1 0 2668 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_23
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_38
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_38
timestamp 1586364061
transform 1 0 4600 0 -1 24480
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_52
timestamp 1586364061
transform 1 0 5888 0 -1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_69
timestamp 1586364061
transform 1 0 7452 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_71
timestamp 1586364061
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_75
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_86
timestamp 1586364061
transform 1 0 9016 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_88
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_92
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_105
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_109
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_102
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_106
timestamp 1586364061
transform 1 0 10856 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_113
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_113
timestamp 1586364061
transform 1 0 11500 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_137
timestamp 1586364061
transform 1 0 13708 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_21
timestamp 1586364061
transform 1 0 3036 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_25
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3956 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_29
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_36
timestamp 1586364061
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_40
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_71
timestamp 1586364061
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_75
timestamp 1586364061
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_79
timestamp 1586364061
transform 1 0 8372 0 1 24480
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8832 0 1 24480
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_41_95
timestamp 1586364061
transform 1 0 9844 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_99
timestamp 1586364061
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_112
timestamp 1586364061
transform 1 0 11408 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_116
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_120
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_1  _148_
timestamp 1586364061
transform 1 0 4416 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_4  FILLER_42_39
timestamp 1586364061
transform 1 0 4692 0 -1 25568
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 5060 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_45
timestamp 1586364061
transform 1 0 5244 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_49
timestamp 1586364061
transform 1 0 5612 0 -1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 7176 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_60
timestamp 1586364061
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_64
timestamp 1586364061
transform 1 0 6992 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 8372 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_77
timestamp 1586364061
transform 1 0 8188 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_81
timestamp 1586364061
transform 1 0 8556 0 -1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_85
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_42_91
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_104
timestamp 1586364061
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_108
timestamp 1586364061
transform 1 0 11040 0 -1 25568
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_12  FILLER_42_121
timestamp 1586364061
transform 1 0 12236 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_133
timestamp 1586364061
transform 1 0 13340 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_145
timestamp 1586364061
transform 1 0 14444 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 2944 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_19
timestamp 1586364061
transform 1 0 2852 0 1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_43_22
timestamp 1586364061
transform 1 0 3128 0 1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 4876 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 3864 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_35
timestamp 1586364061
transform 1 0 4324 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_39
timestamp 1586364061
transform 1 0 4692 0 1 25568
box -38 -48 222 592
use scs8hd_buf_1  _071_
timestamp 1586364061
transform 1 0 5060 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 5612 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 5980 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_46
timestamp 1586364061
transform 1 0 5336 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_43_55
timestamp 1586364061
transform 1 0 6164 0 1 25568
box -38 -48 590 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 7176 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 6992 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8740 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 8188 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_75
timestamp 1586364061
transform 1 0 8004 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_79
timestamp 1586364061
transform 1 0 8372 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 9936 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_94
timestamp 1586364061
transform 1 0 9752 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 10304 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_98
timestamp 1586364061
transform 1 0 10120 0 1 25568
box -38 -48 222 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_111
timestamp 1586364061
transform 1 0 11316 0 1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_43_115
timestamp 1586364061
transform 1 0 11684 0 1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_43_121
timestamp 1586364061
transform 1 0 12236 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_126
timestamp 1586364061
transform 1 0 12696 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_138
timestamp 1586364061
transform 1 0 13800 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_8  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  FILLER_44_11
timestamp 1586364061
transform 1 0 2116 0 -1 26656
box -38 -48 314 592
use scs8hd_buf_1  _130_
timestamp 1586364061
transform 1 0 2944 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 2392 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 3404 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_16
timestamp 1586364061
transform 1 0 2576 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_44_23
timestamp 1586364061
transform 1 0 3220 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_41
timestamp 1586364061
transform 1 0 4876 0 -1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 5612 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_45
timestamp 1586364061
transform 1 0 5244 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 7268 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_58
timestamp 1586364061
transform 1 0 6440 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_1  FILLER_44_66
timestamp 1586364061
transform 1 0 7176 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_69
timestamp 1586364061
transform 1 0 7452 0 -1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 7820 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 7636 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_82
timestamp 1586364061
transform 1 0 8648 0 -1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 8832 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_86
timestamp 1586364061
transform 1 0 9016 0 -1 26656
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_102
timestamp 1586364061
transform 1 0 10488 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_106
timestamp 1586364061
transform 1 0 10856 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_113
timestamp 1586364061
transform 1 0 11500 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_125
timestamp 1586364061
transform 1 0 12604 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_44_137
timestamp 1586364061
transform 1 0 13708 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_1  FILLER_44_145
timestamp 1586364061
transform 1 0 14444 0 -1 26656
box -38 -48 130 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 2116 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 1932 0 1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 590 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 3128 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 2944 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 2576 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_14
timestamp 1586364061
transform 1 0 2392 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_18
timestamp 1586364061
transform 1 0 2760 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_31
timestamp 1586364061
transform 1 0 3956 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_35
timestamp 1586364061
transform 1 0 4324 0 1 26656
box -38 -48 130 592
use scs8hd_fill_1  FILLER_45_38
timestamp 1586364061
transform 1 0 4600 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5704 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_48
timestamp 1586364061
transform 1 0 5520 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_52
timestamp 1586364061
transform 1 0 5888 0 1 26656
box -38 -48 314 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 7268 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 7084 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_57
timestamp 1586364061
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 8648 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 8280 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_76
timestamp 1586364061
transform 1 0 8096 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_80
timestamp 1586364061
transform 1 0 8464 0 1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 8832 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_93
timestamp 1586364061
transform 1 0 9660 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_97
timestamp 1586364061
transform 1 0 10028 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_104
timestamp 1586364061
transform 1 0 10672 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_108
timestamp 1586364061
transform 1 0 11040 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_120
timestamp 1586364061
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_135
timestamp 1586364061
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_143
timestamp 1586364061
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2116 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 774 592
use scs8hd_decap_3  FILLER_46_11
timestamp 1586364061
transform 1 0 2116 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 774 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 2392 0 -1 27744
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_23
timestamp 1586364061
transform 1 0 3220 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_14
timestamp 1586364061
transform 1 0 2392 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_18
timestamp 1586364061
transform 1 0 2760 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_25
timestamp 1586364061
transform 1 0 3404 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 27744
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4140 0 1 27744
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_29
timestamp 1586364061
transform 1 0 3772 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_47
timestamp 1586364061
transform 1 0 5428 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_44
timestamp 1586364061
transform 1 0 5152 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_48
timestamp 1586364061
transform 1 0 5520 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_52
timestamp 1586364061
transform 1 0 5888 0 1 27744
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_46_64
timestamp 1586364061
transform 1 0 6992 0 -1 27744
box -38 -48 590 592
use scs8hd_fill_2  FILLER_47_57
timestamp 1586364061
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_65
timestamp 1586364061
transform 1 0 7084 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_47_69
timestamp 1586364061
transform 1 0 7452 0 1 27744
box -38 -48 406 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 7728 0 -1 27744
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8096 0 1 27744
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_81
timestamp 1586364061
transform 1 0 8556 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_73
timestamp 1586364061
transform 1 0 7820 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_87
timestamp 1586364061
transform 1 0 9108 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_89
timestamp 1586364061
transform 1 0 9292 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_85
timestamp 1586364061
transform 1 0 8924 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_91
timestamp 1586364061
transform 1 0 9476 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9844 0 1 27744
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_102
timestamp 1586364061
transform 1 0 10488 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_47_106
timestamp 1586364061
transform 1 0 10856 0 1 27744
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_114
timestamp 1586364061
transform 1 0 11592 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_112
timestamp 1586364061
transform 1 0 11408 0 1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_120
timestamp 1586364061
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_126
timestamp 1586364061
transform 1 0 12696 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_46_138
timestamp 1586364061
transform 1 0 13800 0 -1 27744
box -38 -48 774 592
use scs8hd_decap_12  FILLER_47_127
timestamp 1586364061
transform 1 0 12788 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_decap_6  FILLER_47_139
timestamp 1586364061
transform 1 0 13892 0 1 27744
box -38 -48 590 592
use scs8hd_fill_1  FILLER_47_145
timestamp 1586364061
transform 1 0 14444 0 1 27744
box -38 -48 130 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_4  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_19
timestamp 1586364061
transform 1 0 2852 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_23
timestamp 1586364061
transform 1 0 3220 0 -1 28832
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_6  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6164 0 -1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_47
timestamp 1586364061
transform 1 0 5428 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_51
timestamp 1586364061
transform 1 0 5796 0 -1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_66
timestamp 1586364061
transform 1 0 7176 0 -1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_70
timestamp 1586364061
transform 1 0 7544 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_83
timestamp 1586364061
transform 1 0 8740 0 -1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_87
timestamp 1586364061
transform 1 0 9108 0 -1 28832
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_102
timestamp 1586364061
transform 1 0 10488 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_106
timestamp 1586364061
transform 1 0 10856 0 -1 28832
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_48_113
timestamp 1586364061
transform 1 0 11500 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_12  FILLER_48_124
timestamp 1586364061
transform 1 0 12512 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_48_136
timestamp 1586364061
transform 1 0 13616 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_144
timestamp 1586364061
transform 1 0 14352 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 1564 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_7
timestamp 1586364061
transform 1 0 1748 0 1 28832
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_19
timestamp 1586364061
transform 1 0 2852 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_25
timestamp 1586364061
transform 1 0 3404 0 1 28832
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_29
timestamp 1586364061
transform 1 0 3772 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_36
timestamp 1586364061
transform 1 0 4416 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_40
timestamp 1586364061
transform 1 0 4784 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_53
timestamp 1586364061
transform 1 0 5980 0 1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_57
timestamp 1586364061
transform 1 0 6348 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_73
timestamp 1586364061
transform 1 0 7820 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_77
timestamp 1586364061
transform 1 0 8188 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_90
timestamp 1586364061
transform 1 0 9384 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_94
timestamp 1586364061
transform 1 0 9752 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_107
timestamp 1586364061
transform 1 0 10948 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 12052 0 1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_49_111
timestamp 1586364061
transform 1 0 11316 0 1 28832
box -38 -48 774 592
use scs8hd_fill_1  FILLER_49_121
timestamp 1586364061
transform 1 0 12236 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_143
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_7
timestamp 1586364061
transform 1 0 1748 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_19
timestamp 1586364061
transform 1 0 2852 0 -1 29920
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_50_38
timestamp 1586364061
transform 1 0 4600 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_50_50
timestamp 1586364061
transform 1 0 5704 0 -1 29920
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6440 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_60
timestamp 1586364061
transform 1 0 6624 0 -1 29920
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_73
timestamp 1586364061
transform 1 0 7820 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_77
timestamp 1586364061
transform 1 0 8188 0 -1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_50_84
timestamp 1586364061
transform 1 0 8832 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_12  FILLER_50_102
timestamp 1586364061
transform 1 0 10488 0 -1 29920
box -38 -48 1142 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 12052 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_4  FILLER_50_114
timestamp 1586364061
transform 1 0 11592 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_50_118
timestamp 1586364061
transform 1 0 11960 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_123
timestamp 1586364061
transform 1 0 12420 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_135
timestamp 1586364061
transform 1 0 13524 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_50_143
timestamp 1586364061
transform 1 0 14260 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 4600 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_33
timestamp 1586364061
transform 1 0 4140 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_36
timestamp 1586364061
transform 1 0 4416 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_40
timestamp 1586364061
transform 1 0 4784 0 1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 5152 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 4968 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_53
timestamp 1586364061
transform 1 0 5980 0 1 29920
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 6440 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_57
timestamp 1586364061
transform 1 0 6348 0 1 29920
box -38 -48 130 592
use scs8hd_fill_1  FILLER_51_60
timestamp 1586364061
transform 1 0 6624 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_65
timestamp 1586364061
transform 1 0 7084 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_69
timestamp 1586364061
transform 1 0 7452 0 1 29920
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 29920
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_85
timestamp 1586364061
transform 1 0 8924 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_89
timestamp 1586364061
transform 1 0 9292 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_96
timestamp 1586364061
transform 1 0 9936 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_100
timestamp 1586364061
transform 1 0 10304 0 1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_51_104
timestamp 1586364061
transform 1 0 10672 0 1 29920
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_51_112
timestamp 1586364061
transform 1 0 11408 0 1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_51_120
timestamp 1586364061
transform 1 0 12144 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_53_18
timestamp 1586364061
transform 1 0 2760 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 2576 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_22
timestamp 1586364061
transform 1 0 3128 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_52_23
timestamp 1586364061
transform 1 0 3220 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 3404 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 3220 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 774 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 3404 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_34
timestamp 1586364061
transform 1 0 4232 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_38
timestamp 1586364061
transform 1 0 4600 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_37
timestamp 1586364061
transform 1 0 4508 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4324 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4784 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_50
timestamp 1586364061
transform 1 0 5704 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_4  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 406 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 6440 0 -1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_67
timestamp 1586364061
transform 1 0 7268 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_57
timestamp 1586364061
transform 1 0 6348 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 31008
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_71
timestamp 1586364061
transform 1 0 7636 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_71
timestamp 1586364061
transform 1 0 7636 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_75
timestamp 1586364061
transform 1 0 8004 0 1 31008
box -38 -48 406 592
use scs8hd_decap_3  FILLER_53_88
timestamp 1586364061
transform 1 0 9200 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_84
timestamp 1586364061
transform 1 0 8832 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_88
timestamp 1586364061
transform 1 0 9200 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_84
timestamp 1586364061
transform 1 0 8832 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 11224 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_102
timestamp 1586364061
transform 1 0 10488 0 -1 31008
box -38 -48 774 592
use scs8hd_fill_2  FILLER_53_102
timestamp 1586364061
transform 1 0 10488 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_106
timestamp 1586364061
transform 1 0 10856 0 1 31008
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_113
timestamp 1586364061
transform 1 0 11500 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_112
timestamp 1586364061
transform 1 0 11408 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_53_116
timestamp 1586364061
transform 1 0 11776 0 1 31008
box -38 -48 590 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_125
timestamp 1586364061
transform 1 0 12604 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_52_137
timestamp 1586364061
transform 1 0 13708 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_8  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_145
timestamp 1586364061
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_143
timestamp 1586364061
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 2576 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_20
timestamp 1586364061
transform 1 0 2944 0 -1 32096
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4232 0 -1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  FILLER_54_28
timestamp 1586364061
transform 1 0 3680 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_45
timestamp 1586364061
transform 1 0 5244 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_49
timestamp 1586364061
transform 1 0 5612 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_53
timestamp 1586364061
transform 1 0 5980 0 -1 32096
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 32096
box -38 -48 866 592
use scs8hd_fill_1  FILLER_54_61
timestamp 1586364061
transform 1 0 6716 0 -1 32096
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_71
timestamp 1586364061
transform 1 0 7636 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_75
timestamp 1586364061
transform 1 0 8004 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_82
timestamp 1586364061
transform 1 0 8648 0 -1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_86
timestamp 1586364061
transform 1 0 9016 0 -1 32096
box -38 -48 406 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 11224 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_102
timestamp 1586364061
transform 1 0 10488 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_106
timestamp 1586364061
transform 1 0 10856 0 -1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 12420 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_119
timestamp 1586364061
transform 1 0 12052 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_125
timestamp 1586364061
transform 1 0 12604 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_54_137
timestamp 1586364061
transform 1 0 13708 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_8  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 774 592
use scs8hd_decap_3  FILLER_55_11
timestamp 1586364061
transform 1 0 2116 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 2392 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 2760 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_16
timestamp 1586364061
transform 1 0 2576 0 1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_55_20
timestamp 1586364061
transform 1 0 2944 0 1 32096
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4324 0 1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_55_28
timestamp 1586364061
transform 1 0 3680 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_31
timestamp 1586364061
transform 1 0 3956 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_46
timestamp 1586364061
transform 1 0 5336 0 1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_55_50
timestamp 1586364061
transform 1 0 5704 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_53
timestamp 1586364061
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_57
timestamp 1586364061
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8648 0 1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_74
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_78
timestamp 1586364061
transform 1 0 8280 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_93
timestamp 1586364061
transform 1 0 9660 0 1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10396 0 1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_97
timestamp 1586364061
transform 1 0 10028 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 11592 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_112
timestamp 1586364061
transform 1 0 11408 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_116
timestamp 1586364061
transform 1 0 11776 0 1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_55_132
timestamp 1586364061
transform 1 0 13248 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_144
timestamp 1586364061
transform 1 0 14352 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_3  FILLER_56_11
timestamp 1586364061
transform 1 0 2116 0 -1 33184
box -38 -48 314 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 2392 0 -1 33184
box -38 -48 866 592
use scs8hd_decap_8  FILLER_56_23
timestamp 1586364061
transform 1 0 3220 0 -1 33184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 4600 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_36
timestamp 1586364061
transform 1 0 4416 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_40
timestamp 1586364061
transform 1 0 4784 0 -1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_53
timestamp 1586364061
transform 1 0 5980 0 -1 33184
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 -1 33184
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_56_72
timestamp 1586364061
transform 1 0 7728 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_56_83
timestamp 1586364061
transform 1 0 8740 0 -1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8924 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 9384 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_87
timestamp 1586364061
transform 1 0 9108 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_1  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 11132 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_103
timestamp 1586364061
transform 1 0 10580 0 -1 33184
box -38 -48 590 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 11316 0 -1 33184
box -38 -48 866 592
use scs8hd_decap_8  FILLER_56_120
timestamp 1586364061
transform 1 0 12144 0 -1 33184
box -38 -48 774 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 12880 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_131
timestamp 1586364061
transform 1 0 13156 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_56_143
timestamp 1586364061
transform 1 0 14260 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 3220 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 3036 0 1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4784 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 4232 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_32
timestamp 1586364061
transform 1 0 4048 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_36
timestamp 1586364061
transform 1 0 4416 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_57
timestamp 1586364061
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8740 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 8372 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_73
timestamp 1586364061
transform 1 0 7820 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_77
timestamp 1586364061
transform 1 0 8188 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_81
timestamp 1586364061
transform 1 0 8556 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 9936 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_94
timestamp 1586364061
transform 1 0 9752 0 1 33184
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 10488 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 10304 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_111
timestamp 1586364061
transform 1 0 11316 0 1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_57_115
timestamp 1586364061
transform 1 0 11684 0 1 33184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_57_121
timestamp 1586364061
transform 1 0 12236 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_135
timestamp 1586364061
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_143
timestamp 1586364061
transform 1 0 14260 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 3220 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_6  FILLER_58_25
timestamp 1586364061
transform 1 0 3404 0 -1 34272
box -38 -48 590 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 4600 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_6  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_47
timestamp 1586364061
transform 1 0 5428 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_51
timestamp 1586364061
transform 1 0 5796 0 -1 34272
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 34272
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_58_57
timestamp 1586364061
transform 1 0 6348 0 -1 34272
box -38 -48 130 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 8372 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_8  FILLER_58_71
timestamp 1586364061
transform 1 0 7636 0 -1 34272
box -38 -48 774 592
use scs8hd_fill_2  FILLER_58_83
timestamp 1586364061
transform 1 0 8740 0 -1 34272
box -38 -48 222 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_87
timestamp 1586364061
transform 1 0 9108 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_58_91
timestamp 1586364061
transform 1 0 9476 0 -1 34272
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 10672 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_102
timestamp 1586364061
transform 1 0 10488 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_106
timestamp 1586364061
transform 1 0 10856 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_113
timestamp 1586364061
transform 1 0 11500 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_125
timestamp 1586364061
transform 1 0 12604 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_58_137
timestamp 1586364061
transform 1 0 13708 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_58_145
timestamp 1586364061
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3496 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 774 592
use scs8hd_decap_3  FILLER_59_23
timestamp 1586364061
transform 1 0 3220 0 1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_32
timestamp 1586364061
transform 1 0 4048 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 4232 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 314 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 3680 0 1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_60_39
timestamp 1586364061
transform 1 0 4692 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_4  FILLER_60_35
timestamp 1586364061
transform 1 0 4324 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_36
timestamp 1586364061
transform 1 0 4416 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4784 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4784 0 1 34272
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 -1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_55
timestamp 1586364061
transform 1 0 6164 0 1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_60_42
timestamp 1586364061
transform 1 0 4968 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_60_52
timestamp 1586364061
transform 1 0 5888 0 -1 35360
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6716 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_60
timestamp 1586364061
transform 1 0 6624 0 -1 35360
box -38 -48 130 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 8372 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_73
timestamp 1586364061
transform 1 0 7820 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_77
timestamp 1586364061
transform 1 0 8188 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_60_72
timestamp 1586364061
transform 1 0 7728 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_76
timestamp 1586364061
transform 1 0 8096 0 -1 35360
box -38 -48 406 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_90
timestamp 1586364061
transform 1 0 9384 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  FILLER_59_95
timestamp 1586364061
transform 1 0 9844 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_84
timestamp 1586364061
transform 1 0 8832 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_88
timestamp 1586364061
transform 1 0 9200 0 -1 35360
box -38 -48 406 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 10120 0 1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_101
timestamp 1586364061
transform 1 0 10396 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_97
timestamp 1586364061
transform 1 0 10028 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_109
timestamp 1586364061
transform 1 0 11132 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 12512 0 1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_113
timestamp 1586364061
transform 1 0 11500 0 1 34272
box -38 -48 774 592
use scs8hd_fill_1  FILLER_59_121
timestamp 1586364061
transform 1 0 12236 0 1 34272
box -38 -48 130 592
use scs8hd_fill_1  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_60_121
timestamp 1586364061
transform 1 0 12236 0 -1 35360
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 13064 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_128
timestamp 1586364061
transform 1 0 12880 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_132
timestamp 1586364061
transform 1 0 13248 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_133
timestamp 1586364061
transform 1 0 13340 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_144
timestamp 1586364061
transform 1 0 14352 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_145
timestamp 1586364061
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 4876 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_44
timestamp 1586364061
transform 1 0 5152 0 1 35360
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_56
timestamp 1586364061
transform 1 0 6256 0 1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_61_60
timestamp 1586364061
transform 1 0 6624 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_65
timestamp 1586364061
transform 1 0 7084 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_69
timestamp 1586364061
transform 1 0 7452 0 1 35360
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 1 35360
box -38 -48 222 592
use scs8hd_decap_8  FILLER_61_83
timestamp 1586364061
transform 1 0 8740 0 1 35360
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9476 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_94
timestamp 1586364061
transform 1 0 9752 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_98
timestamp 1586364061
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_110
timestamp 1586364061
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_105
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_117
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_129
timestamp 1586364061
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_4  FILLER_62_141
timestamp 1586364061
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 1232 480 1352 6 address[0]
port 0 nsew default input
rlabel metal2 s 2318 0 2374 480 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 3680 480 3800 6 address[2]
port 2 nsew default input
rlabel metal2 s 662 39520 718 40000 6 address[3]
port 3 nsew default input
rlabel metal2 s 3238 0 3294 480 6 address[4]
port 4 nsew default input
rlabel metal3 s 15520 1776 16000 1896 6 address[5]
port 5 nsew default input
rlabel metal3 s 15520 5312 16000 5432 6 address[6]
port 6 nsew default input
rlabel metal2 s 1950 39520 2006 40000 6 chany_bottom_in[0]
port 7 nsew default input
rlabel metal2 s 3330 39520 3386 40000 6 chany_bottom_in[1]
port 8 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[2]
port 9 nsew default input
rlabel metal2 s 5170 0 5226 480 6 chany_bottom_in[3]
port 10 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chany_bottom_in[4]
port 11 nsew default input
rlabel metal3 s 15520 8984 16000 9104 6 chany_bottom_in[5]
port 12 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chany_bottom_in[6]
port 13 nsew default input
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_in[7]
port 14 nsew default input
rlabel metal2 s 4618 39520 4674 40000 6 chany_bottom_in[8]
port 15 nsew default input
rlabel metal2 s 7010 0 7066 480 6 chany_bottom_out[0]
port 16 nsew default tristate
rlabel metal3 s 0 11160 480 11280 6 chany_bottom_out[1]
port 17 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chany_bottom_out[2]
port 18 nsew default tristate
rlabel metal2 s 7930 0 7986 480 6 chany_bottom_out[3]
port 19 nsew default tristate
rlabel metal2 s 5998 39520 6054 40000 6 chany_bottom_out[4]
port 20 nsew default tristate
rlabel metal2 s 7286 39520 7342 40000 6 chany_bottom_out[5]
port 21 nsew default tristate
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_out[6]
port 22 nsew default tristate
rlabel metal2 s 8666 39520 8722 40000 6 chany_bottom_out[7]
port 23 nsew default tristate
rlabel metal3 s 15520 12656 16000 12776 6 chany_bottom_out[8]
port 24 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 chany_top_in[0]
port 25 nsew default input
rlabel metal2 s 9862 0 9918 480 6 chany_top_in[1]
port 26 nsew default input
rlabel metal3 s 0 18640 480 18760 6 chany_top_in[2]
port 27 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chany_top_in[3]
port 28 nsew default input
rlabel metal3 s 0 23672 480 23792 6 chany_top_in[4]
port 29 nsew default input
rlabel metal2 s 9954 39520 10010 40000 6 chany_top_in[5]
port 30 nsew default input
rlabel metal3 s 0 26120 480 26240 6 chany_top_in[6]
port 31 nsew default input
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_in[7]
port 32 nsew default input
rlabel metal3 s 0 28704 480 28824 6 chany_top_in[8]
port 33 nsew default input
rlabel metal3 s 15520 16192 16000 16312 6 chany_top_out[0]
port 34 nsew default tristate
rlabel metal3 s 0 31152 480 31272 6 chany_top_out[1]
port 35 nsew default tristate
rlabel metal3 s 0 33600 480 33720 6 chany_top_out[2]
port 36 nsew default tristate
rlabel metal3 s 0 36184 480 36304 6 chany_top_out[3]
port 37 nsew default tristate
rlabel metal2 s 10782 0 10838 480 6 chany_top_out[4]
port 38 nsew default tristate
rlabel metal2 s 12622 39520 12678 40000 6 chany_top_out[5]
port 39 nsew default tristate
rlabel metal2 s 14002 39520 14058 40000 6 chany_top_out[6]
port 40 nsew default tristate
rlabel metal2 s 15290 39520 15346 40000 6 chany_top_out[7]
port 41 nsew default tristate
rlabel metal2 s 11702 0 11758 480 6 chany_top_out[8]
port 42 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 data_in
port 43 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 44 nsew default input
rlabel metal3 s 0 38632 480 38752 6 left_grid_pin_1_
port 45 nsew default tristate
rlabel metal2 s 12714 0 12770 480 6 left_grid_pin_5_
port 46 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 left_grid_pin_9_
port 47 nsew default tristate
rlabel metal3 s 15520 19864 16000 19984 6 right_grid_pin_0_
port 48 nsew default tristate
rlabel metal3 s 15520 30744 16000 30864 6 right_grid_pin_10_
port 49 nsew default tristate
rlabel metal3 s 15520 34416 16000 34536 6 right_grid_pin_12_
port 50 nsew default tristate
rlabel metal3 s 15520 38088 16000 38208 6 right_grid_pin_14_
port 51 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 right_grid_pin_2_
port 52 nsew default tristate
rlabel metal3 s 15520 23536 16000 23656 6 right_grid_pin_4_
port 53 nsew default tristate
rlabel metal3 s 15520 27208 16000 27328 6 right_grid_pin_6_
port 54 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 right_grid_pin_8_
port 55 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 56 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 57 nsew default input
<< end >>
