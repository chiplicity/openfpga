VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 138.600 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.000 2.400 68.600 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.920 2.400 115.520 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 2.720 140.000 3.320 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 31.280 140.000 31.880 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 34.000 140.000 34.600 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 36.720 140.000 37.320 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 39.440 140.000 40.040 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 42.840 140.000 43.440 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 45.560 140.000 46.160 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 48.280 140.000 48.880 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 51.000 140.000 51.600 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 53.720 140.000 54.320 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 57.120 140.000 57.720 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 5.440 140.000 6.040 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 8.160 140.000 8.760 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 10.880 140.000 11.480 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 14.280 140.000 14.880 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 17.000 140.000 17.600 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 19.720 140.000 20.320 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 22.440 140.000 23.040 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 25.160 140.000 25.760 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 28.560 140.000 29.160 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 59.840 140.000 60.440 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 88.400 140.000 89.000 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 91.120 140.000 91.720 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 93.840 140.000 94.440 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 96.560 140.000 97.160 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 99.960 140.000 100.560 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 102.680 140.000 103.280 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 105.400 140.000 106.000 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 108.120 140.000 108.720 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 110.840 140.000 111.440 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 114.240 140.000 114.840 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 62.560 140.000 63.160 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 65.280 140.000 65.880 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 68.000 140.000 68.600 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 71.400 140.000 72.000 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 74.120 140.000 74.720 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 76.840 140.000 77.440 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 79.560 140.000 80.160 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 82.280 140.000 82.880 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 85.680 140.000 86.280 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 136.200 4.970 138.600 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 136.200 39.010 138.600 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 136.200 42.230 138.600 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 136.200 45.910 138.600 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 136.200 49.130 138.600 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 136.200 52.810 138.600 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 136.200 56.030 138.600 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 136.200 59.710 138.600 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 136.200 62.930 138.600 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 136.200 66.150 138.600 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 136.200 69.830 138.600 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 136.200 8.190 138.600 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 136.200 11.870 138.600 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 136.200 15.090 138.600 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 136.200 18.770 138.600 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 136.200 21.990 138.600 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 136.200 25.210 138.600 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 136.200 28.890 138.600 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 136.200 32.110 138.600 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 136.200 35.790 138.600 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 136.200 73.050 138.600 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 136.200 107.090 138.600 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 136.200 110.770 138.600 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 136.200 113.990 138.600 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.390 136.200 117.670 138.600 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 136.200 120.890 138.600 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 136.200 124.110 138.600 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.510 136.200 127.790 138.600 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 136.200 131.010 138.600 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.410 136.200 134.690 138.600 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 136.200 137.910 138.600 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 136.200 76.730 138.600 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.670 136.200 79.950 138.600 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 136.200 83.170 138.600 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 136.200 86.850 138.600 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 136.200 90.070 138.600 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 136.200 93.750 138.600 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 136.200 96.970 138.600 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 136.200 100.650 138.600 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 136.200 103.870 138.600 ;
    END
  END chany_top_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.760 2.400 22.360 ;
    END
  END prog_clk
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 0.000 140.000 0.600 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_top_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 116.960 140.000 117.560 ;
    END
  END right_top_grid_pin_42_
  PIN right_top_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 119.680 140.000 120.280 ;
    END
  END right_top_grid_pin_43_
  PIN right_top_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 122.400 140.000 123.000 ;
    END
  END right_top_grid_pin_44_
  PIN right_top_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 125.120 140.000 125.720 ;
    END
  END right_top_grid_pin_45_
  PIN right_top_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 128.520 140.000 129.120 ;
    END
  END right_top_grid_pin_46_
  PIN right_top_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 131.240 140.000 131.840 ;
    END
  END right_top_grid_pin_47_
  PIN right_top_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 133.960 140.000 134.560 ;
    END
  END right_top_grid_pin_48_
  PIN right_top_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.680 140.000 137.280 ;
    END
  END right_top_grid_pin_49_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 136.200 1.750 138.600 ;
    END
  END top_left_grid_pin_1_
  PIN vpwr
    USE POWER ; 
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 9.240 29.655 126.680 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ; 
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 9.240 52.985 126.680 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 9.395 134.320 126.525 ;
      LAYER met1 ;
        RECT 5.520 9.240 137.930 131.500 ;
      LAYER met2 ;
        RECT 2.030 135.920 4.410 137.165 ;
        RECT 5.250 135.920 7.630 137.165 ;
        RECT 8.470 135.920 11.310 137.165 ;
        RECT 12.150 135.920 14.530 137.165 ;
        RECT 15.370 135.920 18.210 137.165 ;
        RECT 19.050 135.920 21.430 137.165 ;
        RECT 22.270 135.920 24.650 137.165 ;
        RECT 25.490 135.920 28.330 137.165 ;
        RECT 29.170 135.920 31.550 137.165 ;
        RECT 32.390 135.920 35.230 137.165 ;
        RECT 36.070 135.920 38.450 137.165 ;
        RECT 39.290 135.920 41.670 137.165 ;
        RECT 42.510 135.920 45.350 137.165 ;
        RECT 46.190 135.920 48.570 137.165 ;
        RECT 49.410 135.920 52.250 137.165 ;
        RECT 53.090 135.920 55.470 137.165 ;
        RECT 56.310 135.920 59.150 137.165 ;
        RECT 59.990 135.920 62.370 137.165 ;
        RECT 63.210 135.920 65.590 137.165 ;
        RECT 66.430 135.920 69.270 137.165 ;
        RECT 70.110 135.920 72.490 137.165 ;
        RECT 73.330 135.920 76.170 137.165 ;
        RECT 77.010 135.920 79.390 137.165 ;
        RECT 80.230 135.920 82.610 137.165 ;
        RECT 83.450 135.920 86.290 137.165 ;
        RECT 87.130 135.920 89.510 137.165 ;
        RECT 90.350 135.920 93.190 137.165 ;
        RECT 94.030 135.920 96.410 137.165 ;
        RECT 97.250 135.920 100.090 137.165 ;
        RECT 100.930 135.920 103.310 137.165 ;
        RECT 104.150 135.920 106.530 137.165 ;
        RECT 107.370 135.920 110.210 137.165 ;
        RECT 111.050 135.920 113.430 137.165 ;
        RECT 114.270 135.920 117.110 137.165 ;
        RECT 117.950 135.920 120.330 137.165 ;
        RECT 121.170 135.920 123.550 137.165 ;
        RECT 124.390 135.920 127.230 137.165 ;
        RECT 128.070 135.920 130.450 137.165 ;
        RECT 131.290 135.920 134.130 137.165 ;
        RECT 134.970 135.920 137.350 137.165 ;
        RECT 1.540 0.115 137.900 135.920 ;
      LAYER met3 ;
        RECT 1.905 136.280 137.200 137.145 ;
        RECT 1.905 134.960 137.600 136.280 ;
        RECT 1.905 133.560 137.200 134.960 ;
        RECT 1.905 132.240 137.600 133.560 ;
        RECT 1.905 130.840 137.200 132.240 ;
        RECT 1.905 129.520 137.600 130.840 ;
        RECT 1.905 128.120 137.200 129.520 ;
        RECT 1.905 126.120 137.600 128.120 ;
        RECT 1.905 124.720 137.200 126.120 ;
        RECT 1.905 123.400 137.600 124.720 ;
        RECT 1.905 122.000 137.200 123.400 ;
        RECT 1.905 120.680 137.600 122.000 ;
        RECT 1.905 119.280 137.200 120.680 ;
        RECT 1.905 117.960 137.600 119.280 ;
        RECT 1.905 116.560 137.200 117.960 ;
        RECT 1.905 115.920 137.600 116.560 ;
        RECT 2.800 115.240 137.600 115.920 ;
        RECT 2.800 114.520 137.200 115.240 ;
        RECT 1.905 113.840 137.200 114.520 ;
        RECT 1.905 111.840 137.600 113.840 ;
        RECT 1.905 110.440 137.200 111.840 ;
        RECT 1.905 109.120 137.600 110.440 ;
        RECT 1.905 107.720 137.200 109.120 ;
        RECT 1.905 106.400 137.600 107.720 ;
        RECT 1.905 105.000 137.200 106.400 ;
        RECT 1.905 103.680 137.600 105.000 ;
        RECT 1.905 102.280 137.200 103.680 ;
        RECT 1.905 100.960 137.600 102.280 ;
        RECT 1.905 99.560 137.200 100.960 ;
        RECT 1.905 97.560 137.600 99.560 ;
        RECT 1.905 96.160 137.200 97.560 ;
        RECT 1.905 94.840 137.600 96.160 ;
        RECT 1.905 93.440 137.200 94.840 ;
        RECT 1.905 92.120 137.600 93.440 ;
        RECT 1.905 90.720 137.200 92.120 ;
        RECT 1.905 89.400 137.600 90.720 ;
        RECT 1.905 88.000 137.200 89.400 ;
        RECT 1.905 86.680 137.600 88.000 ;
        RECT 1.905 85.280 137.200 86.680 ;
        RECT 1.905 83.280 137.600 85.280 ;
        RECT 1.905 81.880 137.200 83.280 ;
        RECT 1.905 80.560 137.600 81.880 ;
        RECT 1.905 79.160 137.200 80.560 ;
        RECT 1.905 77.840 137.600 79.160 ;
        RECT 1.905 76.440 137.200 77.840 ;
        RECT 1.905 75.120 137.600 76.440 ;
        RECT 1.905 73.720 137.200 75.120 ;
        RECT 1.905 72.400 137.600 73.720 ;
        RECT 1.905 71.000 137.200 72.400 ;
        RECT 1.905 69.000 137.600 71.000 ;
        RECT 2.800 67.600 137.200 69.000 ;
        RECT 1.905 66.280 137.600 67.600 ;
        RECT 1.905 64.880 137.200 66.280 ;
        RECT 1.905 63.560 137.600 64.880 ;
        RECT 1.905 62.160 137.200 63.560 ;
        RECT 1.905 60.840 137.600 62.160 ;
        RECT 1.905 59.440 137.200 60.840 ;
        RECT 1.905 58.120 137.600 59.440 ;
        RECT 1.905 56.720 137.200 58.120 ;
        RECT 1.905 54.720 137.600 56.720 ;
        RECT 1.905 53.320 137.200 54.720 ;
        RECT 1.905 52.000 137.600 53.320 ;
        RECT 1.905 50.600 137.200 52.000 ;
        RECT 1.905 49.280 137.600 50.600 ;
        RECT 1.905 47.880 137.200 49.280 ;
        RECT 1.905 46.560 137.600 47.880 ;
        RECT 1.905 45.160 137.200 46.560 ;
        RECT 1.905 43.840 137.600 45.160 ;
        RECT 1.905 42.440 137.200 43.840 ;
        RECT 1.905 40.440 137.600 42.440 ;
        RECT 1.905 39.040 137.200 40.440 ;
        RECT 1.905 37.720 137.600 39.040 ;
        RECT 1.905 36.320 137.200 37.720 ;
        RECT 1.905 35.000 137.600 36.320 ;
        RECT 1.905 33.600 137.200 35.000 ;
        RECT 1.905 32.280 137.600 33.600 ;
        RECT 1.905 30.880 137.200 32.280 ;
        RECT 1.905 29.560 137.600 30.880 ;
        RECT 1.905 28.160 137.200 29.560 ;
        RECT 1.905 26.160 137.600 28.160 ;
        RECT 1.905 24.760 137.200 26.160 ;
        RECT 1.905 23.440 137.600 24.760 ;
        RECT 1.905 22.760 137.200 23.440 ;
        RECT 2.800 22.040 137.200 22.760 ;
        RECT 2.800 21.360 137.600 22.040 ;
        RECT 1.905 20.720 137.600 21.360 ;
        RECT 1.905 19.320 137.200 20.720 ;
        RECT 1.905 18.000 137.600 19.320 ;
        RECT 1.905 16.600 137.200 18.000 ;
        RECT 1.905 15.280 137.600 16.600 ;
        RECT 1.905 13.880 137.200 15.280 ;
        RECT 1.905 11.880 137.600 13.880 ;
        RECT 1.905 10.480 137.200 11.880 ;
        RECT 1.905 9.160 137.600 10.480 ;
        RECT 1.905 7.760 137.200 9.160 ;
        RECT 1.905 6.440 137.600 7.760 ;
        RECT 1.905 5.040 137.200 6.440 ;
        RECT 1.905 3.720 137.600 5.040 ;
        RECT 1.905 2.320 137.200 3.720 ;
        RECT 1.905 1.000 137.600 2.320 ;
        RECT 1.905 0.135 137.200 1.000 ;
      LAYER met4 ;
        RECT 30.055 9.240 50.985 126.680 ;
        RECT 53.385 9.240 122.985 126.680 ;
      LAYER met5 ;
        RECT 30.020 101.500 120.860 106.500 ;
  END
END sb_0__0_
END LIBRARY

