//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: FPGA Verilog Testbench for Top-level netlist of Design: and2
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Oct  7 01:24:55 2020
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

module and2_autocheck_top_tb;
// ----- Local wires for global ports of FPGA fabric -----
wire [0:0] set;
wire [0:0] reset;
wire [0:0] clk;

// ----- Local wires for I/Os of FPGA fabric -----
wire [0:95] gfpga_pad_GPIO_PAD;



reg [0:0] config_done;
wire [0:0] prog_clock;
reg [0:0] prog_clock_reg;
wire [0:0] op_clock;
reg [0:0] op_clock_reg;
reg [0:0] prog_reset;
reg [0:0] prog_set;
reg [0:0] greset;
reg [0:0] gset;
// ---- Address port for frame-based decoder -----
reg [0:15] address;
// ---- Data input port for frame-based decoder -----
reg [0:0] data_in;
// ---- Wire enable port of frame-based decoders  -----
wire [0:0] enable;
reg [0:0] enable_reg;
	assign enable[0]= ~enable_reg[0] & ~config_done[0];
// ----- Shared inputs -------
	reg [0:0] a;
	reg [0:0] b;

// ----- FPGA fabric outputs -------
	wire [0:0] out_c_fpga;

`ifdef AUTOCHECKED_SIMULATION

// ----- Benchmark outputs -------
	wire [0:0] out_c_benchmark;

// ----- Output vectors checking flags -------
	reg [0:0] out_c_flag;

`endif

// ----- Error counter: Deposit an error for config_done signal is not raised at the beginning -----
	integer nb_error= 1;
// ----- Number of clock cycles in configuration phase: 3807 -----
// ----- Begin configuration done signal generation -----
initial
	begin
		config_done[0] = 1'b0;
	end

// ----- End configuration done signal generation -----

// ----- Begin raw programming clock signal generation -----
initial
	begin
		prog_clock_reg[0] = 1'b0;
	end
always
	begin
		#5	prog_clock_reg[0] = ~prog_clock_reg[0];
	end

// ----- End raw programming clock signal generation -----

// ----- Actual programming clock is triggered only when config_done and prog_reset are disabled -----
	assign prog_clock[0] = prog_clock_reg[0] & (~config_done[0]) & (~prog_reset[0]);

// ----- Begin raw operating clock signal generation -----
initial
	begin
		op_clock_reg[0] = 1'b0;
	end
always wait(~greset)
	begin
		#0.4885859489	op_clock_reg[0] = ~op_clock_reg[0];
	end

// ----- End raw operating clock signal generation -----
// ----- Actual operating clock is triggered only when config_done is enabled -----
	assign op_clock[0] = op_clock_reg[0] & config_done[0];

// ----- Begin programming reset signal generation -----
initial
	begin
		prog_reset[0] = 1'b1;
	#10	prog_reset[0] = 1'b0;
	end

// ----- End programming reset signal generation -----

// ----- Begin programming set signal generation -----
initial
	begin
		prog_set[0] = 1'b1;
	#10	prog_set[0] = 1'b0;
	end

// ----- End programming set signal generation -----

// ----- Begin operating reset signal generation -----
// ----- Reset signal is enabled until the first clock cycle in operation phase -----
initial
	begin
		greset[0] = 1'b1;
	wait(config_done)
	#0.9771718979	greset[0] = 1'b1;
	#1.954343796	greset[0] = 1'b0;
	end

// ----- End operating reset signal generation -----
// ----- Begin operating set signal generation: always disabled -----
initial
	begin
		gset[0] = 1'b0;
	end

// ----- End operating set signal generation: always disabled -----

// ---- Generate enable signal waveform  -----
initial
	begin
		enable_reg[0] = 1'b0;
		#2.5;
		forever enable_reg[0] = #5 ~enable_reg[0];
	end

// ----- Begin connecting global ports of FPGA fabric to stimuli -----
	assign clk[0] = op_clock[0];
	assign reset[0] = greset[0];
	assign set[0] = gset[0];
// ----- End connecting global ports of FPGA fabric to stimuli -----
// ----- FPGA top-level module to be capsulated -----
	fpga_top FPGA_DUT (
		.set(set[0]),
		.reset(reset[0]),
		.clk(clk[0]),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:95]),
		.enable(enable[0]),
		.address(address[0:15]),
		.data_in(data_in[0]));

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input a is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[50] -----
	assign gfpga_pad_GPIO_PAD[50] = a[0];
// ----- Blif Benchmark input b is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[53] -----
	assign gfpga_pad_GPIO_PAD[53] = b[0];
// ----- Blif Benchmark output out_c is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[54] -----
	assign out_c_fpga[0] = gfpga_pad_GPIO_PAD[54];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_GPIO_PAD[0] = 1'b0;
	assign gfpga_pad_GPIO_PAD[1] = 1'b0;
	assign gfpga_pad_GPIO_PAD[2] = 1'b0;
	assign gfpga_pad_GPIO_PAD[3] = 1'b0;
	assign gfpga_pad_GPIO_PAD[4] = 1'b0;
	assign gfpga_pad_GPIO_PAD[5] = 1'b0;
	assign gfpga_pad_GPIO_PAD[6] = 1'b0;
	assign gfpga_pad_GPIO_PAD[7] = 1'b0;
	assign gfpga_pad_GPIO_PAD[8] = 1'b0;
	assign gfpga_pad_GPIO_PAD[9] = 1'b0;
	assign gfpga_pad_GPIO_PAD[10] = 1'b0;
	assign gfpga_pad_GPIO_PAD[11] = 1'b0;
	assign gfpga_pad_GPIO_PAD[12] = 1'b0;
	assign gfpga_pad_GPIO_PAD[13] = 1'b0;
	assign gfpga_pad_GPIO_PAD[14] = 1'b0;
	assign gfpga_pad_GPIO_PAD[15] = 1'b0;
	assign gfpga_pad_GPIO_PAD[16] = 1'b0;
	assign gfpga_pad_GPIO_PAD[17] = 1'b0;
	assign gfpga_pad_GPIO_PAD[18] = 1'b0;
	assign gfpga_pad_GPIO_PAD[19] = 1'b0;
	assign gfpga_pad_GPIO_PAD[20] = 1'b0;
	assign gfpga_pad_GPIO_PAD[21] = 1'b0;
	assign gfpga_pad_GPIO_PAD[22] = 1'b0;
	assign gfpga_pad_GPIO_PAD[23] = 1'b0;
	assign gfpga_pad_GPIO_PAD[24] = 1'b0;
	assign gfpga_pad_GPIO_PAD[25] = 1'b0;
	assign gfpga_pad_GPIO_PAD[26] = 1'b0;
	assign gfpga_pad_GPIO_PAD[27] = 1'b0;
	assign gfpga_pad_GPIO_PAD[28] = 1'b0;
	assign gfpga_pad_GPIO_PAD[29] = 1'b0;
	assign gfpga_pad_GPIO_PAD[30] = 1'b0;
	assign gfpga_pad_GPIO_PAD[31] = 1'b0;
	assign gfpga_pad_GPIO_PAD[32] = 1'b0;
	assign gfpga_pad_GPIO_PAD[33] = 1'b0;
	assign gfpga_pad_GPIO_PAD[34] = 1'b0;
	assign gfpga_pad_GPIO_PAD[35] = 1'b0;
	assign gfpga_pad_GPIO_PAD[36] = 1'b0;
	assign gfpga_pad_GPIO_PAD[37] = 1'b0;
	assign gfpga_pad_GPIO_PAD[38] = 1'b0;
	assign gfpga_pad_GPIO_PAD[39] = 1'b0;
	assign gfpga_pad_GPIO_PAD[40] = 1'b0;
	assign gfpga_pad_GPIO_PAD[41] = 1'b0;
	assign gfpga_pad_GPIO_PAD[42] = 1'b0;
	assign gfpga_pad_GPIO_PAD[43] = 1'b0;
	assign gfpga_pad_GPIO_PAD[44] = 1'b0;
	assign gfpga_pad_GPIO_PAD[45] = 1'b0;
	assign gfpga_pad_GPIO_PAD[46] = 1'b0;
	assign gfpga_pad_GPIO_PAD[47] = 1'b0;
	assign gfpga_pad_GPIO_PAD[48] = 1'b0;
	assign gfpga_pad_GPIO_PAD[49] = 1'b0;
	assign gfpga_pad_GPIO_PAD[51] = 1'b0;
	assign gfpga_pad_GPIO_PAD[52] = 1'b0;
	assign gfpga_pad_GPIO_PAD[55] = 1'b0;
	assign gfpga_pad_GPIO_PAD[56] = 1'b0;
	assign gfpga_pad_GPIO_PAD[57] = 1'b0;
	assign gfpga_pad_GPIO_PAD[58] = 1'b0;
	assign gfpga_pad_GPIO_PAD[59] = 1'b0;
	assign gfpga_pad_GPIO_PAD[60] = 1'b0;
	assign gfpga_pad_GPIO_PAD[61] = 1'b0;
	assign gfpga_pad_GPIO_PAD[62] = 1'b0;
	assign gfpga_pad_GPIO_PAD[63] = 1'b0;
	assign gfpga_pad_GPIO_PAD[64] = 1'b0;
	assign gfpga_pad_GPIO_PAD[65] = 1'b0;
	assign gfpga_pad_GPIO_PAD[66] = 1'b0;
	assign gfpga_pad_GPIO_PAD[67] = 1'b0;
	assign gfpga_pad_GPIO_PAD[68] = 1'b0;
	assign gfpga_pad_GPIO_PAD[69] = 1'b0;
	assign gfpga_pad_GPIO_PAD[70] = 1'b0;
	assign gfpga_pad_GPIO_PAD[71] = 1'b0;
	assign gfpga_pad_GPIO_PAD[72] = 1'b0;
	assign gfpga_pad_GPIO_PAD[73] = 1'b0;
	assign gfpga_pad_GPIO_PAD[74] = 1'b0;
	assign gfpga_pad_GPIO_PAD[75] = 1'b0;
	assign gfpga_pad_GPIO_PAD[76] = 1'b0;
	assign gfpga_pad_GPIO_PAD[77] = 1'b0;
	assign gfpga_pad_GPIO_PAD[78] = 1'b0;
	assign gfpga_pad_GPIO_PAD[79] = 1'b0;
	assign gfpga_pad_GPIO_PAD[80] = 1'b0;
	assign gfpga_pad_GPIO_PAD[81] = 1'b0;
	assign gfpga_pad_GPIO_PAD[82] = 1'b0;
	assign gfpga_pad_GPIO_PAD[83] = 1'b0;
	assign gfpga_pad_GPIO_PAD[84] = 1'b0;
	assign gfpga_pad_GPIO_PAD[85] = 1'b0;
	assign gfpga_pad_GPIO_PAD[86] = 1'b0;
	assign gfpga_pad_GPIO_PAD[87] = 1'b0;
	assign gfpga_pad_GPIO_PAD[88] = 1'b0;
	assign gfpga_pad_GPIO_PAD[89] = 1'b0;
	assign gfpga_pad_GPIO_PAD[90] = 1'b0;
	assign gfpga_pad_GPIO_PAD[91] = 1'b0;
	assign gfpga_pad_GPIO_PAD[92] = 1'b0;
	assign gfpga_pad_GPIO_PAD[93] = 1'b0;
	assign gfpga_pad_GPIO_PAD[94] = 1'b0;
	assign gfpga_pad_GPIO_PAD[95] = 1'b0;

`ifdef AUTOCHECKED_SIMULATION
// ----- Reference Benchmark Instanication -------
	and2 REF_DUT(
		.a(a),
		.b(b),
		.c(out_c_benchmark)	);
// ----- End reference Benchmark Instanication -------

`endif


// ----- Task: assign address and data values at rising edge of enable signal -----
task prog_cycle_task;
input [0:15] address_val;
input [0:0] data_in_val;
	begin
		@(negedge prog_clock[0]);
			address[0:15] = address_val[0:15];

			data_in[0] = data_in_val[0];

	end
endtask

// ----- Begin bitstream loading during configuration phase -----
initial
	begin
// ----- Address port default input -----
		address[0:15] = {16{1'b0}};
// ----- Data-input port default input -----
		data_in[0] = 1'b0;
		prog_cycle_task(16'b0000000000000000, 1'b1);
		prog_cycle_task(16'b0100000000000000, 1'b1);
		prog_cycle_task(16'b0010000000000000, 1'b1);
		prog_cycle_task(16'b0110000000000000, 1'b1);
		prog_cycle_task(16'b0001000000000000, 1'b1);
		prog_cycle_task(16'b0101000000000000, 1'b1);
		prog_cycle_task(16'b0011000000000000, 1'b0);
		prog_cycle_task(16'b0111000000000000, 1'b1);
		prog_cycle_task(16'b0000000000100000, 1'b1);
		prog_cycle_task(16'b0100000000100000, 1'b1);
		prog_cycle_task(16'b0010000000100000, 1'b1);
		prog_cycle_task(16'b0110000000100000, 1'b1);
		prog_cycle_task(16'b0001000000100000, 1'b1);
		prog_cycle_task(16'b0101000000100000, 1'b1);
		prog_cycle_task(16'b0011000000100000, 1'b1);
		prog_cycle_task(16'b0111000000100000, 1'b1);
		prog_cycle_task(16'b0000000000010000, 1'b1);
		prog_cycle_task(16'b0100000000010000, 1'b1);
		prog_cycle_task(16'b0010000000010000, 1'b1);
		prog_cycle_task(16'b0110000000010000, 1'b1);
		prog_cycle_task(16'b0001000000010000, 1'b1);
		prog_cycle_task(16'b0101000000010000, 1'b1);
		prog_cycle_task(16'b0011000000010000, 1'b1);
		prog_cycle_task(16'b0111000000010000, 1'b1);
		prog_cycle_task(16'b0000000000110000, 1'b1);
		prog_cycle_task(16'b0100000000110000, 1'b1);
		prog_cycle_task(16'b0010000000110000, 1'b1);
		prog_cycle_task(16'b0110000000110000, 1'b1);
		prog_cycle_task(16'b0001000000110000, 1'b1);
		prog_cycle_task(16'b0101000000110000, 1'b1);
		prog_cycle_task(16'b0011000000110000, 1'b1);
		prog_cycle_task(16'b0111000000110000, 1'b1);
		prog_cycle_task(16'b0000000000001000, 1'b1);
		prog_cycle_task(16'b0100000000001000, 1'b1);
		prog_cycle_task(16'b0010000000001000, 1'b1);
		prog_cycle_task(16'b0110000000001000, 1'b1);
		prog_cycle_task(16'b0001000000001000, 1'b1);
		prog_cycle_task(16'b0101000000001000, 1'b1);
		prog_cycle_task(16'b0011000000001000, 1'b1);
		prog_cycle_task(16'b0111000000001000, 1'b1);
		prog_cycle_task(16'b0000000000101000, 1'b1);
		prog_cycle_task(16'b0100000000101000, 1'b1);
		prog_cycle_task(16'b0010000000101000, 1'b1);
		prog_cycle_task(16'b0110000000101000, 1'b1);
		prog_cycle_task(16'b0001000000101000, 1'b1);
		prog_cycle_task(16'b0101000000101000, 1'b1);
		prog_cycle_task(16'b0011000000101000, 1'b1);
		prog_cycle_task(16'b0111000000101000, 1'b1);
		prog_cycle_task(16'b0000000000011000, 1'b0);
		prog_cycle_task(16'b1000000000011000, 1'b0);
		prog_cycle_task(16'b0100000000011000, 1'b0);
		prog_cycle_task(16'b1100000000011000, 1'b0);
		prog_cycle_task(16'b0010000000011000, 1'b0);
		prog_cycle_task(16'b1010000000011000, 1'b0);
		prog_cycle_task(16'b0110000000011000, 1'b0);
		prog_cycle_task(16'b1110000000011000, 1'b0);
		prog_cycle_task(16'b0001000000011000, 1'b0);
		prog_cycle_task(16'b1001000000011000, 1'b0);
		prog_cycle_task(16'b0101000000011000, 1'b0);
		prog_cycle_task(16'b1101000000011000, 1'b0);
		prog_cycle_task(16'b0011000000011000, 1'b0);
		prog_cycle_task(16'b1011000000011000, 1'b0);
		prog_cycle_task(16'b0111000000011000, 1'b0);
		prog_cycle_task(16'b1111000000011000, 1'b0);
		prog_cycle_task(16'b0000100000011000, 1'b0);
		prog_cycle_task(16'b1000100000011000, 1'b0);
		prog_cycle_task(16'b0100100000011000, 1'b0);
		prog_cycle_task(16'b1100100000011000, 1'b0);
		prog_cycle_task(16'b0010100000011000, 1'b0);
		prog_cycle_task(16'b1010100000011000, 1'b0);
		prog_cycle_task(16'b0110100000011000, 1'b0);
		prog_cycle_task(16'b1110100000011000, 1'b0);
		prog_cycle_task(16'b0001100000011000, 1'b0);
		prog_cycle_task(16'b1001100000011000, 1'b0);
		prog_cycle_task(16'b0101100000011000, 1'b0);
		prog_cycle_task(16'b1101100000011000, 1'b0);
		prog_cycle_task(16'b0011100000011000, 1'b0);
		prog_cycle_task(16'b1011100000011000, 1'b0);
		prog_cycle_task(16'b0111100000011000, 1'b0);
		prog_cycle_task(16'b1111100000011000, 1'b0);
		prog_cycle_task(16'b0000010000011000, 1'b0);
		prog_cycle_task(16'b1000010000011000, 1'b0);
		prog_cycle_task(16'b0100010000011000, 1'b0);
		prog_cycle_task(16'b1100010000011000, 1'b0);
		prog_cycle_task(16'b0000000000111000, 1'b0);
		prog_cycle_task(16'b1000000000111000, 1'b0);
		prog_cycle_task(16'b0100000000111000, 1'b0);
		prog_cycle_task(16'b1100000000111000, 1'b0);
		prog_cycle_task(16'b0010000000111000, 1'b0);
		prog_cycle_task(16'b1010000000111000, 1'b1);
		prog_cycle_task(16'b0001000000111000, 1'b0);
		prog_cycle_task(16'b1001000000111000, 1'b0);
		prog_cycle_task(16'b0101000000111000, 1'b0);
		prog_cycle_task(16'b1101000000111000, 1'b0);
		prog_cycle_task(16'b0011000000111000, 1'b0);
		prog_cycle_task(16'b1011000000111000, 1'b1);
		prog_cycle_task(16'b0000100000111000, 1'b0);
		prog_cycle_task(16'b1000100000111000, 1'b0);
		prog_cycle_task(16'b0100100000111000, 1'b0);
		prog_cycle_task(16'b1100100000111000, 1'b0);
		prog_cycle_task(16'b0010100000111000, 1'b0);
		prog_cycle_task(16'b1010100000111000, 1'b1);
		prog_cycle_task(16'b0001100000111000, 1'b0);
		prog_cycle_task(16'b1001100000111000, 1'b0);
		prog_cycle_task(16'b0101100000111000, 1'b0);
		prog_cycle_task(16'b1101100000111000, 1'b0);
		prog_cycle_task(16'b0011100000111000, 1'b0);
		prog_cycle_task(16'b1011100000111000, 1'b1);
		prog_cycle_task(16'b0000010000111000, 1'b0);
		prog_cycle_task(16'b1000010000111000, 1'b0);
		prog_cycle_task(16'b0100010000111000, 1'b0);
		prog_cycle_task(16'b1100010000111000, 1'b0);
		prog_cycle_task(16'b0010010000111000, 1'b0);
		prog_cycle_task(16'b1010010000111000, 1'b1);
		prog_cycle_task(16'b0001010000111000, 1'b0);
		prog_cycle_task(16'b1001010000111000, 1'b0);
		prog_cycle_task(16'b0101010000111000, 1'b0);
		prog_cycle_task(16'b1101010000111000, 1'b0);
		prog_cycle_task(16'b0011010000111000, 1'b0);
		prog_cycle_task(16'b1011010000111000, 1'b1);
		prog_cycle_task(16'b0000110000111000, 1'b0);
		prog_cycle_task(16'b1000110000111000, 1'b0);
		prog_cycle_task(16'b0100110000111000, 1'b0);
		prog_cycle_task(16'b1100110000111000, 1'b0);
		prog_cycle_task(16'b0010110000111000, 1'b0);
		prog_cycle_task(16'b1010110000111000, 1'b1);
		prog_cycle_task(16'b0001110000111000, 1'b0);
		prog_cycle_task(16'b1001110000111000, 1'b0);
		prog_cycle_task(16'b0101110000111000, 1'b0);
		prog_cycle_task(16'b1101110000111000, 1'b0);
		prog_cycle_task(16'b0011110000111000, 1'b0);
		prog_cycle_task(16'b1011110000111000, 1'b1);
		prog_cycle_task(16'b0000001000111000, 1'b0);
		prog_cycle_task(16'b1000001000111000, 1'b0);
		prog_cycle_task(16'b0100001000111000, 1'b0);
		prog_cycle_task(16'b1100001000111000, 1'b0);
		prog_cycle_task(16'b0010001000111000, 1'b0);
		prog_cycle_task(16'b1010001000111000, 1'b1);
		prog_cycle_task(16'b0001001000111000, 1'b0);
		prog_cycle_task(16'b1001001000111000, 1'b0);
		prog_cycle_task(16'b0000101000111000, 1'b0);
		prog_cycle_task(16'b1000101000111000, 1'b0);
		prog_cycle_task(16'b0000000000000100, 1'b1);
		prog_cycle_task(16'b0100000000000100, 1'b1);
		prog_cycle_task(16'b0010000000000100, 1'b1);
		prog_cycle_task(16'b0110000000000100, 1'b1);
		prog_cycle_task(16'b0001000000000100, 1'b1);
		prog_cycle_task(16'b0101000000000100, 1'b1);
		prog_cycle_task(16'b0011000000000100, 1'b1);
		prog_cycle_task(16'b0111000000000100, 1'b1);
		prog_cycle_task(16'b0000000000100100, 1'b0);
		prog_cycle_task(16'b1000000000100100, 1'b0);
		prog_cycle_task(16'b0100000000100100, 1'b1);
		prog_cycle_task(16'b1100000000100100, 1'b0);
		prog_cycle_task(16'b0010000000100100, 1'b0);
		prog_cycle_task(16'b1010000000100100, 1'b1);
		prog_cycle_task(16'b0001000000100100, 1'b0);
		prog_cycle_task(16'b1001000000100100, 1'b0);
		prog_cycle_task(16'b0101000000100100, 1'b1);
		prog_cycle_task(16'b1101000000100100, 1'b0);
		prog_cycle_task(16'b0011000000100100, 1'b0);
		prog_cycle_task(16'b1011000000100100, 1'b1);
		prog_cycle_task(16'b0000100000100100, 1'b0);
		prog_cycle_task(16'b1000100000100100, 1'b0);
		prog_cycle_task(16'b0100100000100100, 1'b1);
		prog_cycle_task(16'b1100100000100100, 1'b0);
		prog_cycle_task(16'b0010100000100100, 1'b0);
		prog_cycle_task(16'b1010100000100100, 1'b1);
		prog_cycle_task(16'b0001100000100100, 1'b0);
		prog_cycle_task(16'b1001100000100100, 1'b0);
		prog_cycle_task(16'b0000010000100100, 1'b0);
		prog_cycle_task(16'b1000010000100100, 1'b0);
		prog_cycle_task(16'b0001010000100100, 1'b0);
		prog_cycle_task(16'b1001010000100100, 1'b0);
		prog_cycle_task(16'b0000110000100100, 1'b0);
		prog_cycle_task(16'b1000110000100100, 1'b0);
		prog_cycle_task(16'b0001110000100100, 1'b0);
		prog_cycle_task(16'b1001110000100100, 1'b0);
		prog_cycle_task(16'b0000001000100100, 1'b0);
		prog_cycle_task(16'b1000001000100100, 1'b0);
		prog_cycle_task(16'b0001001000100100, 1'b0);
		prog_cycle_task(16'b1001001000100100, 1'b0);
		prog_cycle_task(16'b0000101000100100, 1'b0);
		prog_cycle_task(16'b1000101000100100, 1'b0);
		prog_cycle_task(16'b0001101000100100, 1'b0);
		prog_cycle_task(16'b1001101000100100, 1'b0);
		prog_cycle_task(16'b0000011000100100, 1'b0);
		prog_cycle_task(16'b1000011000100100, 1'b0);
		prog_cycle_task(16'b0100011000100100, 1'b1);
		prog_cycle_task(16'b1100011000100100, 1'b0);
		prog_cycle_task(16'b0010011000100100, 1'b0);
		prog_cycle_task(16'b1010011000100100, 1'b1);
		prog_cycle_task(16'b0001011000100100, 1'b0);
		prog_cycle_task(16'b1001011000100100, 1'b0);
		prog_cycle_task(16'b0101011000100100, 1'b1);
		prog_cycle_task(16'b1101011000100100, 1'b0);
		prog_cycle_task(16'b0011011000100100, 1'b0);
		prog_cycle_task(16'b1011011000100100, 1'b1);
		prog_cycle_task(16'b0000111000100100, 1'b0);
		prog_cycle_task(16'b1000111000100100, 1'b0);
		prog_cycle_task(16'b0100111000100100, 1'b1);
		prog_cycle_task(16'b1100111000100100, 1'b0);
		prog_cycle_task(16'b0010111000100100, 1'b0);
		prog_cycle_task(16'b1010111000100100, 1'b1);
		prog_cycle_task(16'b0000000000010100, 1'b0);
		prog_cycle_task(16'b1000000000010100, 1'b0);
		prog_cycle_task(16'b0100000000010100, 1'b0);
		prog_cycle_task(16'b1100000000010100, 1'b0);
		prog_cycle_task(16'b0010000000010100, 1'b0);
		prog_cycle_task(16'b1010000000010100, 1'b1);
		prog_cycle_task(16'b0001000000010100, 1'b0);
		prog_cycle_task(16'b1001000000010100, 1'b0);
		prog_cycle_task(16'b0101000000010100, 1'b0);
		prog_cycle_task(16'b1101000000010100, 1'b0);
		prog_cycle_task(16'b0011000000010100, 1'b0);
		prog_cycle_task(16'b1011000000010100, 1'b1);
		prog_cycle_task(16'b0000100000010100, 1'b0);
		prog_cycle_task(16'b1000100000010100, 1'b0);
		prog_cycle_task(16'b0100100000010100, 1'b0);
		prog_cycle_task(16'b1100100000010100, 1'b0);
		prog_cycle_task(16'b0010100000010100, 1'b0);
		prog_cycle_task(16'b1010100000010100, 1'b1);
		prog_cycle_task(16'b0001100000010100, 1'b0);
		prog_cycle_task(16'b1001100000010100, 1'b0);
		prog_cycle_task(16'b0101100000010100, 1'b0);
		prog_cycle_task(16'b1101100000010100, 1'b0);
		prog_cycle_task(16'b0011100000010100, 1'b0);
		prog_cycle_task(16'b1011100000010100, 1'b1);
		prog_cycle_task(16'b0000010000010100, 1'b0);
		prog_cycle_task(16'b1000010000010100, 1'b0);
		prog_cycle_task(16'b0100010000010100, 1'b0);
		prog_cycle_task(16'b1100010000010100, 1'b0);
		prog_cycle_task(16'b0010010000010100, 1'b0);
		prog_cycle_task(16'b1010010000010100, 1'b1);
		prog_cycle_task(16'b0001010000010100, 1'b0);
		prog_cycle_task(16'b1001010000010100, 1'b0);
		prog_cycle_task(16'b0101010000010100, 1'b0);
		prog_cycle_task(16'b1101010000010100, 1'b0);
		prog_cycle_task(16'b0011010000010100, 1'b0);
		prog_cycle_task(16'b1011010000010100, 1'b1);
		prog_cycle_task(16'b0000110000010100, 1'b0);
		prog_cycle_task(16'b1000110000010100, 1'b0);
		prog_cycle_task(16'b0100110000010100, 1'b0);
		prog_cycle_task(16'b1100110000010100, 1'b0);
		prog_cycle_task(16'b0010110000010100, 1'b0);
		prog_cycle_task(16'b1010110000010100, 1'b1);
		prog_cycle_task(16'b0001110000010100, 1'b0);
		prog_cycle_task(16'b1001110000010100, 1'b0);
		prog_cycle_task(16'b0101110000010100, 1'b0);
		prog_cycle_task(16'b1101110000010100, 1'b0);
		prog_cycle_task(16'b0011110000010100, 1'b0);
		prog_cycle_task(16'b1011110000010100, 1'b1);
		prog_cycle_task(16'b0000001000010100, 1'b0);
		prog_cycle_task(16'b1000001000010100, 1'b0);
		prog_cycle_task(16'b0100001000010100, 1'b0);
		prog_cycle_task(16'b1100001000010100, 1'b0);
		prog_cycle_task(16'b0010001000010100, 1'b0);
		prog_cycle_task(16'b1010001000010100, 1'b1);
		prog_cycle_task(16'b0001001000010100, 1'b0);
		prog_cycle_task(16'b1001001000010100, 1'b0);
		prog_cycle_task(16'b0000101000010100, 1'b0);
		prog_cycle_task(16'b1000101000010100, 1'b0);
		prog_cycle_task(16'b0000000000110100, 1'b1);
		prog_cycle_task(16'b0100000000110100, 1'b1);
		prog_cycle_task(16'b0010000000110100, 1'b1);
		prog_cycle_task(16'b0110000000110100, 1'b1);
		prog_cycle_task(16'b0001000000110100, 1'b1);
		prog_cycle_task(16'b0101000000110100, 1'b1);
		prog_cycle_task(16'b0011000000110100, 1'b1);
		prog_cycle_task(16'b0111000000110100, 1'b1);
		prog_cycle_task(16'b0000000000001100, 1'b0);
		prog_cycle_task(16'b1000000000001100, 1'b0);
		prog_cycle_task(16'b0100000000001100, 1'b1);
		prog_cycle_task(16'b1100000000001100, 1'b0);
		prog_cycle_task(16'b0010000000001100, 1'b0);
		prog_cycle_task(16'b1010000000001100, 1'b1);
		prog_cycle_task(16'b0001000000001100, 1'b0);
		prog_cycle_task(16'b1001000000001100, 1'b0);
		prog_cycle_task(16'b0101000000001100, 1'b1);
		prog_cycle_task(16'b1101000000001100, 1'b0);
		prog_cycle_task(16'b0011000000001100, 1'b0);
		prog_cycle_task(16'b1011000000001100, 1'b1);
		prog_cycle_task(16'b0000100000001100, 1'b0);
		prog_cycle_task(16'b1000100000001100, 1'b0);
		prog_cycle_task(16'b0100100000001100, 1'b1);
		prog_cycle_task(16'b1100100000001100, 1'b0);
		prog_cycle_task(16'b0010100000001100, 1'b0);
		prog_cycle_task(16'b1010100000001100, 1'b1);
		prog_cycle_task(16'b0001100000001100, 1'b0);
		prog_cycle_task(16'b1001100000001100, 1'b0);
		prog_cycle_task(16'b0000010000001100, 1'b0);
		prog_cycle_task(16'b1000010000001100, 1'b0);
		prog_cycle_task(16'b0001010000001100, 1'b0);
		prog_cycle_task(16'b1001010000001100, 1'b0);
		prog_cycle_task(16'b0000110000001100, 1'b0);
		prog_cycle_task(16'b1000110000001100, 1'b0);
		prog_cycle_task(16'b0001110000001100, 1'b0);
		prog_cycle_task(16'b1001110000001100, 1'b0);
		prog_cycle_task(16'b0000001000001100, 1'b0);
		prog_cycle_task(16'b1000001000001100, 1'b0);
		prog_cycle_task(16'b0001001000001100, 1'b0);
		prog_cycle_task(16'b1001001000001100, 1'b0);
		prog_cycle_task(16'b0000101000001100, 1'b0);
		prog_cycle_task(16'b1000101000001100, 1'b0);
		prog_cycle_task(16'b0001101000001100, 1'b0);
		prog_cycle_task(16'b1001101000001100, 1'b0);
		prog_cycle_task(16'b0000011000001100, 1'b0);
		prog_cycle_task(16'b1000011000001100, 1'b0);
		prog_cycle_task(16'b0100011000001100, 1'b1);
		prog_cycle_task(16'b1100011000001100, 1'b0);
		prog_cycle_task(16'b0010011000001100, 1'b0);
		prog_cycle_task(16'b1010011000001100, 1'b1);
		prog_cycle_task(16'b0001011000001100, 1'b0);
		prog_cycle_task(16'b1001011000001100, 1'b0);
		prog_cycle_task(16'b0101011000001100, 1'b1);
		prog_cycle_task(16'b1101011000001100, 1'b0);
		prog_cycle_task(16'b0011011000001100, 1'b0);
		prog_cycle_task(16'b1011011000001100, 1'b1);
		prog_cycle_task(16'b0000111000001100, 1'b0);
		prog_cycle_task(16'b1000111000001100, 1'b0);
		prog_cycle_task(16'b0100111000001100, 1'b1);
		prog_cycle_task(16'b1100111000001100, 1'b0);
		prog_cycle_task(16'b0010111000001100, 1'b0);
		prog_cycle_task(16'b1010111000001100, 1'b1);
		prog_cycle_task(16'b0000000000101100, 1'b0);
		prog_cycle_task(16'b1000000000101100, 1'b0);
		prog_cycle_task(16'b0100000000101100, 1'b0);
		prog_cycle_task(16'b1100000000101100, 1'b0);
		prog_cycle_task(16'b0010000000101100, 1'b0);
		prog_cycle_task(16'b1010000000101100, 1'b1);
		prog_cycle_task(16'b0001000000101100, 1'b0);
		prog_cycle_task(16'b1001000000101100, 1'b0);
		prog_cycle_task(16'b0101000000101100, 1'b0);
		prog_cycle_task(16'b1101000000101100, 1'b0);
		prog_cycle_task(16'b0011000000101100, 1'b0);
		prog_cycle_task(16'b1011000000101100, 1'b1);
		prog_cycle_task(16'b0000100000101100, 1'b0);
		prog_cycle_task(16'b1000100000101100, 1'b0);
		prog_cycle_task(16'b0100100000101100, 1'b0);
		prog_cycle_task(16'b1100100000101100, 1'b0);
		prog_cycle_task(16'b0010100000101100, 1'b0);
		prog_cycle_task(16'b1010100000101100, 1'b1);
		prog_cycle_task(16'b0001100000101100, 1'b0);
		prog_cycle_task(16'b1001100000101100, 1'b0);
		prog_cycle_task(16'b0101100000101100, 1'b0);
		prog_cycle_task(16'b1101100000101100, 1'b0);
		prog_cycle_task(16'b0011100000101100, 1'b0);
		prog_cycle_task(16'b1011100000101100, 1'b1);
		prog_cycle_task(16'b0000010000101100, 1'b0);
		prog_cycle_task(16'b1000010000101100, 1'b0);
		prog_cycle_task(16'b0100010000101100, 1'b0);
		prog_cycle_task(16'b1100010000101100, 1'b0);
		prog_cycle_task(16'b0010010000101100, 1'b0);
		prog_cycle_task(16'b1010010000101100, 1'b1);
		prog_cycle_task(16'b0001010000101100, 1'b0);
		prog_cycle_task(16'b1001010000101100, 1'b0);
		prog_cycle_task(16'b0101010000101100, 1'b0);
		prog_cycle_task(16'b1101010000101100, 1'b0);
		prog_cycle_task(16'b0011010000101100, 1'b0);
		prog_cycle_task(16'b1011010000101100, 1'b1);
		prog_cycle_task(16'b0000110000101100, 1'b0);
		prog_cycle_task(16'b1000110000101100, 1'b0);
		prog_cycle_task(16'b0100110000101100, 1'b0);
		prog_cycle_task(16'b1100110000101100, 1'b0);
		prog_cycle_task(16'b0010110000101100, 1'b0);
		prog_cycle_task(16'b1010110000101100, 1'b1);
		prog_cycle_task(16'b0001110000101100, 1'b0);
		prog_cycle_task(16'b1001110000101100, 1'b0);
		prog_cycle_task(16'b0101110000101100, 1'b0);
		prog_cycle_task(16'b1101110000101100, 1'b0);
		prog_cycle_task(16'b0011110000101100, 1'b0);
		prog_cycle_task(16'b1011110000101100, 1'b1);
		prog_cycle_task(16'b0000001000101100, 1'b0);
		prog_cycle_task(16'b1000001000101100, 1'b0);
		prog_cycle_task(16'b0100001000101100, 1'b0);
		prog_cycle_task(16'b1100001000101100, 1'b0);
		prog_cycle_task(16'b0010001000101100, 1'b0);
		prog_cycle_task(16'b1010001000101100, 1'b1);
		prog_cycle_task(16'b0001001000101100, 1'b0);
		prog_cycle_task(16'b1001001000101100, 1'b0);
		prog_cycle_task(16'b0000101000101100, 1'b0);
		prog_cycle_task(16'b1000101000101100, 1'b0);
		prog_cycle_task(16'b0000000000011100, 1'b1);
		prog_cycle_task(16'b0100000000011100, 1'b1);
		prog_cycle_task(16'b0010000000011100, 1'b1);
		prog_cycle_task(16'b0110000000011100, 1'b1);
		prog_cycle_task(16'b0001000000011100, 1'b1);
		prog_cycle_task(16'b0101000000011100, 1'b1);
		prog_cycle_task(16'b0011000000011100, 1'b1);
		prog_cycle_task(16'b0111000000011100, 1'b1);
		prog_cycle_task(16'b0000000000111100, 1'b0);
		prog_cycle_task(16'b1000000000111100, 1'b0);
		prog_cycle_task(16'b0100000000111100, 1'b0);
		prog_cycle_task(16'b1100000000111100, 1'b0);
		prog_cycle_task(16'b0010000000111100, 1'b0);
		prog_cycle_task(16'b1010000000111100, 1'b0);
		prog_cycle_task(16'b0110000000111100, 1'b0);
		prog_cycle_task(16'b1110000000111100, 1'b0);
		prog_cycle_task(16'b0001000000111100, 1'b0);
		prog_cycle_task(16'b1001000000111100, 1'b0);
		prog_cycle_task(16'b0101000000111100, 1'b0);
		prog_cycle_task(16'b1101000000111100, 1'b0);
		prog_cycle_task(16'b0011000000111100, 1'b0);
		prog_cycle_task(16'b1011000000111100, 1'b0);
		prog_cycle_task(16'b0111000000111100, 1'b0);
		prog_cycle_task(16'b1111000000111100, 1'b0);
		prog_cycle_task(16'b0000100000111100, 1'b0);
		prog_cycle_task(16'b1000100000111100, 1'b0);
		prog_cycle_task(16'b0100100000111100, 1'b0);
		prog_cycle_task(16'b1100100000111100, 1'b0);
		prog_cycle_task(16'b0010100000111100, 1'b0);
		prog_cycle_task(16'b1010100000111100, 1'b0);
		prog_cycle_task(16'b0110100000111100, 1'b0);
		prog_cycle_task(16'b1110100000111100, 1'b0);
		prog_cycle_task(16'b0001100000111100, 1'b0);
		prog_cycle_task(16'b1001100000111100, 1'b0);
		prog_cycle_task(16'b0101100000111100, 1'b0);
		prog_cycle_task(16'b1101100000111100, 1'b0);
		prog_cycle_task(16'b0011100000111100, 1'b0);
		prog_cycle_task(16'b1011100000111100, 1'b0);
		prog_cycle_task(16'b0111100000111100, 1'b0);
		prog_cycle_task(16'b1111100000111100, 1'b0);
		prog_cycle_task(16'b0000010000111100, 1'b0);
		prog_cycle_task(16'b1000010000111100, 1'b0);
		prog_cycle_task(16'b0100010000111100, 1'b0);
		prog_cycle_task(16'b1100010000111100, 1'b0);
		prog_cycle_task(16'b0000000000000010, 1'b0);
		prog_cycle_task(16'b1000000000000010, 1'b0);
		prog_cycle_task(16'b0100000000000010, 1'b1);
		prog_cycle_task(16'b1100000000000010, 1'b0);
		prog_cycle_task(16'b0010000000000010, 1'b0);
		prog_cycle_task(16'b1010000000000010, 1'b1);
		prog_cycle_task(16'b0001000000000010, 1'b0);
		prog_cycle_task(16'b1001000000000010, 1'b0);
		prog_cycle_task(16'b0101000000000010, 1'b1);
		prog_cycle_task(16'b1101000000000010, 1'b0);
		prog_cycle_task(16'b0011000000000010, 1'b0);
		prog_cycle_task(16'b1011000000000010, 1'b1);
		prog_cycle_task(16'b0000100000000010, 1'b0);
		prog_cycle_task(16'b1000100000000010, 1'b0);
		prog_cycle_task(16'b0100100000000010, 1'b1);
		prog_cycle_task(16'b1100100000000010, 1'b0);
		prog_cycle_task(16'b0010100000000010, 1'b0);
		prog_cycle_task(16'b1010100000000010, 1'b1);
		prog_cycle_task(16'b0001100000000010, 1'b0);
		prog_cycle_task(16'b1001100000000010, 1'b0);
		prog_cycle_task(16'b0000010000000010, 1'b0);
		prog_cycle_task(16'b1000010000000010, 1'b0);
		prog_cycle_task(16'b0001010000000010, 1'b0);
		prog_cycle_task(16'b1001010000000010, 1'b0);
		prog_cycle_task(16'b0000110000000010, 1'b0);
		prog_cycle_task(16'b1000110000000010, 1'b0);
		prog_cycle_task(16'b0001110000000010, 1'b0);
		prog_cycle_task(16'b1001110000000010, 1'b0);
		prog_cycle_task(16'b0000001000000010, 1'b0);
		prog_cycle_task(16'b1000001000000010, 1'b0);
		prog_cycle_task(16'b0001001000000010, 1'b0);
		prog_cycle_task(16'b1001001000000010, 1'b0);
		prog_cycle_task(16'b0000101000000010, 1'b0);
		prog_cycle_task(16'b1000101000000010, 1'b0);
		prog_cycle_task(16'b0100101000000010, 1'b1);
		prog_cycle_task(16'b1100101000000010, 1'b0);
		prog_cycle_task(16'b0010101000000010, 1'b0);
		prog_cycle_task(16'b1010101000000010, 1'b1);
		prog_cycle_task(16'b0001101000000010, 1'b0);
		prog_cycle_task(16'b1001101000000010, 1'b0);
		prog_cycle_task(16'b0101101000000010, 1'b1);
		prog_cycle_task(16'b1101101000000010, 1'b0);
		prog_cycle_task(16'b0011101000000010, 1'b0);
		prog_cycle_task(16'b1011101000000010, 1'b1);
		prog_cycle_task(16'b0000011000000010, 1'b0);
		prog_cycle_task(16'b1000011000000010, 1'b0);
		prog_cycle_task(16'b0100011000000010, 1'b1);
		prog_cycle_task(16'b1100011000000010, 1'b0);
		prog_cycle_task(16'b0010011000000010, 1'b0);
		prog_cycle_task(16'b1010011000000010, 1'b1);
		prog_cycle_task(16'b0000000000100010, 1'b0);
		prog_cycle_task(16'b1000000000100010, 1'b0);
		prog_cycle_task(16'b0100000000100010, 1'b0);
		prog_cycle_task(16'b1100000000100010, 1'b0);
		prog_cycle_task(16'b0010000000100010, 1'b0);
		prog_cycle_task(16'b1010000000100010, 1'b1);
		prog_cycle_task(16'b0001000000100010, 1'b0);
		prog_cycle_task(16'b1001000000100010, 1'b0);
		prog_cycle_task(16'b0000100000100010, 1'b0);
		prog_cycle_task(16'b1000100000100010, 1'b0);
		prog_cycle_task(16'b0100100000100010, 1'b0);
		prog_cycle_task(16'b1100100000100010, 1'b0);
		prog_cycle_task(16'b0010100000100010, 1'b0);
		prog_cycle_task(16'b1010100000100010, 1'b1);
		prog_cycle_task(16'b0001100000100010, 1'b0);
		prog_cycle_task(16'b1001100000100010, 1'b0);
		prog_cycle_task(16'b0101100000100010, 1'b0);
		prog_cycle_task(16'b1101100000100010, 1'b0);
		prog_cycle_task(16'b0011100000100010, 1'b0);
		prog_cycle_task(16'b1011100000100010, 1'b1);
		prog_cycle_task(16'b0000010000100010, 1'b0);
		prog_cycle_task(16'b1000010000100010, 1'b0);
		prog_cycle_task(16'b0100010000100010, 1'b0);
		prog_cycle_task(16'b1100010000100010, 1'b0);
		prog_cycle_task(16'b0010010000100010, 1'b0);
		prog_cycle_task(16'b1010010000100010, 1'b1);
		prog_cycle_task(16'b0001010000100010, 1'b0);
		prog_cycle_task(16'b1001010000100010, 1'b0);
		prog_cycle_task(16'b0101010000100010, 1'b0);
		prog_cycle_task(16'b1101010000100010, 1'b0);
		prog_cycle_task(16'b0011010000100010, 1'b0);
		prog_cycle_task(16'b1011010000100010, 1'b1);
		prog_cycle_task(16'b0000110000100010, 1'b0);
		prog_cycle_task(16'b1000110000100010, 1'b0);
		prog_cycle_task(16'b0100110000100010, 1'b0);
		prog_cycle_task(16'b1100110000100010, 1'b0);
		prog_cycle_task(16'b0010110000100010, 1'b0);
		prog_cycle_task(16'b1010110000100010, 1'b1);
		prog_cycle_task(16'b0001110000100010, 1'b0);
		prog_cycle_task(16'b1001110000100010, 1'b0);
		prog_cycle_task(16'b0101110000100010, 1'b0);
		prog_cycle_task(16'b1101110000100010, 1'b0);
		prog_cycle_task(16'b0011110000100010, 1'b0);
		prog_cycle_task(16'b1011110000100010, 1'b1);
		prog_cycle_task(16'b0000001000100010, 1'b0);
		prog_cycle_task(16'b1000001000100010, 1'b0);
		prog_cycle_task(16'b0100001000100010, 1'b0);
		prog_cycle_task(16'b1100001000100010, 1'b0);
		prog_cycle_task(16'b0010001000100010, 1'b0);
		prog_cycle_task(16'b1010001000100010, 1'b1);
		prog_cycle_task(16'b0001001000100010, 1'b0);
		prog_cycle_task(16'b1001001000100010, 1'b0);
		prog_cycle_task(16'b0101001000100010, 1'b0);
		prog_cycle_task(16'b1101001000100010, 1'b0);
		prog_cycle_task(16'b0011001000100010, 1'b0);
		prog_cycle_task(16'b1011001000100010, 1'b1);
		prog_cycle_task(16'b0000000000010010, 1'b1);
		prog_cycle_task(16'b0100000000010010, 1'b1);
		prog_cycle_task(16'b0010000000010010, 1'b1);
		prog_cycle_task(16'b0110000000010010, 1'b1);
		prog_cycle_task(16'b0001000000010010, 1'b1);
		prog_cycle_task(16'b0101000000010010, 1'b1);
		prog_cycle_task(16'b0011000000010010, 1'b1);
		prog_cycle_task(16'b0111000000010010, 1'b1);
		prog_cycle_task(16'b0000000000110010, 1'b0);
		prog_cycle_task(16'b1000000000110010, 1'b0);
		prog_cycle_task(16'b0100000000110010, 1'b1);
		prog_cycle_task(16'b1100000000110010, 1'b0);
		prog_cycle_task(16'b0010000000110010, 1'b0);
		prog_cycle_task(16'b1010000000110010, 1'b1);
		prog_cycle_task(16'b0001000000110010, 1'b0);
		prog_cycle_task(16'b1001000000110010, 1'b0);
		prog_cycle_task(16'b0101000000110010, 1'b1);
		prog_cycle_task(16'b1101000000110010, 1'b0);
		prog_cycle_task(16'b0011000000110010, 1'b0);
		prog_cycle_task(16'b1011000000110010, 1'b1);
		prog_cycle_task(16'b0000100000110010, 1'b0);
		prog_cycle_task(16'b1000100000110010, 1'b0);
		prog_cycle_task(16'b0100100000110010, 1'b1);
		prog_cycle_task(16'b1100100000110010, 1'b0);
		prog_cycle_task(16'b0010100000110010, 1'b0);
		prog_cycle_task(16'b1010100000110010, 1'b1);
		prog_cycle_task(16'b0001100000110010, 1'b0);
		prog_cycle_task(16'b1001100000110010, 1'b0);
		prog_cycle_task(16'b0000010000110010, 1'b0);
		prog_cycle_task(16'b1000010000110010, 1'b0);
		prog_cycle_task(16'b0001010000110010, 1'b0);
		prog_cycle_task(16'b1001010000110010, 1'b0);
		prog_cycle_task(16'b0000110000110010, 1'b0);
		prog_cycle_task(16'b1000110000110010, 1'b0);
		prog_cycle_task(16'b0001110000110010, 1'b0);
		prog_cycle_task(16'b1001110000110010, 1'b0);
		prog_cycle_task(16'b0000001000110010, 1'b0);
		prog_cycle_task(16'b1000001000110010, 1'b0);
		prog_cycle_task(16'b0001001000110010, 1'b0);
		prog_cycle_task(16'b1001001000110010, 1'b0);
		prog_cycle_task(16'b0000101000110010, 1'b0);
		prog_cycle_task(16'b1000101000110010, 1'b0);
		prog_cycle_task(16'b0100101000110010, 1'b1);
		prog_cycle_task(16'b1100101000110010, 1'b0);
		prog_cycle_task(16'b0010101000110010, 1'b0);
		prog_cycle_task(16'b1010101000110010, 1'b1);
		prog_cycle_task(16'b0001101000110010, 1'b0);
		prog_cycle_task(16'b1001101000110010, 1'b0);
		prog_cycle_task(16'b0101101000110010, 1'b1);
		prog_cycle_task(16'b1101101000110010, 1'b0);
		prog_cycle_task(16'b0011101000110010, 1'b0);
		prog_cycle_task(16'b1011101000110010, 1'b1);
		prog_cycle_task(16'b0000011000110010, 1'b0);
		prog_cycle_task(16'b1000011000110010, 1'b0);
		prog_cycle_task(16'b0100011000110010, 1'b1);
		prog_cycle_task(16'b1100011000110010, 1'b0);
		prog_cycle_task(16'b0010011000110010, 1'b0);
		prog_cycle_task(16'b1010011000110010, 1'b1);
		prog_cycle_task(16'b0000000000001010, 1'b0);
		prog_cycle_task(16'b1000000000001010, 1'b0);
		prog_cycle_task(16'b0100000000001010, 1'b0);
		prog_cycle_task(16'b1100000000001010, 1'b0);
		prog_cycle_task(16'b0010000000001010, 1'b0);
		prog_cycle_task(16'b1010000000001010, 1'b1);
		prog_cycle_task(16'b0001000000001010, 1'b0);
		prog_cycle_task(16'b1001000000001010, 1'b0);
		prog_cycle_task(16'b0000100000001010, 1'b0);
		prog_cycle_task(16'b1000100000001010, 1'b0);
		prog_cycle_task(16'b0100100000001010, 1'b0);
		prog_cycle_task(16'b1100100000001010, 1'b0);
		prog_cycle_task(16'b0010100000001010, 1'b0);
		prog_cycle_task(16'b1010100000001010, 1'b1);
		prog_cycle_task(16'b0001100000001010, 1'b0);
		prog_cycle_task(16'b1001100000001010, 1'b0);
		prog_cycle_task(16'b0101100000001010, 1'b0);
		prog_cycle_task(16'b1101100000001010, 1'b0);
		prog_cycle_task(16'b0011100000001010, 1'b0);
		prog_cycle_task(16'b1011100000001010, 1'b1);
		prog_cycle_task(16'b0000010000001010, 1'b0);
		prog_cycle_task(16'b1000010000001010, 1'b0);
		prog_cycle_task(16'b0100010000001010, 1'b0);
		prog_cycle_task(16'b1100010000001010, 1'b0);
		prog_cycle_task(16'b0010010000001010, 1'b0);
		prog_cycle_task(16'b1010010000001010, 1'b1);
		prog_cycle_task(16'b0001010000001010, 1'b0);
		prog_cycle_task(16'b1001010000001010, 1'b0);
		prog_cycle_task(16'b0101010000001010, 1'b0);
		prog_cycle_task(16'b1101010000001010, 1'b0);
		prog_cycle_task(16'b0011010000001010, 1'b0);
		prog_cycle_task(16'b1011010000001010, 1'b1);
		prog_cycle_task(16'b0000110000001010, 1'b0);
		prog_cycle_task(16'b1000110000001010, 1'b0);
		prog_cycle_task(16'b0100110000001010, 1'b0);
		prog_cycle_task(16'b1100110000001010, 1'b0);
		prog_cycle_task(16'b0010110000001010, 1'b0);
		prog_cycle_task(16'b1010110000001010, 1'b1);
		prog_cycle_task(16'b0001110000001010, 1'b0);
		prog_cycle_task(16'b1001110000001010, 1'b0);
		prog_cycle_task(16'b0101110000001010, 1'b0);
		prog_cycle_task(16'b1101110000001010, 1'b0);
		prog_cycle_task(16'b0011110000001010, 1'b0);
		prog_cycle_task(16'b1011110000001010, 1'b1);
		prog_cycle_task(16'b0000001000001010, 1'b0);
		prog_cycle_task(16'b1000001000001010, 1'b0);
		prog_cycle_task(16'b0100001000001010, 1'b0);
		prog_cycle_task(16'b1100001000001010, 1'b0);
		prog_cycle_task(16'b0010001000001010, 1'b0);
		prog_cycle_task(16'b1010001000001010, 1'b1);
		prog_cycle_task(16'b0001001000001010, 1'b0);
		prog_cycle_task(16'b1001001000001010, 1'b0);
		prog_cycle_task(16'b0101001000001010, 1'b0);
		prog_cycle_task(16'b1101001000001010, 1'b0);
		prog_cycle_task(16'b0011001000001010, 1'b0);
		prog_cycle_task(16'b1011001000001010, 1'b1);
		prog_cycle_task(16'b0000000000101010, 1'b1);
		prog_cycle_task(16'b0100000000101010, 1'b1);
		prog_cycle_task(16'b0010000000101010, 1'b1);
		prog_cycle_task(16'b0110000000101010, 1'b1);
		prog_cycle_task(16'b0001000000101010, 1'b1);
		prog_cycle_task(16'b0101000000101010, 1'b1);
		prog_cycle_task(16'b0011000000101010, 1'b1);
		prog_cycle_task(16'b0111000000101010, 1'b1);
		prog_cycle_task(16'b0000000000011010, 1'b0);
		prog_cycle_task(16'b1000000000011010, 1'b0);
		prog_cycle_task(16'b0100000000011010, 1'b0);
		prog_cycle_task(16'b1100000000011010, 1'b0);
		prog_cycle_task(16'b0010000000011010, 1'b0);
		prog_cycle_task(16'b1010000000011010, 1'b0);
		prog_cycle_task(16'b0110000000011010, 1'b0);
		prog_cycle_task(16'b1110000000011010, 1'b0);
		prog_cycle_task(16'b0001000000011010, 1'b0);
		prog_cycle_task(16'b1001000000011010, 1'b0);
		prog_cycle_task(16'b0101000000011010, 1'b0);
		prog_cycle_task(16'b1101000000011010, 1'b0);
		prog_cycle_task(16'b0011000000011010, 1'b0);
		prog_cycle_task(16'b1011000000011010, 1'b0);
		prog_cycle_task(16'b0111000000011010, 1'b0);
		prog_cycle_task(16'b1111000000011010, 1'b0);
		prog_cycle_task(16'b0000100000011010, 1'b0);
		prog_cycle_task(16'b1000100000011010, 1'b0);
		prog_cycle_task(16'b0100100000011010, 1'b0);
		prog_cycle_task(16'b1100100000011010, 1'b0);
		prog_cycle_task(16'b0010100000011010, 1'b0);
		prog_cycle_task(16'b1010100000011010, 1'b0);
		prog_cycle_task(16'b0110100000011010, 1'b0);
		prog_cycle_task(16'b1110100000011010, 1'b0);
		prog_cycle_task(16'b0001100000011010, 1'b0);
		prog_cycle_task(16'b1001100000011010, 1'b0);
		prog_cycle_task(16'b0101100000011010, 1'b0);
		prog_cycle_task(16'b1101100000011010, 1'b0);
		prog_cycle_task(16'b0011100000011010, 1'b0);
		prog_cycle_task(16'b1011100000011010, 1'b0);
		prog_cycle_task(16'b0111100000011010, 1'b0);
		prog_cycle_task(16'b1111100000011010, 1'b1);
		prog_cycle_task(16'b0000010000011010, 1'b0);
		prog_cycle_task(16'b1000010000011010, 1'b0);
		prog_cycle_task(16'b0100010000011010, 1'b0);
		prog_cycle_task(16'b1100010000011010, 1'b0);
		prog_cycle_task(16'b0000000000111010, 1'b0);
		prog_cycle_task(16'b1000000000111010, 1'b0);
		prog_cycle_task(16'b0100000000111010, 1'b0);
		prog_cycle_task(16'b1100000000111010, 1'b0);
		prog_cycle_task(16'b0010000000111010, 1'b0);
		prog_cycle_task(16'b1010000000111010, 1'b1);
		prog_cycle_task(16'b0001000000111010, 1'b0);
		prog_cycle_task(16'b1001000000111010, 1'b0);
		prog_cycle_task(16'b0000100000111010, 1'b0);
		prog_cycle_task(16'b1000100000111010, 1'b0);
		prog_cycle_task(16'b0100100000111010, 1'b0);
		prog_cycle_task(16'b1100100000111010, 1'b0);
		prog_cycle_task(16'b0010100000111010, 1'b0);
		prog_cycle_task(16'b1010100000111010, 1'b1);
		prog_cycle_task(16'b0001100000111010, 1'b0);
		prog_cycle_task(16'b1001100000111010, 1'b0);
		prog_cycle_task(16'b0101100000111010, 1'b0);
		prog_cycle_task(16'b1101100000111010, 1'b0);
		prog_cycle_task(16'b0011100000111010, 1'b0);
		prog_cycle_task(16'b1011100000111010, 1'b1);
		prog_cycle_task(16'b0000010000111010, 1'b0);
		prog_cycle_task(16'b1000010000111010, 1'b0);
		prog_cycle_task(16'b0100010000111010, 1'b0);
		prog_cycle_task(16'b1100010000111010, 1'b0);
		prog_cycle_task(16'b0010010000111010, 1'b0);
		prog_cycle_task(16'b1010010000111010, 1'b1);
		prog_cycle_task(16'b0001010000111010, 1'b0);
		prog_cycle_task(16'b1001010000111010, 1'b0);
		prog_cycle_task(16'b0101010000111010, 1'b0);
		prog_cycle_task(16'b1101010000111010, 1'b0);
		prog_cycle_task(16'b0011010000111010, 1'b0);
		prog_cycle_task(16'b1011010000111010, 1'b1);
		prog_cycle_task(16'b0000110000111010, 1'b0);
		prog_cycle_task(16'b1000110000111010, 1'b0);
		prog_cycle_task(16'b0100110000111010, 1'b0);
		prog_cycle_task(16'b1100110000111010, 1'b0);
		prog_cycle_task(16'b0010110000111010, 1'b0);
		prog_cycle_task(16'b1010110000111010, 1'b1);
		prog_cycle_task(16'b0001110000111010, 1'b0);
		prog_cycle_task(16'b1001110000111010, 1'b0);
		prog_cycle_task(16'b0101110000111010, 1'b0);
		prog_cycle_task(16'b1101110000111010, 1'b0);
		prog_cycle_task(16'b0011110000111010, 1'b0);
		prog_cycle_task(16'b1011110000111010, 1'b1);
		prog_cycle_task(16'b0000001000111010, 1'b0);
		prog_cycle_task(16'b1000001000111010, 1'b0);
		prog_cycle_task(16'b0100001000111010, 1'b0);
		prog_cycle_task(16'b1100001000111010, 1'b0);
		prog_cycle_task(16'b0010001000111010, 1'b0);
		prog_cycle_task(16'b1010001000111010, 1'b1);
		prog_cycle_task(16'b0001001000111010, 1'b0);
		prog_cycle_task(16'b1001001000111010, 1'b0);
		prog_cycle_task(16'b0101001000111010, 1'b0);
		prog_cycle_task(16'b1101001000111010, 1'b0);
		prog_cycle_task(16'b0011001000111010, 1'b0);
		prog_cycle_task(16'b1011001000111010, 1'b1);
		prog_cycle_task(16'b0000000000000110, 1'b1);
		prog_cycle_task(16'b0100000000000110, 1'b1);
		prog_cycle_task(16'b0010000000000110, 1'b1);
		prog_cycle_task(16'b0110000000000110, 1'b1);
		prog_cycle_task(16'b0001000000000110, 1'b1);
		prog_cycle_task(16'b0101000000000110, 1'b1);
		prog_cycle_task(16'b0011000000000110, 1'b1);
		prog_cycle_task(16'b0111000000000110, 1'b1);
		prog_cycle_task(16'b0000000000100110, 1'b0);
		prog_cycle_task(16'b1000000000100110, 1'b0);
		prog_cycle_task(16'b0100000000100110, 1'b0);
		prog_cycle_task(16'b1100000000100110, 1'b0);
		prog_cycle_task(16'b0010000000100110, 1'b0);
		prog_cycle_task(16'b1010000000100110, 1'b1);
		prog_cycle_task(16'b0001000000100110, 1'b0);
		prog_cycle_task(16'b1001000000100110, 1'b0);
		prog_cycle_task(16'b0000100000100110, 1'b0);
		prog_cycle_task(16'b1000100000100110, 1'b1);
		prog_cycle_task(16'b0001100000100110, 1'b0);
		prog_cycle_task(16'b1001100000100110, 1'b0);
		prog_cycle_task(16'b0000010000100110, 1'b0);
		prog_cycle_task(16'b1000010000100110, 1'b0);
		prog_cycle_task(16'b0100010000100110, 1'b0);
		prog_cycle_task(16'b1100010000100110, 1'b0);
		prog_cycle_task(16'b0010010000100110, 1'b0);
		prog_cycle_task(16'b1010010000100110, 1'b1);
		prog_cycle_task(16'b0001010000100110, 1'b0);
		prog_cycle_task(16'b1001010000100110, 1'b0);
		prog_cycle_task(16'b0101010000100110, 1'b1);
		prog_cycle_task(16'b1101010000100110, 1'b0);
		prog_cycle_task(16'b0011010000100110, 1'b0);
		prog_cycle_task(16'b1011010000100110, 1'b1);
		prog_cycle_task(16'b0000110000100110, 1'b0);
		prog_cycle_task(16'b1000110000100110, 1'b0);
		prog_cycle_task(16'b0100110000100110, 1'b1);
		prog_cycle_task(16'b1100110000100110, 1'b0);
		prog_cycle_task(16'b0010110000100110, 1'b0);
		prog_cycle_task(16'b1010110000100110, 1'b1);
		prog_cycle_task(16'b0001110000100110, 1'b0);
		prog_cycle_task(16'b1001110000100110, 1'b0);
		prog_cycle_task(16'b0101110000100110, 1'b1);
		prog_cycle_task(16'b1101110000100110, 1'b0);
		prog_cycle_task(16'b0011110000100110, 1'b0);
		prog_cycle_task(16'b1011110000100110, 1'b1);
		prog_cycle_task(16'b0000001000100110, 1'b1);
		prog_cycle_task(16'b1000001000100110, 1'b0);
		prog_cycle_task(16'b0100001000100110, 1'b0);
		prog_cycle_task(16'b1100001000100110, 1'b0);
		prog_cycle_task(16'b0010001000100110, 1'b0);
		prog_cycle_task(16'b1010001000100110, 1'b1);
		prog_cycle_task(16'b0001001000100110, 1'b0);
		prog_cycle_task(16'b1001001000100110, 1'b0);
		prog_cycle_task(16'b0101001000100110, 1'b1);
		prog_cycle_task(16'b1101001000100110, 1'b0);
		prog_cycle_task(16'b0011001000100110, 1'b0);
		prog_cycle_task(16'b1011001000100110, 1'b1);
		prog_cycle_task(16'b0000101000100110, 1'b0);
		prog_cycle_task(16'b1000101000100110, 1'b1);
		prog_cycle_task(16'b0100101000100110, 1'b0);
		prog_cycle_task(16'b1100101000100110, 1'b1);
		prog_cycle_task(16'b0010101000100110, 1'b0);
		prog_cycle_task(16'b1010101000100110, 1'b0);
		prog_cycle_task(16'b0000000000010110, 1'b0);
		prog_cycle_task(16'b1000000000010110, 1'b1);
		prog_cycle_task(16'b0100000000010110, 1'b0);
		prog_cycle_task(16'b1100000000010110, 1'b1);
		prog_cycle_task(16'b0010000000010110, 1'b0);
		prog_cycle_task(16'b1010000000010110, 1'b0);
		prog_cycle_task(16'b0001000000010110, 1'b0);
		prog_cycle_task(16'b1001000000010110, 1'b0);
		prog_cycle_task(16'b0000100000010110, 1'b0);
		prog_cycle_task(16'b1000100000010110, 1'b0);
		prog_cycle_task(16'b0100100000010110, 1'b0);
		prog_cycle_task(16'b1100100000010110, 1'b0);
		prog_cycle_task(16'b0010100000010110, 1'b0);
		prog_cycle_task(16'b1010100000010110, 1'b1);
		prog_cycle_task(16'b0001100000010110, 1'b0);
		prog_cycle_task(16'b1001100000010110, 1'b0);
		prog_cycle_task(16'b0101100000010110, 1'b0);
		prog_cycle_task(16'b1101100000010110, 1'b0);
		prog_cycle_task(16'b0011100000010110, 1'b0);
		prog_cycle_task(16'b1011100000010110, 1'b1);
		prog_cycle_task(16'b0000010000010110, 1'b0);
		prog_cycle_task(16'b1000010000010110, 1'b0);
		prog_cycle_task(16'b0100010000010110, 1'b0);
		prog_cycle_task(16'b1100010000010110, 1'b0);
		prog_cycle_task(16'b0010010000010110, 1'b0);
		prog_cycle_task(16'b1010010000010110, 1'b1);
		prog_cycle_task(16'b0001010000010110, 1'b0);
		prog_cycle_task(16'b1001010000010110, 1'b0);
		prog_cycle_task(16'b0101010000010110, 1'b0);
		prog_cycle_task(16'b1101010000010110, 1'b0);
		prog_cycle_task(16'b0011010000010110, 1'b0);
		prog_cycle_task(16'b1011010000010110, 1'b1);
		prog_cycle_task(16'b0000110000010110, 1'b0);
		prog_cycle_task(16'b1000110000010110, 1'b0);
		prog_cycle_task(16'b0100110000010110, 1'b0);
		prog_cycle_task(16'b1100110000010110, 1'b0);
		prog_cycle_task(16'b0010110000010110, 1'b0);
		prog_cycle_task(16'b1010110000010110, 1'b1);
		prog_cycle_task(16'b0001110000010110, 1'b0);
		prog_cycle_task(16'b1001110000010110, 1'b0);
		prog_cycle_task(16'b0101110000010110, 1'b0);
		prog_cycle_task(16'b1101110000010110, 1'b0);
		prog_cycle_task(16'b0011110000010110, 1'b0);
		prog_cycle_task(16'b1011110000010110, 1'b1);
		prog_cycle_task(16'b0000001000010110, 1'b0);
		prog_cycle_task(16'b1000001000010110, 1'b0);
		prog_cycle_task(16'b0100001000010110, 1'b0);
		prog_cycle_task(16'b1100001000010110, 1'b0);
		prog_cycle_task(16'b0010001000010110, 1'b0);
		prog_cycle_task(16'b1010001000010110, 1'b1);
		prog_cycle_task(16'b0001001000010110, 1'b0);
		prog_cycle_task(16'b1001001000010110, 1'b0);
		prog_cycle_task(16'b0101001000010110, 1'b1);
		prog_cycle_task(16'b1101001000010110, 1'b0);
		prog_cycle_task(16'b0011001000010110, 1'b1);
		prog_cycle_task(16'b1011001000010110, 1'b0);
		prog_cycle_task(16'b0000101000010110, 1'b0);
		prog_cycle_task(16'b1000101000010110, 1'b0);
		prog_cycle_task(16'b0100101000010110, 1'b0);
		prog_cycle_task(16'b1100101000010110, 1'b0);
		prog_cycle_task(16'b0010101000010110, 1'b0);
		prog_cycle_task(16'b1010101000010110, 1'b1);
		prog_cycle_task(16'b0000000000110110, 1'b0);
		prog_cycle_task(16'b1000000000110110, 1'b0);
		prog_cycle_task(16'b0100000000110110, 1'b0);
		prog_cycle_task(16'b1100000000110110, 1'b0);
		prog_cycle_task(16'b0010000000110110, 1'b0);
		prog_cycle_task(16'b1010000000110110, 1'b1);
		prog_cycle_task(16'b0001000000110110, 1'b0);
		prog_cycle_task(16'b1001000000110110, 1'b0);
		prog_cycle_task(16'b0000100000110110, 1'b0);
		prog_cycle_task(16'b1000100000110110, 1'b0);
		prog_cycle_task(16'b0100100000110110, 1'b0);
		prog_cycle_task(16'b1100100000110110, 1'b0);
		prog_cycle_task(16'b0010100000110110, 1'b0);
		prog_cycle_task(16'b1010100000110110, 1'b1);
		prog_cycle_task(16'b0001100000110110, 1'b0);
		prog_cycle_task(16'b1001100000110110, 1'b0);
		prog_cycle_task(16'b0000010000110110, 1'b1);
		prog_cycle_task(16'b1000010000110110, 1'b1);
		prog_cycle_task(16'b0000000000001110, 1'b0);
		prog_cycle_task(16'b1000000000001110, 1'b0);
		prog_cycle_task(16'b0100000000001110, 1'b0);
		prog_cycle_task(16'b1100000000001110, 1'b0);
		prog_cycle_task(16'b0010000000001110, 1'b0);
		prog_cycle_task(16'b1010000000001110, 1'b0);
		prog_cycle_task(16'b0110000000001110, 1'b0);
		prog_cycle_task(16'b1110000000001110, 1'b0);
		prog_cycle_task(16'b0001000000001110, 1'b0);
		prog_cycle_task(16'b1001000000001110, 1'b0);
		prog_cycle_task(16'b0101000000001110, 1'b0);
		prog_cycle_task(16'b1101000000001110, 1'b0);
		prog_cycle_task(16'b0011000000001110, 1'b0);
		prog_cycle_task(16'b1011000000001110, 1'b0);
		prog_cycle_task(16'b0111000000001110, 1'b0);
		prog_cycle_task(16'b1111000000001110, 1'b0);
		prog_cycle_task(16'b0000100000001110, 1'b0);
		prog_cycle_task(16'b1000100000001110, 1'b0);
		prog_cycle_task(16'b0100100000001110, 1'b1);
		prog_cycle_task(16'b0000010000001110, 1'b0);
		prog_cycle_task(16'b1000010000001110, 1'b0);
		prog_cycle_task(16'b0100010000001110, 1'b0);
		prog_cycle_task(16'b1100010000001110, 1'b0);
		prog_cycle_task(16'b0010010000001110, 1'b0);
		prog_cycle_task(16'b1010010000001110, 1'b0);
		prog_cycle_task(16'b0110010000001110, 1'b0);
		prog_cycle_task(16'b1110010000001110, 1'b0);
		prog_cycle_task(16'b0001010000001110, 1'b0);
		prog_cycle_task(16'b1001010000001110, 1'b0);
		prog_cycle_task(16'b0101010000001110, 1'b0);
		prog_cycle_task(16'b1101010000001110, 1'b0);
		prog_cycle_task(16'b0011010000001110, 1'b0);
		prog_cycle_task(16'b1011010000001110, 1'b0);
		prog_cycle_task(16'b0111010000001110, 1'b0);
		prog_cycle_task(16'b1111010000001110, 1'b0);
		prog_cycle_task(16'b0000110000001110, 1'b0);
		prog_cycle_task(16'b1000110000001110, 1'b0);
		prog_cycle_task(16'b0100110000001110, 1'b1);
		prog_cycle_task(16'b0000001000001110, 1'b0);
		prog_cycle_task(16'b1000001000001110, 1'b0);
		prog_cycle_task(16'b0100001000001110, 1'b0);
		prog_cycle_task(16'b1100001000001110, 1'b0);
		prog_cycle_task(16'b0010001000001110, 1'b0);
		prog_cycle_task(16'b1010001000001110, 1'b0);
		prog_cycle_task(16'b0110001000001110, 1'b0);
		prog_cycle_task(16'b1110001000001110, 1'b0);
		prog_cycle_task(16'b0001001000001110, 1'b0);
		prog_cycle_task(16'b1001001000001110, 1'b0);
		prog_cycle_task(16'b0101001000001110, 1'b0);
		prog_cycle_task(16'b1101001000001110, 1'b0);
		prog_cycle_task(16'b0011001000001110, 1'b0);
		prog_cycle_task(16'b1011001000001110, 1'b0);
		prog_cycle_task(16'b0111001000001110, 1'b0);
		prog_cycle_task(16'b1111001000001110, 1'b0);
		prog_cycle_task(16'b0000101000001110, 1'b0);
		prog_cycle_task(16'b1000101000001110, 1'b0);
		prog_cycle_task(16'b0100101000001110, 1'b1);
		prog_cycle_task(16'b0000011000001110, 1'b1);
		prog_cycle_task(16'b1000011000001110, 1'b0);
		prog_cycle_task(16'b0100011000001110, 1'b1);
		prog_cycle_task(16'b1100011000001110, 1'b0);
		prog_cycle_task(16'b0010011000001110, 1'b1);
		prog_cycle_task(16'b1010011000001110, 1'b0);
		prog_cycle_task(16'b0110011000001110, 1'b1);
		prog_cycle_task(16'b1110011000001110, 1'b0);
		prog_cycle_task(16'b0001011000001110, 1'b0);
		prog_cycle_task(16'b1001011000001110, 1'b0);
		prog_cycle_task(16'b0101011000001110, 1'b0);
		prog_cycle_task(16'b1101011000001110, 1'b0);
		prog_cycle_task(16'b0011011000001110, 1'b0);
		prog_cycle_task(16'b1011011000001110, 1'b0);
		prog_cycle_task(16'b0111011000001110, 1'b0);
		prog_cycle_task(16'b1111011000001110, 1'b0);
		prog_cycle_task(16'b0000111000001110, 1'b0);
		prog_cycle_task(16'b1000111000001110, 1'b1);
		prog_cycle_task(16'b0100111000001110, 1'b0);
		prog_cycle_task(16'b0000000100001110, 1'b0);
		prog_cycle_task(16'b1000000100001110, 1'b0);
		prog_cycle_task(16'b0100000100001110, 1'b1);
		prog_cycle_task(16'b1100000100001110, 1'b0);
		prog_cycle_task(16'b0010000100001110, 1'b0);
		prog_cycle_task(16'b1010000100001110, 1'b0);
		prog_cycle_task(16'b0110000100001110, 1'b0);
		prog_cycle_task(16'b1110000100001110, 1'b1);
		prog_cycle_task(16'b0000010100001110, 1'b0);
		prog_cycle_task(16'b1000010100001110, 1'b0);
		prog_cycle_task(16'b0100010100001110, 1'b1);
		prog_cycle_task(16'b1100010100001110, 1'b0);
		prog_cycle_task(16'b0010010100001110, 1'b0);
		prog_cycle_task(16'b1010010100001110, 1'b0);
		prog_cycle_task(16'b0110010100001110, 1'b0);
		prog_cycle_task(16'b1110010100001110, 1'b1);
		prog_cycle_task(16'b0000001100001110, 1'b0);
		prog_cycle_task(16'b1000001100001110, 1'b0);
		prog_cycle_task(16'b0100001100001110, 1'b1);
		prog_cycle_task(16'b1100001100001110, 1'b0);
		prog_cycle_task(16'b0010001100001110, 1'b0);
		prog_cycle_task(16'b1010001100001110, 1'b0);
		prog_cycle_task(16'b0110001100001110, 1'b0);
		prog_cycle_task(16'b1110001100001110, 1'b1);
		prog_cycle_task(16'b0000011100001110, 1'b0);
		prog_cycle_task(16'b1000011100001110, 1'b0);
		prog_cycle_task(16'b0100011100001110, 1'b1);
		prog_cycle_task(16'b1100011100001110, 1'b0);
		prog_cycle_task(16'b0010011100001110, 1'b0);
		prog_cycle_task(16'b1010011100001110, 1'b0);
		prog_cycle_task(16'b0110011100001110, 1'b0);
		prog_cycle_task(16'b1110011100001110, 1'b1);
		prog_cycle_task(16'b0000000010001110, 1'b0);
		prog_cycle_task(16'b1000000010001110, 1'b0);
		prog_cycle_task(16'b0100000010001110, 1'b1);
		prog_cycle_task(16'b1100000010001110, 1'b0);
		prog_cycle_task(16'b0010000010001110, 1'b0);
		prog_cycle_task(16'b1010000010001110, 1'b0);
		prog_cycle_task(16'b0110000010001110, 1'b0);
		prog_cycle_task(16'b1110000010001110, 1'b1);
		prog_cycle_task(16'b0000010010001110, 1'b0);
		prog_cycle_task(16'b1000010010001110, 1'b0);
		prog_cycle_task(16'b0100010010001110, 1'b1);
		prog_cycle_task(16'b1100010010001110, 1'b0);
		prog_cycle_task(16'b0010010010001110, 1'b0);
		prog_cycle_task(16'b1010010010001110, 1'b0);
		prog_cycle_task(16'b0110010010001110, 1'b0);
		prog_cycle_task(16'b1110010010001110, 1'b1);
		prog_cycle_task(16'b0000001010001110, 1'b0);
		prog_cycle_task(16'b1000001010001110, 1'b0);
		prog_cycle_task(16'b0100001010001110, 1'b1);
		prog_cycle_task(16'b1100001010001110, 1'b0);
		prog_cycle_task(16'b0010001010001110, 1'b0);
		prog_cycle_task(16'b1010001010001110, 1'b0);
		prog_cycle_task(16'b0110001010001110, 1'b0);
		prog_cycle_task(16'b1110001010001110, 1'b1);
		prog_cycle_task(16'b0000011010001110, 1'b0);
		prog_cycle_task(16'b1000011010001110, 1'b0);
		prog_cycle_task(16'b0100011010001110, 1'b1);
		prog_cycle_task(16'b1100011010001110, 1'b0);
		prog_cycle_task(16'b0010011010001110, 1'b0);
		prog_cycle_task(16'b1010011010001110, 1'b0);
		prog_cycle_task(16'b0110011010001110, 1'b0);
		prog_cycle_task(16'b1110011010001110, 1'b1);
		prog_cycle_task(16'b0000000110001110, 1'b0);
		prog_cycle_task(16'b1000000110001110, 1'b0);
		prog_cycle_task(16'b0100000110001110, 1'b1);
		prog_cycle_task(16'b1100000110001110, 1'b0);
		prog_cycle_task(16'b0010000110001110, 1'b0);
		prog_cycle_task(16'b1010000110001110, 1'b0);
		prog_cycle_task(16'b0110000110001110, 1'b0);
		prog_cycle_task(16'b1110000110001110, 1'b1);
		prog_cycle_task(16'b0000010110001110, 1'b0);
		prog_cycle_task(16'b1000010110001110, 1'b0);
		prog_cycle_task(16'b0100010110001110, 1'b1);
		prog_cycle_task(16'b1100010110001110, 1'b0);
		prog_cycle_task(16'b0010010110001110, 1'b0);
		prog_cycle_task(16'b1010010110001110, 1'b0);
		prog_cycle_task(16'b0110010110001110, 1'b0);
		prog_cycle_task(16'b1110010110001110, 1'b1);
		prog_cycle_task(16'b0000001110001110, 1'b0);
		prog_cycle_task(16'b1000001110001110, 1'b0);
		prog_cycle_task(16'b0100001110001110, 1'b1);
		prog_cycle_task(16'b1100001110001110, 1'b0);
		prog_cycle_task(16'b0010001110001110, 1'b0);
		prog_cycle_task(16'b1010001110001110, 1'b0);
		prog_cycle_task(16'b0110001110001110, 1'b0);
		prog_cycle_task(16'b1110001110001110, 1'b1);
		prog_cycle_task(16'b0000011110001110, 1'b0);
		prog_cycle_task(16'b1000011110001110, 1'b0);
		prog_cycle_task(16'b0100011110001110, 1'b1);
		prog_cycle_task(16'b1100011110001110, 1'b0);
		prog_cycle_task(16'b0010011110001110, 1'b0);
		prog_cycle_task(16'b1010011110001110, 1'b0);
		prog_cycle_task(16'b0110011110001110, 1'b0);
		prog_cycle_task(16'b1110011110001110, 1'b1);
		prog_cycle_task(16'b0000000001001110, 1'b0);
		prog_cycle_task(16'b1000000001001110, 1'b1);
		prog_cycle_task(16'b0100000001001110, 1'b0);
		prog_cycle_task(16'b1100000001001110, 1'b0);
		prog_cycle_task(16'b0010000001001110, 1'b0);
		prog_cycle_task(16'b1010000001001110, 1'b0);
		prog_cycle_task(16'b0110000001001110, 1'b1);
		prog_cycle_task(16'b1110000001001110, 1'b0);
		prog_cycle_task(16'b0000010001001110, 1'b0);
		prog_cycle_task(16'b1000010001001110, 1'b0);
		prog_cycle_task(16'b0100010001001110, 1'b1);
		prog_cycle_task(16'b1100010001001110, 1'b0);
		prog_cycle_task(16'b0010010001001110, 1'b0);
		prog_cycle_task(16'b1010010001001110, 1'b0);
		prog_cycle_task(16'b0110010001001110, 1'b0);
		prog_cycle_task(16'b1110010001001110, 1'b1);
		prog_cycle_task(16'b0000001001001110, 1'b0);
		prog_cycle_task(16'b1000001001001110, 1'b0);
		prog_cycle_task(16'b0100001001001110, 1'b1);
		prog_cycle_task(16'b1100001001001110, 1'b0);
		prog_cycle_task(16'b0010001001001110, 1'b0);
		prog_cycle_task(16'b1010001001001110, 1'b0);
		prog_cycle_task(16'b0110001001001110, 1'b0);
		prog_cycle_task(16'b1110001001001110, 1'b1);
		prog_cycle_task(16'b0000011001001110, 1'b0);
		prog_cycle_task(16'b1000011001001110, 1'b0);
		prog_cycle_task(16'b0100011001001110, 1'b1);
		prog_cycle_task(16'b1100011001001110, 1'b0);
		prog_cycle_task(16'b0010011001001110, 1'b1);
		prog_cycle_task(16'b1010011001001110, 1'b0);
		prog_cycle_task(16'b0110011001001110, 1'b0);
		prog_cycle_task(16'b1110011001001110, 1'b0);
		prog_cycle_task(16'b0000000000101110, 1'b0);
		prog_cycle_task(16'b1000000000101110, 1'b0);
		prog_cycle_task(16'b0100000000101110, 1'b0);
		prog_cycle_task(16'b1100000000101110, 1'b0);
		prog_cycle_task(16'b0010000000101110, 1'b0);
		prog_cycle_task(16'b1010000000101110, 1'b1);
		prog_cycle_task(16'b0001000000101110, 1'b0);
		prog_cycle_task(16'b1001000000101110, 1'b0);
		prog_cycle_task(16'b0000100000101110, 1'b0);
		prog_cycle_task(16'b1000100000101110, 1'b0);
		prog_cycle_task(16'b0001100000101110, 1'b0);
		prog_cycle_task(16'b1001100000101110, 1'b0);
		prog_cycle_task(16'b0000010000101110, 1'b0);
		prog_cycle_task(16'b1000010000101110, 1'b0);
		prog_cycle_task(16'b0100010000101110, 1'b0);
		prog_cycle_task(16'b1100010000101110, 1'b0);
		prog_cycle_task(16'b0010010000101110, 1'b0);
		prog_cycle_task(16'b1010010000101110, 1'b1);
		prog_cycle_task(16'b0001010000101110, 1'b0);
		prog_cycle_task(16'b1001010000101110, 1'b0);
		prog_cycle_task(16'b0101010000101110, 1'b1);
		prog_cycle_task(16'b1101010000101110, 1'b0);
		prog_cycle_task(16'b0011010000101110, 1'b0);
		prog_cycle_task(16'b1011010000101110, 1'b1);
		prog_cycle_task(16'b0000110000101110, 1'b0);
		prog_cycle_task(16'b1000110000101110, 1'b0);
		prog_cycle_task(16'b0100110000101110, 1'b1);
		prog_cycle_task(16'b1100110000101110, 1'b0);
		prog_cycle_task(16'b0010110000101110, 1'b0);
		prog_cycle_task(16'b1010110000101110, 1'b1);
		prog_cycle_task(16'b0001110000101110, 1'b0);
		prog_cycle_task(16'b1001110000101110, 1'b0);
		prog_cycle_task(16'b0101110000101110, 1'b1);
		prog_cycle_task(16'b1101110000101110, 1'b0);
		prog_cycle_task(16'b0011110000101110, 1'b0);
		prog_cycle_task(16'b1011110000101110, 1'b1);
		prog_cycle_task(16'b0000001000101110, 1'b0);
		prog_cycle_task(16'b1000001000101110, 1'b0);
		prog_cycle_task(16'b0100001000101110, 1'b1);
		prog_cycle_task(16'b1100001000101110, 1'b0);
		prog_cycle_task(16'b0010001000101110, 1'b0);
		prog_cycle_task(16'b1010001000101110, 1'b1);
		prog_cycle_task(16'b0001001000101110, 1'b0);
		prog_cycle_task(16'b1001001000101110, 1'b0);
		prog_cycle_task(16'b0101001000101110, 1'b1);
		prog_cycle_task(16'b1101001000101110, 1'b0);
		prog_cycle_task(16'b0011001000101110, 1'b0);
		prog_cycle_task(16'b1011001000101110, 1'b1);
		prog_cycle_task(16'b0000101000101110, 1'b0);
		prog_cycle_task(16'b1000101000101110, 1'b0);
		prog_cycle_task(16'b0100101000101110, 1'b1);
		prog_cycle_task(16'b1100101000101110, 1'b0);
		prog_cycle_task(16'b0010101000101110, 1'b0);
		prog_cycle_task(16'b1010101000101110, 1'b1);
		prog_cycle_task(16'b0000000000011110, 1'b0);
		prog_cycle_task(16'b1000000000011110, 1'b0);
		prog_cycle_task(16'b0100000000011110, 1'b0);
		prog_cycle_task(16'b1100000000011110, 1'b0);
		prog_cycle_task(16'b0010000000011110, 1'b0);
		prog_cycle_task(16'b1010000000011110, 1'b1);
		prog_cycle_task(16'b0001000000011110, 1'b0);
		prog_cycle_task(16'b1001000000011110, 1'b0);
		prog_cycle_task(16'b0000100000011110, 1'b0);
		prog_cycle_task(16'b1000100000011110, 1'b0);
		prog_cycle_task(16'b0100100000011110, 1'b0);
		prog_cycle_task(16'b1100100000011110, 1'b0);
		prog_cycle_task(16'b0010100000011110, 1'b0);
		prog_cycle_task(16'b1010100000011110, 1'b1);
		prog_cycle_task(16'b0001100000011110, 1'b0);
		prog_cycle_task(16'b1001100000011110, 1'b0);
		prog_cycle_task(16'b0101100000011110, 1'b0);
		prog_cycle_task(16'b1101100000011110, 1'b0);
		prog_cycle_task(16'b0011100000011110, 1'b0);
		prog_cycle_task(16'b1011100000011110, 1'b1);
		prog_cycle_task(16'b0000010000011110, 1'b0);
		prog_cycle_task(16'b1000010000011110, 1'b0);
		prog_cycle_task(16'b0100010000011110, 1'b0);
		prog_cycle_task(16'b1100010000011110, 1'b0);
		prog_cycle_task(16'b0010010000011110, 1'b0);
		prog_cycle_task(16'b1010010000011110, 1'b1);
		prog_cycle_task(16'b0001010000011110, 1'b0);
		prog_cycle_task(16'b1001010000011110, 1'b0);
		prog_cycle_task(16'b0101010000011110, 1'b0);
		prog_cycle_task(16'b1101010000011110, 1'b0);
		prog_cycle_task(16'b0011010000011110, 1'b0);
		prog_cycle_task(16'b1011010000011110, 1'b1);
		prog_cycle_task(16'b0000110000011110, 1'b0);
		prog_cycle_task(16'b1000110000011110, 1'b0);
		prog_cycle_task(16'b0100110000011110, 1'b0);
		prog_cycle_task(16'b1100110000011110, 1'b0);
		prog_cycle_task(16'b0010110000011110, 1'b0);
		prog_cycle_task(16'b1010110000011110, 1'b1);
		prog_cycle_task(16'b0001110000011110, 1'b0);
		prog_cycle_task(16'b1001110000011110, 1'b0);
		prog_cycle_task(16'b0101110000011110, 1'b0);
		prog_cycle_task(16'b1101110000011110, 1'b0);
		prog_cycle_task(16'b0011110000011110, 1'b0);
		prog_cycle_task(16'b1011110000011110, 1'b1);
		prog_cycle_task(16'b0000001000011110, 1'b0);
		prog_cycle_task(16'b1000001000011110, 1'b0);
		prog_cycle_task(16'b0100001000011110, 1'b0);
		prog_cycle_task(16'b1100001000011110, 1'b0);
		prog_cycle_task(16'b0010001000011110, 1'b0);
		prog_cycle_task(16'b1010001000011110, 1'b1);
		prog_cycle_task(16'b0001001000011110, 1'b0);
		prog_cycle_task(16'b1001001000011110, 1'b0);
		prog_cycle_task(16'b0101001000011110, 1'b0);
		prog_cycle_task(16'b1101001000011110, 1'b0);
		prog_cycle_task(16'b0011001000011110, 1'b0);
		prog_cycle_task(16'b1011001000011110, 1'b1);
		prog_cycle_task(16'b0000101000011110, 1'b0);
		prog_cycle_task(16'b1000101000011110, 1'b0);
		prog_cycle_task(16'b0100101000011110, 1'b0);
		prog_cycle_task(16'b1100101000011110, 1'b0);
		prog_cycle_task(16'b0010101000011110, 1'b0);
		prog_cycle_task(16'b1010101000011110, 1'b1);
		prog_cycle_task(16'b0000000000111110, 1'b0);
		prog_cycle_task(16'b1000000000111110, 1'b0);
		prog_cycle_task(16'b0100000000111110, 1'b0);
		prog_cycle_task(16'b1100000000111110, 1'b0);
		prog_cycle_task(16'b0010000000111110, 1'b0);
		prog_cycle_task(16'b1010000000111110, 1'b1);
		prog_cycle_task(16'b0001000000111110, 1'b0);
		prog_cycle_task(16'b1001000000111110, 1'b0);
		prog_cycle_task(16'b0000100000111110, 1'b0);
		prog_cycle_task(16'b1000100000111110, 1'b0);
		prog_cycle_task(16'b0100100000111110, 1'b0);
		prog_cycle_task(16'b1100100000111110, 1'b0);
		prog_cycle_task(16'b0010100000111110, 1'b0);
		prog_cycle_task(16'b1010100000111110, 1'b1);
		prog_cycle_task(16'b0001100000111110, 1'b0);
		prog_cycle_task(16'b1001100000111110, 1'b0);
		prog_cycle_task(16'b0000010000111110, 1'b0);
		prog_cycle_task(16'b1000010000111110, 1'b0);
		prog_cycle_task(16'b0000000000000001, 1'b0);
		prog_cycle_task(16'b1000000000000001, 1'b0);
		prog_cycle_task(16'b0100000000000001, 1'b0);
		prog_cycle_task(16'b1100000000000001, 1'b0);
		prog_cycle_task(16'b0010000000000001, 1'b0);
		prog_cycle_task(16'b1010000000000001, 1'b0);
		prog_cycle_task(16'b0110000000000001, 1'b0);
		prog_cycle_task(16'b1110000000000001, 1'b0);
		prog_cycle_task(16'b0001000000000001, 1'b0);
		prog_cycle_task(16'b1001000000000001, 1'b0);
		prog_cycle_task(16'b0101000000000001, 1'b0);
		prog_cycle_task(16'b1101000000000001, 1'b0);
		prog_cycle_task(16'b0011000000000001, 1'b0);
		prog_cycle_task(16'b1011000000000001, 1'b0);
		prog_cycle_task(16'b0111000000000001, 1'b0);
		prog_cycle_task(16'b1111000000000001, 1'b0);
		prog_cycle_task(16'b0000100000000001, 1'b0);
		prog_cycle_task(16'b1000100000000001, 1'b0);
		prog_cycle_task(16'b0100100000000001, 1'b1);
		prog_cycle_task(16'b0000010000000001, 1'b0);
		prog_cycle_task(16'b1000010000000001, 1'b0);
		prog_cycle_task(16'b0100010000000001, 1'b0);
		prog_cycle_task(16'b1100010000000001, 1'b0);
		prog_cycle_task(16'b0010010000000001, 1'b0);
		prog_cycle_task(16'b1010010000000001, 1'b0);
		prog_cycle_task(16'b0110010000000001, 1'b0);
		prog_cycle_task(16'b1110010000000001, 1'b0);
		prog_cycle_task(16'b0001010000000001, 1'b0);
		prog_cycle_task(16'b1001010000000001, 1'b0);
		prog_cycle_task(16'b0101010000000001, 1'b0);
		prog_cycle_task(16'b1101010000000001, 1'b0);
		prog_cycle_task(16'b0011010000000001, 1'b0);
		prog_cycle_task(16'b1011010000000001, 1'b0);
		prog_cycle_task(16'b0111010000000001, 1'b0);
		prog_cycle_task(16'b1111010000000001, 1'b0);
		prog_cycle_task(16'b0000110000000001, 1'b0);
		prog_cycle_task(16'b1000110000000001, 1'b0);
		prog_cycle_task(16'b0100110000000001, 1'b1);
		prog_cycle_task(16'b0000001000000001, 1'b0);
		prog_cycle_task(16'b1000001000000001, 1'b0);
		prog_cycle_task(16'b0100001000000001, 1'b0);
		prog_cycle_task(16'b1100001000000001, 1'b0);
		prog_cycle_task(16'b0010001000000001, 1'b0);
		prog_cycle_task(16'b1010001000000001, 1'b0);
		prog_cycle_task(16'b0110001000000001, 1'b0);
		prog_cycle_task(16'b1110001000000001, 1'b0);
		prog_cycle_task(16'b0001001000000001, 1'b0);
		prog_cycle_task(16'b1001001000000001, 1'b0);
		prog_cycle_task(16'b0101001000000001, 1'b0);
		prog_cycle_task(16'b1101001000000001, 1'b0);
		prog_cycle_task(16'b0011001000000001, 1'b0);
		prog_cycle_task(16'b1011001000000001, 1'b0);
		prog_cycle_task(16'b0111001000000001, 1'b0);
		prog_cycle_task(16'b1111001000000001, 1'b0);
		prog_cycle_task(16'b0000101000000001, 1'b0);
		prog_cycle_task(16'b1000101000000001, 1'b0);
		prog_cycle_task(16'b0100101000000001, 1'b1);
		prog_cycle_task(16'b0000011000000001, 1'b0);
		prog_cycle_task(16'b1000011000000001, 1'b0);
		prog_cycle_task(16'b0100011000000001, 1'b0);
		prog_cycle_task(16'b1100011000000001, 1'b0);
		prog_cycle_task(16'b0010011000000001, 1'b0);
		prog_cycle_task(16'b1010011000000001, 1'b0);
		prog_cycle_task(16'b0110011000000001, 1'b0);
		prog_cycle_task(16'b1110011000000001, 1'b0);
		prog_cycle_task(16'b0001011000000001, 1'b0);
		prog_cycle_task(16'b1001011000000001, 1'b0);
		prog_cycle_task(16'b0101011000000001, 1'b0);
		prog_cycle_task(16'b1101011000000001, 1'b0);
		prog_cycle_task(16'b0011011000000001, 1'b0);
		prog_cycle_task(16'b1011011000000001, 1'b0);
		prog_cycle_task(16'b0111011000000001, 1'b0);
		prog_cycle_task(16'b1111011000000001, 1'b0);
		prog_cycle_task(16'b0000111000000001, 1'b0);
		prog_cycle_task(16'b1000111000000001, 1'b0);
		prog_cycle_task(16'b0100111000000001, 1'b1);
		prog_cycle_task(16'b0000000100000001, 1'b0);
		prog_cycle_task(16'b1000000100000001, 1'b0);
		prog_cycle_task(16'b0100000100000001, 1'b1);
		prog_cycle_task(16'b1100000100000001, 1'b0);
		prog_cycle_task(16'b0010000100000001, 1'b0);
		prog_cycle_task(16'b1010000100000001, 1'b0);
		prog_cycle_task(16'b0110000100000001, 1'b0);
		prog_cycle_task(16'b1110000100000001, 1'b1);
		prog_cycle_task(16'b0000010100000001, 1'b0);
		prog_cycle_task(16'b1000010100000001, 1'b0);
		prog_cycle_task(16'b0100010100000001, 1'b1);
		prog_cycle_task(16'b1100010100000001, 1'b0);
		prog_cycle_task(16'b0010010100000001, 1'b0);
		prog_cycle_task(16'b1010010100000001, 1'b0);
		prog_cycle_task(16'b0110010100000001, 1'b0);
		prog_cycle_task(16'b1110010100000001, 1'b1);
		prog_cycle_task(16'b0000001100000001, 1'b0);
		prog_cycle_task(16'b1000001100000001, 1'b0);
		prog_cycle_task(16'b0100001100000001, 1'b1);
		prog_cycle_task(16'b1100001100000001, 1'b0);
		prog_cycle_task(16'b0010001100000001, 1'b0);
		prog_cycle_task(16'b1010001100000001, 1'b0);
		prog_cycle_task(16'b0110001100000001, 1'b0);
		prog_cycle_task(16'b1110001100000001, 1'b1);
		prog_cycle_task(16'b0000011100000001, 1'b0);
		prog_cycle_task(16'b1000011100000001, 1'b0);
		prog_cycle_task(16'b0100011100000001, 1'b1);
		prog_cycle_task(16'b1100011100000001, 1'b0);
		prog_cycle_task(16'b0010011100000001, 1'b0);
		prog_cycle_task(16'b1010011100000001, 1'b0);
		prog_cycle_task(16'b0110011100000001, 1'b0);
		prog_cycle_task(16'b1110011100000001, 1'b1);
		prog_cycle_task(16'b0000000010000001, 1'b0);
		prog_cycle_task(16'b1000000010000001, 1'b0);
		prog_cycle_task(16'b0100000010000001, 1'b1);
		prog_cycle_task(16'b1100000010000001, 1'b0);
		prog_cycle_task(16'b0010000010000001, 1'b0);
		prog_cycle_task(16'b1010000010000001, 1'b0);
		prog_cycle_task(16'b0110000010000001, 1'b0);
		prog_cycle_task(16'b1110000010000001, 1'b1);
		prog_cycle_task(16'b0000010010000001, 1'b0);
		prog_cycle_task(16'b1000010010000001, 1'b0);
		prog_cycle_task(16'b0100010010000001, 1'b1);
		prog_cycle_task(16'b1100010010000001, 1'b0);
		prog_cycle_task(16'b0010010010000001, 1'b0);
		prog_cycle_task(16'b1010010010000001, 1'b0);
		prog_cycle_task(16'b0110010010000001, 1'b0);
		prog_cycle_task(16'b1110010010000001, 1'b1);
		prog_cycle_task(16'b0000001010000001, 1'b0);
		prog_cycle_task(16'b1000001010000001, 1'b0);
		prog_cycle_task(16'b0100001010000001, 1'b1);
		prog_cycle_task(16'b1100001010000001, 1'b0);
		prog_cycle_task(16'b0010001010000001, 1'b0);
		prog_cycle_task(16'b1010001010000001, 1'b0);
		prog_cycle_task(16'b0110001010000001, 1'b0);
		prog_cycle_task(16'b1110001010000001, 1'b1);
		prog_cycle_task(16'b0000011010000001, 1'b0);
		prog_cycle_task(16'b1000011010000001, 1'b0);
		prog_cycle_task(16'b0100011010000001, 1'b1);
		prog_cycle_task(16'b1100011010000001, 1'b0);
		prog_cycle_task(16'b0010011010000001, 1'b0);
		prog_cycle_task(16'b1010011010000001, 1'b0);
		prog_cycle_task(16'b0110011010000001, 1'b0);
		prog_cycle_task(16'b1110011010000001, 1'b1);
		prog_cycle_task(16'b0000000110000001, 1'b0);
		prog_cycle_task(16'b1000000110000001, 1'b0);
		prog_cycle_task(16'b0100000110000001, 1'b1);
		prog_cycle_task(16'b1100000110000001, 1'b0);
		prog_cycle_task(16'b0010000110000001, 1'b0);
		prog_cycle_task(16'b1010000110000001, 1'b0);
		prog_cycle_task(16'b0110000110000001, 1'b0);
		prog_cycle_task(16'b1110000110000001, 1'b1);
		prog_cycle_task(16'b0000010110000001, 1'b0);
		prog_cycle_task(16'b1000010110000001, 1'b0);
		prog_cycle_task(16'b0100010110000001, 1'b1);
		prog_cycle_task(16'b1100010110000001, 1'b0);
		prog_cycle_task(16'b0010010110000001, 1'b0);
		prog_cycle_task(16'b1010010110000001, 1'b0);
		prog_cycle_task(16'b0110010110000001, 1'b0);
		prog_cycle_task(16'b1110010110000001, 1'b1);
		prog_cycle_task(16'b0000001110000001, 1'b0);
		prog_cycle_task(16'b1000001110000001, 1'b0);
		prog_cycle_task(16'b0100001110000001, 1'b1);
		prog_cycle_task(16'b1100001110000001, 1'b0);
		prog_cycle_task(16'b0010001110000001, 1'b0);
		prog_cycle_task(16'b1010001110000001, 1'b0);
		prog_cycle_task(16'b0110001110000001, 1'b0);
		prog_cycle_task(16'b1110001110000001, 1'b1);
		prog_cycle_task(16'b0000011110000001, 1'b0);
		prog_cycle_task(16'b1000011110000001, 1'b0);
		prog_cycle_task(16'b0100011110000001, 1'b1);
		prog_cycle_task(16'b1100011110000001, 1'b0);
		prog_cycle_task(16'b0010011110000001, 1'b0);
		prog_cycle_task(16'b1010011110000001, 1'b0);
		prog_cycle_task(16'b0110011110000001, 1'b0);
		prog_cycle_task(16'b1110011110000001, 1'b1);
		prog_cycle_task(16'b0000000001000001, 1'b0);
		prog_cycle_task(16'b1000000001000001, 1'b0);
		prog_cycle_task(16'b0100000001000001, 1'b1);
		prog_cycle_task(16'b1100000001000001, 1'b0);
		prog_cycle_task(16'b0010000001000001, 1'b0);
		prog_cycle_task(16'b1010000001000001, 1'b0);
		prog_cycle_task(16'b0110000001000001, 1'b0);
		prog_cycle_task(16'b1110000001000001, 1'b1);
		prog_cycle_task(16'b0000010001000001, 1'b0);
		prog_cycle_task(16'b1000010001000001, 1'b0);
		prog_cycle_task(16'b0100010001000001, 1'b1);
		prog_cycle_task(16'b1100010001000001, 1'b0);
		prog_cycle_task(16'b0010010001000001, 1'b0);
		prog_cycle_task(16'b1010010001000001, 1'b0);
		prog_cycle_task(16'b0110010001000001, 1'b0);
		prog_cycle_task(16'b1110010001000001, 1'b1);
		prog_cycle_task(16'b0000001001000001, 1'b0);
		prog_cycle_task(16'b1000001001000001, 1'b0);
		prog_cycle_task(16'b0100001001000001, 1'b1);
		prog_cycle_task(16'b1100001001000001, 1'b0);
		prog_cycle_task(16'b0010001001000001, 1'b0);
		prog_cycle_task(16'b1010001001000001, 1'b0);
		prog_cycle_task(16'b0110001001000001, 1'b0);
		prog_cycle_task(16'b1110001001000001, 1'b1);
		prog_cycle_task(16'b0000011001000001, 1'b0);
		prog_cycle_task(16'b1000011001000001, 1'b0);
		prog_cycle_task(16'b0100011001000001, 1'b1);
		prog_cycle_task(16'b1100011001000001, 1'b0);
		prog_cycle_task(16'b0010011001000001, 1'b0);
		prog_cycle_task(16'b1010011001000001, 1'b0);
		prog_cycle_task(16'b0110011001000001, 1'b0);
		prog_cycle_task(16'b1110011001000001, 1'b1);
		prog_cycle_task(16'b0000000000100001, 1'b0);
		prog_cycle_task(16'b1000000000100001, 1'b0);
		prog_cycle_task(16'b0100000000100001, 1'b0);
		prog_cycle_task(16'b1100000000100001, 1'b0);
		prog_cycle_task(16'b0010000000100001, 1'b0);
		prog_cycle_task(16'b1010000000100001, 1'b0);
		prog_cycle_task(16'b0110000000100001, 1'b0);
		prog_cycle_task(16'b1110000000100001, 1'b0);
		prog_cycle_task(16'b0001000000100001, 1'b0);
		prog_cycle_task(16'b1001000000100001, 1'b0);
		prog_cycle_task(16'b0101000000100001, 1'b0);
		prog_cycle_task(16'b1101000000100001, 1'b0);
		prog_cycle_task(16'b0011000000100001, 1'b0);
		prog_cycle_task(16'b1011000000100001, 1'b0);
		prog_cycle_task(16'b0111000000100001, 1'b0);
		prog_cycle_task(16'b1111000000100001, 1'b0);
		prog_cycle_task(16'b0000100000100001, 1'b0);
		prog_cycle_task(16'b1000100000100001, 1'b0);
		prog_cycle_task(16'b0100100000100001, 1'b0);
		prog_cycle_task(16'b1100100000100001, 1'b0);
		prog_cycle_task(16'b0010100000100001, 1'b0);
		prog_cycle_task(16'b1010100000100001, 1'b0);
		prog_cycle_task(16'b0110100000100001, 1'b0);
		prog_cycle_task(16'b1110100000100001, 1'b0);
		prog_cycle_task(16'b0001100000100001, 1'b0);
		prog_cycle_task(16'b1001100000100001, 1'b0);
		prog_cycle_task(16'b0101100000100001, 1'b0);
		prog_cycle_task(16'b1101100000100001, 1'b0);
		prog_cycle_task(16'b0011100000100001, 1'b0);
		prog_cycle_task(16'b1011100000100001, 1'b0);
		prog_cycle_task(16'b0111100000100001, 1'b0);
		prog_cycle_task(16'b1111100000100001, 1'b0);
		prog_cycle_task(16'b0000010000100001, 1'b0);
		prog_cycle_task(16'b1000010000100001, 1'b0);
		prog_cycle_task(16'b0100010000100001, 1'b0);
		prog_cycle_task(16'b1100010000100001, 1'b0);
		prog_cycle_task(16'b0000000000010001, 1'b0);
		prog_cycle_task(16'b1000000000010001, 1'b0);
		prog_cycle_task(16'b0100000000010001, 1'b0);
		prog_cycle_task(16'b1100000000010001, 1'b0);
		prog_cycle_task(16'b0010000000010001, 1'b0);
		prog_cycle_task(16'b1010000000010001, 1'b1);
		prog_cycle_task(16'b0001000000010001, 1'b0);
		prog_cycle_task(16'b1001000000010001, 1'b0);
		prog_cycle_task(16'b0000100000010001, 1'b0);
		prog_cycle_task(16'b1000100000010001, 1'b0);
		prog_cycle_task(16'b0100100000010001, 1'b0);
		prog_cycle_task(16'b1100100000010001, 1'b0);
		prog_cycle_task(16'b0010100000010001, 1'b0);
		prog_cycle_task(16'b1010100000010001, 1'b1);
		prog_cycle_task(16'b0001100000010001, 1'b0);
		prog_cycle_task(16'b1001100000010001, 1'b0);
		prog_cycle_task(16'b0101100000010001, 1'b0);
		prog_cycle_task(16'b1101100000010001, 1'b0);
		prog_cycle_task(16'b0011100000010001, 1'b0);
		prog_cycle_task(16'b1011100000010001, 1'b1);
		prog_cycle_task(16'b0000010000010001, 1'b0);
		prog_cycle_task(16'b1000010000010001, 1'b0);
		prog_cycle_task(16'b0100010000010001, 1'b0);
		prog_cycle_task(16'b1100010000010001, 1'b0);
		prog_cycle_task(16'b0010010000010001, 1'b0);
		prog_cycle_task(16'b1010010000010001, 1'b1);
		prog_cycle_task(16'b0001010000010001, 1'b0);
		prog_cycle_task(16'b1001010000010001, 1'b0);
		prog_cycle_task(16'b0101010000010001, 1'b0);
		prog_cycle_task(16'b1101010000010001, 1'b0);
		prog_cycle_task(16'b0011010000010001, 1'b0);
		prog_cycle_task(16'b1011010000010001, 1'b1);
		prog_cycle_task(16'b0000110000010001, 1'b0);
		prog_cycle_task(16'b1000110000010001, 1'b0);
		prog_cycle_task(16'b0100110000010001, 1'b0);
		prog_cycle_task(16'b1100110000010001, 1'b0);
		prog_cycle_task(16'b0010110000010001, 1'b0);
		prog_cycle_task(16'b1010110000010001, 1'b1);
		prog_cycle_task(16'b0001110000010001, 1'b0);
		prog_cycle_task(16'b1001110000010001, 1'b0);
		prog_cycle_task(16'b0101110000010001, 1'b0);
		prog_cycle_task(16'b1101110000010001, 1'b0);
		prog_cycle_task(16'b0011110000010001, 1'b0);
		prog_cycle_task(16'b1011110000010001, 1'b1);
		prog_cycle_task(16'b0000001000010001, 1'b0);
		prog_cycle_task(16'b1000001000010001, 1'b0);
		prog_cycle_task(16'b0100001000010001, 1'b0);
		prog_cycle_task(16'b1100001000010001, 1'b0);
		prog_cycle_task(16'b0010001000010001, 1'b0);
		prog_cycle_task(16'b1010001000010001, 1'b1);
		prog_cycle_task(16'b0001001000010001, 1'b0);
		prog_cycle_task(16'b1001001000010001, 1'b0);
		prog_cycle_task(16'b0101001000010001, 1'b0);
		prog_cycle_task(16'b1101001000010001, 1'b0);
		prog_cycle_task(16'b0011001000010001, 1'b0);
		prog_cycle_task(16'b1011001000010001, 1'b1);
		prog_cycle_task(16'b0000101000010001, 1'b0);
		prog_cycle_task(16'b1000101000010001, 1'b0);
		prog_cycle_task(16'b0100101000010001, 1'b0);
		prog_cycle_task(16'b1100101000010001, 1'b0);
		prog_cycle_task(16'b0010101000010001, 1'b0);
		prog_cycle_task(16'b1010101000010001, 1'b1);
		prog_cycle_task(16'b0000000000110001, 1'b0);
		prog_cycle_task(16'b1000000000110001, 1'b0);
		prog_cycle_task(16'b0100000000110001, 1'b0);
		prog_cycle_task(16'b1100000000110001, 1'b0);
		prog_cycle_task(16'b0010000000110001, 1'b0);
		prog_cycle_task(16'b1010000000110001, 1'b1);
		prog_cycle_task(16'b0001000000110001, 1'b0);
		prog_cycle_task(16'b1001000000110001, 1'b0);
		prog_cycle_task(16'b0101000000110001, 1'b0);
		prog_cycle_task(16'b1101000000110001, 1'b0);
		prog_cycle_task(16'b0011000000110001, 1'b0);
		prog_cycle_task(16'b1011000000110001, 1'b1);
		prog_cycle_task(16'b0000100000110001, 1'b0);
		prog_cycle_task(16'b1000100000110001, 1'b0);
		prog_cycle_task(16'b0100100000110001, 1'b0);
		prog_cycle_task(16'b1100100000110001, 1'b0);
		prog_cycle_task(16'b0010100000110001, 1'b0);
		prog_cycle_task(16'b1010100000110001, 1'b1);
		prog_cycle_task(16'b0001100000110001, 1'b0);
		prog_cycle_task(16'b1001100000110001, 1'b0);
		prog_cycle_task(16'b0101100000110001, 1'b0);
		prog_cycle_task(16'b1101100000110001, 1'b0);
		prog_cycle_task(16'b0011100000110001, 1'b0);
		prog_cycle_task(16'b1011100000110001, 1'b1);
		prog_cycle_task(16'b0000010000110001, 1'b0);
		prog_cycle_task(16'b1000010000110001, 1'b0);
		prog_cycle_task(16'b0100010000110001, 1'b0);
		prog_cycle_task(16'b1100010000110001, 1'b0);
		prog_cycle_task(16'b0010010000110001, 1'b0);
		prog_cycle_task(16'b1010010000110001, 1'b1);
		prog_cycle_task(16'b0001010000110001, 1'b0);
		prog_cycle_task(16'b1001010000110001, 1'b0);
		prog_cycle_task(16'b0101010000110001, 1'b0);
		prog_cycle_task(16'b1101010000110001, 1'b0);
		prog_cycle_task(16'b0011010000110001, 1'b0);
		prog_cycle_task(16'b1011010000110001, 1'b1);
		prog_cycle_task(16'b0000110000110001, 1'b0);
		prog_cycle_task(16'b1000110000110001, 1'b0);
		prog_cycle_task(16'b0100110000110001, 1'b0);
		prog_cycle_task(16'b1100110000110001, 1'b0);
		prog_cycle_task(16'b0010110000110001, 1'b0);
		prog_cycle_task(16'b1010110000110001, 1'b1);
		prog_cycle_task(16'b0001110000110001, 1'b0);
		prog_cycle_task(16'b1001110000110001, 1'b0);
		prog_cycle_task(16'b0101110000110001, 1'b0);
		prog_cycle_task(16'b1101110000110001, 1'b0);
		prog_cycle_task(16'b0011110000110001, 1'b0);
		prog_cycle_task(16'b1011110000110001, 1'b1);
		prog_cycle_task(16'b0000001000110001, 1'b0);
		prog_cycle_task(16'b1000001000110001, 1'b0);
		prog_cycle_task(16'b0100001000110001, 1'b0);
		prog_cycle_task(16'b1100001000110001, 1'b0);
		prog_cycle_task(16'b0010001000110001, 1'b0);
		prog_cycle_task(16'b1010001000110001, 1'b1);
		prog_cycle_task(16'b0001001000110001, 1'b0);
		prog_cycle_task(16'b1001001000110001, 1'b0);
		prog_cycle_task(16'b0000101000110001, 1'b0);
		prog_cycle_task(16'b1000101000110001, 1'b0);
		prog_cycle_task(16'b0000000000001001, 1'b0);
		prog_cycle_task(16'b1000000000001001, 1'b0);
		prog_cycle_task(16'b0100000000001001, 1'b0);
		prog_cycle_task(16'b1100000000001001, 1'b0);
		prog_cycle_task(16'b0010000000001001, 1'b0);
		prog_cycle_task(16'b1010000000001001, 1'b0);
		prog_cycle_task(16'b0110000000001001, 1'b0);
		prog_cycle_task(16'b1110000000001001, 1'b0);
		prog_cycle_task(16'b0001000000001001, 1'b0);
		prog_cycle_task(16'b1001000000001001, 1'b0);
		prog_cycle_task(16'b0101000000001001, 1'b0);
		prog_cycle_task(16'b1101000000001001, 1'b0);
		prog_cycle_task(16'b0011000000001001, 1'b0);
		prog_cycle_task(16'b1011000000001001, 1'b0);
		prog_cycle_task(16'b0111000000001001, 1'b0);
		prog_cycle_task(16'b1111000000001001, 1'b0);
		prog_cycle_task(16'b0000100000001001, 1'b0);
		prog_cycle_task(16'b1000100000001001, 1'b0);
		prog_cycle_task(16'b0100100000001001, 1'b1);
		prog_cycle_task(16'b0000010000001001, 1'b0);
		prog_cycle_task(16'b1000010000001001, 1'b0);
		prog_cycle_task(16'b0100010000001001, 1'b0);
		prog_cycle_task(16'b1100010000001001, 1'b0);
		prog_cycle_task(16'b0010010000001001, 1'b0);
		prog_cycle_task(16'b1010010000001001, 1'b0);
		prog_cycle_task(16'b0110010000001001, 1'b0);
		prog_cycle_task(16'b1110010000001001, 1'b0);
		prog_cycle_task(16'b0001010000001001, 1'b0);
		prog_cycle_task(16'b1001010000001001, 1'b0);
		prog_cycle_task(16'b0101010000001001, 1'b0);
		prog_cycle_task(16'b1101010000001001, 1'b0);
		prog_cycle_task(16'b0011010000001001, 1'b0);
		prog_cycle_task(16'b1011010000001001, 1'b0);
		prog_cycle_task(16'b0111010000001001, 1'b0);
		prog_cycle_task(16'b1111010000001001, 1'b0);
		prog_cycle_task(16'b0000110000001001, 1'b0);
		prog_cycle_task(16'b1000110000001001, 1'b0);
		prog_cycle_task(16'b0100110000001001, 1'b1);
		prog_cycle_task(16'b0000001000001001, 1'b0);
		prog_cycle_task(16'b1000001000001001, 1'b0);
		prog_cycle_task(16'b0100001000001001, 1'b0);
		prog_cycle_task(16'b1100001000001001, 1'b0);
		prog_cycle_task(16'b0010001000001001, 1'b0);
		prog_cycle_task(16'b1010001000001001, 1'b0);
		prog_cycle_task(16'b0110001000001001, 1'b0);
		prog_cycle_task(16'b1110001000001001, 1'b0);
		prog_cycle_task(16'b0001001000001001, 1'b0);
		prog_cycle_task(16'b1001001000001001, 1'b0);
		prog_cycle_task(16'b0101001000001001, 1'b0);
		prog_cycle_task(16'b1101001000001001, 1'b0);
		prog_cycle_task(16'b0011001000001001, 1'b0);
		prog_cycle_task(16'b1011001000001001, 1'b0);
		prog_cycle_task(16'b0111001000001001, 1'b0);
		prog_cycle_task(16'b1111001000001001, 1'b0);
		prog_cycle_task(16'b0000101000001001, 1'b0);
		prog_cycle_task(16'b1000101000001001, 1'b0);
		prog_cycle_task(16'b0100101000001001, 1'b1);
		prog_cycle_task(16'b0000011000001001, 1'b0);
		prog_cycle_task(16'b1000011000001001, 1'b0);
		prog_cycle_task(16'b0100011000001001, 1'b0);
		prog_cycle_task(16'b1100011000001001, 1'b0);
		prog_cycle_task(16'b0010011000001001, 1'b0);
		prog_cycle_task(16'b1010011000001001, 1'b0);
		prog_cycle_task(16'b0110011000001001, 1'b0);
		prog_cycle_task(16'b1110011000001001, 1'b0);
		prog_cycle_task(16'b0001011000001001, 1'b0);
		prog_cycle_task(16'b1001011000001001, 1'b0);
		prog_cycle_task(16'b0101011000001001, 1'b0);
		prog_cycle_task(16'b1101011000001001, 1'b0);
		prog_cycle_task(16'b0011011000001001, 1'b0);
		prog_cycle_task(16'b1011011000001001, 1'b0);
		prog_cycle_task(16'b0111011000001001, 1'b0);
		prog_cycle_task(16'b1111011000001001, 1'b0);
		prog_cycle_task(16'b0000111000001001, 1'b0);
		prog_cycle_task(16'b1000111000001001, 1'b0);
		prog_cycle_task(16'b0100111000001001, 1'b1);
		prog_cycle_task(16'b0000000100001001, 1'b0);
		prog_cycle_task(16'b1000000100001001, 1'b0);
		prog_cycle_task(16'b0100000100001001, 1'b1);
		prog_cycle_task(16'b1100000100001001, 1'b0);
		prog_cycle_task(16'b0010000100001001, 1'b0);
		prog_cycle_task(16'b1010000100001001, 1'b0);
		prog_cycle_task(16'b0110000100001001, 1'b0);
		prog_cycle_task(16'b1110000100001001, 1'b1);
		prog_cycle_task(16'b0000010100001001, 1'b0);
		prog_cycle_task(16'b1000010100001001, 1'b0);
		prog_cycle_task(16'b0100010100001001, 1'b1);
		prog_cycle_task(16'b1100010100001001, 1'b0);
		prog_cycle_task(16'b0010010100001001, 1'b0);
		prog_cycle_task(16'b1010010100001001, 1'b0);
		prog_cycle_task(16'b0110010100001001, 1'b0);
		prog_cycle_task(16'b1110010100001001, 1'b1);
		prog_cycle_task(16'b0000001100001001, 1'b0);
		prog_cycle_task(16'b1000001100001001, 1'b0);
		prog_cycle_task(16'b0100001100001001, 1'b1);
		prog_cycle_task(16'b1100001100001001, 1'b0);
		prog_cycle_task(16'b0010001100001001, 1'b0);
		prog_cycle_task(16'b1010001100001001, 1'b0);
		prog_cycle_task(16'b0110001100001001, 1'b0);
		prog_cycle_task(16'b1110001100001001, 1'b1);
		prog_cycle_task(16'b0000011100001001, 1'b0);
		prog_cycle_task(16'b1000011100001001, 1'b0);
		prog_cycle_task(16'b0100011100001001, 1'b1);
		prog_cycle_task(16'b1100011100001001, 1'b0);
		prog_cycle_task(16'b0010011100001001, 1'b0);
		prog_cycle_task(16'b1010011100001001, 1'b0);
		prog_cycle_task(16'b0110011100001001, 1'b0);
		prog_cycle_task(16'b1110011100001001, 1'b1);
		prog_cycle_task(16'b0000000010001001, 1'b0);
		prog_cycle_task(16'b1000000010001001, 1'b0);
		prog_cycle_task(16'b0100000010001001, 1'b1);
		prog_cycle_task(16'b1100000010001001, 1'b0);
		prog_cycle_task(16'b0010000010001001, 1'b0);
		prog_cycle_task(16'b1010000010001001, 1'b0);
		prog_cycle_task(16'b0110000010001001, 1'b0);
		prog_cycle_task(16'b1110000010001001, 1'b1);
		prog_cycle_task(16'b0000010010001001, 1'b0);
		prog_cycle_task(16'b1000010010001001, 1'b0);
		prog_cycle_task(16'b0100010010001001, 1'b1);
		prog_cycle_task(16'b1100010010001001, 1'b0);
		prog_cycle_task(16'b0010010010001001, 1'b0);
		prog_cycle_task(16'b1010010010001001, 1'b0);
		prog_cycle_task(16'b0110010010001001, 1'b0);
		prog_cycle_task(16'b1110010010001001, 1'b1);
		prog_cycle_task(16'b0000001010001001, 1'b0);
		prog_cycle_task(16'b1000001010001001, 1'b0);
		prog_cycle_task(16'b0100001010001001, 1'b1);
		prog_cycle_task(16'b1100001010001001, 1'b0);
		prog_cycle_task(16'b0010001010001001, 1'b0);
		prog_cycle_task(16'b1010001010001001, 1'b0);
		prog_cycle_task(16'b0110001010001001, 1'b0);
		prog_cycle_task(16'b1110001010001001, 1'b1);
		prog_cycle_task(16'b0000011010001001, 1'b0);
		prog_cycle_task(16'b1000011010001001, 1'b0);
		prog_cycle_task(16'b0100011010001001, 1'b1);
		prog_cycle_task(16'b1100011010001001, 1'b0);
		prog_cycle_task(16'b0010011010001001, 1'b0);
		prog_cycle_task(16'b1010011010001001, 1'b0);
		prog_cycle_task(16'b0110011010001001, 1'b0);
		prog_cycle_task(16'b1110011010001001, 1'b1);
		prog_cycle_task(16'b0000000110001001, 1'b0);
		prog_cycle_task(16'b1000000110001001, 1'b0);
		prog_cycle_task(16'b0100000110001001, 1'b1);
		prog_cycle_task(16'b1100000110001001, 1'b0);
		prog_cycle_task(16'b0010000110001001, 1'b0);
		prog_cycle_task(16'b1010000110001001, 1'b0);
		prog_cycle_task(16'b0110000110001001, 1'b0);
		prog_cycle_task(16'b1110000110001001, 1'b1);
		prog_cycle_task(16'b0000010110001001, 1'b0);
		prog_cycle_task(16'b1000010110001001, 1'b0);
		prog_cycle_task(16'b0100010110001001, 1'b1);
		prog_cycle_task(16'b1100010110001001, 1'b0);
		prog_cycle_task(16'b0010010110001001, 1'b0);
		prog_cycle_task(16'b1010010110001001, 1'b0);
		prog_cycle_task(16'b0110010110001001, 1'b0);
		prog_cycle_task(16'b1110010110001001, 1'b1);
		prog_cycle_task(16'b0000001110001001, 1'b0);
		prog_cycle_task(16'b1000001110001001, 1'b0);
		prog_cycle_task(16'b0100001110001001, 1'b1);
		prog_cycle_task(16'b1100001110001001, 1'b0);
		prog_cycle_task(16'b0010001110001001, 1'b0);
		prog_cycle_task(16'b1010001110001001, 1'b0);
		prog_cycle_task(16'b0110001110001001, 1'b0);
		prog_cycle_task(16'b1110001110001001, 1'b1);
		prog_cycle_task(16'b0000011110001001, 1'b0);
		prog_cycle_task(16'b1000011110001001, 1'b0);
		prog_cycle_task(16'b0100011110001001, 1'b1);
		prog_cycle_task(16'b1100011110001001, 1'b0);
		prog_cycle_task(16'b0010011110001001, 1'b0);
		prog_cycle_task(16'b1010011110001001, 1'b0);
		prog_cycle_task(16'b0110011110001001, 1'b0);
		prog_cycle_task(16'b1110011110001001, 1'b1);
		prog_cycle_task(16'b0000000001001001, 1'b0);
		prog_cycle_task(16'b1000000001001001, 1'b0);
		prog_cycle_task(16'b0100000001001001, 1'b1);
		prog_cycle_task(16'b1100000001001001, 1'b0);
		prog_cycle_task(16'b0010000001001001, 1'b0);
		prog_cycle_task(16'b1010000001001001, 1'b0);
		prog_cycle_task(16'b0110000001001001, 1'b0);
		prog_cycle_task(16'b1110000001001001, 1'b1);
		prog_cycle_task(16'b0000010001001001, 1'b0);
		prog_cycle_task(16'b1000010001001001, 1'b0);
		prog_cycle_task(16'b0100010001001001, 1'b1);
		prog_cycle_task(16'b1100010001001001, 1'b0);
		prog_cycle_task(16'b0010010001001001, 1'b0);
		prog_cycle_task(16'b1010010001001001, 1'b0);
		prog_cycle_task(16'b0110010001001001, 1'b0);
		prog_cycle_task(16'b1110010001001001, 1'b1);
		prog_cycle_task(16'b0000001001001001, 1'b0);
		prog_cycle_task(16'b1000001001001001, 1'b0);
		prog_cycle_task(16'b0100001001001001, 1'b1);
		prog_cycle_task(16'b1100001001001001, 1'b0);
		prog_cycle_task(16'b0010001001001001, 1'b0);
		prog_cycle_task(16'b1010001001001001, 1'b0);
		prog_cycle_task(16'b0110001001001001, 1'b0);
		prog_cycle_task(16'b1110001001001001, 1'b1);
		prog_cycle_task(16'b0000011001001001, 1'b0);
		prog_cycle_task(16'b1000011001001001, 1'b0);
		prog_cycle_task(16'b0100011001001001, 1'b1);
		prog_cycle_task(16'b1100011001001001, 1'b0);
		prog_cycle_task(16'b0010011001001001, 1'b0);
		prog_cycle_task(16'b1010011001001001, 1'b0);
		prog_cycle_task(16'b0110011001001001, 1'b0);
		prog_cycle_task(16'b1110011001001001, 1'b1);
		prog_cycle_task(16'b0000000000101001, 1'b0);
		prog_cycle_task(16'b1000000000101001, 1'b0);
		prog_cycle_task(16'b0100000000101001, 1'b1);
		prog_cycle_task(16'b1100000000101001, 1'b0);
		prog_cycle_task(16'b0010000000101001, 1'b0);
		prog_cycle_task(16'b1010000000101001, 1'b1);
		prog_cycle_task(16'b0001000000101001, 1'b0);
		prog_cycle_task(16'b1001000000101001, 1'b0);
		prog_cycle_task(16'b0101000000101001, 1'b1);
		prog_cycle_task(16'b1101000000101001, 1'b0);
		prog_cycle_task(16'b0011000000101001, 1'b0);
		prog_cycle_task(16'b1011000000101001, 1'b1);
		prog_cycle_task(16'b0000100000101001, 1'b0);
		prog_cycle_task(16'b1000100000101001, 1'b0);
		prog_cycle_task(16'b0100100000101001, 1'b1);
		prog_cycle_task(16'b1100100000101001, 1'b0);
		prog_cycle_task(16'b0010100000101001, 1'b0);
		prog_cycle_task(16'b1010100000101001, 1'b1);
		prog_cycle_task(16'b0001100000101001, 1'b0);
		prog_cycle_task(16'b1001100000101001, 1'b0);
		prog_cycle_task(16'b0101100000101001, 1'b1);
		prog_cycle_task(16'b1101100000101001, 1'b0);
		prog_cycle_task(16'b0011100000101001, 1'b0);
		prog_cycle_task(16'b1011100000101001, 1'b1);
		prog_cycle_task(16'b0000010000101001, 1'b0);
		prog_cycle_task(16'b1000010000101001, 1'b0);
		prog_cycle_task(16'b0100010000101001, 1'b1);
		prog_cycle_task(16'b1100010000101001, 1'b0);
		prog_cycle_task(16'b0010010000101001, 1'b0);
		prog_cycle_task(16'b1010010000101001, 1'b1);
		prog_cycle_task(16'b0001010000101001, 1'b0);
		prog_cycle_task(16'b1001010000101001, 1'b0);
		prog_cycle_task(16'b0101010000101001, 1'b1);
		prog_cycle_task(16'b1101010000101001, 1'b0);
		prog_cycle_task(16'b0011010000101001, 1'b0);
		prog_cycle_task(16'b1011010000101001, 1'b1);
		prog_cycle_task(16'b0000110000101001, 1'b0);
		prog_cycle_task(16'b1000110000101001, 1'b0);
		prog_cycle_task(16'b0001110000101001, 1'b0);
		prog_cycle_task(16'b1001110000101001, 1'b0);
		prog_cycle_task(16'b0000001000101001, 1'b0);
		prog_cycle_task(16'b1000001000101001, 1'b0);
		prog_cycle_task(16'b0001001000101001, 1'b0);
		prog_cycle_task(16'b1001001000101001, 1'b0);
		prog_cycle_task(16'b0000101000101001, 1'b0);
		prog_cycle_task(16'b1000101000101001, 1'b0);
		prog_cycle_task(16'b0001101000101001, 1'b0);
		prog_cycle_task(16'b1001101000101001, 1'b0);
		prog_cycle_task(16'b0000011000101001, 1'b0);
		prog_cycle_task(16'b1000011000101001, 1'b0);
		prog_cycle_task(16'b0001011000101001, 1'b0);
		prog_cycle_task(16'b1001011000101001, 1'b0);
		prog_cycle_task(16'b0000111000101001, 1'b0);
		prog_cycle_task(16'b1000111000101001, 1'b0);
		prog_cycle_task(16'b0000000000011001, 1'b0);
		prog_cycle_task(16'b1000000000011001, 1'b0);
		prog_cycle_task(16'b0100000000011001, 1'b0);
		prog_cycle_task(16'b1100000000011001, 1'b0);
		prog_cycle_task(16'b0010000000011001, 1'b0);
		prog_cycle_task(16'b1010000000011001, 1'b1);
		prog_cycle_task(16'b0001000000011001, 1'b0);
		prog_cycle_task(16'b1001000000011001, 1'b0);
		prog_cycle_task(16'b0000100000011001, 1'b0);
		prog_cycle_task(16'b1000100000011001, 1'b0);
		prog_cycle_task(16'b0100100000011001, 1'b0);
		prog_cycle_task(16'b1100100000011001, 1'b0);
		prog_cycle_task(16'b0010100000011001, 1'b0);
		prog_cycle_task(16'b1010100000011001, 1'b1);
		prog_cycle_task(16'b0001100000011001, 1'b0);
		prog_cycle_task(16'b1001100000011001, 1'b0);
		prog_cycle_task(16'b0101100000011001, 1'b0);
		prog_cycle_task(16'b1101100000011001, 1'b0);
		prog_cycle_task(16'b0011100000011001, 1'b0);
		prog_cycle_task(16'b1011100000011001, 1'b1);
		prog_cycle_task(16'b0000010000011001, 1'b0);
		prog_cycle_task(16'b1000010000011001, 1'b0);
		prog_cycle_task(16'b0001010000011001, 1'b0);
		prog_cycle_task(16'b1001010000011001, 1'b0);
		prog_cycle_task(16'b0000000000111001, 1'b0);
		prog_cycle_task(16'b1000000000111001, 1'b0);
		prog_cycle_task(16'b0100000000111001, 1'b0);
		prog_cycle_task(16'b1100000000111001, 1'b0);
		prog_cycle_task(16'b0010000000111001, 1'b0);
		prog_cycle_task(16'b1010000000111001, 1'b1);
		prog_cycle_task(16'b0001000000111001, 1'b0);
		prog_cycle_task(16'b1001000000111001, 1'b0);
		prog_cycle_task(16'b0101000000111001, 1'b0);
		prog_cycle_task(16'b1101000000111001, 1'b0);
		prog_cycle_task(16'b0011000000111001, 1'b0);
		prog_cycle_task(16'b1011000000111001, 1'b1);
		prog_cycle_task(16'b0000100000111001, 1'b0);
		prog_cycle_task(16'b1000100000111001, 1'b0);
		prog_cycle_task(16'b0100100000111001, 1'b0);
		prog_cycle_task(16'b1100100000111001, 1'b0);
		prog_cycle_task(16'b0010100000111001, 1'b0);
		prog_cycle_task(16'b1010100000111001, 1'b1);
		prog_cycle_task(16'b0001100000111001, 1'b0);
		prog_cycle_task(16'b1001100000111001, 1'b0);
		prog_cycle_task(16'b0101100000111001, 1'b0);
		prog_cycle_task(16'b1101100000111001, 1'b0);
		prog_cycle_task(16'b0011100000111001, 1'b0);
		prog_cycle_task(16'b1011100000111001, 1'b1);
		prog_cycle_task(16'b0000010000111001, 1'b0);
		prog_cycle_task(16'b1000010000111001, 1'b0);
		prog_cycle_task(16'b0100010000111001, 1'b0);
		prog_cycle_task(16'b1100010000111001, 1'b0);
		prog_cycle_task(16'b0010010000111001, 1'b0);
		prog_cycle_task(16'b1010010000111001, 1'b1);
		prog_cycle_task(16'b0001010000111001, 1'b0);
		prog_cycle_task(16'b1001010000111001, 1'b0);
		prog_cycle_task(16'b0101010000111001, 1'b0);
		prog_cycle_task(16'b1101010000111001, 1'b0);
		prog_cycle_task(16'b0011010000111001, 1'b0);
		prog_cycle_task(16'b1011010000111001, 1'b1);
		prog_cycle_task(16'b0000110000111001, 1'b0);
		prog_cycle_task(16'b1000110000111001, 1'b0);
		prog_cycle_task(16'b0100110000111001, 1'b0);
		prog_cycle_task(16'b1100110000111001, 1'b0);
		prog_cycle_task(16'b0010110000111001, 1'b0);
		prog_cycle_task(16'b1010110000111001, 1'b1);
		prog_cycle_task(16'b0001110000111001, 1'b0);
		prog_cycle_task(16'b1001110000111001, 1'b0);
		prog_cycle_task(16'b0101110000111001, 1'b0);
		prog_cycle_task(16'b1101110000111001, 1'b0);
		prog_cycle_task(16'b0011110000111001, 1'b0);
		prog_cycle_task(16'b1011110000111001, 1'b1);
		prog_cycle_task(16'b0000001000111001, 1'b0);
		prog_cycle_task(16'b1000001000111001, 1'b0);
		prog_cycle_task(16'b0100001000111001, 1'b0);
		prog_cycle_task(16'b1100001000111001, 1'b0);
		prog_cycle_task(16'b0010001000111001, 1'b0);
		prog_cycle_task(16'b1010001000111001, 1'b1);
		prog_cycle_task(16'b0001001000111001, 1'b0);
		prog_cycle_task(16'b1001001000111001, 1'b0);
		prog_cycle_task(16'b0000101000111001, 1'b0);
		prog_cycle_task(16'b1000101000111001, 1'b0);
		prog_cycle_task(16'b0000000000000101, 1'b0);
		prog_cycle_task(16'b1000000000000101, 1'b0);
		prog_cycle_task(16'b0100000000000101, 1'b0);
		prog_cycle_task(16'b1100000000000101, 1'b0);
		prog_cycle_task(16'b0010000000000101, 1'b0);
		prog_cycle_task(16'b1010000000000101, 1'b0);
		prog_cycle_task(16'b0110000000000101, 1'b0);
		prog_cycle_task(16'b1110000000000101, 1'b0);
		prog_cycle_task(16'b0001000000000101, 1'b0);
		prog_cycle_task(16'b1001000000000101, 1'b0);
		prog_cycle_task(16'b0101000000000101, 1'b0);
		prog_cycle_task(16'b1101000000000101, 1'b0);
		prog_cycle_task(16'b0011000000000101, 1'b0);
		prog_cycle_task(16'b1011000000000101, 1'b0);
		prog_cycle_task(16'b0111000000000101, 1'b0);
		prog_cycle_task(16'b1111000000000101, 1'b0);
		prog_cycle_task(16'b0000100000000101, 1'b0);
		prog_cycle_task(16'b1000100000000101, 1'b0);
		prog_cycle_task(16'b0100100000000101, 1'b1);
		prog_cycle_task(16'b0000010000000101, 1'b0);
		prog_cycle_task(16'b1000010000000101, 1'b0);
		prog_cycle_task(16'b0100010000000101, 1'b0);
		prog_cycle_task(16'b1100010000000101, 1'b0);
		prog_cycle_task(16'b0010010000000101, 1'b0);
		prog_cycle_task(16'b1010010000000101, 1'b0);
		prog_cycle_task(16'b0110010000000101, 1'b0);
		prog_cycle_task(16'b1110010000000101, 1'b0);
		prog_cycle_task(16'b0001010000000101, 1'b0);
		prog_cycle_task(16'b1001010000000101, 1'b0);
		prog_cycle_task(16'b0101010000000101, 1'b0);
		prog_cycle_task(16'b1101010000000101, 1'b0);
		prog_cycle_task(16'b0011010000000101, 1'b0);
		prog_cycle_task(16'b1011010000000101, 1'b0);
		prog_cycle_task(16'b0111010000000101, 1'b0);
		prog_cycle_task(16'b1111010000000101, 1'b0);
		prog_cycle_task(16'b0000110000000101, 1'b0);
		prog_cycle_task(16'b1000110000000101, 1'b0);
		prog_cycle_task(16'b0100110000000101, 1'b1);
		prog_cycle_task(16'b0000001000000101, 1'b0);
		prog_cycle_task(16'b1000001000000101, 1'b0);
		prog_cycle_task(16'b0100001000000101, 1'b0);
		prog_cycle_task(16'b1100001000000101, 1'b0);
		prog_cycle_task(16'b0010001000000101, 1'b0);
		prog_cycle_task(16'b1010001000000101, 1'b0);
		prog_cycle_task(16'b0110001000000101, 1'b0);
		prog_cycle_task(16'b1110001000000101, 1'b0);
		prog_cycle_task(16'b0001001000000101, 1'b0);
		prog_cycle_task(16'b1001001000000101, 1'b0);
		prog_cycle_task(16'b0101001000000101, 1'b0);
		prog_cycle_task(16'b1101001000000101, 1'b0);
		prog_cycle_task(16'b0011001000000101, 1'b0);
		prog_cycle_task(16'b1011001000000101, 1'b0);
		prog_cycle_task(16'b0111001000000101, 1'b0);
		prog_cycle_task(16'b1111001000000101, 1'b0);
		prog_cycle_task(16'b0000101000000101, 1'b0);
		prog_cycle_task(16'b1000101000000101, 1'b0);
		prog_cycle_task(16'b0100101000000101, 1'b1);
		prog_cycle_task(16'b0000011000000101, 1'b0);
		prog_cycle_task(16'b1000011000000101, 1'b0);
		prog_cycle_task(16'b0100011000000101, 1'b0);
		prog_cycle_task(16'b1100011000000101, 1'b0);
		prog_cycle_task(16'b0010011000000101, 1'b0);
		prog_cycle_task(16'b1010011000000101, 1'b0);
		prog_cycle_task(16'b0110011000000101, 1'b0);
		prog_cycle_task(16'b1110011000000101, 1'b0);
		prog_cycle_task(16'b0001011000000101, 1'b0);
		prog_cycle_task(16'b1001011000000101, 1'b0);
		prog_cycle_task(16'b0101011000000101, 1'b0);
		prog_cycle_task(16'b1101011000000101, 1'b0);
		prog_cycle_task(16'b0011011000000101, 1'b0);
		prog_cycle_task(16'b1011011000000101, 1'b0);
		prog_cycle_task(16'b0111011000000101, 1'b0);
		prog_cycle_task(16'b1111011000000101, 1'b0);
		prog_cycle_task(16'b0000111000000101, 1'b0);
		prog_cycle_task(16'b1000111000000101, 1'b0);
		prog_cycle_task(16'b0100111000000101, 1'b1);
		prog_cycle_task(16'b0000000100000101, 1'b0);
		prog_cycle_task(16'b1000000100000101, 1'b0);
		prog_cycle_task(16'b0100000100000101, 1'b1);
		prog_cycle_task(16'b1100000100000101, 1'b0);
		prog_cycle_task(16'b0010000100000101, 1'b0);
		prog_cycle_task(16'b1010000100000101, 1'b0);
		prog_cycle_task(16'b0110000100000101, 1'b0);
		prog_cycle_task(16'b1110000100000101, 1'b1);
		prog_cycle_task(16'b0000010100000101, 1'b0);
		prog_cycle_task(16'b1000010100000101, 1'b0);
		prog_cycle_task(16'b0100010100000101, 1'b1);
		prog_cycle_task(16'b1100010100000101, 1'b0);
		prog_cycle_task(16'b0010010100000101, 1'b0);
		prog_cycle_task(16'b1010010100000101, 1'b0);
		prog_cycle_task(16'b0110010100000101, 1'b0);
		prog_cycle_task(16'b1110010100000101, 1'b1);
		prog_cycle_task(16'b0000001100000101, 1'b0);
		prog_cycle_task(16'b1000001100000101, 1'b0);
		prog_cycle_task(16'b0100001100000101, 1'b1);
		prog_cycle_task(16'b1100001100000101, 1'b0);
		prog_cycle_task(16'b0010001100000101, 1'b0);
		prog_cycle_task(16'b1010001100000101, 1'b0);
		prog_cycle_task(16'b0110001100000101, 1'b0);
		prog_cycle_task(16'b1110001100000101, 1'b1);
		prog_cycle_task(16'b0000011100000101, 1'b0);
		prog_cycle_task(16'b1000011100000101, 1'b0);
		prog_cycle_task(16'b0100011100000101, 1'b1);
		prog_cycle_task(16'b1100011100000101, 1'b0);
		prog_cycle_task(16'b0010011100000101, 1'b0);
		prog_cycle_task(16'b1010011100000101, 1'b0);
		prog_cycle_task(16'b0110011100000101, 1'b0);
		prog_cycle_task(16'b1110011100000101, 1'b1);
		prog_cycle_task(16'b0000000010000101, 1'b0);
		prog_cycle_task(16'b1000000010000101, 1'b0);
		prog_cycle_task(16'b0100000010000101, 1'b1);
		prog_cycle_task(16'b1100000010000101, 1'b0);
		prog_cycle_task(16'b0010000010000101, 1'b0);
		prog_cycle_task(16'b1010000010000101, 1'b0);
		prog_cycle_task(16'b0110000010000101, 1'b0);
		prog_cycle_task(16'b1110000010000101, 1'b1);
		prog_cycle_task(16'b0000010010000101, 1'b0);
		prog_cycle_task(16'b1000010010000101, 1'b0);
		prog_cycle_task(16'b0100010010000101, 1'b1);
		prog_cycle_task(16'b1100010010000101, 1'b0);
		prog_cycle_task(16'b0010010010000101, 1'b0);
		prog_cycle_task(16'b1010010010000101, 1'b0);
		prog_cycle_task(16'b0110010010000101, 1'b0);
		prog_cycle_task(16'b1110010010000101, 1'b1);
		prog_cycle_task(16'b0000001010000101, 1'b0);
		prog_cycle_task(16'b1000001010000101, 1'b0);
		prog_cycle_task(16'b0100001010000101, 1'b1);
		prog_cycle_task(16'b1100001010000101, 1'b0);
		prog_cycle_task(16'b0010001010000101, 1'b0);
		prog_cycle_task(16'b1010001010000101, 1'b0);
		prog_cycle_task(16'b0110001010000101, 1'b0);
		prog_cycle_task(16'b1110001010000101, 1'b1);
		prog_cycle_task(16'b0000011010000101, 1'b0);
		prog_cycle_task(16'b1000011010000101, 1'b0);
		prog_cycle_task(16'b0100011010000101, 1'b1);
		prog_cycle_task(16'b1100011010000101, 1'b0);
		prog_cycle_task(16'b0010011010000101, 1'b0);
		prog_cycle_task(16'b1010011010000101, 1'b0);
		prog_cycle_task(16'b0110011010000101, 1'b0);
		prog_cycle_task(16'b1110011010000101, 1'b1);
		prog_cycle_task(16'b0000000110000101, 1'b0);
		prog_cycle_task(16'b1000000110000101, 1'b0);
		prog_cycle_task(16'b0100000110000101, 1'b1);
		prog_cycle_task(16'b1100000110000101, 1'b0);
		prog_cycle_task(16'b0010000110000101, 1'b0);
		prog_cycle_task(16'b1010000110000101, 1'b0);
		prog_cycle_task(16'b0110000110000101, 1'b0);
		prog_cycle_task(16'b1110000110000101, 1'b1);
		prog_cycle_task(16'b0000010110000101, 1'b0);
		prog_cycle_task(16'b1000010110000101, 1'b0);
		prog_cycle_task(16'b0100010110000101, 1'b1);
		prog_cycle_task(16'b1100010110000101, 1'b0);
		prog_cycle_task(16'b0010010110000101, 1'b0);
		prog_cycle_task(16'b1010010110000101, 1'b0);
		prog_cycle_task(16'b0110010110000101, 1'b0);
		prog_cycle_task(16'b1110010110000101, 1'b1);
		prog_cycle_task(16'b0000001110000101, 1'b0);
		prog_cycle_task(16'b1000001110000101, 1'b0);
		prog_cycle_task(16'b0100001110000101, 1'b1);
		prog_cycle_task(16'b1100001110000101, 1'b0);
		prog_cycle_task(16'b0010001110000101, 1'b0);
		prog_cycle_task(16'b1010001110000101, 1'b0);
		prog_cycle_task(16'b0110001110000101, 1'b0);
		prog_cycle_task(16'b1110001110000101, 1'b1);
		prog_cycle_task(16'b0000011110000101, 1'b0);
		prog_cycle_task(16'b1000011110000101, 1'b0);
		prog_cycle_task(16'b0100011110000101, 1'b1);
		prog_cycle_task(16'b1100011110000101, 1'b0);
		prog_cycle_task(16'b0010011110000101, 1'b0);
		prog_cycle_task(16'b1010011110000101, 1'b0);
		prog_cycle_task(16'b0110011110000101, 1'b0);
		prog_cycle_task(16'b1110011110000101, 1'b1);
		prog_cycle_task(16'b0000000001000101, 1'b0);
		prog_cycle_task(16'b1000000001000101, 1'b0);
		prog_cycle_task(16'b0100000001000101, 1'b1);
		prog_cycle_task(16'b1100000001000101, 1'b0);
		prog_cycle_task(16'b0010000001000101, 1'b0);
		prog_cycle_task(16'b1010000001000101, 1'b0);
		prog_cycle_task(16'b0110000001000101, 1'b0);
		prog_cycle_task(16'b1110000001000101, 1'b1);
		prog_cycle_task(16'b0000010001000101, 1'b0);
		prog_cycle_task(16'b1000010001000101, 1'b0);
		prog_cycle_task(16'b0100010001000101, 1'b1);
		prog_cycle_task(16'b1100010001000101, 1'b0);
		prog_cycle_task(16'b0010010001000101, 1'b0);
		prog_cycle_task(16'b1010010001000101, 1'b0);
		prog_cycle_task(16'b0110010001000101, 1'b0);
		prog_cycle_task(16'b1110010001000101, 1'b1);
		prog_cycle_task(16'b0000001001000101, 1'b0);
		prog_cycle_task(16'b1000001001000101, 1'b0);
		prog_cycle_task(16'b0100001001000101, 1'b1);
		prog_cycle_task(16'b1100001001000101, 1'b0);
		prog_cycle_task(16'b0010001001000101, 1'b0);
		prog_cycle_task(16'b1010001001000101, 1'b0);
		prog_cycle_task(16'b0110001001000101, 1'b0);
		prog_cycle_task(16'b1110001001000101, 1'b1);
		prog_cycle_task(16'b0000011001000101, 1'b0);
		prog_cycle_task(16'b1000011001000101, 1'b0);
		prog_cycle_task(16'b0100011001000101, 1'b1);
		prog_cycle_task(16'b1100011001000101, 1'b0);
		prog_cycle_task(16'b0010011001000101, 1'b0);
		prog_cycle_task(16'b1010011001000101, 1'b0);
		prog_cycle_task(16'b0110011001000101, 1'b0);
		prog_cycle_task(16'b1110011001000101, 1'b1);
		prog_cycle_task(16'b0000000000100101, 1'b0);
		prog_cycle_task(16'b1000000000100101, 1'b0);
		prog_cycle_task(16'b0100000000100101, 1'b0);
		prog_cycle_task(16'b1100000000100101, 1'b0);
		prog_cycle_task(16'b0010000000100101, 1'b0);
		prog_cycle_task(16'b1010000000100101, 1'b0);
		prog_cycle_task(16'b0110000000100101, 1'b0);
		prog_cycle_task(16'b1110000000100101, 1'b1);
		prog_cycle_task(16'b0001000000100101, 1'b0);
		prog_cycle_task(16'b1001000000100101, 1'b0);
		prog_cycle_task(16'b0101000000100101, 1'b0);
		prog_cycle_task(16'b1101000000100101, 1'b0);
		prog_cycle_task(16'b0011000000100101, 1'b0);
		prog_cycle_task(16'b1011000000100101, 1'b0);
		prog_cycle_task(16'b0111000000100101, 1'b0);
		prog_cycle_task(16'b1111000000100101, 1'b1);
		prog_cycle_task(16'b0000100000100101, 1'b0);
		prog_cycle_task(16'b1000100000100101, 1'b0);
		prog_cycle_task(16'b0100100000100101, 1'b1);
		prog_cycle_task(16'b1100100000100101, 1'b0);
		prog_cycle_task(16'b0010100000100101, 1'b0);
		prog_cycle_task(16'b1010100000100101, 1'b1);
		prog_cycle_task(16'b0001100000100101, 1'b0);
		prog_cycle_task(16'b1001100000100101, 1'b0);
		prog_cycle_task(16'b0101100000100101, 1'b0);
		prog_cycle_task(16'b1101100000100101, 1'b0);
		prog_cycle_task(16'b0011100000100101, 1'b0);
		prog_cycle_task(16'b1011100000100101, 1'b0);
		prog_cycle_task(16'b0111100000100101, 1'b0);
		prog_cycle_task(16'b1111100000100101, 1'b1);
		prog_cycle_task(16'b0000010000100101, 1'b0);
		prog_cycle_task(16'b1000010000100101, 1'b0);
		prog_cycle_task(16'b0100010000100101, 1'b0);
		prog_cycle_task(16'b1100010000100101, 1'b0);
		prog_cycle_task(16'b0010010000100101, 1'b0);
		prog_cycle_task(16'b1010010000100101, 1'b0);
		prog_cycle_task(16'b0110010000100101, 1'b0);
		prog_cycle_task(16'b1110010000100101, 1'b1);
		prog_cycle_task(16'b0001010000100101, 1'b0);
		prog_cycle_task(16'b1001010000100101, 1'b0);
		prog_cycle_task(16'b0101010000100101, 1'b1);
		prog_cycle_task(16'b1101010000100101, 1'b0);
		prog_cycle_task(16'b0011010000100101, 1'b0);
		prog_cycle_task(16'b1011010000100101, 1'b1);
		prog_cycle_task(16'b0000110000100101, 1'b0);
		prog_cycle_task(16'b1000110000100101, 1'b0);
		prog_cycle_task(16'b0100110000100101, 1'b0);
		prog_cycle_task(16'b1100110000100101, 1'b0);
		prog_cycle_task(16'b0010110000100101, 1'b0);
		prog_cycle_task(16'b1010110000100101, 1'b0);
		prog_cycle_task(16'b0110110000100101, 1'b0);
		prog_cycle_task(16'b1110110000100101, 1'b1);
		prog_cycle_task(16'b0001110000100101, 1'b0);
		prog_cycle_task(16'b1001110000100101, 1'b0);
		prog_cycle_task(16'b0101110000100101, 1'b0);
		prog_cycle_task(16'b1101110000100101, 1'b0);
		prog_cycle_task(16'b0011110000100101, 1'b0);
		prog_cycle_task(16'b1011110000100101, 1'b0);
		prog_cycle_task(16'b0111110000100101, 1'b0);
		prog_cycle_task(16'b1111110000100101, 1'b1);
		prog_cycle_task(16'b0000001000100101, 1'b0);
		prog_cycle_task(16'b1000001000100101, 1'b0);
		prog_cycle_task(16'b0100001000100101, 1'b1);
		prog_cycle_task(16'b1100001000100101, 1'b0);
		prog_cycle_task(16'b0010001000100101, 1'b0);
		prog_cycle_task(16'b1010001000100101, 1'b1);
		prog_cycle_task(16'b0001001000100101, 1'b0);
		prog_cycle_task(16'b1001001000100101, 1'b0);
		prog_cycle_task(16'b0101001000100101, 1'b0);
		prog_cycle_task(16'b1101001000100101, 1'b0);
		prog_cycle_task(16'b0011001000100101, 1'b0);
		prog_cycle_task(16'b1011001000100101, 1'b0);
		prog_cycle_task(16'b0111001000100101, 1'b0);
		prog_cycle_task(16'b1111001000100101, 1'b1);
		prog_cycle_task(16'b0000101000100101, 1'b0);
		prog_cycle_task(16'b1000101000100101, 1'b0);
		prog_cycle_task(16'b0100101000100101, 1'b0);
		prog_cycle_task(16'b1100101000100101, 1'b0);
		prog_cycle_task(16'b0010101000100101, 1'b0);
		prog_cycle_task(16'b1010101000100101, 1'b0);
		prog_cycle_task(16'b0110101000100101, 1'b0);
		prog_cycle_task(16'b1110101000100101, 1'b1);
		prog_cycle_task(16'b0001101000100101, 1'b0);
		prog_cycle_task(16'b1001101000100101, 1'b0);
		prog_cycle_task(16'b0101101000100101, 1'b1);
		prog_cycle_task(16'b1101101000100101, 1'b0);
		prog_cycle_task(16'b0011101000100101, 1'b0);
		prog_cycle_task(16'b1011101000100101, 1'b1);
		prog_cycle_task(16'b0000000000010101, 1'b0);
		prog_cycle_task(16'b1000000000010101, 1'b0);
		prog_cycle_task(16'b0100000000010101, 1'b0);
		prog_cycle_task(16'b1100000000010101, 1'b0);
		prog_cycle_task(16'b0010000000010101, 1'b0);
		prog_cycle_task(16'b1010000000010101, 1'b1);
		prog_cycle_task(16'b0001000000010101, 1'b0);
		prog_cycle_task(16'b1001000000010101, 1'b0);
		prog_cycle_task(16'b0000100000010101, 1'b0);
		prog_cycle_task(16'b1000100000010101, 1'b0);
		prog_cycle_task(16'b0100100000010101, 1'b0);
		prog_cycle_task(16'b1100100000010101, 1'b0);
		prog_cycle_task(16'b0010100000010101, 1'b0);
		prog_cycle_task(16'b1010100000010101, 1'b1);
		prog_cycle_task(16'b0001100000010101, 1'b0);
		prog_cycle_task(16'b1001100000010101, 1'b0);
		prog_cycle_task(16'b0101100000010101, 1'b0);
		prog_cycle_task(16'b1101100000010101, 1'b0);
		prog_cycle_task(16'b0011100000010101, 1'b0);
		prog_cycle_task(16'b1011100000010101, 1'b1);
		prog_cycle_task(16'b0000010000010101, 1'b0);
		prog_cycle_task(16'b1000010000010101, 1'b0);
		prog_cycle_task(16'b0001010000010101, 1'b0);
		prog_cycle_task(16'b1001010000010101, 1'b0);
		prog_cycle_task(16'b0000000000110101, 1'b0);
		prog_cycle_task(16'b1000000000110101, 1'b0);
		prog_cycle_task(16'b0100000000110101, 1'b0);
		prog_cycle_task(16'b1100000000110101, 1'b0);
		prog_cycle_task(16'b0010000000110101, 1'b0);
		prog_cycle_task(16'b1010000000110101, 1'b1);
		prog_cycle_task(16'b0001000000110101, 1'b0);
		prog_cycle_task(16'b1001000000110101, 1'b0);
		prog_cycle_task(16'b0000100000110101, 1'b0);
		prog_cycle_task(16'b1000100000110101, 1'b0);
		prog_cycle_task(16'b0100100000110101, 1'b0);
		prog_cycle_task(16'b1100100000110101, 1'b0);
		prog_cycle_task(16'b0010100000110101, 1'b0);
		prog_cycle_task(16'b1010100000110101, 1'b1);
		prog_cycle_task(16'b0001100000110101, 1'b0);
		prog_cycle_task(16'b1001100000110101, 1'b0);
		prog_cycle_task(16'b0000010000110101, 1'b0);
		prog_cycle_task(16'b1000010000110101, 1'b0);
		prog_cycle_task(16'b0000000000001101, 1'b0);
		prog_cycle_task(16'b1000000000001101, 1'b0);
		prog_cycle_task(16'b0100000000001101, 1'b0);
		prog_cycle_task(16'b1100000000001101, 1'b0);
		prog_cycle_task(16'b0010000000001101, 1'b0);
		prog_cycle_task(16'b1010000000001101, 1'b0);
		prog_cycle_task(16'b0110000000001101, 1'b0);
		prog_cycle_task(16'b1110000000001101, 1'b0);
		prog_cycle_task(16'b0001000000001101, 1'b0);
		prog_cycle_task(16'b1001000000001101, 1'b0);
		prog_cycle_task(16'b0101000000001101, 1'b0);
		prog_cycle_task(16'b1101000000001101, 1'b0);
		prog_cycle_task(16'b0011000000001101, 1'b0);
		prog_cycle_task(16'b1011000000001101, 1'b0);
		prog_cycle_task(16'b0111000000001101, 1'b0);
		prog_cycle_task(16'b1111000000001101, 1'b0);
		prog_cycle_task(16'b0000100000001101, 1'b0);
		prog_cycle_task(16'b1000100000001101, 1'b0);
		prog_cycle_task(16'b0100100000001101, 1'b1);
		prog_cycle_task(16'b0000010000001101, 1'b0);
		prog_cycle_task(16'b1000010000001101, 1'b0);
		prog_cycle_task(16'b0100010000001101, 1'b0);
		prog_cycle_task(16'b1100010000001101, 1'b0);
		prog_cycle_task(16'b0010010000001101, 1'b0);
		prog_cycle_task(16'b1010010000001101, 1'b0);
		prog_cycle_task(16'b0110010000001101, 1'b0);
		prog_cycle_task(16'b1110010000001101, 1'b0);
		prog_cycle_task(16'b0001010000001101, 1'b0);
		prog_cycle_task(16'b1001010000001101, 1'b0);
		prog_cycle_task(16'b0101010000001101, 1'b0);
		prog_cycle_task(16'b1101010000001101, 1'b0);
		prog_cycle_task(16'b0011010000001101, 1'b0);
		prog_cycle_task(16'b1011010000001101, 1'b0);
		prog_cycle_task(16'b0111010000001101, 1'b0);
		prog_cycle_task(16'b1111010000001101, 1'b0);
		prog_cycle_task(16'b0000110000001101, 1'b0);
		prog_cycle_task(16'b1000110000001101, 1'b0);
		prog_cycle_task(16'b0100110000001101, 1'b1);
		prog_cycle_task(16'b0000001000001101, 1'b0);
		prog_cycle_task(16'b1000001000001101, 1'b0);
		prog_cycle_task(16'b0100001000001101, 1'b0);
		prog_cycle_task(16'b1100001000001101, 1'b0);
		prog_cycle_task(16'b0010001000001101, 1'b0);
		prog_cycle_task(16'b1010001000001101, 1'b0);
		prog_cycle_task(16'b0110001000001101, 1'b0);
		prog_cycle_task(16'b1110001000001101, 1'b0);
		prog_cycle_task(16'b0001001000001101, 1'b0);
		prog_cycle_task(16'b1001001000001101, 1'b0);
		prog_cycle_task(16'b0101001000001101, 1'b0);
		prog_cycle_task(16'b1101001000001101, 1'b0);
		prog_cycle_task(16'b0011001000001101, 1'b0);
		prog_cycle_task(16'b1011001000001101, 1'b0);
		prog_cycle_task(16'b0111001000001101, 1'b0);
		prog_cycle_task(16'b1111001000001101, 1'b0);
		prog_cycle_task(16'b0000101000001101, 1'b0);
		prog_cycle_task(16'b1000101000001101, 1'b0);
		prog_cycle_task(16'b0100101000001101, 1'b1);
		prog_cycle_task(16'b0000011000001101, 1'b0);
		prog_cycle_task(16'b1000011000001101, 1'b0);
		prog_cycle_task(16'b0100011000001101, 1'b0);
		prog_cycle_task(16'b1100011000001101, 1'b0);
		prog_cycle_task(16'b0010011000001101, 1'b0);
		prog_cycle_task(16'b1010011000001101, 1'b0);
		prog_cycle_task(16'b0110011000001101, 1'b0);
		prog_cycle_task(16'b1110011000001101, 1'b0);
		prog_cycle_task(16'b0001011000001101, 1'b0);
		prog_cycle_task(16'b1001011000001101, 1'b0);
		prog_cycle_task(16'b0101011000001101, 1'b0);
		prog_cycle_task(16'b1101011000001101, 1'b0);
		prog_cycle_task(16'b0011011000001101, 1'b0);
		prog_cycle_task(16'b1011011000001101, 1'b0);
		prog_cycle_task(16'b0111011000001101, 1'b0);
		prog_cycle_task(16'b1111011000001101, 1'b0);
		prog_cycle_task(16'b0000111000001101, 1'b0);
		prog_cycle_task(16'b1000111000001101, 1'b0);
		prog_cycle_task(16'b0100111000001101, 1'b1);
		prog_cycle_task(16'b0000000100001101, 1'b0);
		prog_cycle_task(16'b1000000100001101, 1'b0);
		prog_cycle_task(16'b0100000100001101, 1'b1);
		prog_cycle_task(16'b1100000100001101, 1'b0);
		prog_cycle_task(16'b0010000100001101, 1'b0);
		prog_cycle_task(16'b1010000100001101, 1'b0);
		prog_cycle_task(16'b0110000100001101, 1'b0);
		prog_cycle_task(16'b1110000100001101, 1'b1);
		prog_cycle_task(16'b0000010100001101, 1'b0);
		prog_cycle_task(16'b1000010100001101, 1'b0);
		prog_cycle_task(16'b0100010100001101, 1'b1);
		prog_cycle_task(16'b1100010100001101, 1'b0);
		prog_cycle_task(16'b0010010100001101, 1'b0);
		prog_cycle_task(16'b1010010100001101, 1'b0);
		prog_cycle_task(16'b0110010100001101, 1'b0);
		prog_cycle_task(16'b1110010100001101, 1'b1);
		prog_cycle_task(16'b0000001100001101, 1'b0);
		prog_cycle_task(16'b1000001100001101, 1'b0);
		prog_cycle_task(16'b0100001100001101, 1'b1);
		prog_cycle_task(16'b1100001100001101, 1'b0);
		prog_cycle_task(16'b0010001100001101, 1'b0);
		prog_cycle_task(16'b1010001100001101, 1'b0);
		prog_cycle_task(16'b0110001100001101, 1'b0);
		prog_cycle_task(16'b1110001100001101, 1'b1);
		prog_cycle_task(16'b0000011100001101, 1'b0);
		prog_cycle_task(16'b1000011100001101, 1'b0);
		prog_cycle_task(16'b0100011100001101, 1'b1);
		prog_cycle_task(16'b1100011100001101, 1'b0);
		prog_cycle_task(16'b0010011100001101, 1'b0);
		prog_cycle_task(16'b1010011100001101, 1'b0);
		prog_cycle_task(16'b0110011100001101, 1'b0);
		prog_cycle_task(16'b1110011100001101, 1'b1);
		prog_cycle_task(16'b0000000010001101, 1'b0);
		prog_cycle_task(16'b1000000010001101, 1'b0);
		prog_cycle_task(16'b0100000010001101, 1'b1);
		prog_cycle_task(16'b1100000010001101, 1'b0);
		prog_cycle_task(16'b0010000010001101, 1'b0);
		prog_cycle_task(16'b1010000010001101, 1'b0);
		prog_cycle_task(16'b0110000010001101, 1'b0);
		prog_cycle_task(16'b1110000010001101, 1'b1);
		prog_cycle_task(16'b0000010010001101, 1'b0);
		prog_cycle_task(16'b1000010010001101, 1'b0);
		prog_cycle_task(16'b0100010010001101, 1'b1);
		prog_cycle_task(16'b1100010010001101, 1'b0);
		prog_cycle_task(16'b0010010010001101, 1'b0);
		prog_cycle_task(16'b1010010010001101, 1'b0);
		prog_cycle_task(16'b0110010010001101, 1'b0);
		prog_cycle_task(16'b1110010010001101, 1'b1);
		prog_cycle_task(16'b0000001010001101, 1'b0);
		prog_cycle_task(16'b1000001010001101, 1'b0);
		prog_cycle_task(16'b0100001010001101, 1'b1);
		prog_cycle_task(16'b1100001010001101, 1'b0);
		prog_cycle_task(16'b0010001010001101, 1'b0);
		prog_cycle_task(16'b1010001010001101, 1'b0);
		prog_cycle_task(16'b0110001010001101, 1'b0);
		prog_cycle_task(16'b1110001010001101, 1'b1);
		prog_cycle_task(16'b0000011010001101, 1'b0);
		prog_cycle_task(16'b1000011010001101, 1'b0);
		prog_cycle_task(16'b0100011010001101, 1'b1);
		prog_cycle_task(16'b1100011010001101, 1'b0);
		prog_cycle_task(16'b0010011010001101, 1'b0);
		prog_cycle_task(16'b1010011010001101, 1'b0);
		prog_cycle_task(16'b0110011010001101, 1'b0);
		prog_cycle_task(16'b1110011010001101, 1'b1);
		prog_cycle_task(16'b0000000110001101, 1'b0);
		prog_cycle_task(16'b1000000110001101, 1'b0);
		prog_cycle_task(16'b0100000110001101, 1'b1);
		prog_cycle_task(16'b1100000110001101, 1'b0);
		prog_cycle_task(16'b0010000110001101, 1'b0);
		prog_cycle_task(16'b1010000110001101, 1'b0);
		prog_cycle_task(16'b0110000110001101, 1'b0);
		prog_cycle_task(16'b1110000110001101, 1'b1);
		prog_cycle_task(16'b0000010110001101, 1'b0);
		prog_cycle_task(16'b1000010110001101, 1'b0);
		prog_cycle_task(16'b0100010110001101, 1'b1);
		prog_cycle_task(16'b1100010110001101, 1'b0);
		prog_cycle_task(16'b0010010110001101, 1'b0);
		prog_cycle_task(16'b1010010110001101, 1'b0);
		prog_cycle_task(16'b0110010110001101, 1'b0);
		prog_cycle_task(16'b1110010110001101, 1'b1);
		prog_cycle_task(16'b0000001110001101, 1'b0);
		prog_cycle_task(16'b1000001110001101, 1'b0);
		prog_cycle_task(16'b0100001110001101, 1'b1);
		prog_cycle_task(16'b1100001110001101, 1'b0);
		prog_cycle_task(16'b0010001110001101, 1'b0);
		prog_cycle_task(16'b1010001110001101, 1'b0);
		prog_cycle_task(16'b0110001110001101, 1'b0);
		prog_cycle_task(16'b1110001110001101, 1'b1);
		prog_cycle_task(16'b0000011110001101, 1'b0);
		prog_cycle_task(16'b1000011110001101, 1'b0);
		prog_cycle_task(16'b0100011110001101, 1'b1);
		prog_cycle_task(16'b1100011110001101, 1'b0);
		prog_cycle_task(16'b0010011110001101, 1'b0);
		prog_cycle_task(16'b1010011110001101, 1'b0);
		prog_cycle_task(16'b0110011110001101, 1'b0);
		prog_cycle_task(16'b1110011110001101, 1'b1);
		prog_cycle_task(16'b0000000001001101, 1'b0);
		prog_cycle_task(16'b1000000001001101, 1'b0);
		prog_cycle_task(16'b0100000001001101, 1'b1);
		prog_cycle_task(16'b1100000001001101, 1'b0);
		prog_cycle_task(16'b0010000001001101, 1'b0);
		prog_cycle_task(16'b1010000001001101, 1'b0);
		prog_cycle_task(16'b0110000001001101, 1'b0);
		prog_cycle_task(16'b1110000001001101, 1'b1);
		prog_cycle_task(16'b0000010001001101, 1'b0);
		prog_cycle_task(16'b1000010001001101, 1'b0);
		prog_cycle_task(16'b0100010001001101, 1'b1);
		prog_cycle_task(16'b1100010001001101, 1'b0);
		prog_cycle_task(16'b0010010001001101, 1'b0);
		prog_cycle_task(16'b1010010001001101, 1'b0);
		prog_cycle_task(16'b0110010001001101, 1'b0);
		prog_cycle_task(16'b1110010001001101, 1'b1);
		prog_cycle_task(16'b0000001001001101, 1'b0);
		prog_cycle_task(16'b1000001001001101, 1'b0);
		prog_cycle_task(16'b0100001001001101, 1'b1);
		prog_cycle_task(16'b1100001001001101, 1'b0);
		prog_cycle_task(16'b0010001001001101, 1'b0);
		prog_cycle_task(16'b1010001001001101, 1'b0);
		prog_cycle_task(16'b0110001001001101, 1'b0);
		prog_cycle_task(16'b1110001001001101, 1'b1);
		prog_cycle_task(16'b0000011001001101, 1'b0);
		prog_cycle_task(16'b1000011001001101, 1'b0);
		prog_cycle_task(16'b0100011001001101, 1'b1);
		prog_cycle_task(16'b1100011001001101, 1'b0);
		prog_cycle_task(16'b0010011001001101, 1'b0);
		prog_cycle_task(16'b1010011001001101, 1'b0);
		prog_cycle_task(16'b0110011001001101, 1'b0);
		prog_cycle_task(16'b1110011001001101, 1'b1);
		prog_cycle_task(16'b0000000000101101, 1'b0);
		prog_cycle_task(16'b1000000000101101, 1'b0);
		prog_cycle_task(16'b0100000000101101, 1'b0);
		prog_cycle_task(16'b1100000000101101, 1'b0);
		prog_cycle_task(16'b0010000000101101, 1'b0);
		prog_cycle_task(16'b1010000000101101, 1'b0);
		prog_cycle_task(16'b0110000000101101, 1'b0);
		prog_cycle_task(16'b1110000000101101, 1'b1);
		prog_cycle_task(16'b0001000000101101, 1'b0);
		prog_cycle_task(16'b1001000000101101, 1'b0);
		prog_cycle_task(16'b0101000000101101, 1'b0);
		prog_cycle_task(16'b1101000000101101, 1'b0);
		prog_cycle_task(16'b0011000000101101, 1'b0);
		prog_cycle_task(16'b1011000000101101, 1'b0);
		prog_cycle_task(16'b0111000000101101, 1'b0);
		prog_cycle_task(16'b1111000000101101, 1'b1);
		prog_cycle_task(16'b0000100000101101, 1'b0);
		prog_cycle_task(16'b1000100000101101, 1'b0);
		prog_cycle_task(16'b0100100000101101, 1'b1);
		prog_cycle_task(16'b1100100000101101, 1'b0);
		prog_cycle_task(16'b0010100000101101, 1'b0);
		prog_cycle_task(16'b1010100000101101, 1'b1);
		prog_cycle_task(16'b0001100000101101, 1'b0);
		prog_cycle_task(16'b1001100000101101, 1'b0);
		prog_cycle_task(16'b0101100000101101, 1'b0);
		prog_cycle_task(16'b1101100000101101, 1'b0);
		prog_cycle_task(16'b0011100000101101, 1'b0);
		prog_cycle_task(16'b1011100000101101, 1'b0);
		prog_cycle_task(16'b0111100000101101, 1'b0);
		prog_cycle_task(16'b1111100000101101, 1'b1);
		prog_cycle_task(16'b0000010000101101, 1'b0);
		prog_cycle_task(16'b1000010000101101, 1'b0);
		prog_cycle_task(16'b0100010000101101, 1'b0);
		prog_cycle_task(16'b1100010000101101, 1'b0);
		prog_cycle_task(16'b0010010000101101, 1'b0);
		prog_cycle_task(16'b1010010000101101, 1'b0);
		prog_cycle_task(16'b0110010000101101, 1'b0);
		prog_cycle_task(16'b1110010000101101, 1'b1);
		prog_cycle_task(16'b0001010000101101, 1'b0);
		prog_cycle_task(16'b1001010000101101, 1'b0);
		prog_cycle_task(16'b0101010000101101, 1'b1);
		prog_cycle_task(16'b1101010000101101, 1'b0);
		prog_cycle_task(16'b0011010000101101, 1'b0);
		prog_cycle_task(16'b1011010000101101, 1'b1);
		prog_cycle_task(16'b0000110000101101, 1'b0);
		prog_cycle_task(16'b1000110000101101, 1'b0);
		prog_cycle_task(16'b0100110000101101, 1'b0);
		prog_cycle_task(16'b1100110000101101, 1'b0);
		prog_cycle_task(16'b0010110000101101, 1'b0);
		prog_cycle_task(16'b1010110000101101, 1'b0);
		prog_cycle_task(16'b0110110000101101, 1'b0);
		prog_cycle_task(16'b1110110000101101, 1'b1);
		prog_cycle_task(16'b0001110000101101, 1'b0);
		prog_cycle_task(16'b1001110000101101, 1'b1);
		prog_cycle_task(16'b0101110000101101, 1'b0);
		prog_cycle_task(16'b1101110000101101, 1'b0);
		prog_cycle_task(16'b0011110000101101, 1'b0);
		prog_cycle_task(16'b1011110000101101, 1'b1);
		prog_cycle_task(16'b0111110000101101, 1'b0);
		prog_cycle_task(16'b1111110000101101, 1'b0);
		prog_cycle_task(16'b0000001000101101, 1'b0);
		prog_cycle_task(16'b1000001000101101, 1'b0);
		prog_cycle_task(16'b0100001000101101, 1'b1);
		prog_cycle_task(16'b1100001000101101, 1'b0);
		prog_cycle_task(16'b0010001000101101, 1'b0);
		prog_cycle_task(16'b1010001000101101, 1'b1);
		prog_cycle_task(16'b0001001000101101, 1'b0);
		prog_cycle_task(16'b1001001000101101, 1'b0);
		prog_cycle_task(16'b0101001000101101, 1'b0);
		prog_cycle_task(16'b1101001000101101, 1'b0);
		prog_cycle_task(16'b0011001000101101, 1'b0);
		prog_cycle_task(16'b1011001000101101, 1'b0);
		prog_cycle_task(16'b0111001000101101, 1'b0);
		prog_cycle_task(16'b1111001000101101, 1'b1);
		prog_cycle_task(16'b0000101000101101, 1'b0);
		prog_cycle_task(16'b1000101000101101, 1'b0);
		prog_cycle_task(16'b0100101000101101, 1'b0);
		prog_cycle_task(16'b1100101000101101, 1'b0);
		prog_cycle_task(16'b0010101000101101, 1'b0);
		prog_cycle_task(16'b1010101000101101, 1'b0);
		prog_cycle_task(16'b0110101000101101, 1'b0);
		prog_cycle_task(16'b1110101000101101, 1'b1);
		prog_cycle_task(16'b0001101000101101, 1'b0);
		prog_cycle_task(16'b1001101000101101, 1'b0);
		prog_cycle_task(16'b0101101000101101, 1'b1);
		prog_cycle_task(16'b1101101000101101, 1'b0);
		prog_cycle_task(16'b0011101000101101, 1'b0);
		prog_cycle_task(16'b1011101000101101, 1'b1);
		prog_cycle_task(16'b0000000000011101, 1'b0);
		prog_cycle_task(16'b1000000000011101, 1'b0);
		prog_cycle_task(16'b0100000000011101, 1'b0);
		prog_cycle_task(16'b1100000000011101, 1'b0);
		prog_cycle_task(16'b0010000000011101, 1'b0);
		prog_cycle_task(16'b1010000000011101, 1'b1);
		prog_cycle_task(16'b0001000000011101, 1'b0);
		prog_cycle_task(16'b1001000000011101, 1'b0);
		prog_cycle_task(16'b0000100000011101, 1'b0);
		prog_cycle_task(16'b1000100000011101, 1'b0);
		prog_cycle_task(16'b0100100000011101, 1'b0);
		prog_cycle_task(16'b1100100000011101, 1'b0);
		prog_cycle_task(16'b0010100000011101, 1'b0);
		prog_cycle_task(16'b1010100000011101, 1'b1);
		prog_cycle_task(16'b0001100000011101, 1'b0);
		prog_cycle_task(16'b1001100000011101, 1'b0);
		prog_cycle_task(16'b0101100000011101, 1'b0);
		prog_cycle_task(16'b1101100000011101, 1'b0);
		prog_cycle_task(16'b0011100000011101, 1'b0);
		prog_cycle_task(16'b1011100000011101, 1'b1);
		prog_cycle_task(16'b0000010000011101, 1'b0);
		prog_cycle_task(16'b1000010000011101, 1'b0);
		prog_cycle_task(16'b0001010000011101, 1'b0);
		prog_cycle_task(16'b1001010000011101, 1'b0);
		prog_cycle_task(16'b0000000000111101, 1'b0);
		prog_cycle_task(16'b1000000000111101, 1'b0);
		prog_cycle_task(16'b0100000000111101, 1'b0);
		prog_cycle_task(16'b1100000000111101, 1'b0);
		prog_cycle_task(16'b0010000000111101, 1'b0);
		prog_cycle_task(16'b1010000000111101, 1'b1);
		prog_cycle_task(16'b0001000000111101, 1'b0);
		prog_cycle_task(16'b1001000000111101, 1'b0);
		prog_cycle_task(16'b0000100000111101, 1'b0);
		prog_cycle_task(16'b1000100000111101, 1'b0);
		prog_cycle_task(16'b0100100000111101, 1'b0);
		prog_cycle_task(16'b1100100000111101, 1'b0);
		prog_cycle_task(16'b0010100000111101, 1'b0);
		prog_cycle_task(16'b1010100000111101, 1'b1);
		prog_cycle_task(16'b0001100000111101, 1'b0);
		prog_cycle_task(16'b1001100000111101, 1'b0);
		prog_cycle_task(16'b0000010000111101, 1'b0);
		prog_cycle_task(16'b1000010000111101, 1'b0);
		prog_cycle_task(16'b0000000000000011, 1'b0);
		prog_cycle_task(16'b1000000000000011, 1'b0);
		prog_cycle_task(16'b0100000000000011, 1'b0);
		prog_cycle_task(16'b1100000000000011, 1'b0);
		prog_cycle_task(16'b0010000000000011, 1'b0);
		prog_cycle_task(16'b1010000000000011, 1'b0);
		prog_cycle_task(16'b0110000000000011, 1'b0);
		prog_cycle_task(16'b1110000000000011, 1'b0);
		prog_cycle_task(16'b0001000000000011, 1'b0);
		prog_cycle_task(16'b1001000000000011, 1'b0);
		prog_cycle_task(16'b0101000000000011, 1'b0);
		prog_cycle_task(16'b1101000000000011, 1'b0);
		prog_cycle_task(16'b0011000000000011, 1'b0);
		prog_cycle_task(16'b1011000000000011, 1'b0);
		prog_cycle_task(16'b0111000000000011, 1'b0);
		prog_cycle_task(16'b1111000000000011, 1'b0);
		prog_cycle_task(16'b0000100000000011, 1'b0);
		prog_cycle_task(16'b1000100000000011, 1'b0);
		prog_cycle_task(16'b0100100000000011, 1'b1);
		prog_cycle_task(16'b0000010000000011, 1'b0);
		prog_cycle_task(16'b1000010000000011, 1'b0);
		prog_cycle_task(16'b0100010000000011, 1'b0);
		prog_cycle_task(16'b1100010000000011, 1'b0);
		prog_cycle_task(16'b0010010000000011, 1'b0);
		prog_cycle_task(16'b1010010000000011, 1'b0);
		prog_cycle_task(16'b0110010000000011, 1'b0);
		prog_cycle_task(16'b1110010000000011, 1'b0);
		prog_cycle_task(16'b0001010000000011, 1'b0);
		prog_cycle_task(16'b1001010000000011, 1'b0);
		prog_cycle_task(16'b0101010000000011, 1'b0);
		prog_cycle_task(16'b1101010000000011, 1'b0);
		prog_cycle_task(16'b0011010000000011, 1'b0);
		prog_cycle_task(16'b1011010000000011, 1'b0);
		prog_cycle_task(16'b0111010000000011, 1'b0);
		prog_cycle_task(16'b1111010000000011, 1'b0);
		prog_cycle_task(16'b0000110000000011, 1'b0);
		prog_cycle_task(16'b1000110000000011, 1'b0);
		prog_cycle_task(16'b0100110000000011, 1'b1);
		prog_cycle_task(16'b0000001000000011, 1'b0);
		prog_cycle_task(16'b1000001000000011, 1'b0);
		prog_cycle_task(16'b0100001000000011, 1'b0);
		prog_cycle_task(16'b1100001000000011, 1'b0);
		prog_cycle_task(16'b0010001000000011, 1'b0);
		prog_cycle_task(16'b1010001000000011, 1'b0);
		prog_cycle_task(16'b0110001000000011, 1'b0);
		prog_cycle_task(16'b1110001000000011, 1'b0);
		prog_cycle_task(16'b0001001000000011, 1'b0);
		prog_cycle_task(16'b1001001000000011, 1'b0);
		prog_cycle_task(16'b0101001000000011, 1'b0);
		prog_cycle_task(16'b1101001000000011, 1'b0);
		prog_cycle_task(16'b0011001000000011, 1'b0);
		prog_cycle_task(16'b1011001000000011, 1'b0);
		prog_cycle_task(16'b0111001000000011, 1'b0);
		prog_cycle_task(16'b1111001000000011, 1'b0);
		prog_cycle_task(16'b0000101000000011, 1'b0);
		prog_cycle_task(16'b1000101000000011, 1'b0);
		prog_cycle_task(16'b0100101000000011, 1'b1);
		prog_cycle_task(16'b0000011000000011, 1'b0);
		prog_cycle_task(16'b1000011000000011, 1'b0);
		prog_cycle_task(16'b0100011000000011, 1'b0);
		prog_cycle_task(16'b1100011000000011, 1'b0);
		prog_cycle_task(16'b0010011000000011, 1'b0);
		prog_cycle_task(16'b1010011000000011, 1'b0);
		prog_cycle_task(16'b0110011000000011, 1'b0);
		prog_cycle_task(16'b1110011000000011, 1'b0);
		prog_cycle_task(16'b0001011000000011, 1'b0);
		prog_cycle_task(16'b1001011000000011, 1'b0);
		prog_cycle_task(16'b0101011000000011, 1'b0);
		prog_cycle_task(16'b1101011000000011, 1'b0);
		prog_cycle_task(16'b0011011000000011, 1'b0);
		prog_cycle_task(16'b1011011000000011, 1'b0);
		prog_cycle_task(16'b0111011000000011, 1'b0);
		prog_cycle_task(16'b1111011000000011, 1'b0);
		prog_cycle_task(16'b0000111000000011, 1'b0);
		prog_cycle_task(16'b1000111000000011, 1'b0);
		prog_cycle_task(16'b0100111000000011, 1'b1);
		prog_cycle_task(16'b0000000100000011, 1'b0);
		prog_cycle_task(16'b1000000100000011, 1'b0);
		prog_cycle_task(16'b0100000100000011, 1'b1);
		prog_cycle_task(16'b1100000100000011, 1'b0);
		prog_cycle_task(16'b0010000100000011, 1'b0);
		prog_cycle_task(16'b1010000100000011, 1'b0);
		prog_cycle_task(16'b0110000100000011, 1'b0);
		prog_cycle_task(16'b1110000100000011, 1'b1);
		prog_cycle_task(16'b0000010100000011, 1'b0);
		prog_cycle_task(16'b1000010100000011, 1'b0);
		prog_cycle_task(16'b0100010100000011, 1'b1);
		prog_cycle_task(16'b1100010100000011, 1'b0);
		prog_cycle_task(16'b0010010100000011, 1'b0);
		prog_cycle_task(16'b1010010100000011, 1'b0);
		prog_cycle_task(16'b0110010100000011, 1'b0);
		prog_cycle_task(16'b1110010100000011, 1'b1);
		prog_cycle_task(16'b0000001100000011, 1'b0);
		prog_cycle_task(16'b1000001100000011, 1'b0);
		prog_cycle_task(16'b0100001100000011, 1'b1);
		prog_cycle_task(16'b1100001100000011, 1'b0);
		prog_cycle_task(16'b0010001100000011, 1'b0);
		prog_cycle_task(16'b1010001100000011, 1'b0);
		prog_cycle_task(16'b0110001100000011, 1'b0);
		prog_cycle_task(16'b1110001100000011, 1'b1);
		prog_cycle_task(16'b0000011100000011, 1'b0);
		prog_cycle_task(16'b1000011100000011, 1'b0);
		prog_cycle_task(16'b0100011100000011, 1'b1);
		prog_cycle_task(16'b1100011100000011, 1'b0);
		prog_cycle_task(16'b0010011100000011, 1'b0);
		prog_cycle_task(16'b1010011100000011, 1'b0);
		prog_cycle_task(16'b0110011100000011, 1'b0);
		prog_cycle_task(16'b1110011100000011, 1'b1);
		prog_cycle_task(16'b0000000010000011, 1'b0);
		prog_cycle_task(16'b1000000010000011, 1'b0);
		prog_cycle_task(16'b0100000010000011, 1'b1);
		prog_cycle_task(16'b1100000010000011, 1'b0);
		prog_cycle_task(16'b0010000010000011, 1'b0);
		prog_cycle_task(16'b1010000010000011, 1'b0);
		prog_cycle_task(16'b0110000010000011, 1'b0);
		prog_cycle_task(16'b1110000010000011, 1'b1);
		prog_cycle_task(16'b0000010010000011, 1'b0);
		prog_cycle_task(16'b1000010010000011, 1'b0);
		prog_cycle_task(16'b0100010010000011, 1'b1);
		prog_cycle_task(16'b1100010010000011, 1'b0);
		prog_cycle_task(16'b0010010010000011, 1'b0);
		prog_cycle_task(16'b1010010010000011, 1'b0);
		prog_cycle_task(16'b0110010010000011, 1'b0);
		prog_cycle_task(16'b1110010010000011, 1'b1);
		prog_cycle_task(16'b0000001010000011, 1'b0);
		prog_cycle_task(16'b1000001010000011, 1'b0);
		prog_cycle_task(16'b0100001010000011, 1'b1);
		prog_cycle_task(16'b1100001010000011, 1'b0);
		prog_cycle_task(16'b0010001010000011, 1'b0);
		prog_cycle_task(16'b1010001010000011, 1'b0);
		prog_cycle_task(16'b0110001010000011, 1'b0);
		prog_cycle_task(16'b1110001010000011, 1'b1);
		prog_cycle_task(16'b0000011010000011, 1'b0);
		prog_cycle_task(16'b1000011010000011, 1'b0);
		prog_cycle_task(16'b0100011010000011, 1'b1);
		prog_cycle_task(16'b1100011010000011, 1'b0);
		prog_cycle_task(16'b0010011010000011, 1'b0);
		prog_cycle_task(16'b1010011010000011, 1'b0);
		prog_cycle_task(16'b0110011010000011, 1'b0);
		prog_cycle_task(16'b1110011010000011, 1'b1);
		prog_cycle_task(16'b0000000110000011, 1'b0);
		prog_cycle_task(16'b1000000110000011, 1'b0);
		prog_cycle_task(16'b0100000110000011, 1'b1);
		prog_cycle_task(16'b1100000110000011, 1'b0);
		prog_cycle_task(16'b0010000110000011, 1'b0);
		prog_cycle_task(16'b1010000110000011, 1'b0);
		prog_cycle_task(16'b0110000110000011, 1'b0);
		prog_cycle_task(16'b1110000110000011, 1'b1);
		prog_cycle_task(16'b0000010110000011, 1'b0);
		prog_cycle_task(16'b1000010110000011, 1'b0);
		prog_cycle_task(16'b0100010110000011, 1'b1);
		prog_cycle_task(16'b1100010110000011, 1'b0);
		prog_cycle_task(16'b0010010110000011, 1'b0);
		prog_cycle_task(16'b1010010110000011, 1'b0);
		prog_cycle_task(16'b0110010110000011, 1'b0);
		prog_cycle_task(16'b1110010110000011, 1'b1);
		prog_cycle_task(16'b0000001110000011, 1'b0);
		prog_cycle_task(16'b1000001110000011, 1'b0);
		prog_cycle_task(16'b0100001110000011, 1'b1);
		prog_cycle_task(16'b1100001110000011, 1'b0);
		prog_cycle_task(16'b0010001110000011, 1'b0);
		prog_cycle_task(16'b1010001110000011, 1'b0);
		prog_cycle_task(16'b0110001110000011, 1'b0);
		prog_cycle_task(16'b1110001110000011, 1'b1);
		prog_cycle_task(16'b0000011110000011, 1'b0);
		prog_cycle_task(16'b1000011110000011, 1'b0);
		prog_cycle_task(16'b0100011110000011, 1'b1);
		prog_cycle_task(16'b1100011110000011, 1'b0);
		prog_cycle_task(16'b0010011110000011, 1'b0);
		prog_cycle_task(16'b1010011110000011, 1'b0);
		prog_cycle_task(16'b0110011110000011, 1'b0);
		prog_cycle_task(16'b1110011110000011, 1'b1);
		prog_cycle_task(16'b0000000001000011, 1'b0);
		prog_cycle_task(16'b1000000001000011, 1'b0);
		prog_cycle_task(16'b0100000001000011, 1'b1);
		prog_cycle_task(16'b1100000001000011, 1'b0);
		prog_cycle_task(16'b0010000001000011, 1'b0);
		prog_cycle_task(16'b1010000001000011, 1'b0);
		prog_cycle_task(16'b0110000001000011, 1'b0);
		prog_cycle_task(16'b1110000001000011, 1'b1);
		prog_cycle_task(16'b0000010001000011, 1'b0);
		prog_cycle_task(16'b1000010001000011, 1'b0);
		prog_cycle_task(16'b0100010001000011, 1'b1);
		prog_cycle_task(16'b1100010001000011, 1'b0);
		prog_cycle_task(16'b0010010001000011, 1'b0);
		prog_cycle_task(16'b1010010001000011, 1'b0);
		prog_cycle_task(16'b0110010001000011, 1'b0);
		prog_cycle_task(16'b1110010001000011, 1'b1);
		prog_cycle_task(16'b0000001001000011, 1'b0);
		prog_cycle_task(16'b1000001001000011, 1'b0);
		prog_cycle_task(16'b0100001001000011, 1'b1);
		prog_cycle_task(16'b1100001001000011, 1'b0);
		prog_cycle_task(16'b0010001001000011, 1'b0);
		prog_cycle_task(16'b1010001001000011, 1'b0);
		prog_cycle_task(16'b0110001001000011, 1'b0);
		prog_cycle_task(16'b1110001001000011, 1'b1);
		prog_cycle_task(16'b0000011001000011, 1'b0);
		prog_cycle_task(16'b1000011001000011, 1'b0);
		prog_cycle_task(16'b0100011001000011, 1'b1);
		prog_cycle_task(16'b1100011001000011, 1'b0);
		prog_cycle_task(16'b0010011001000011, 1'b0);
		prog_cycle_task(16'b1010011001000011, 1'b0);
		prog_cycle_task(16'b0110011001000011, 1'b0);
		prog_cycle_task(16'b1110011001000011, 1'b1);
		prog_cycle_task(16'b0000000000100011, 1'b0);
		prog_cycle_task(16'b1000000000100011, 1'b0);
		prog_cycle_task(16'b0100000000100011, 1'b0);
		prog_cycle_task(16'b1100000000100011, 1'b0);
		prog_cycle_task(16'b0010000000100011, 1'b0);
		prog_cycle_task(16'b1010000000100011, 1'b0);
		prog_cycle_task(16'b0110000000100011, 1'b0);
		prog_cycle_task(16'b1110000000100011, 1'b1);
		prog_cycle_task(16'b0001000000100011, 1'b0);
		prog_cycle_task(16'b1001000000100011, 1'b0);
		prog_cycle_task(16'b0101000000100011, 1'b0);
		prog_cycle_task(16'b1101000000100011, 1'b0);
		prog_cycle_task(16'b0011000000100011, 1'b0);
		prog_cycle_task(16'b1011000000100011, 1'b0);
		prog_cycle_task(16'b0111000000100011, 1'b0);
		prog_cycle_task(16'b1111000000100011, 1'b1);
		prog_cycle_task(16'b0000100000100011, 1'b0);
		prog_cycle_task(16'b1000100000100011, 1'b0);
		prog_cycle_task(16'b0100100000100011, 1'b1);
		prog_cycle_task(16'b1100100000100011, 1'b0);
		prog_cycle_task(16'b0010100000100011, 1'b0);
		prog_cycle_task(16'b1010100000100011, 1'b1);
		prog_cycle_task(16'b0001100000100011, 1'b0);
		prog_cycle_task(16'b1001100000100011, 1'b0);
		prog_cycle_task(16'b0101100000100011, 1'b0);
		prog_cycle_task(16'b1101100000100011, 1'b0);
		prog_cycle_task(16'b0011100000100011, 1'b0);
		prog_cycle_task(16'b1011100000100011, 1'b0);
		prog_cycle_task(16'b0111100000100011, 1'b0);
		prog_cycle_task(16'b1111100000100011, 1'b1);
		prog_cycle_task(16'b0000010000100011, 1'b0);
		prog_cycle_task(16'b1000010000100011, 1'b0);
		prog_cycle_task(16'b0100010000100011, 1'b0);
		prog_cycle_task(16'b1100010000100011, 1'b0);
		prog_cycle_task(16'b0010010000100011, 1'b0);
		prog_cycle_task(16'b1010010000100011, 1'b0);
		prog_cycle_task(16'b0110010000100011, 1'b0);
		prog_cycle_task(16'b1110010000100011, 1'b1);
		prog_cycle_task(16'b0001010000100011, 1'b0);
		prog_cycle_task(16'b1001010000100011, 1'b0);
		prog_cycle_task(16'b0101010000100011, 1'b1);
		prog_cycle_task(16'b1101010000100011, 1'b0);
		prog_cycle_task(16'b0011010000100011, 1'b0);
		prog_cycle_task(16'b1011010000100011, 1'b1);
		prog_cycle_task(16'b0000110000100011, 1'b0);
		prog_cycle_task(16'b1000110000100011, 1'b0);
		prog_cycle_task(16'b0100110000100011, 1'b0);
		prog_cycle_task(16'b1100110000100011, 1'b0);
		prog_cycle_task(16'b0010110000100011, 1'b0);
		prog_cycle_task(16'b1010110000100011, 1'b0);
		prog_cycle_task(16'b0110110000100011, 1'b0);
		prog_cycle_task(16'b1110110000100011, 1'b1);
		prog_cycle_task(16'b0001110000100011, 1'b0);
		prog_cycle_task(16'b1001110000100011, 1'b0);
		prog_cycle_task(16'b0101110000100011, 1'b0);
		prog_cycle_task(16'b1101110000100011, 1'b0);
		prog_cycle_task(16'b0011110000100011, 1'b0);
		prog_cycle_task(16'b1011110000100011, 1'b0);
		prog_cycle_task(16'b0111110000100011, 1'b0);
		prog_cycle_task(16'b1111110000100011, 1'b1);
		prog_cycle_task(16'b0000001000100011, 1'b0);
		prog_cycle_task(16'b1000001000100011, 1'b0);
		prog_cycle_task(16'b0100001000100011, 1'b1);
		prog_cycle_task(16'b1100001000100011, 1'b0);
		prog_cycle_task(16'b0010001000100011, 1'b0);
		prog_cycle_task(16'b1010001000100011, 1'b1);
		prog_cycle_task(16'b0001001000100011, 1'b0);
		prog_cycle_task(16'b1001001000100011, 1'b0);
		prog_cycle_task(16'b0101001000100011, 1'b0);
		prog_cycle_task(16'b1101001000100011, 1'b0);
		prog_cycle_task(16'b0011001000100011, 1'b0);
		prog_cycle_task(16'b1011001000100011, 1'b0);
		prog_cycle_task(16'b0111001000100011, 1'b0);
		prog_cycle_task(16'b1111001000100011, 1'b1);
		prog_cycle_task(16'b0000101000100011, 1'b0);
		prog_cycle_task(16'b1000101000100011, 1'b0);
		prog_cycle_task(16'b0100101000100011, 1'b0);
		prog_cycle_task(16'b1100101000100011, 1'b0);
		prog_cycle_task(16'b0010101000100011, 1'b0);
		prog_cycle_task(16'b1010101000100011, 1'b0);
		prog_cycle_task(16'b0110101000100011, 1'b0);
		prog_cycle_task(16'b1110101000100011, 1'b1);
		prog_cycle_task(16'b0001101000100011, 1'b0);
		prog_cycle_task(16'b1001101000100011, 1'b0);
		prog_cycle_task(16'b0101101000100011, 1'b1);
		prog_cycle_task(16'b1101101000100011, 1'b0);
		prog_cycle_task(16'b0011101000100011, 1'b0);
		prog_cycle_task(16'b1011101000100011, 1'b1);
		prog_cycle_task(16'b0000000000010011, 1'b0);
		prog_cycle_task(16'b1000000000010011, 1'b0);
		prog_cycle_task(16'b0100000000010011, 1'b0);
		prog_cycle_task(16'b1100000000010011, 1'b0);
		prog_cycle_task(16'b0010000000010011, 1'b0);
		prog_cycle_task(16'b1010000000010011, 1'b1);
		prog_cycle_task(16'b0001000000010011, 1'b0);
		prog_cycle_task(16'b1001000000010011, 1'b0);
		prog_cycle_task(16'b0000100000010011, 1'b0);
		prog_cycle_task(16'b1000100000010011, 1'b0);
		prog_cycle_task(16'b0100100000010011, 1'b0);
		prog_cycle_task(16'b1100100000010011, 1'b0);
		prog_cycle_task(16'b0010100000010011, 1'b0);
		prog_cycle_task(16'b1010100000010011, 1'b1);
		prog_cycle_task(16'b0001100000010011, 1'b0);
		prog_cycle_task(16'b1001100000010011, 1'b0);
		prog_cycle_task(16'b0101100000010011, 1'b0);
		prog_cycle_task(16'b1101100000010011, 1'b0);
		prog_cycle_task(16'b0011100000010011, 1'b0);
		prog_cycle_task(16'b1011100000010011, 1'b1);
		prog_cycle_task(16'b0000010000010011, 1'b0);
		prog_cycle_task(16'b1000010000010011, 1'b0);
		prog_cycle_task(16'b0001010000010011, 1'b0);
		prog_cycle_task(16'b1001010000010011, 1'b0);
		prog_cycle_task(16'b0000000000110011, 1'b0);
		prog_cycle_task(16'b1000000000110011, 1'b0);
		prog_cycle_task(16'b0100000000110011, 1'b0);
		prog_cycle_task(16'b1100000000110011, 1'b0);
		prog_cycle_task(16'b0010000000110011, 1'b0);
		prog_cycle_task(16'b1010000000110011, 1'b1);
		prog_cycle_task(16'b0001000000110011, 1'b0);
		prog_cycle_task(16'b1001000000110011, 1'b0);
		prog_cycle_task(16'b0000100000110011, 1'b0);
		prog_cycle_task(16'b1000100000110011, 1'b0);
		prog_cycle_task(16'b0100100000110011, 1'b0);
		prog_cycle_task(16'b1100100000110011, 1'b0);
		prog_cycle_task(16'b0010100000110011, 1'b0);
		prog_cycle_task(16'b1010100000110011, 1'b1);
		prog_cycle_task(16'b0001100000110011, 1'b0);
		prog_cycle_task(16'b1001100000110011, 1'b0);
		prog_cycle_task(16'b0000010000110011, 1'b0);
		prog_cycle_task(16'b1000010000110011, 1'b0);
		prog_cycle_task(16'b0000000000001011, 1'b0);
		prog_cycle_task(16'b1000000000001011, 1'b0);
		prog_cycle_task(16'b0100000000001011, 1'b0);
		prog_cycle_task(16'b1100000000001011, 1'b0);
		prog_cycle_task(16'b0010000000001011, 1'b0);
		prog_cycle_task(16'b1010000000001011, 1'b0);
		prog_cycle_task(16'b0110000000001011, 1'b0);
		prog_cycle_task(16'b1110000000001011, 1'b0);
		prog_cycle_task(16'b0001000000001011, 1'b0);
		prog_cycle_task(16'b1001000000001011, 1'b0);
		prog_cycle_task(16'b0101000000001011, 1'b0);
		prog_cycle_task(16'b1101000000001011, 1'b0);
		prog_cycle_task(16'b0011000000001011, 1'b0);
		prog_cycle_task(16'b1011000000001011, 1'b0);
		prog_cycle_task(16'b0111000000001011, 1'b0);
		prog_cycle_task(16'b1111000000001011, 1'b0);
		prog_cycle_task(16'b0000100000001011, 1'b0);
		prog_cycle_task(16'b1000100000001011, 1'b0);
		prog_cycle_task(16'b0100100000001011, 1'b1);
		prog_cycle_task(16'b0000010000001011, 1'b0);
		prog_cycle_task(16'b1000010000001011, 1'b0);
		prog_cycle_task(16'b0100010000001011, 1'b0);
		prog_cycle_task(16'b1100010000001011, 1'b0);
		prog_cycle_task(16'b0010010000001011, 1'b0);
		prog_cycle_task(16'b1010010000001011, 1'b0);
		prog_cycle_task(16'b0110010000001011, 1'b0);
		prog_cycle_task(16'b1110010000001011, 1'b0);
		prog_cycle_task(16'b0001010000001011, 1'b0);
		prog_cycle_task(16'b1001010000001011, 1'b0);
		prog_cycle_task(16'b0101010000001011, 1'b0);
		prog_cycle_task(16'b1101010000001011, 1'b0);
		prog_cycle_task(16'b0011010000001011, 1'b0);
		prog_cycle_task(16'b1011010000001011, 1'b0);
		prog_cycle_task(16'b0111010000001011, 1'b0);
		prog_cycle_task(16'b1111010000001011, 1'b0);
		prog_cycle_task(16'b0000110000001011, 1'b0);
		prog_cycle_task(16'b1000110000001011, 1'b0);
		prog_cycle_task(16'b0100110000001011, 1'b1);
		prog_cycle_task(16'b0000001000001011, 1'b0);
		prog_cycle_task(16'b1000001000001011, 1'b0);
		prog_cycle_task(16'b0100001000001011, 1'b0);
		prog_cycle_task(16'b1100001000001011, 1'b0);
		prog_cycle_task(16'b0010001000001011, 1'b0);
		prog_cycle_task(16'b1010001000001011, 1'b0);
		prog_cycle_task(16'b0110001000001011, 1'b0);
		prog_cycle_task(16'b1110001000001011, 1'b0);
		prog_cycle_task(16'b0001001000001011, 1'b0);
		prog_cycle_task(16'b1001001000001011, 1'b0);
		prog_cycle_task(16'b0101001000001011, 1'b0);
		prog_cycle_task(16'b1101001000001011, 1'b0);
		prog_cycle_task(16'b0011001000001011, 1'b0);
		prog_cycle_task(16'b1011001000001011, 1'b0);
		prog_cycle_task(16'b0111001000001011, 1'b0);
		prog_cycle_task(16'b1111001000001011, 1'b0);
		prog_cycle_task(16'b0000101000001011, 1'b0);
		prog_cycle_task(16'b1000101000001011, 1'b0);
		prog_cycle_task(16'b0100101000001011, 1'b1);
		prog_cycle_task(16'b0000011000001011, 1'b0);
		prog_cycle_task(16'b1000011000001011, 1'b0);
		prog_cycle_task(16'b0100011000001011, 1'b0);
		prog_cycle_task(16'b1100011000001011, 1'b0);
		prog_cycle_task(16'b0010011000001011, 1'b0);
		prog_cycle_task(16'b1010011000001011, 1'b0);
		prog_cycle_task(16'b0110011000001011, 1'b0);
		prog_cycle_task(16'b1110011000001011, 1'b0);
		prog_cycle_task(16'b0001011000001011, 1'b0);
		prog_cycle_task(16'b1001011000001011, 1'b0);
		prog_cycle_task(16'b0101011000001011, 1'b0);
		prog_cycle_task(16'b1101011000001011, 1'b0);
		prog_cycle_task(16'b0011011000001011, 1'b0);
		prog_cycle_task(16'b1011011000001011, 1'b0);
		prog_cycle_task(16'b0111011000001011, 1'b0);
		prog_cycle_task(16'b1111011000001011, 1'b0);
		prog_cycle_task(16'b0000111000001011, 1'b0);
		prog_cycle_task(16'b1000111000001011, 1'b0);
		prog_cycle_task(16'b0100111000001011, 1'b1);
		prog_cycle_task(16'b0000000100001011, 1'b0);
		prog_cycle_task(16'b1000000100001011, 1'b0);
		prog_cycle_task(16'b0100000100001011, 1'b1);
		prog_cycle_task(16'b1100000100001011, 1'b0);
		prog_cycle_task(16'b0010000100001011, 1'b0);
		prog_cycle_task(16'b1010000100001011, 1'b0);
		prog_cycle_task(16'b0110000100001011, 1'b0);
		prog_cycle_task(16'b1110000100001011, 1'b1);
		prog_cycle_task(16'b0000010100001011, 1'b0);
		prog_cycle_task(16'b1000010100001011, 1'b0);
		prog_cycle_task(16'b0100010100001011, 1'b1);
		prog_cycle_task(16'b1100010100001011, 1'b0);
		prog_cycle_task(16'b0010010100001011, 1'b0);
		prog_cycle_task(16'b1010010100001011, 1'b0);
		prog_cycle_task(16'b0110010100001011, 1'b0);
		prog_cycle_task(16'b1110010100001011, 1'b1);
		prog_cycle_task(16'b0000001100001011, 1'b0);
		prog_cycle_task(16'b1000001100001011, 1'b0);
		prog_cycle_task(16'b0100001100001011, 1'b1);
		prog_cycle_task(16'b1100001100001011, 1'b0);
		prog_cycle_task(16'b0010001100001011, 1'b0);
		prog_cycle_task(16'b1010001100001011, 1'b0);
		prog_cycle_task(16'b0110001100001011, 1'b0);
		prog_cycle_task(16'b1110001100001011, 1'b1);
		prog_cycle_task(16'b0000011100001011, 1'b0);
		prog_cycle_task(16'b1000011100001011, 1'b0);
		prog_cycle_task(16'b0100011100001011, 1'b1);
		prog_cycle_task(16'b1100011100001011, 1'b0);
		prog_cycle_task(16'b0010011100001011, 1'b0);
		prog_cycle_task(16'b1010011100001011, 1'b0);
		prog_cycle_task(16'b0110011100001011, 1'b0);
		prog_cycle_task(16'b1110011100001011, 1'b1);
		prog_cycle_task(16'b0000000010001011, 1'b0);
		prog_cycle_task(16'b1000000010001011, 1'b0);
		prog_cycle_task(16'b0100000010001011, 1'b1);
		prog_cycle_task(16'b1100000010001011, 1'b0);
		prog_cycle_task(16'b0010000010001011, 1'b0);
		prog_cycle_task(16'b1010000010001011, 1'b0);
		prog_cycle_task(16'b0110000010001011, 1'b0);
		prog_cycle_task(16'b1110000010001011, 1'b1);
		prog_cycle_task(16'b0000010010001011, 1'b0);
		prog_cycle_task(16'b1000010010001011, 1'b0);
		prog_cycle_task(16'b0100010010001011, 1'b1);
		prog_cycle_task(16'b1100010010001011, 1'b0);
		prog_cycle_task(16'b0010010010001011, 1'b0);
		prog_cycle_task(16'b1010010010001011, 1'b0);
		prog_cycle_task(16'b0110010010001011, 1'b0);
		prog_cycle_task(16'b1110010010001011, 1'b1);
		prog_cycle_task(16'b0000001010001011, 1'b0);
		prog_cycle_task(16'b1000001010001011, 1'b0);
		prog_cycle_task(16'b0100001010001011, 1'b1);
		prog_cycle_task(16'b1100001010001011, 1'b0);
		prog_cycle_task(16'b0010001010001011, 1'b0);
		prog_cycle_task(16'b1010001010001011, 1'b0);
		prog_cycle_task(16'b0110001010001011, 1'b0);
		prog_cycle_task(16'b1110001010001011, 1'b1);
		prog_cycle_task(16'b0000011010001011, 1'b0);
		prog_cycle_task(16'b1000011010001011, 1'b0);
		prog_cycle_task(16'b0100011010001011, 1'b1);
		prog_cycle_task(16'b1100011010001011, 1'b0);
		prog_cycle_task(16'b0010011010001011, 1'b0);
		prog_cycle_task(16'b1010011010001011, 1'b0);
		prog_cycle_task(16'b0110011010001011, 1'b0);
		prog_cycle_task(16'b1110011010001011, 1'b1);
		prog_cycle_task(16'b0000000110001011, 1'b0);
		prog_cycle_task(16'b1000000110001011, 1'b0);
		prog_cycle_task(16'b0100000110001011, 1'b1);
		prog_cycle_task(16'b1100000110001011, 1'b0);
		prog_cycle_task(16'b0010000110001011, 1'b0);
		prog_cycle_task(16'b1010000110001011, 1'b0);
		prog_cycle_task(16'b0110000110001011, 1'b0);
		prog_cycle_task(16'b1110000110001011, 1'b1);
		prog_cycle_task(16'b0000010110001011, 1'b0);
		prog_cycle_task(16'b1000010110001011, 1'b0);
		prog_cycle_task(16'b0100010110001011, 1'b1);
		prog_cycle_task(16'b1100010110001011, 1'b0);
		prog_cycle_task(16'b0010010110001011, 1'b0);
		prog_cycle_task(16'b1010010110001011, 1'b0);
		prog_cycle_task(16'b0110010110001011, 1'b0);
		prog_cycle_task(16'b1110010110001011, 1'b1);
		prog_cycle_task(16'b0000001110001011, 1'b0);
		prog_cycle_task(16'b1000001110001011, 1'b0);
		prog_cycle_task(16'b0100001110001011, 1'b1);
		prog_cycle_task(16'b1100001110001011, 1'b0);
		prog_cycle_task(16'b0010001110001011, 1'b0);
		prog_cycle_task(16'b1010001110001011, 1'b0);
		prog_cycle_task(16'b0110001110001011, 1'b0);
		prog_cycle_task(16'b1110001110001011, 1'b1);
		prog_cycle_task(16'b0000011110001011, 1'b0);
		prog_cycle_task(16'b1000011110001011, 1'b0);
		prog_cycle_task(16'b0100011110001011, 1'b1);
		prog_cycle_task(16'b1100011110001011, 1'b0);
		prog_cycle_task(16'b0010011110001011, 1'b0);
		prog_cycle_task(16'b1010011110001011, 1'b0);
		prog_cycle_task(16'b0110011110001011, 1'b0);
		prog_cycle_task(16'b1110011110001011, 1'b1);
		prog_cycle_task(16'b0000000001001011, 1'b0);
		prog_cycle_task(16'b1000000001001011, 1'b0);
		prog_cycle_task(16'b0100000001001011, 1'b1);
		prog_cycle_task(16'b1100000001001011, 1'b0);
		prog_cycle_task(16'b0010000001001011, 1'b0);
		prog_cycle_task(16'b1010000001001011, 1'b0);
		prog_cycle_task(16'b0110000001001011, 1'b0);
		prog_cycle_task(16'b1110000001001011, 1'b1);
		prog_cycle_task(16'b0000010001001011, 1'b0);
		prog_cycle_task(16'b1000010001001011, 1'b0);
		prog_cycle_task(16'b0100010001001011, 1'b1);
		prog_cycle_task(16'b1100010001001011, 1'b0);
		prog_cycle_task(16'b0010010001001011, 1'b0);
		prog_cycle_task(16'b1010010001001011, 1'b0);
		prog_cycle_task(16'b0110010001001011, 1'b0);
		prog_cycle_task(16'b1110010001001011, 1'b1);
		prog_cycle_task(16'b0000001001001011, 1'b0);
		prog_cycle_task(16'b1000001001001011, 1'b0);
		prog_cycle_task(16'b0100001001001011, 1'b1);
		prog_cycle_task(16'b1100001001001011, 1'b0);
		prog_cycle_task(16'b0010001001001011, 1'b0);
		prog_cycle_task(16'b1010001001001011, 1'b0);
		prog_cycle_task(16'b0110001001001011, 1'b0);
		prog_cycle_task(16'b1110001001001011, 1'b1);
		prog_cycle_task(16'b0000011001001011, 1'b0);
		prog_cycle_task(16'b1000011001001011, 1'b0);
		prog_cycle_task(16'b0100011001001011, 1'b1);
		prog_cycle_task(16'b1100011001001011, 1'b0);
		prog_cycle_task(16'b0010011001001011, 1'b0);
		prog_cycle_task(16'b1010011001001011, 1'b0);
		prog_cycle_task(16'b0110011001001011, 1'b0);
		prog_cycle_task(16'b1110011001001011, 1'b1);
		prog_cycle_task(16'b0000000000101011, 1'b0);
		prog_cycle_task(16'b1000000000101011, 1'b0);
		prog_cycle_task(16'b0100000000101011, 1'b0);
		prog_cycle_task(16'b1100000000101011, 1'b0);
		prog_cycle_task(16'b0010000000101011, 1'b0);
		prog_cycle_task(16'b1010000000101011, 1'b0);
		prog_cycle_task(16'b0110000000101011, 1'b0);
		prog_cycle_task(16'b1110000000101011, 1'b1);
		prog_cycle_task(16'b0001000000101011, 1'b0);
		prog_cycle_task(16'b1001000000101011, 1'b0);
		prog_cycle_task(16'b0101000000101011, 1'b0);
		prog_cycle_task(16'b1101000000101011, 1'b0);
		prog_cycle_task(16'b0011000000101011, 1'b0);
		prog_cycle_task(16'b1011000000101011, 1'b0);
		prog_cycle_task(16'b0111000000101011, 1'b0);
		prog_cycle_task(16'b1111000000101011, 1'b1);
		prog_cycle_task(16'b0000100000101011, 1'b0);
		prog_cycle_task(16'b1000100000101011, 1'b0);
		prog_cycle_task(16'b0100100000101011, 1'b1);
		prog_cycle_task(16'b1100100000101011, 1'b0);
		prog_cycle_task(16'b0010100000101011, 1'b0);
		prog_cycle_task(16'b1010100000101011, 1'b1);
		prog_cycle_task(16'b0001100000101011, 1'b0);
		prog_cycle_task(16'b1001100000101011, 1'b0);
		prog_cycle_task(16'b0101100000101011, 1'b0);
		prog_cycle_task(16'b1101100000101011, 1'b0);
		prog_cycle_task(16'b0011100000101011, 1'b0);
		prog_cycle_task(16'b1011100000101011, 1'b0);
		prog_cycle_task(16'b0111100000101011, 1'b0);
		prog_cycle_task(16'b1111100000101011, 1'b1);
		prog_cycle_task(16'b0000010000101011, 1'b0);
		prog_cycle_task(16'b1000010000101011, 1'b0);
		prog_cycle_task(16'b0100010000101011, 1'b0);
		prog_cycle_task(16'b1100010000101011, 1'b0);
		prog_cycle_task(16'b0010010000101011, 1'b0);
		prog_cycle_task(16'b1010010000101011, 1'b0);
		prog_cycle_task(16'b0110010000101011, 1'b0);
		prog_cycle_task(16'b1110010000101011, 1'b1);
		prog_cycle_task(16'b0001010000101011, 1'b0);
		prog_cycle_task(16'b1001010000101011, 1'b0);
		prog_cycle_task(16'b0101010000101011, 1'b1);
		prog_cycle_task(16'b1101010000101011, 1'b0);
		prog_cycle_task(16'b0011010000101011, 1'b0);
		prog_cycle_task(16'b1011010000101011, 1'b1);
		prog_cycle_task(16'b0000110000101011, 1'b0);
		prog_cycle_task(16'b1000110000101011, 1'b0);
		prog_cycle_task(16'b0100110000101011, 1'b0);
		prog_cycle_task(16'b1100110000101011, 1'b0);
		prog_cycle_task(16'b0010110000101011, 1'b0);
		prog_cycle_task(16'b1010110000101011, 1'b0);
		prog_cycle_task(16'b0110110000101011, 1'b0);
		prog_cycle_task(16'b1110110000101011, 1'b1);
		prog_cycle_task(16'b0001110000101011, 1'b0);
		prog_cycle_task(16'b1001110000101011, 1'b0);
		prog_cycle_task(16'b0101110000101011, 1'b0);
		prog_cycle_task(16'b1101110000101011, 1'b0);
		prog_cycle_task(16'b0011110000101011, 1'b0);
		prog_cycle_task(16'b1011110000101011, 1'b0);
		prog_cycle_task(16'b0111110000101011, 1'b0);
		prog_cycle_task(16'b1111110000101011, 1'b1);
		prog_cycle_task(16'b0000001000101011, 1'b0);
		prog_cycle_task(16'b1000001000101011, 1'b0);
		prog_cycle_task(16'b0100001000101011, 1'b1);
		prog_cycle_task(16'b1100001000101011, 1'b0);
		prog_cycle_task(16'b0010001000101011, 1'b0);
		prog_cycle_task(16'b1010001000101011, 1'b1);
		prog_cycle_task(16'b0001001000101011, 1'b0);
		prog_cycle_task(16'b1001001000101011, 1'b0);
		prog_cycle_task(16'b0101001000101011, 1'b0);
		prog_cycle_task(16'b1101001000101011, 1'b0);
		prog_cycle_task(16'b0011001000101011, 1'b0);
		prog_cycle_task(16'b1011001000101011, 1'b0);
		prog_cycle_task(16'b0111001000101011, 1'b0);
		prog_cycle_task(16'b1111001000101011, 1'b1);
		prog_cycle_task(16'b0000101000101011, 1'b0);
		prog_cycle_task(16'b1000101000101011, 1'b0);
		prog_cycle_task(16'b0100101000101011, 1'b0);
		prog_cycle_task(16'b1100101000101011, 1'b0);
		prog_cycle_task(16'b0010101000101011, 1'b0);
		prog_cycle_task(16'b1010101000101011, 1'b0);
		prog_cycle_task(16'b0110101000101011, 1'b0);
		prog_cycle_task(16'b1110101000101011, 1'b1);
		prog_cycle_task(16'b0001101000101011, 1'b0);
		prog_cycle_task(16'b1001101000101011, 1'b0);
		prog_cycle_task(16'b0101101000101011, 1'b1);
		prog_cycle_task(16'b1101101000101011, 1'b0);
		prog_cycle_task(16'b0011101000101011, 1'b0);
		prog_cycle_task(16'b1011101000101011, 1'b1);
		prog_cycle_task(16'b0000000000011011, 1'b0);
		prog_cycle_task(16'b1000000000011011, 1'b0);
		prog_cycle_task(16'b0100000000011011, 1'b0);
		prog_cycle_task(16'b1100000000011011, 1'b0);
		prog_cycle_task(16'b0010000000011011, 1'b0);
		prog_cycle_task(16'b1010000000011011, 1'b1);
		prog_cycle_task(16'b0001000000011011, 1'b0);
		prog_cycle_task(16'b1001000000011011, 1'b0);
		prog_cycle_task(16'b0000100000011011, 1'b0);
		prog_cycle_task(16'b1000100000011011, 1'b0);
		prog_cycle_task(16'b0100100000011011, 1'b0);
		prog_cycle_task(16'b1100100000011011, 1'b0);
		prog_cycle_task(16'b0010100000011011, 1'b0);
		prog_cycle_task(16'b1010100000011011, 1'b1);
		prog_cycle_task(16'b0001100000011011, 1'b0);
		prog_cycle_task(16'b1001100000011011, 1'b0);
		prog_cycle_task(16'b0101100000011011, 1'b0);
		prog_cycle_task(16'b1101100000011011, 1'b0);
		prog_cycle_task(16'b0011100000011011, 1'b0);
		prog_cycle_task(16'b1011100000011011, 1'b1);
		prog_cycle_task(16'b0000010000011011, 1'b0);
		prog_cycle_task(16'b1000010000011011, 1'b0);
		prog_cycle_task(16'b0001010000011011, 1'b0);
		prog_cycle_task(16'b1001010000011011, 1'b0);
		prog_cycle_task(16'b0000000000111011, 1'b0);
		prog_cycle_task(16'b1000000000111011, 1'b0);
		prog_cycle_task(16'b0100000000111011, 1'b0);
		prog_cycle_task(16'b1100000000111011, 1'b0);
		prog_cycle_task(16'b0010000000111011, 1'b0);
		prog_cycle_task(16'b1010000000111011, 1'b1);
		prog_cycle_task(16'b0001000000111011, 1'b0);
		prog_cycle_task(16'b1001000000111011, 1'b0);
		prog_cycle_task(16'b0000100000111011, 1'b0);
		prog_cycle_task(16'b1000100000111011, 1'b0);
		prog_cycle_task(16'b0100100000111011, 1'b0);
		prog_cycle_task(16'b1100100000111011, 1'b0);
		prog_cycle_task(16'b0010100000111011, 1'b0);
		prog_cycle_task(16'b1010100000111011, 1'b1);
		prog_cycle_task(16'b0001100000111011, 1'b0);
		prog_cycle_task(16'b1001100000111011, 1'b0);
		prog_cycle_task(16'b0000010000111011, 1'b0);
		prog_cycle_task(16'b1000010000111011, 1'b0);
		prog_cycle_task(16'b0000000000000111, 1'b0);
		prog_cycle_task(16'b1000000000000111, 1'b0);
		prog_cycle_task(16'b0100000000000111, 1'b0);
		prog_cycle_task(16'b1100000000000111, 1'b0);
		prog_cycle_task(16'b0010000000000111, 1'b0);
		prog_cycle_task(16'b1010000000000111, 1'b0);
		prog_cycle_task(16'b0110000000000111, 1'b0);
		prog_cycle_task(16'b1110000000000111, 1'b0);
		prog_cycle_task(16'b0001000000000111, 1'b0);
		prog_cycle_task(16'b1001000000000111, 1'b0);
		prog_cycle_task(16'b0101000000000111, 1'b0);
		prog_cycle_task(16'b1101000000000111, 1'b0);
		prog_cycle_task(16'b0011000000000111, 1'b0);
		prog_cycle_task(16'b1011000000000111, 1'b0);
		prog_cycle_task(16'b0111000000000111, 1'b0);
		prog_cycle_task(16'b1111000000000111, 1'b0);
		prog_cycle_task(16'b0000100000000111, 1'b0);
		prog_cycle_task(16'b1000100000000111, 1'b0);
		prog_cycle_task(16'b0100100000000111, 1'b1);
		prog_cycle_task(16'b0000010000000111, 1'b0);
		prog_cycle_task(16'b1000010000000111, 1'b0);
		prog_cycle_task(16'b0100010000000111, 1'b0);
		prog_cycle_task(16'b1100010000000111, 1'b0);
		prog_cycle_task(16'b0010010000000111, 1'b0);
		prog_cycle_task(16'b1010010000000111, 1'b0);
		prog_cycle_task(16'b0110010000000111, 1'b0);
		prog_cycle_task(16'b1110010000000111, 1'b0);
		prog_cycle_task(16'b0001010000000111, 1'b0);
		prog_cycle_task(16'b1001010000000111, 1'b0);
		prog_cycle_task(16'b0101010000000111, 1'b0);
		prog_cycle_task(16'b1101010000000111, 1'b0);
		prog_cycle_task(16'b0011010000000111, 1'b0);
		prog_cycle_task(16'b1011010000000111, 1'b0);
		prog_cycle_task(16'b0111010000000111, 1'b0);
		prog_cycle_task(16'b1111010000000111, 1'b0);
		prog_cycle_task(16'b0000110000000111, 1'b0);
		prog_cycle_task(16'b1000110000000111, 1'b0);
		prog_cycle_task(16'b0100110000000111, 1'b1);
		prog_cycle_task(16'b0000001000000111, 1'b0);
		prog_cycle_task(16'b1000001000000111, 1'b0);
		prog_cycle_task(16'b0100001000000111, 1'b0);
		prog_cycle_task(16'b1100001000000111, 1'b0);
		prog_cycle_task(16'b0010001000000111, 1'b0);
		prog_cycle_task(16'b1010001000000111, 1'b0);
		prog_cycle_task(16'b0110001000000111, 1'b0);
		prog_cycle_task(16'b1110001000000111, 1'b0);
		prog_cycle_task(16'b0001001000000111, 1'b0);
		prog_cycle_task(16'b1001001000000111, 1'b0);
		prog_cycle_task(16'b0101001000000111, 1'b0);
		prog_cycle_task(16'b1101001000000111, 1'b0);
		prog_cycle_task(16'b0011001000000111, 1'b0);
		prog_cycle_task(16'b1011001000000111, 1'b0);
		prog_cycle_task(16'b0111001000000111, 1'b0);
		prog_cycle_task(16'b1111001000000111, 1'b0);
		prog_cycle_task(16'b0000101000000111, 1'b0);
		prog_cycle_task(16'b1000101000000111, 1'b0);
		prog_cycle_task(16'b0100101000000111, 1'b1);
		prog_cycle_task(16'b0000011000000111, 1'b0);
		prog_cycle_task(16'b1000011000000111, 1'b0);
		prog_cycle_task(16'b0100011000000111, 1'b0);
		prog_cycle_task(16'b1100011000000111, 1'b0);
		prog_cycle_task(16'b0010011000000111, 1'b0);
		prog_cycle_task(16'b1010011000000111, 1'b0);
		prog_cycle_task(16'b0110011000000111, 1'b0);
		prog_cycle_task(16'b1110011000000111, 1'b0);
		prog_cycle_task(16'b0001011000000111, 1'b0);
		prog_cycle_task(16'b1001011000000111, 1'b0);
		prog_cycle_task(16'b0101011000000111, 1'b0);
		prog_cycle_task(16'b1101011000000111, 1'b0);
		prog_cycle_task(16'b0011011000000111, 1'b0);
		prog_cycle_task(16'b1011011000000111, 1'b0);
		prog_cycle_task(16'b0111011000000111, 1'b0);
		prog_cycle_task(16'b1111011000000111, 1'b0);
		prog_cycle_task(16'b0000111000000111, 1'b0);
		prog_cycle_task(16'b1000111000000111, 1'b0);
		prog_cycle_task(16'b0100111000000111, 1'b1);
		prog_cycle_task(16'b0000000100000111, 1'b0);
		prog_cycle_task(16'b1000000100000111, 1'b0);
		prog_cycle_task(16'b0100000100000111, 1'b1);
		prog_cycle_task(16'b1100000100000111, 1'b0);
		prog_cycle_task(16'b0010000100000111, 1'b0);
		prog_cycle_task(16'b1010000100000111, 1'b0);
		prog_cycle_task(16'b0110000100000111, 1'b0);
		prog_cycle_task(16'b1110000100000111, 1'b1);
		prog_cycle_task(16'b0000010100000111, 1'b0);
		prog_cycle_task(16'b1000010100000111, 1'b0);
		prog_cycle_task(16'b0100010100000111, 1'b1);
		prog_cycle_task(16'b1100010100000111, 1'b0);
		prog_cycle_task(16'b0010010100000111, 1'b0);
		prog_cycle_task(16'b1010010100000111, 1'b0);
		prog_cycle_task(16'b0110010100000111, 1'b0);
		prog_cycle_task(16'b1110010100000111, 1'b1);
		prog_cycle_task(16'b0000001100000111, 1'b0);
		prog_cycle_task(16'b1000001100000111, 1'b0);
		prog_cycle_task(16'b0100001100000111, 1'b1);
		prog_cycle_task(16'b1100001100000111, 1'b0);
		prog_cycle_task(16'b0010001100000111, 1'b0);
		prog_cycle_task(16'b1010001100000111, 1'b0);
		prog_cycle_task(16'b0110001100000111, 1'b0);
		prog_cycle_task(16'b1110001100000111, 1'b1);
		prog_cycle_task(16'b0000011100000111, 1'b0);
		prog_cycle_task(16'b1000011100000111, 1'b0);
		prog_cycle_task(16'b0100011100000111, 1'b1);
		prog_cycle_task(16'b1100011100000111, 1'b0);
		prog_cycle_task(16'b0010011100000111, 1'b0);
		prog_cycle_task(16'b1010011100000111, 1'b0);
		prog_cycle_task(16'b0110011100000111, 1'b0);
		prog_cycle_task(16'b1110011100000111, 1'b1);
		prog_cycle_task(16'b0000000010000111, 1'b0);
		prog_cycle_task(16'b1000000010000111, 1'b0);
		prog_cycle_task(16'b0100000010000111, 1'b1);
		prog_cycle_task(16'b1100000010000111, 1'b0);
		prog_cycle_task(16'b0010000010000111, 1'b0);
		prog_cycle_task(16'b1010000010000111, 1'b0);
		prog_cycle_task(16'b0110000010000111, 1'b0);
		prog_cycle_task(16'b1110000010000111, 1'b1);
		prog_cycle_task(16'b0000010010000111, 1'b0);
		prog_cycle_task(16'b1000010010000111, 1'b0);
		prog_cycle_task(16'b0100010010000111, 1'b1);
		prog_cycle_task(16'b1100010010000111, 1'b0);
		prog_cycle_task(16'b0010010010000111, 1'b0);
		prog_cycle_task(16'b1010010010000111, 1'b0);
		prog_cycle_task(16'b0110010010000111, 1'b0);
		prog_cycle_task(16'b1110010010000111, 1'b1);
		prog_cycle_task(16'b0000001010000111, 1'b0);
		prog_cycle_task(16'b1000001010000111, 1'b0);
		prog_cycle_task(16'b0100001010000111, 1'b1);
		prog_cycle_task(16'b1100001010000111, 1'b0);
		prog_cycle_task(16'b0010001010000111, 1'b0);
		prog_cycle_task(16'b1010001010000111, 1'b0);
		prog_cycle_task(16'b0110001010000111, 1'b0);
		prog_cycle_task(16'b1110001010000111, 1'b1);
		prog_cycle_task(16'b0000011010000111, 1'b0);
		prog_cycle_task(16'b1000011010000111, 1'b0);
		prog_cycle_task(16'b0100011010000111, 1'b1);
		prog_cycle_task(16'b1100011010000111, 1'b0);
		prog_cycle_task(16'b0010011010000111, 1'b0);
		prog_cycle_task(16'b1010011010000111, 1'b0);
		prog_cycle_task(16'b0110011010000111, 1'b0);
		prog_cycle_task(16'b1110011010000111, 1'b1);
		prog_cycle_task(16'b0000000110000111, 1'b0);
		prog_cycle_task(16'b1000000110000111, 1'b0);
		prog_cycle_task(16'b0100000110000111, 1'b1);
		prog_cycle_task(16'b1100000110000111, 1'b0);
		prog_cycle_task(16'b0010000110000111, 1'b0);
		prog_cycle_task(16'b1010000110000111, 1'b0);
		prog_cycle_task(16'b0110000110000111, 1'b0);
		prog_cycle_task(16'b1110000110000111, 1'b1);
		prog_cycle_task(16'b0000010110000111, 1'b0);
		prog_cycle_task(16'b1000010110000111, 1'b0);
		prog_cycle_task(16'b0100010110000111, 1'b1);
		prog_cycle_task(16'b1100010110000111, 1'b0);
		prog_cycle_task(16'b0010010110000111, 1'b0);
		prog_cycle_task(16'b1010010110000111, 1'b0);
		prog_cycle_task(16'b0110010110000111, 1'b0);
		prog_cycle_task(16'b1110010110000111, 1'b1);
		prog_cycle_task(16'b0000001110000111, 1'b0);
		prog_cycle_task(16'b1000001110000111, 1'b0);
		prog_cycle_task(16'b0100001110000111, 1'b1);
		prog_cycle_task(16'b1100001110000111, 1'b0);
		prog_cycle_task(16'b0010001110000111, 1'b0);
		prog_cycle_task(16'b1010001110000111, 1'b0);
		prog_cycle_task(16'b0110001110000111, 1'b0);
		prog_cycle_task(16'b1110001110000111, 1'b1);
		prog_cycle_task(16'b0000011110000111, 1'b0);
		prog_cycle_task(16'b1000011110000111, 1'b0);
		prog_cycle_task(16'b0100011110000111, 1'b1);
		prog_cycle_task(16'b1100011110000111, 1'b0);
		prog_cycle_task(16'b0010011110000111, 1'b0);
		prog_cycle_task(16'b1010011110000111, 1'b0);
		prog_cycle_task(16'b0110011110000111, 1'b0);
		prog_cycle_task(16'b1110011110000111, 1'b1);
		prog_cycle_task(16'b0000000001000111, 1'b0);
		prog_cycle_task(16'b1000000001000111, 1'b0);
		prog_cycle_task(16'b0100000001000111, 1'b1);
		prog_cycle_task(16'b1100000001000111, 1'b0);
		prog_cycle_task(16'b0010000001000111, 1'b0);
		prog_cycle_task(16'b1010000001000111, 1'b0);
		prog_cycle_task(16'b0110000001000111, 1'b0);
		prog_cycle_task(16'b1110000001000111, 1'b1);
		prog_cycle_task(16'b0000010001000111, 1'b0);
		prog_cycle_task(16'b1000010001000111, 1'b0);
		prog_cycle_task(16'b0100010001000111, 1'b1);
		prog_cycle_task(16'b1100010001000111, 1'b0);
		prog_cycle_task(16'b0010010001000111, 1'b0);
		prog_cycle_task(16'b1010010001000111, 1'b0);
		prog_cycle_task(16'b0110010001000111, 1'b0);
		prog_cycle_task(16'b1110010001000111, 1'b1);
		prog_cycle_task(16'b0000001001000111, 1'b0);
		prog_cycle_task(16'b1000001001000111, 1'b0);
		prog_cycle_task(16'b0100001001000111, 1'b1);
		prog_cycle_task(16'b1100001001000111, 1'b0);
		prog_cycle_task(16'b0010001001000111, 1'b0);
		prog_cycle_task(16'b1010001001000111, 1'b0);
		prog_cycle_task(16'b0110001001000111, 1'b0);
		prog_cycle_task(16'b1110001001000111, 1'b1);
		prog_cycle_task(16'b0000011001000111, 1'b0);
		prog_cycle_task(16'b1000011001000111, 1'b0);
		prog_cycle_task(16'b0100011001000111, 1'b1);
		prog_cycle_task(16'b1100011001000111, 1'b0);
		prog_cycle_task(16'b0010011001000111, 1'b0);
		prog_cycle_task(16'b1010011001000111, 1'b0);
		prog_cycle_task(16'b0110011001000111, 1'b0);
		prog_cycle_task(16'b1110011001000111, 1'b1);
		prog_cycle_task(16'b0000000000100111, 1'b0);
		prog_cycle_task(16'b1000000000100111, 1'b0);
		prog_cycle_task(16'b0100000000100111, 1'b1);
		prog_cycle_task(16'b1100000000100111, 1'b0);
		prog_cycle_task(16'b0010000000100111, 1'b0);
		prog_cycle_task(16'b1010000000100111, 1'b1);
		prog_cycle_task(16'b0001000000100111, 1'b0);
		prog_cycle_task(16'b1001000000100111, 1'b0);
		prog_cycle_task(16'b0101000000100111, 1'b1);
		prog_cycle_task(16'b1101000000100111, 1'b0);
		prog_cycle_task(16'b0011000000100111, 1'b0);
		prog_cycle_task(16'b1011000000100111, 1'b1);
		prog_cycle_task(16'b0000100000100111, 1'b0);
		prog_cycle_task(16'b1000100000100111, 1'b0);
		prog_cycle_task(16'b0100100000100111, 1'b1);
		prog_cycle_task(16'b1100100000100111, 1'b0);
		prog_cycle_task(16'b0010100000100111, 1'b0);
		prog_cycle_task(16'b1010100000100111, 1'b1);
		prog_cycle_task(16'b0001100000100111, 1'b0);
		prog_cycle_task(16'b1001100000100111, 1'b0);
		prog_cycle_task(16'b0101100000100111, 1'b1);
		prog_cycle_task(16'b1101100000100111, 1'b0);
		prog_cycle_task(16'b0011100000100111, 1'b0);
		prog_cycle_task(16'b1011100000100111, 1'b1);
		prog_cycle_task(16'b0000010000100111, 1'b0);
		prog_cycle_task(16'b1000010000100111, 1'b0);
		prog_cycle_task(16'b0100010000100111, 1'b1);
		prog_cycle_task(16'b1100010000100111, 1'b0);
		prog_cycle_task(16'b0010010000100111, 1'b0);
		prog_cycle_task(16'b1010010000100111, 1'b1);
		prog_cycle_task(16'b0001010000100111, 1'b0);
		prog_cycle_task(16'b1001010000100111, 1'b0);
		prog_cycle_task(16'b0101010000100111, 1'b1);
		prog_cycle_task(16'b1101010000100111, 1'b0);
		prog_cycle_task(16'b0011010000100111, 1'b0);
		prog_cycle_task(16'b1011010000100111, 1'b1);
		prog_cycle_task(16'b0000110000100111, 1'b0);
		prog_cycle_task(16'b1000110000100111, 1'b0);
		prog_cycle_task(16'b0001110000100111, 1'b0);
		prog_cycle_task(16'b1001110000100111, 1'b0);
		prog_cycle_task(16'b0000001000100111, 1'b0);
		prog_cycle_task(16'b1000001000100111, 1'b0);
		prog_cycle_task(16'b0001001000100111, 1'b0);
		prog_cycle_task(16'b1001001000100111, 1'b0);
		prog_cycle_task(16'b0000101000100111, 1'b0);
		prog_cycle_task(16'b1000101000100111, 1'b0);
		prog_cycle_task(16'b0001101000100111, 1'b0);
		prog_cycle_task(16'b1001101000100111, 1'b0);
		prog_cycle_task(16'b0000011000100111, 1'b0);
		prog_cycle_task(16'b1000011000100111, 1'b0);
		prog_cycle_task(16'b0001011000100111, 1'b0);
		prog_cycle_task(16'b1001011000100111, 1'b0);
		prog_cycle_task(16'b0000111000100111, 1'b0);
		prog_cycle_task(16'b1000111000100111, 1'b0);
		prog_cycle_task(16'b0000000000010111, 1'b0);
		prog_cycle_task(16'b1000000000010111, 1'b0);
		prog_cycle_task(16'b0100000000010111, 1'b0);
		prog_cycle_task(16'b1100000000010111, 1'b0);
		prog_cycle_task(16'b0010000000010111, 1'b0);
		prog_cycle_task(16'b1010000000010111, 1'b1);
		prog_cycle_task(16'b0001000000010111, 1'b0);
		prog_cycle_task(16'b1001000000010111, 1'b0);
		prog_cycle_task(16'b0000100000010111, 1'b0);
		prog_cycle_task(16'b1000100000010111, 1'b0);
		prog_cycle_task(16'b0100100000010111, 1'b0);
		prog_cycle_task(16'b1100100000010111, 1'b0);
		prog_cycle_task(16'b0010100000010111, 1'b0);
		prog_cycle_task(16'b1010100000010111, 1'b1);
		prog_cycle_task(16'b0001100000010111, 1'b0);
		prog_cycle_task(16'b1001100000010111, 1'b0);
		prog_cycle_task(16'b0101100000010111, 1'b0);
		prog_cycle_task(16'b1101100000010111, 1'b0);
		prog_cycle_task(16'b0011100000010111, 1'b0);
		prog_cycle_task(16'b1011100000010111, 1'b1);
		prog_cycle_task(16'b0000010000010111, 1'b0);
		prog_cycle_task(16'b1000010000010111, 1'b0);
		prog_cycle_task(16'b0001010000010111, 1'b0);
		prog_cycle_task(16'b1001010000010111, 1'b0);
		prog_cycle_task(16'b0000000000110111, 1'b0);
		prog_cycle_task(16'b1000000000110111, 1'b0);
		prog_cycle_task(16'b0100000000110111, 1'b0);
		prog_cycle_task(16'b1100000000110111, 1'b0);
		prog_cycle_task(16'b0010000000110111, 1'b0);
		prog_cycle_task(16'b1010000000110111, 1'b1);
		prog_cycle_task(16'b0001000000110111, 1'b0);
		prog_cycle_task(16'b1001000000110111, 1'b0);
		prog_cycle_task(16'b0101000000110111, 1'b0);
		prog_cycle_task(16'b1101000000110111, 1'b0);
		prog_cycle_task(16'b0011000000110111, 1'b0);
		prog_cycle_task(16'b1011000000110111, 1'b1);
		prog_cycle_task(16'b0000100000110111, 1'b0);
		prog_cycle_task(16'b1000100000110111, 1'b0);
		prog_cycle_task(16'b0100100000110111, 1'b0);
		prog_cycle_task(16'b1100100000110111, 1'b0);
		prog_cycle_task(16'b0010100000110111, 1'b0);
		prog_cycle_task(16'b1010100000110111, 1'b1);
		prog_cycle_task(16'b0001100000110111, 1'b0);
		prog_cycle_task(16'b1001100000110111, 1'b0);
		prog_cycle_task(16'b0101100000110111, 1'b0);
		prog_cycle_task(16'b1101100000110111, 1'b0);
		prog_cycle_task(16'b0011100000110111, 1'b0);
		prog_cycle_task(16'b1011100000110111, 1'b1);
		prog_cycle_task(16'b0000010000110111, 1'b0);
		prog_cycle_task(16'b1000010000110111, 1'b0);
		prog_cycle_task(16'b0100010000110111, 1'b0);
		prog_cycle_task(16'b1100010000110111, 1'b0);
		prog_cycle_task(16'b0010010000110111, 1'b0);
		prog_cycle_task(16'b1010010000110111, 1'b1);
		prog_cycle_task(16'b0001010000110111, 1'b0);
		prog_cycle_task(16'b1001010000110111, 1'b0);
		prog_cycle_task(16'b0101010000110111, 1'b0);
		prog_cycle_task(16'b1101010000110111, 1'b0);
		prog_cycle_task(16'b0011010000110111, 1'b0);
		prog_cycle_task(16'b1011010000110111, 1'b1);
		prog_cycle_task(16'b0000110000110111, 1'b0);
		prog_cycle_task(16'b1000110000110111, 1'b0);
		prog_cycle_task(16'b0100110000110111, 1'b0);
		prog_cycle_task(16'b1100110000110111, 1'b0);
		prog_cycle_task(16'b0010110000110111, 1'b0);
		prog_cycle_task(16'b1010110000110111, 1'b1);
		prog_cycle_task(16'b0001110000110111, 1'b0);
		prog_cycle_task(16'b1001110000110111, 1'b0);
		prog_cycle_task(16'b0101110000110111, 1'b0);
		prog_cycle_task(16'b1101110000110111, 1'b0);
		prog_cycle_task(16'b0011110000110111, 1'b0);
		prog_cycle_task(16'b1011110000110111, 1'b1);
		prog_cycle_task(16'b0000001000110111, 1'b0);
		prog_cycle_task(16'b1000001000110111, 1'b0);
		prog_cycle_task(16'b0100001000110111, 1'b0);
		prog_cycle_task(16'b1100001000110111, 1'b0);
		prog_cycle_task(16'b0010001000110111, 1'b0);
		prog_cycle_task(16'b1010001000110111, 1'b1);
		prog_cycle_task(16'b0001001000110111, 1'b0);
		prog_cycle_task(16'b1001001000110111, 1'b0);
		prog_cycle_task(16'b0000101000110111, 1'b0);
		prog_cycle_task(16'b1000101000110111, 1'b0);
		prog_cycle_task(16'b0000000000001111, 1'b0);
		prog_cycle_task(16'b1000000000001111, 1'b0);
		prog_cycle_task(16'b0100000000001111, 1'b0);
		prog_cycle_task(16'b1100000000001111, 1'b0);
		prog_cycle_task(16'b0010000000001111, 1'b0);
		prog_cycle_task(16'b1010000000001111, 1'b0);
		prog_cycle_task(16'b0110000000001111, 1'b0);
		prog_cycle_task(16'b1110000000001111, 1'b0);
		prog_cycle_task(16'b0001000000001111, 1'b0);
		prog_cycle_task(16'b1001000000001111, 1'b0);
		prog_cycle_task(16'b0101000000001111, 1'b0);
		prog_cycle_task(16'b1101000000001111, 1'b0);
		prog_cycle_task(16'b0011000000001111, 1'b0);
		prog_cycle_task(16'b1011000000001111, 1'b0);
		prog_cycle_task(16'b0111000000001111, 1'b0);
		prog_cycle_task(16'b1111000000001111, 1'b0);
		prog_cycle_task(16'b0000100000001111, 1'b0);
		prog_cycle_task(16'b1000100000001111, 1'b0);
		prog_cycle_task(16'b0100100000001111, 1'b1);
		prog_cycle_task(16'b0000010000001111, 1'b0);
		prog_cycle_task(16'b1000010000001111, 1'b0);
		prog_cycle_task(16'b0100010000001111, 1'b0);
		prog_cycle_task(16'b1100010000001111, 1'b0);
		prog_cycle_task(16'b0010010000001111, 1'b0);
		prog_cycle_task(16'b1010010000001111, 1'b0);
		prog_cycle_task(16'b0110010000001111, 1'b0);
		prog_cycle_task(16'b1110010000001111, 1'b0);
		prog_cycle_task(16'b0001010000001111, 1'b0);
		prog_cycle_task(16'b1001010000001111, 1'b0);
		prog_cycle_task(16'b0101010000001111, 1'b0);
		prog_cycle_task(16'b1101010000001111, 1'b0);
		prog_cycle_task(16'b0011010000001111, 1'b0);
		prog_cycle_task(16'b1011010000001111, 1'b0);
		prog_cycle_task(16'b0111010000001111, 1'b0);
		prog_cycle_task(16'b1111010000001111, 1'b0);
		prog_cycle_task(16'b0000110000001111, 1'b0);
		prog_cycle_task(16'b1000110000001111, 1'b0);
		prog_cycle_task(16'b0100110000001111, 1'b1);
		prog_cycle_task(16'b0000001000001111, 1'b0);
		prog_cycle_task(16'b1000001000001111, 1'b0);
		prog_cycle_task(16'b0100001000001111, 1'b0);
		prog_cycle_task(16'b1100001000001111, 1'b0);
		prog_cycle_task(16'b0010001000001111, 1'b0);
		prog_cycle_task(16'b1010001000001111, 1'b0);
		prog_cycle_task(16'b0110001000001111, 1'b0);
		prog_cycle_task(16'b1110001000001111, 1'b0);
		prog_cycle_task(16'b0001001000001111, 1'b0);
		prog_cycle_task(16'b1001001000001111, 1'b0);
		prog_cycle_task(16'b0101001000001111, 1'b0);
		prog_cycle_task(16'b1101001000001111, 1'b0);
		prog_cycle_task(16'b0011001000001111, 1'b0);
		prog_cycle_task(16'b1011001000001111, 1'b0);
		prog_cycle_task(16'b0111001000001111, 1'b0);
		prog_cycle_task(16'b1111001000001111, 1'b0);
		prog_cycle_task(16'b0000101000001111, 1'b0);
		prog_cycle_task(16'b1000101000001111, 1'b0);
		prog_cycle_task(16'b0100101000001111, 1'b1);
		prog_cycle_task(16'b0000011000001111, 1'b0);
		prog_cycle_task(16'b1000011000001111, 1'b0);
		prog_cycle_task(16'b0100011000001111, 1'b0);
		prog_cycle_task(16'b1100011000001111, 1'b0);
		prog_cycle_task(16'b0010011000001111, 1'b0);
		prog_cycle_task(16'b1010011000001111, 1'b0);
		prog_cycle_task(16'b0110011000001111, 1'b0);
		prog_cycle_task(16'b1110011000001111, 1'b0);
		prog_cycle_task(16'b0001011000001111, 1'b0);
		prog_cycle_task(16'b1001011000001111, 1'b0);
		prog_cycle_task(16'b0101011000001111, 1'b0);
		prog_cycle_task(16'b1101011000001111, 1'b0);
		prog_cycle_task(16'b0011011000001111, 1'b0);
		prog_cycle_task(16'b1011011000001111, 1'b0);
		prog_cycle_task(16'b0111011000001111, 1'b0);
		prog_cycle_task(16'b1111011000001111, 1'b0);
		prog_cycle_task(16'b0000111000001111, 1'b0);
		prog_cycle_task(16'b1000111000001111, 1'b0);
		prog_cycle_task(16'b0100111000001111, 1'b1);
		prog_cycle_task(16'b0000000100001111, 1'b0);
		prog_cycle_task(16'b1000000100001111, 1'b0);
		prog_cycle_task(16'b0100000100001111, 1'b1);
		prog_cycle_task(16'b1100000100001111, 1'b0);
		prog_cycle_task(16'b0010000100001111, 1'b0);
		prog_cycle_task(16'b1010000100001111, 1'b0);
		prog_cycle_task(16'b0110000100001111, 1'b0);
		prog_cycle_task(16'b1110000100001111, 1'b1);
		prog_cycle_task(16'b0000010100001111, 1'b0);
		prog_cycle_task(16'b1000010100001111, 1'b0);
		prog_cycle_task(16'b0100010100001111, 1'b1);
		prog_cycle_task(16'b1100010100001111, 1'b0);
		prog_cycle_task(16'b0010010100001111, 1'b0);
		prog_cycle_task(16'b1010010100001111, 1'b0);
		prog_cycle_task(16'b0110010100001111, 1'b0);
		prog_cycle_task(16'b1110010100001111, 1'b1);
		prog_cycle_task(16'b0000001100001111, 1'b0);
		prog_cycle_task(16'b1000001100001111, 1'b0);
		prog_cycle_task(16'b0100001100001111, 1'b1);
		prog_cycle_task(16'b1100001100001111, 1'b0);
		prog_cycle_task(16'b0010001100001111, 1'b0);
		prog_cycle_task(16'b1010001100001111, 1'b0);
		prog_cycle_task(16'b0110001100001111, 1'b0);
		prog_cycle_task(16'b1110001100001111, 1'b1);
		prog_cycle_task(16'b0000011100001111, 1'b0);
		prog_cycle_task(16'b1000011100001111, 1'b0);
		prog_cycle_task(16'b0100011100001111, 1'b1);
		prog_cycle_task(16'b1100011100001111, 1'b0);
		prog_cycle_task(16'b0010011100001111, 1'b0);
		prog_cycle_task(16'b1010011100001111, 1'b0);
		prog_cycle_task(16'b0110011100001111, 1'b0);
		prog_cycle_task(16'b1110011100001111, 1'b1);
		prog_cycle_task(16'b0000000010001111, 1'b0);
		prog_cycle_task(16'b1000000010001111, 1'b0);
		prog_cycle_task(16'b0100000010001111, 1'b1);
		prog_cycle_task(16'b1100000010001111, 1'b0);
		prog_cycle_task(16'b0010000010001111, 1'b0);
		prog_cycle_task(16'b1010000010001111, 1'b0);
		prog_cycle_task(16'b0110000010001111, 1'b0);
		prog_cycle_task(16'b1110000010001111, 1'b1);
		prog_cycle_task(16'b0000010010001111, 1'b0);
		prog_cycle_task(16'b1000010010001111, 1'b0);
		prog_cycle_task(16'b0100010010001111, 1'b1);
		prog_cycle_task(16'b1100010010001111, 1'b0);
		prog_cycle_task(16'b0010010010001111, 1'b0);
		prog_cycle_task(16'b1010010010001111, 1'b0);
		prog_cycle_task(16'b0110010010001111, 1'b0);
		prog_cycle_task(16'b1110010010001111, 1'b1);
		prog_cycle_task(16'b0000001010001111, 1'b0);
		prog_cycle_task(16'b1000001010001111, 1'b0);
		prog_cycle_task(16'b0100001010001111, 1'b1);
		prog_cycle_task(16'b1100001010001111, 1'b0);
		prog_cycle_task(16'b0010001010001111, 1'b0);
		prog_cycle_task(16'b1010001010001111, 1'b0);
		prog_cycle_task(16'b0110001010001111, 1'b0);
		prog_cycle_task(16'b1110001010001111, 1'b1);
		prog_cycle_task(16'b0000011010001111, 1'b0);
		prog_cycle_task(16'b1000011010001111, 1'b0);
		prog_cycle_task(16'b0100011010001111, 1'b1);
		prog_cycle_task(16'b1100011010001111, 1'b0);
		prog_cycle_task(16'b0010011010001111, 1'b0);
		prog_cycle_task(16'b1010011010001111, 1'b0);
		prog_cycle_task(16'b0110011010001111, 1'b0);
		prog_cycle_task(16'b1110011010001111, 1'b1);
		prog_cycle_task(16'b0000000110001111, 1'b0);
		prog_cycle_task(16'b1000000110001111, 1'b0);
		prog_cycle_task(16'b0100000110001111, 1'b1);
		prog_cycle_task(16'b1100000110001111, 1'b0);
		prog_cycle_task(16'b0010000110001111, 1'b0);
		prog_cycle_task(16'b1010000110001111, 1'b0);
		prog_cycle_task(16'b0110000110001111, 1'b0);
		prog_cycle_task(16'b1110000110001111, 1'b1);
		prog_cycle_task(16'b0000010110001111, 1'b0);
		prog_cycle_task(16'b1000010110001111, 1'b0);
		prog_cycle_task(16'b0100010110001111, 1'b1);
		prog_cycle_task(16'b1100010110001111, 1'b0);
		prog_cycle_task(16'b0010010110001111, 1'b0);
		prog_cycle_task(16'b1010010110001111, 1'b0);
		prog_cycle_task(16'b0110010110001111, 1'b0);
		prog_cycle_task(16'b1110010110001111, 1'b1);
		prog_cycle_task(16'b0000001110001111, 1'b0);
		prog_cycle_task(16'b1000001110001111, 1'b0);
		prog_cycle_task(16'b0100001110001111, 1'b1);
		prog_cycle_task(16'b1100001110001111, 1'b0);
		prog_cycle_task(16'b0010001110001111, 1'b0);
		prog_cycle_task(16'b1010001110001111, 1'b0);
		prog_cycle_task(16'b0110001110001111, 1'b0);
		prog_cycle_task(16'b1110001110001111, 1'b1);
		prog_cycle_task(16'b0000011110001111, 1'b0);
		prog_cycle_task(16'b1000011110001111, 1'b0);
		prog_cycle_task(16'b0100011110001111, 1'b1);
		prog_cycle_task(16'b1100011110001111, 1'b0);
		prog_cycle_task(16'b0010011110001111, 1'b0);
		prog_cycle_task(16'b1010011110001111, 1'b0);
		prog_cycle_task(16'b0110011110001111, 1'b0);
		prog_cycle_task(16'b1110011110001111, 1'b1);
		prog_cycle_task(16'b0000000001001111, 1'b0);
		prog_cycle_task(16'b1000000001001111, 1'b0);
		prog_cycle_task(16'b0100000001001111, 1'b1);
		prog_cycle_task(16'b1100000001001111, 1'b0);
		prog_cycle_task(16'b0010000001001111, 1'b0);
		prog_cycle_task(16'b1010000001001111, 1'b0);
		prog_cycle_task(16'b0110000001001111, 1'b0);
		prog_cycle_task(16'b1110000001001111, 1'b1);
		prog_cycle_task(16'b0000010001001111, 1'b0);
		prog_cycle_task(16'b1000010001001111, 1'b0);
		prog_cycle_task(16'b0100010001001111, 1'b1);
		prog_cycle_task(16'b1100010001001111, 1'b0);
		prog_cycle_task(16'b0010010001001111, 1'b0);
		prog_cycle_task(16'b1010010001001111, 1'b0);
		prog_cycle_task(16'b0110010001001111, 1'b0);
		prog_cycle_task(16'b1110010001001111, 1'b1);
		prog_cycle_task(16'b0000001001001111, 1'b0);
		prog_cycle_task(16'b1000001001001111, 1'b0);
		prog_cycle_task(16'b0100001001001111, 1'b1);
		prog_cycle_task(16'b1100001001001111, 1'b0);
		prog_cycle_task(16'b0010001001001111, 1'b0);
		prog_cycle_task(16'b1010001001001111, 1'b0);
		prog_cycle_task(16'b0110001001001111, 1'b0);
		prog_cycle_task(16'b1110001001001111, 1'b1);
		prog_cycle_task(16'b0000011001001111, 1'b0);
		prog_cycle_task(16'b1000011001001111, 1'b0);
		prog_cycle_task(16'b0100011001001111, 1'b1);
		prog_cycle_task(16'b1100011001001111, 1'b0);
		prog_cycle_task(16'b0010011001001111, 1'b0);
		prog_cycle_task(16'b1010011001001111, 1'b0);
		prog_cycle_task(16'b0110011001001111, 1'b0);
		prog_cycle_task(16'b1110011001001111, 1'b1);
		prog_cycle_task(16'b0000000000000000, 1'b0);
		@(negedge prog_clock[0]);
			config_done[0] <= 1'b1;
	end
// ----- End bitstream loading during configuration phase -----
// ----- Input Initialization -------
	initial begin
		a <= 1'b0;
		b <= 1'b0;

		out_c_flag[0] <= 1'b0;
	end

// ----- Input Stimulus -------
	always@(negedge op_clock[0]) begin
		a <= $random;
		b <= $random;
	end

`ifdef AUTOCHECKED_SIMULATION
// ----- Begin checking output vectors -------
// ----- Skip the first falling edge of clock, it is for initialization -------
	reg [0:0] sim_start;

	always@(negedge op_clock[0]) begin
		if (1'b1 == sim_start[0]) begin
			sim_start[0] <= ~sim_start[0];
		end else begin
			if(!(out_c_fpga === out_c_benchmark) && !(out_c_benchmark === 1'bx)) begin
				out_c_flag <= 1'b1;
			end else begin
				out_c_flag<= 1'b0;
			end
		end
	end

	always@(posedge out_c_flag) begin
		if(out_c_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_c_fpga at time = %t", $realtime);
		end
	end

`endif

`ifdef AUTOCHECKED_SIMULATION
// ----- Configuration done must be raised in the end -------
	always@(posedge config_done[0]) begin
		nb_error = nb_error - 1;
	end
`endif

`ifdef ICARUS_SIMULATOR
// ----- Begin Icarus requirement -------
	initial begin
		$dumpfile("and2_formal.vcd");
		$dumpvars(1, and2_autocheck_top_tb);
	end
`endif
// ----- END Icarus requirement -------

initial begin
	sim_start[0] <= 1'b1;
	$timeformat(-9, 2, "ns", 20);
	$display("Simulation start");
// ----- Can be changed by the user for his/her need -------
	#38091
	if(nb_error == 0) begin
		$display("Simulation Succeed");
	end else begin
		$display("Simulation Failed with %d error(s)", nb_error);
	end
	$finish;
end

endmodule
// ----- END Verilog module for and2_autocheck_top_tb -----

