magic
tech sky130A
magscale 1 2
timestamp 1606226535
<< locali >>
rect 10609 8347 10643 8585
rect 19073 6171 19107 6409
rect 17601 3451 17635 3689
rect 15025 2839 15059 3009
rect 17141 2839 17175 3145
<< viali >>
rect 20729 20009 20763 20043
rect 20545 19873 20579 19907
rect 20177 19465 20211 19499
rect 20729 19465 20763 19499
rect 12449 19261 12483 19295
rect 19993 19261 20027 19295
rect 20545 19261 20579 19295
rect 12633 19125 12667 19159
rect 20453 18921 20487 18955
rect 10149 18853 10183 18887
rect 11713 18853 11747 18887
rect 17386 18853 17420 18887
rect 7757 18785 7791 18819
rect 8677 18785 8711 18819
rect 9873 18785 9907 18819
rect 11437 18785 11471 18819
rect 20269 18785 20303 18819
rect 8033 18717 8067 18751
rect 8953 18717 8987 18751
rect 17141 18717 17175 18751
rect 18521 18581 18555 18615
rect 15301 18377 15335 18411
rect 20729 18309 20763 18343
rect 12725 18241 12759 18275
rect 12449 18173 12483 18207
rect 15117 18173 15151 18207
rect 20545 18173 20579 18207
rect 20453 17833 20487 17867
rect 14565 17765 14599 17799
rect 14289 17697 14323 17731
rect 20269 17697 20303 17731
rect 20729 17289 20763 17323
rect 19993 17153 20027 17187
rect 19717 17085 19751 17119
rect 20545 17085 20579 17119
rect 19993 16677 20027 16711
rect 19717 16609 19751 16643
rect 20177 16201 20211 16235
rect 20729 16201 20763 16235
rect 12725 16065 12759 16099
rect 12449 15997 12483 16031
rect 19993 15997 20027 16031
rect 20545 15997 20579 16031
rect 20453 15657 20487 15691
rect 10517 15521 10551 15555
rect 20269 15521 20303 15555
rect 10793 15453 10827 15487
rect 20177 15113 20211 15147
rect 20729 15045 20763 15079
rect 9873 14909 9907 14943
rect 19993 14909 20027 14943
rect 20545 14909 20579 14943
rect 10149 14841 10183 14875
rect 20453 14569 20487 14603
rect 8217 14501 8251 14535
rect 7941 14433 7975 14467
rect 11621 14433 11655 14467
rect 20269 14433 20303 14467
rect 11805 14365 11839 14399
rect 20729 13957 20763 13991
rect 19993 13889 20027 13923
rect 19717 13821 19751 13855
rect 20545 13821 20579 13855
rect 19349 13481 19383 13515
rect 19993 13413 20027 13447
rect 19165 13345 19199 13379
rect 19717 13345 19751 13379
rect 20729 12937 20763 12971
rect 16681 12801 16715 12835
rect 19809 12801 19843 12835
rect 19625 12733 19659 12767
rect 20545 12733 20579 12767
rect 16129 12597 16163 12631
rect 16497 12597 16531 12631
rect 16589 12597 16623 12631
rect 16037 12393 16071 12427
rect 19441 12325 19475 12359
rect 20177 12325 20211 12359
rect 15945 12257 15979 12291
rect 16856 12257 16890 12291
rect 18613 12257 18647 12291
rect 19165 12257 19199 12291
rect 19901 12257 19935 12291
rect 16221 12189 16255 12223
rect 16589 12189 16623 12223
rect 15577 12053 15611 12087
rect 17969 12053 18003 12087
rect 18797 12053 18831 12087
rect 16865 11849 16899 11883
rect 20729 11849 20763 11883
rect 13645 11713 13679 11747
rect 15025 11713 15059 11747
rect 18061 11713 18095 11747
rect 15485 11645 15519 11679
rect 15752 11645 15786 11679
rect 19809 11645 19843 11679
rect 20545 11645 20579 11679
rect 18306 11577 18340 11611
rect 20085 11577 20119 11611
rect 13093 11509 13127 11543
rect 13461 11509 13495 11543
rect 13553 11509 13587 11543
rect 19441 11509 19475 11543
rect 16681 11305 16715 11339
rect 17693 11305 17727 11339
rect 18245 11305 18279 11339
rect 18705 11305 18739 11339
rect 12725 11237 12759 11271
rect 20177 11237 20211 11271
rect 11989 11169 12023 11203
rect 15117 11169 15151 11203
rect 15301 11169 15335 11203
rect 15568 11169 15602 11203
rect 17601 11169 17635 11203
rect 18613 11169 18647 11203
rect 19349 11169 19383 11203
rect 19901 11169 19935 11203
rect 12265 11101 12299 11135
rect 14381 11101 14415 11135
rect 17877 11101 17911 11135
rect 18797 11101 18831 11135
rect 14933 11033 14967 11067
rect 19533 11033 19567 11067
rect 17233 10965 17267 10999
rect 10977 10761 11011 10795
rect 16405 10761 16439 10795
rect 16681 10761 16715 10795
rect 19441 10761 19475 10795
rect 20913 10761 20947 10795
rect 11621 10625 11655 10659
rect 12909 10625 12943 10659
rect 15025 10625 15059 10659
rect 17233 10625 17267 10659
rect 18061 10625 18095 10659
rect 20269 10625 20303 10659
rect 13369 10557 13403 10591
rect 20085 10557 20119 10591
rect 20729 10557 20763 10591
rect 13636 10489 13670 10523
rect 15270 10489 15304 10523
rect 17141 10489 17175 10523
rect 18328 10489 18362 10523
rect 11345 10421 11379 10455
rect 11437 10421 11471 10455
rect 14749 10421 14783 10455
rect 17049 10421 17083 10455
rect 19717 10421 19751 10455
rect 20177 10421 20211 10455
rect 10793 10217 10827 10251
rect 12633 10217 12667 10251
rect 14289 10217 14323 10251
rect 15301 10217 15335 10251
rect 16313 10217 16347 10251
rect 17877 10217 17911 10251
rect 11520 10149 11554 10183
rect 13154 10149 13188 10183
rect 15761 10149 15795 10183
rect 19064 10149 19098 10183
rect 12909 10081 12943 10115
rect 14749 10081 14783 10115
rect 15669 10081 15703 10115
rect 16865 10081 16899 10115
rect 18797 10081 18831 10115
rect 11253 10013 11287 10047
rect 15853 10013 15887 10047
rect 17049 10013 17083 10047
rect 18337 10013 18371 10047
rect 14565 9877 14599 9911
rect 20177 9877 20211 9911
rect 11621 9673 11655 9707
rect 12725 9605 12759 9639
rect 16497 9605 16531 9639
rect 13277 9537 13311 9571
rect 17049 9537 17083 9571
rect 18797 9537 18831 9571
rect 10241 9469 10275 9503
rect 13093 9469 13127 9503
rect 18245 9469 18279 9503
rect 19064 9469 19098 9503
rect 20545 9469 20579 9503
rect 10508 9401 10542 9435
rect 16865 9401 16899 9435
rect 17509 9401 17543 9435
rect 9597 9333 9631 9367
rect 13185 9333 13219 9367
rect 16957 9333 16991 9367
rect 18429 9333 18463 9367
rect 20177 9333 20211 9367
rect 20729 9333 20763 9367
rect 8585 9129 8619 9163
rect 8953 9129 8987 9163
rect 9045 9129 9079 9163
rect 11069 9129 11103 9163
rect 14197 9129 14231 9163
rect 18521 9129 18555 9163
rect 18613 9129 18647 9163
rect 9956 8993 9990 9027
rect 11989 8993 12023 9027
rect 14565 8993 14599 9027
rect 15669 8993 15703 9027
rect 15936 8993 15970 9027
rect 17417 8993 17451 9027
rect 19432 8993 19466 9027
rect 9229 8925 9263 8959
rect 9689 8925 9723 8959
rect 14657 8925 14691 8959
rect 14749 8925 14783 8959
rect 17601 8925 17635 8959
rect 18797 8925 18831 8959
rect 19165 8925 19199 8959
rect 18153 8857 18187 8891
rect 11805 8789 11839 8823
rect 17049 8789 17083 8823
rect 20545 8789 20579 8823
rect 10609 8585 10643 8619
rect 10701 8585 10735 8619
rect 14749 8585 14783 8619
rect 16405 8585 16439 8619
rect 16681 8585 16715 8619
rect 8585 8449 8619 8483
rect 11253 8449 11287 8483
rect 17233 8449 17267 8483
rect 19625 8449 19659 8483
rect 20545 8449 20579 8483
rect 13369 8381 13403 8415
rect 15025 8381 15059 8415
rect 15281 8381 15315 8415
rect 17049 8381 17083 8415
rect 20361 8381 20395 8415
rect 8852 8313 8886 8347
rect 10609 8313 10643 8347
rect 11069 8313 11103 8347
rect 13636 8313 13670 8347
rect 17141 8313 17175 8347
rect 20453 8313 20487 8347
rect 9965 8245 9999 8279
rect 11161 8245 11195 8279
rect 12449 8245 12483 8279
rect 18981 8245 19015 8279
rect 19349 8245 19383 8279
rect 19441 8245 19475 8279
rect 19993 8245 20027 8279
rect 14013 8041 14047 8075
rect 14657 8041 14691 8075
rect 15485 8041 15519 8075
rect 19165 8041 19199 8075
rect 12878 7973 12912 8007
rect 16580 7973 16614 8007
rect 20269 7973 20303 8007
rect 7941 7905 7975 7939
rect 8208 7905 8242 7939
rect 10701 7905 10735 7939
rect 11244 7905 11278 7939
rect 15669 7905 15703 7939
rect 16313 7905 16347 7939
rect 18429 7905 18463 7939
rect 20177 7905 20211 7939
rect 10977 7837 11011 7871
rect 12633 7837 12667 7871
rect 18705 7837 18739 7871
rect 20361 7837 20395 7871
rect 9321 7701 9355 7735
rect 10517 7701 10551 7735
rect 12357 7701 12391 7735
rect 17693 7701 17727 7735
rect 19809 7701 19843 7735
rect 8677 7497 8711 7531
rect 8953 7497 8987 7531
rect 9965 7497 9999 7531
rect 13461 7497 13495 7531
rect 14473 7497 14507 7531
rect 11069 7429 11103 7463
rect 19625 7429 19659 7463
rect 7297 7361 7331 7395
rect 9505 7361 9539 7395
rect 10517 7361 10551 7395
rect 11621 7361 11655 7395
rect 14013 7361 14047 7395
rect 15025 7361 15059 7395
rect 17141 7361 17175 7395
rect 20361 7361 20395 7395
rect 20453 7361 20487 7395
rect 9321 7293 9355 7327
rect 13921 7293 13955 7327
rect 18245 7293 18279 7327
rect 18512 7293 18546 7327
rect 7564 7225 7598 7259
rect 11437 7225 11471 7259
rect 14933 7225 14967 7259
rect 9413 7157 9447 7191
rect 10333 7157 10367 7191
rect 10425 7157 10459 7191
rect 11529 7157 11563 7191
rect 13277 7157 13311 7191
rect 13829 7157 13863 7191
rect 14841 7157 14875 7191
rect 16497 7157 16531 7191
rect 16865 7157 16899 7191
rect 16957 7157 16991 7191
rect 19901 7157 19935 7191
rect 20269 7157 20303 7191
rect 11437 6953 11471 6987
rect 12449 6953 12483 6987
rect 17877 6953 17911 6987
rect 12541 6885 12575 6919
rect 8217 6817 8251 6851
rect 10324 6817 10358 6851
rect 11989 6817 12023 6851
rect 12909 6817 12943 6851
rect 13176 6817 13210 6851
rect 16017 6817 16051 6851
rect 17785 6817 17819 6851
rect 18613 6817 18647 6851
rect 18880 6817 18914 6851
rect 10057 6749 10091 6783
rect 12633 6749 12667 6783
rect 14565 6749 14599 6783
rect 15761 6749 15795 6783
rect 17969 6749 18003 6783
rect 20269 6749 20303 6783
rect 11805 6681 11839 6715
rect 12081 6681 12115 6715
rect 17141 6681 17175 6715
rect 17417 6681 17451 6715
rect 14289 6613 14323 6647
rect 19993 6613 20027 6647
rect 8401 6409 8435 6443
rect 9873 6409 9907 6443
rect 14013 6409 14047 6443
rect 16957 6409 16991 6443
rect 19073 6409 19107 6443
rect 19257 6409 19291 6443
rect 20269 6409 20303 6443
rect 13001 6341 13035 6375
rect 7021 6273 7055 6307
rect 10517 6273 10551 6307
rect 13645 6273 13679 6307
rect 14565 6273 14599 6307
rect 15025 6273 15059 6307
rect 17509 6273 17543 6307
rect 18889 6273 18923 6307
rect 13369 6205 13403 6239
rect 15292 6205 15326 6239
rect 17325 6205 17359 6239
rect 19717 6273 19751 6307
rect 19809 6273 19843 6307
rect 20821 6273 20855 6307
rect 20729 6205 20763 6239
rect 7288 6137 7322 6171
rect 10241 6137 10275 6171
rect 10885 6137 10919 6171
rect 18613 6137 18647 6171
rect 19073 6137 19107 6171
rect 20637 6137 20671 6171
rect 10333 6069 10367 6103
rect 13461 6069 13495 6103
rect 14381 6069 14415 6103
rect 14473 6069 14507 6103
rect 16405 6069 16439 6103
rect 17417 6069 17451 6103
rect 18245 6069 18279 6103
rect 18705 6069 18739 6103
rect 19625 6069 19659 6103
rect 7757 5865 7791 5899
rect 8033 5865 8067 5899
rect 8401 5865 8435 5899
rect 9045 5865 9079 5899
rect 11069 5865 11103 5899
rect 15853 5865 15887 5899
rect 16957 5865 16991 5899
rect 17325 5865 17359 5899
rect 18981 5865 19015 5899
rect 11612 5797 11646 5831
rect 19441 5797 19475 5831
rect 6377 5729 6411 5763
rect 6644 5729 6678 5763
rect 9956 5729 9990 5763
rect 11345 5729 11379 5763
rect 15393 5729 15427 5763
rect 16221 5729 16255 5763
rect 19349 5729 19383 5763
rect 20269 5729 20303 5763
rect 8493 5661 8527 5695
rect 8585 5661 8619 5695
rect 9689 5661 9723 5695
rect 16313 5661 16347 5695
rect 16497 5661 16531 5695
rect 17417 5661 17451 5695
rect 17509 5661 17543 5695
rect 19533 5661 19567 5695
rect 12725 5525 12759 5559
rect 20453 5525 20487 5559
rect 8217 5321 8251 5355
rect 8493 5321 8527 5355
rect 9597 5321 9631 5355
rect 13277 5321 13311 5355
rect 15853 5321 15887 5355
rect 18613 5321 18647 5355
rect 6837 5185 6871 5219
rect 9045 5185 9079 5219
rect 10241 5185 10275 5219
rect 10701 5185 10735 5219
rect 13829 5185 13863 5219
rect 14841 5185 14875 5219
rect 16497 5185 16531 5219
rect 18981 5185 19015 5219
rect 9965 5117 9999 5151
rect 10057 5117 10091 5151
rect 14749 5117 14783 5151
rect 18429 5117 18463 5151
rect 19248 5117 19282 5151
rect 20637 5117 20671 5151
rect 7104 5049 7138 5083
rect 10968 5049 11002 5083
rect 14657 5049 14691 5083
rect 16313 5049 16347 5083
rect 8861 4981 8895 5015
rect 8953 4981 8987 5015
rect 12081 4981 12115 5015
rect 12449 4981 12483 5015
rect 13645 4981 13679 5015
rect 13737 4981 13771 5015
rect 14289 4981 14323 5015
rect 16221 4981 16255 5015
rect 20361 4981 20395 5015
rect 20821 4981 20855 5015
rect 7021 4777 7055 4811
rect 8585 4777 8619 4811
rect 11069 4777 11103 4811
rect 11621 4777 11655 4811
rect 11989 4777 12023 4811
rect 15301 4777 15335 4811
rect 17877 4777 17911 4811
rect 18245 4777 18279 4811
rect 8953 4709 8987 4743
rect 15761 4709 15795 4743
rect 7389 4641 7423 4675
rect 9945 4641 9979 4675
rect 12081 4641 12115 4675
rect 13093 4641 13127 4675
rect 13360 4641 13394 4675
rect 14749 4641 14783 4675
rect 15669 4641 15703 4675
rect 16764 4641 16798 4675
rect 18613 4641 18647 4675
rect 18705 4641 18739 4675
rect 19901 4641 19935 4675
rect 7481 4573 7515 4607
rect 7665 4573 7699 4607
rect 9045 4573 9079 4607
rect 9229 4573 9263 4607
rect 9689 4573 9723 4607
rect 12173 4573 12207 4607
rect 15853 4573 15887 4607
rect 16497 4573 16531 4607
rect 18797 4573 18831 4607
rect 19993 4573 20027 4607
rect 20177 4573 20211 4607
rect 14473 4437 14507 4471
rect 19533 4437 19567 4471
rect 9873 4233 9907 4267
rect 14657 4233 14691 4267
rect 19717 4233 19751 4267
rect 10977 4165 11011 4199
rect 20913 4165 20947 4199
rect 8033 4097 8067 4131
rect 8493 4097 8527 4131
rect 11529 4097 11563 4131
rect 13277 4097 13311 4131
rect 18061 4097 18095 4131
rect 20177 4097 20211 4131
rect 20361 4097 20395 4131
rect 12449 4029 12483 4063
rect 15485 4029 15519 4063
rect 15752 4029 15786 4063
rect 17417 4029 17451 4063
rect 20729 4029 20763 4063
rect 7849 3961 7883 3995
rect 8760 3961 8794 3995
rect 11437 3961 11471 3995
rect 13544 3961 13578 3995
rect 18328 3961 18362 3995
rect 7389 3893 7423 3927
rect 7757 3893 7791 3927
rect 11345 3893 11379 3927
rect 12633 3893 12667 3927
rect 16865 3893 16899 3927
rect 17601 3893 17635 3927
rect 19441 3893 19475 3927
rect 20085 3893 20119 3927
rect 9321 3689 9355 3723
rect 9689 3689 9723 3723
rect 11989 3689 12023 3723
rect 13185 3689 13219 3723
rect 13645 3689 13679 3723
rect 14197 3689 14231 3723
rect 14657 3689 14691 3723
rect 15301 3689 15335 3723
rect 15669 3689 15703 3723
rect 17601 3689 17635 3723
rect 17693 3689 17727 3723
rect 20545 3689 20579 3723
rect 8208 3621 8242 3655
rect 10600 3621 10634 3655
rect 6285 3553 6319 3587
rect 6552 3553 6586 3587
rect 12357 3553 12391 3587
rect 12449 3553 12483 3587
rect 13553 3553 13587 3587
rect 14565 3553 14599 3587
rect 15761 3553 15795 3587
rect 7941 3485 7975 3519
rect 10333 3485 10367 3519
rect 12633 3485 12667 3519
rect 13829 3485 13863 3519
rect 14841 3485 14875 3519
rect 15945 3485 15979 3519
rect 18061 3553 18095 3587
rect 18705 3553 18739 3587
rect 19432 3553 19466 3587
rect 18153 3485 18187 3519
rect 18337 3485 18371 3519
rect 19165 3485 19199 3519
rect 17601 3417 17635 3451
rect 7665 3349 7699 3383
rect 11713 3349 11747 3383
rect 8217 3145 8251 3179
rect 8677 3145 8711 3179
rect 14105 3145 14139 3179
rect 16957 3145 16991 3179
rect 17141 3145 17175 3179
rect 19533 3145 19567 3179
rect 11805 3077 11839 3111
rect 16497 3077 16531 3111
rect 6837 3009 6871 3043
rect 9137 3009 9171 3043
rect 9321 3009 9355 3043
rect 10425 3009 10459 3043
rect 15025 3009 15059 3043
rect 7104 2941 7138 2975
rect 10692 2941 10726 2975
rect 12725 2941 12759 2975
rect 12992 2873 13026 2907
rect 15117 2941 15151 2975
rect 15384 2941 15418 2975
rect 16773 2941 16807 2975
rect 9045 2805 9079 2839
rect 14381 2805 14415 2839
rect 15025 2805 15059 2839
rect 18797 3077 18831 3111
rect 20177 3009 20211 3043
rect 17325 2941 17359 2975
rect 18061 2941 18095 2975
rect 18613 2941 18647 2975
rect 19901 2941 19935 2975
rect 20545 2941 20579 2975
rect 17141 2805 17175 2839
rect 17509 2805 17543 2839
rect 18245 2805 18279 2839
rect 19993 2805 20027 2839
rect 20729 2805 20763 2839
rect 7297 2601 7331 2635
rect 7757 2601 7791 2635
rect 8309 2601 8343 2635
rect 11069 2601 11103 2635
rect 11529 2601 11563 2635
rect 12081 2601 12115 2635
rect 13001 2601 13035 2635
rect 13369 2601 13403 2635
rect 15485 2601 15519 2635
rect 15853 2601 15887 2635
rect 20729 2601 20763 2635
rect 13461 2533 13495 2567
rect 7665 2465 7699 2499
rect 11437 2465 11471 2499
rect 15945 2465 15979 2499
rect 17417 2465 17451 2499
rect 18705 2465 18739 2499
rect 19441 2465 19475 2499
rect 19993 2465 20027 2499
rect 20545 2465 20579 2499
rect 7849 2397 7883 2431
rect 11713 2397 11747 2431
rect 13645 2397 13679 2431
rect 16037 2397 16071 2431
rect 20177 2329 20211 2363
rect 17601 2261 17635 2295
rect 18889 2261 18923 2295
rect 19625 2261 19659 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 20714 20040 20720 20052
rect 20675 20012 20720 20040
rect 20714 20000 20720 20012
rect 20772 20000 20778 20052
rect 20530 19904 20536 19916
rect 20491 19876 20536 19904
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 20162 19496 20168 19508
rect 20123 19468 20168 19496
rect 20162 19456 20168 19468
rect 20220 19456 20226 19508
rect 20714 19496 20720 19508
rect 20675 19468 20720 19496
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 11698 19252 11704 19304
rect 11756 19292 11762 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 11756 19264 12449 19292
rect 11756 19252 11762 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 19978 19292 19984 19304
rect 19939 19264 19984 19292
rect 12437 19255 12495 19261
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20533 19295 20591 19301
rect 20533 19261 20545 19295
rect 20579 19261 20591 19295
rect 20533 19255 20591 19261
rect 15194 19184 15200 19236
rect 15252 19224 15258 19236
rect 20548 19224 20576 19255
rect 15252 19196 20576 19224
rect 15252 19184 15258 19196
rect 12621 19159 12679 19165
rect 12621 19125 12633 19159
rect 12667 19156 12679 19159
rect 17954 19156 17960 19168
rect 12667 19128 17960 19156
rect 12667 19125 12679 19128
rect 12621 19119 12679 19125
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 19978 18952 19984 18964
rect 10152 18924 19984 18952
rect 10152 18893 10180 18924
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 20438 18952 20444 18964
rect 20399 18924 20444 18952
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 10137 18887 10195 18893
rect 10137 18853 10149 18887
rect 10183 18853 10195 18887
rect 11698 18884 11704 18896
rect 11659 18856 11704 18884
rect 10137 18847 10195 18853
rect 11698 18844 11704 18856
rect 11756 18844 11762 18896
rect 17126 18844 17132 18896
rect 17184 18884 17190 18896
rect 17374 18887 17432 18893
rect 17374 18884 17386 18887
rect 17184 18856 17386 18884
rect 17184 18844 17190 18856
rect 17374 18853 17386 18856
rect 17420 18853 17432 18887
rect 17374 18847 17432 18853
rect 7745 18819 7803 18825
rect 7745 18785 7757 18819
rect 7791 18816 7803 18819
rect 8202 18816 8208 18828
rect 7791 18788 8208 18816
rect 7791 18785 7803 18788
rect 7745 18779 7803 18785
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 8665 18819 8723 18825
rect 8665 18785 8677 18819
rect 8711 18816 8723 18819
rect 8846 18816 8852 18828
rect 8711 18788 8852 18816
rect 8711 18785 8723 18788
rect 8665 18779 8723 18785
rect 8846 18776 8852 18788
rect 8904 18776 8910 18828
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 9861 18819 9919 18825
rect 9861 18816 9873 18819
rect 9732 18788 9873 18816
rect 9732 18776 9738 18788
rect 9861 18785 9873 18788
rect 9907 18785 9919 18819
rect 9861 18779 9919 18785
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 11020 18788 11437 18816
rect 11020 18776 11026 18788
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 11532 18788 12664 18816
rect 8018 18748 8024 18760
rect 7979 18720 8024 18748
rect 8018 18708 8024 18720
rect 8076 18708 8082 18760
rect 8941 18751 8999 18757
rect 8941 18717 8953 18751
rect 8987 18748 8999 18751
rect 11532 18748 11560 18788
rect 8987 18720 11560 18748
rect 8987 18717 8999 18720
rect 8941 18711 8999 18717
rect 5718 18572 5724 18624
rect 5776 18612 5782 18624
rect 12526 18612 12532 18624
rect 5776 18584 12532 18612
rect 5776 18572 5782 18584
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 12636 18612 12664 18788
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 20257 18819 20315 18825
rect 20257 18816 20269 18819
rect 12768 18788 20269 18816
rect 12768 18776 12774 18788
rect 20257 18785 20269 18788
rect 20303 18785 20315 18819
rect 20257 18779 20315 18785
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 17129 18751 17187 18757
rect 17129 18748 17141 18751
rect 17000 18720 17141 18748
rect 17000 18708 17006 18720
rect 17129 18717 17141 18720
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 20530 18680 20536 18692
rect 18064 18652 20536 18680
rect 18064 18612 18092 18652
rect 20530 18640 20536 18652
rect 20588 18640 20594 18692
rect 18506 18612 18512 18624
rect 12636 18584 18092 18612
rect 18467 18584 18512 18612
rect 18506 18572 18512 18584
rect 18564 18572 18570 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 8018 18368 8024 18420
rect 8076 18408 8082 18420
rect 15194 18408 15200 18420
rect 8076 18380 15200 18408
rect 8076 18368 8082 18380
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 15289 18411 15347 18417
rect 15289 18377 15301 18411
rect 15335 18408 15347 18411
rect 17954 18408 17960 18420
rect 15335 18380 17960 18408
rect 15335 18377 15347 18380
rect 15289 18371 15347 18377
rect 17954 18368 17960 18380
rect 18012 18368 18018 18420
rect 20714 18340 20720 18352
rect 20675 18312 20720 18340
rect 20714 18300 20720 18312
rect 20772 18300 20778 18352
rect 12710 18272 12716 18284
rect 12671 18244 12716 18272
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 12434 18204 12440 18216
rect 12395 18176 12440 18204
rect 12434 18164 12440 18176
rect 12492 18164 12498 18216
rect 15102 18204 15108 18216
rect 15063 18176 15108 18204
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20533 18207 20591 18213
rect 20533 18204 20545 18207
rect 20128 18176 20545 18204
rect 20128 18164 20134 18176
rect 20533 18173 20545 18176
rect 20579 18173 20591 18207
rect 20533 18167 20591 18173
rect 12526 18096 12532 18148
rect 12584 18136 12590 18148
rect 12710 18136 12716 18148
rect 12584 18108 12716 18136
rect 12584 18096 12590 18108
rect 12710 18096 12716 18108
rect 12768 18096 12774 18148
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 20438 17864 20444 17876
rect 20399 17836 20444 17864
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 14553 17799 14611 17805
rect 14553 17765 14565 17799
rect 14599 17796 14611 17799
rect 15102 17796 15108 17808
rect 14599 17768 15108 17796
rect 14599 17765 14611 17768
rect 14553 17759 14611 17765
rect 15102 17756 15108 17768
rect 15160 17756 15166 17808
rect 14274 17728 14280 17740
rect 14235 17700 14280 17728
rect 14274 17688 14280 17700
rect 14332 17688 14338 17740
rect 19978 17688 19984 17740
rect 20036 17728 20042 17740
rect 20257 17731 20315 17737
rect 20257 17728 20269 17731
rect 20036 17700 20269 17728
rect 20036 17688 20042 17700
rect 20257 17697 20269 17700
rect 20303 17697 20315 17731
rect 20257 17691 20315 17697
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 20714 17320 20720 17332
rect 20675 17292 20720 17320
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17184 20039 17187
rect 20070 17184 20076 17196
rect 20027 17156 20076 17184
rect 20027 17153 20039 17156
rect 19981 17147 20039 17153
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 19518 17076 19524 17128
rect 19576 17116 19582 17128
rect 19705 17119 19763 17125
rect 19705 17116 19717 17119
rect 19576 17088 19717 17116
rect 19576 17076 19582 17088
rect 19705 17085 19717 17088
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 20533 17119 20591 17125
rect 20533 17085 20545 17119
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 16758 17008 16764 17060
rect 16816 17048 16822 17060
rect 20548 17048 20576 17079
rect 16816 17020 20576 17048
rect 16816 17008 16822 17020
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 19978 16708 19984 16720
rect 19939 16680 19984 16708
rect 19978 16668 19984 16680
rect 20036 16668 20042 16720
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19705 16643 19763 16649
rect 19705 16640 19717 16643
rect 19484 16612 19717 16640
rect 19484 16600 19490 16612
rect 19705 16609 19717 16612
rect 19751 16609 19763 16643
rect 19705 16603 19763 16609
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 20162 16232 20168 16244
rect 20123 16204 20168 16232
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 12713 16099 12771 16105
rect 12713 16065 12725 16099
rect 12759 16096 12771 16099
rect 16758 16096 16764 16108
rect 12759 16068 16764 16096
rect 12759 16065 12771 16068
rect 12713 16059 12771 16065
rect 16758 16056 16764 16068
rect 16816 16056 16822 16108
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 16028 12495 16031
rect 12526 16028 12532 16040
rect 12483 16000 12532 16028
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 19978 16028 19984 16040
rect 19939 16000 19984 16028
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 20070 15988 20076 16040
rect 20128 16028 20134 16040
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20128 16000 20545 16028
rect 20128 15988 20134 16000
rect 20533 15997 20545 16000
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 10042 15512 10048 15564
rect 10100 15552 10106 15564
rect 10505 15555 10563 15561
rect 10505 15552 10517 15555
rect 10100 15524 10517 15552
rect 10100 15512 10106 15524
rect 10505 15521 10517 15524
rect 10551 15521 10563 15555
rect 10505 15515 10563 15521
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 19392 15524 20269 15552
rect 19392 15512 19398 15524
rect 20257 15521 20269 15524
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 10781 15487 10839 15493
rect 10781 15453 10793 15487
rect 10827 15484 10839 15487
rect 19978 15484 19984 15496
rect 10827 15456 19984 15484
rect 10827 15453 10839 15456
rect 10781 15447 10839 15453
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 20162 15144 20168 15156
rect 20123 15116 20168 15144
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 20714 15076 20720 15088
rect 20675 15048 20720 15076
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 9766 14900 9772 14952
rect 9824 14940 9830 14952
rect 9861 14943 9919 14949
rect 9861 14940 9873 14943
rect 9824 14912 9873 14940
rect 9824 14900 9830 14912
rect 9861 14909 9873 14912
rect 9907 14909 9919 14943
rect 9861 14903 9919 14909
rect 16206 14900 16212 14952
rect 16264 14940 16270 14952
rect 19981 14943 20039 14949
rect 19981 14940 19993 14943
rect 16264 14912 19993 14940
rect 16264 14900 16270 14912
rect 19981 14909 19993 14912
rect 20027 14909 20039 14943
rect 19981 14903 20039 14909
rect 20346 14900 20352 14952
rect 20404 14940 20410 14952
rect 20533 14943 20591 14949
rect 20533 14940 20545 14943
rect 20404 14912 20545 14940
rect 20404 14900 20410 14912
rect 20533 14909 20545 14912
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 10137 14875 10195 14881
rect 10137 14841 10149 14875
rect 10183 14872 10195 14875
rect 20070 14872 20076 14884
rect 10183 14844 20076 14872
rect 10183 14841 10195 14844
rect 10137 14835 10195 14841
rect 20070 14832 20076 14844
rect 20128 14832 20134 14884
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 20438 14600 20444 14612
rect 20399 14572 20444 14600
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 8205 14535 8263 14541
rect 8205 14501 8217 14535
rect 8251 14532 8263 14535
rect 19334 14532 19340 14544
rect 8251 14504 19340 14532
rect 8251 14501 8263 14504
rect 8205 14495 8263 14501
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 7374 14424 7380 14476
rect 7432 14464 7438 14476
rect 7929 14467 7987 14473
rect 7929 14464 7941 14467
rect 7432 14436 7941 14464
rect 7432 14424 7438 14436
rect 7929 14433 7941 14436
rect 7975 14433 7987 14467
rect 7929 14427 7987 14433
rect 10870 14424 10876 14476
rect 10928 14464 10934 14476
rect 11609 14467 11667 14473
rect 11609 14464 11621 14467
rect 10928 14436 11621 14464
rect 10928 14424 10934 14436
rect 11609 14433 11621 14436
rect 11655 14433 11667 14467
rect 11609 14427 11667 14433
rect 19978 14424 19984 14476
rect 20036 14464 20042 14476
rect 20257 14467 20315 14473
rect 20257 14464 20269 14467
rect 20036 14436 20269 14464
rect 20036 14424 20042 14436
rect 20257 14433 20269 14436
rect 20303 14433 20315 14467
rect 20257 14427 20315 14433
rect 11793 14399 11851 14405
rect 11793 14365 11805 14399
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11808 14328 11836 14359
rect 16206 14328 16212 14340
rect 11808 14300 16212 14328
rect 16206 14288 16212 14300
rect 16264 14288 16270 14340
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 20622 13948 20628 14000
rect 20680 13988 20686 14000
rect 20717 13991 20775 13997
rect 20717 13988 20729 13991
rect 20680 13960 20729 13988
rect 20680 13948 20686 13960
rect 20717 13957 20729 13960
rect 20763 13957 20775 13991
rect 20717 13951 20775 13957
rect 19981 13923 20039 13929
rect 19981 13889 19993 13923
rect 20027 13920 20039 13923
rect 20346 13920 20352 13932
rect 20027 13892 20352 13920
rect 20027 13889 20039 13892
rect 19981 13883 20039 13889
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 13412 13824 19717 13852
rect 13412 13812 13418 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 19794 13812 19800 13864
rect 19852 13852 19858 13864
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 19852 13824 20545 13852
rect 19852 13812 19858 13824
rect 20533 13821 20545 13824
rect 20579 13821 20591 13855
rect 20533 13815 20591 13821
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 19334 13512 19340 13524
rect 19295 13484 19340 13512
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 19978 13444 19984 13456
rect 19939 13416 19984 13444
rect 19978 13404 19984 13416
rect 20036 13404 20042 13456
rect 19150 13376 19156 13388
rect 19111 13348 19156 13376
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 13262 13268 13268 13320
rect 13320 13308 13326 13320
rect 19720 13308 19748 13339
rect 13320 13280 19748 13308
rect 13320 13268 13326 13280
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 20714 12968 20720 12980
rect 20675 12940 20720 12968
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 16482 12792 16488 12844
rect 16540 12832 16546 12844
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16540 12804 16681 12832
rect 16540 12792 16546 12804
rect 16669 12801 16681 12804
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 19150 12792 19156 12844
rect 19208 12832 19214 12844
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 19208 12804 19809 12832
rect 19208 12792 19214 12804
rect 19797 12801 19809 12804
rect 19843 12801 19855 12835
rect 19797 12795 19855 12801
rect 17402 12724 17408 12776
rect 17460 12764 17466 12776
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 17460 12736 19625 12764
rect 17460 12724 17466 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 20530 12764 20536 12776
rect 20491 12736 20536 12764
rect 19613 12727 19671 12733
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 16114 12628 16120 12640
rect 16075 12600 16120 12628
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 16390 12588 16396 12640
rect 16448 12628 16454 12640
rect 16485 12631 16543 12637
rect 16485 12628 16497 12631
rect 16448 12600 16497 12628
rect 16448 12588 16454 12600
rect 16485 12597 16497 12600
rect 16531 12597 16543 12631
rect 16485 12591 16543 12597
rect 16577 12631 16635 12637
rect 16577 12597 16589 12631
rect 16623 12628 16635 12631
rect 17862 12628 17868 12640
rect 16623 12600 17868 12628
rect 16623 12597 16635 12600
rect 16577 12591 16635 12597
rect 17862 12588 17868 12600
rect 17920 12588 17926 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 16025 12427 16083 12433
rect 16025 12393 16037 12427
rect 16071 12424 16083 12427
rect 16114 12424 16120 12436
rect 16071 12396 16120 12424
rect 16071 12393 16083 12396
rect 16025 12387 16083 12393
rect 16114 12384 16120 12396
rect 16172 12384 16178 12436
rect 19429 12359 19487 12365
rect 19429 12325 19441 12359
rect 19475 12356 19487 12359
rect 19794 12356 19800 12368
rect 19475 12328 19800 12356
rect 19475 12325 19487 12328
rect 19429 12319 19487 12325
rect 19794 12316 19800 12328
rect 19852 12316 19858 12368
rect 20165 12359 20223 12365
rect 20165 12325 20177 12359
rect 20211 12356 20223 12359
rect 20530 12356 20536 12368
rect 20211 12328 20536 12356
rect 20211 12325 20223 12328
rect 20165 12319 20223 12325
rect 20530 12316 20536 12328
rect 20588 12316 20594 12368
rect 15010 12248 15016 12300
rect 15068 12288 15074 12300
rect 16850 12297 16856 12300
rect 15933 12291 15991 12297
rect 15933 12288 15945 12291
rect 15068 12260 15945 12288
rect 15068 12248 15074 12260
rect 15933 12257 15945 12260
rect 15979 12257 15991 12291
rect 16844 12288 16856 12297
rect 15933 12251 15991 12257
rect 16224 12260 16856 12288
rect 16224 12229 16252 12260
rect 16844 12251 16856 12260
rect 16850 12248 16856 12251
rect 16908 12248 16914 12300
rect 18598 12288 18604 12300
rect 18559 12260 18604 12288
rect 18598 12248 18604 12260
rect 18656 12248 18662 12300
rect 18874 12248 18880 12300
rect 18932 12288 18938 12300
rect 19153 12291 19211 12297
rect 19153 12288 19165 12291
rect 18932 12260 19165 12288
rect 18932 12248 18938 12260
rect 19153 12257 19165 12260
rect 19199 12257 19211 12291
rect 19153 12251 19211 12257
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 19889 12291 19947 12297
rect 19889 12288 19901 12291
rect 19300 12260 19901 12288
rect 19300 12248 19306 12260
rect 19889 12257 19901 12260
rect 19935 12257 19947 12291
rect 19889 12251 19947 12257
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 16577 12223 16635 12229
rect 16577 12189 16589 12223
rect 16623 12189 16635 12223
rect 16577 12183 16635 12189
rect 11974 12044 11980 12096
rect 12032 12084 12038 12096
rect 15565 12087 15623 12093
rect 15565 12084 15577 12087
rect 12032 12056 15577 12084
rect 12032 12044 12038 12056
rect 15565 12053 15577 12056
rect 15611 12053 15623 12087
rect 16592 12084 16620 12183
rect 16942 12084 16948 12096
rect 16592 12056 16948 12084
rect 15565 12047 15623 12053
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 17954 12084 17960 12096
rect 17915 12056 17960 12084
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 22462 12084 22468 12096
rect 18831 12056 22468 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 22462 12044 22468 12056
rect 22520 12044 22526 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 16850 11880 16856 11892
rect 16811 11852 16856 11880
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 20717 11883 20775 11889
rect 20717 11849 20729 11883
rect 20763 11880 20775 11883
rect 21082 11880 21088 11892
rect 20763 11852 21088 11880
rect 20763 11849 20775 11852
rect 20717 11843 20775 11849
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 13630 11744 13636 11756
rect 13591 11716 13636 11744
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 15010 11744 15016 11756
rect 14971 11716 15016 11744
rect 15010 11704 15016 11716
rect 15068 11704 15074 11756
rect 16942 11704 16948 11756
rect 17000 11744 17006 11756
rect 17862 11744 17868 11756
rect 17000 11716 17868 11744
rect 17000 11704 17006 11716
rect 17862 11704 17868 11716
rect 17920 11744 17926 11756
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 17920 11716 18061 11744
rect 17920 11704 17926 11716
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 15473 11679 15531 11685
rect 15473 11645 15485 11679
rect 15519 11645 15531 11679
rect 15473 11639 15531 11645
rect 15740 11679 15798 11685
rect 15740 11645 15752 11679
rect 15786 11676 15798 11679
rect 16482 11676 16488 11688
rect 15786 11648 16488 11676
rect 15786 11645 15798 11648
rect 15740 11639 15798 11645
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 15488 11608 15516 11639
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 16960 11608 16988 11704
rect 18782 11636 18788 11688
rect 18840 11676 18846 11688
rect 19797 11679 19855 11685
rect 19797 11676 19809 11679
rect 18840 11648 19809 11676
rect 18840 11636 18846 11648
rect 19797 11645 19809 11648
rect 19843 11645 19855 11679
rect 19797 11639 19855 11645
rect 20162 11636 20168 11688
rect 20220 11676 20226 11688
rect 20533 11679 20591 11685
rect 20533 11676 20545 11679
rect 20220 11648 20545 11676
rect 20220 11636 20226 11648
rect 20533 11645 20545 11648
rect 20579 11645 20591 11679
rect 20533 11639 20591 11645
rect 15344 11580 16988 11608
rect 15344 11568 15350 11580
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 18294 11611 18352 11617
rect 18294 11608 18306 11611
rect 18012 11580 18306 11608
rect 18012 11568 18018 11580
rect 18294 11577 18306 11580
rect 18340 11577 18352 11611
rect 18294 11571 18352 11577
rect 20073 11611 20131 11617
rect 20073 11577 20085 11611
rect 20119 11608 20131 11611
rect 20714 11608 20720 11620
rect 20119 11580 20720 11608
rect 20119 11577 20131 11580
rect 20073 11571 20131 11577
rect 20714 11568 20720 11580
rect 20772 11568 20778 11620
rect 13078 11540 13084 11552
rect 13039 11512 13084 11540
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 13228 11512 13461 11540
rect 13228 11500 13234 11512
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 13449 11503 13507 11509
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 13596 11512 13641 11540
rect 13596 11500 13602 11512
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18506 11540 18512 11552
rect 18104 11512 18512 11540
rect 18104 11500 18110 11512
rect 18506 11500 18512 11512
rect 18564 11540 18570 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 18564 11512 19441 11540
rect 18564 11500 18570 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19429 11503 19487 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 16298 11336 16304 11348
rect 13044 11308 16304 11336
rect 13044 11296 13050 11308
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 16540 11308 16681 11336
rect 16540 11296 16546 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 17681 11339 17739 11345
rect 17681 11305 17693 11339
rect 17727 11336 17739 11339
rect 18233 11339 18291 11345
rect 18233 11336 18245 11339
rect 17727 11308 18245 11336
rect 17727 11305 17739 11308
rect 17681 11299 17739 11305
rect 18233 11305 18245 11308
rect 18279 11305 18291 11339
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18233 11299 18291 11305
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 12710 11268 12716 11280
rect 12671 11240 12716 11268
rect 12710 11228 12716 11240
rect 12768 11228 12774 11280
rect 13078 11228 13084 11280
rect 13136 11268 13142 11280
rect 20162 11268 20168 11280
rect 13136 11240 19932 11268
rect 20123 11240 20168 11268
rect 13136 11228 13142 11240
rect 11974 11200 11980 11212
rect 11935 11172 11980 11200
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 15010 11160 15016 11212
rect 15068 11200 15074 11212
rect 15105 11203 15163 11209
rect 15105 11200 15117 11203
rect 15068 11172 15117 11200
rect 15068 11160 15074 11172
rect 15105 11169 15117 11172
rect 15151 11169 15163 11203
rect 15286 11200 15292 11212
rect 15247 11172 15292 11200
rect 15105 11163 15163 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15556 11203 15614 11209
rect 15556 11169 15568 11203
rect 15602 11200 15614 11203
rect 16390 11200 16396 11212
rect 15602 11172 16396 11200
rect 15602 11169 15614 11172
rect 15556 11163 15614 11169
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 17586 11200 17592 11212
rect 17547 11172 17592 11200
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 18046 11200 18052 11212
rect 17880 11172 18052 11200
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11132 12311 11135
rect 12802 11132 12808 11144
rect 12299 11104 12808 11132
rect 12299 11101 12311 11104
rect 12253 11095 12311 11101
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 14366 11132 14372 11144
rect 14327 11104 14372 11132
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 14918 11064 14924 11076
rect 14831 11036 14924 11064
rect 14918 11024 14924 11036
rect 14976 11064 14982 11076
rect 15304 11064 15332 11160
rect 17880 11141 17908 11172
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 18598 11200 18604 11212
rect 18559 11172 18604 11200
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 19242 11160 19248 11212
rect 19300 11200 19306 11212
rect 19904 11209 19932 11240
rect 20162 11228 20168 11240
rect 20220 11228 20226 11280
rect 19337 11203 19395 11209
rect 19337 11200 19349 11203
rect 19300 11172 19349 11200
rect 19300 11160 19306 11172
rect 19337 11169 19349 11172
rect 19383 11169 19395 11203
rect 19337 11163 19395 11169
rect 19889 11203 19947 11209
rect 19889 11169 19901 11203
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 17865 11135 17923 11141
rect 17865 11101 17877 11135
rect 17911 11101 17923 11135
rect 17865 11095 17923 11101
rect 17954 11092 17960 11144
rect 18012 11132 18018 11144
rect 18785 11135 18843 11141
rect 18785 11132 18797 11135
rect 18012 11104 18797 11132
rect 18012 11092 18018 11104
rect 18785 11101 18797 11104
rect 18831 11101 18843 11135
rect 18785 11095 18843 11101
rect 14976 11036 15332 11064
rect 14976 11024 14982 11036
rect 16298 11024 16304 11076
rect 16356 11064 16362 11076
rect 19521 11067 19579 11073
rect 19521 11064 19533 11067
rect 16356 11036 19533 11064
rect 16356 11024 16362 11036
rect 19521 11033 19533 11036
rect 19567 11033 19579 11067
rect 19521 11027 19579 11033
rect 16850 10956 16856 11008
rect 16908 10996 16914 11008
rect 17221 10999 17279 11005
rect 17221 10996 17233 10999
rect 16908 10968 17233 10996
rect 16908 10956 16914 10968
rect 17221 10965 17233 10968
rect 17267 10965 17279 10999
rect 17221 10959 17279 10965
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 10962 10792 10968 10804
rect 10923 10764 10968 10792
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 16390 10792 16396 10804
rect 16351 10764 16396 10792
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 16669 10795 16727 10801
rect 16669 10761 16681 10795
rect 16715 10792 16727 10795
rect 18782 10792 18788 10804
rect 16715 10764 18788 10792
rect 16715 10761 16727 10764
rect 16669 10755 16727 10761
rect 18782 10752 18788 10764
rect 18840 10752 18846 10804
rect 19426 10792 19432 10804
rect 19339 10764 19432 10792
rect 19426 10752 19432 10764
rect 19484 10792 19490 10804
rect 20898 10792 20904 10804
rect 19484 10764 20300 10792
rect 20859 10764 20904 10792
rect 19484 10752 19490 10764
rect 11606 10656 11612 10668
rect 11567 10628 11612 10656
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 13170 10656 13176 10668
rect 12943 10628 13176 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 14918 10616 14924 10668
rect 14976 10656 14982 10668
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14976 10628 15025 10656
rect 14976 10616 14982 10628
rect 15013 10625 15025 10628
rect 15059 10656 15071 10659
rect 16408 10656 16436 10752
rect 17221 10659 17279 10665
rect 17221 10656 17233 10659
rect 15059 10628 15148 10656
rect 16408 10628 17233 10656
rect 15059 10625 15071 10628
rect 15013 10619 15071 10625
rect 15120 10600 15148 10628
rect 17221 10625 17233 10628
rect 17267 10625 17279 10659
rect 17221 10619 17279 10625
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 20272 10665 20300 10764
rect 20898 10752 20904 10764
rect 20956 10752 20962 10804
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 17920 10628 18061 10656
rect 17920 10616 17926 10628
rect 18049 10625 18061 10628
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10625 20315 10659
rect 20257 10619 20315 10625
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 13446 10588 13452 10600
rect 13403 10560 13452 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 13446 10548 13452 10560
rect 13504 10588 13510 10600
rect 15102 10588 15108 10600
rect 13504 10560 15108 10588
rect 13504 10548 13510 10560
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 16114 10548 16120 10600
rect 16172 10588 16178 10600
rect 18598 10588 18604 10600
rect 16172 10560 18604 10588
rect 16172 10548 16178 10560
rect 18598 10548 18604 10560
rect 18656 10588 18662 10600
rect 20073 10591 20131 10597
rect 20073 10588 20085 10591
rect 18656 10560 20085 10588
rect 18656 10548 18662 10560
rect 20073 10557 20085 10560
rect 20119 10588 20131 10591
rect 20346 10588 20352 10600
rect 20119 10560 20352 10588
rect 20119 10557 20131 10560
rect 20073 10551 20131 10557
rect 20346 10548 20352 10560
rect 20404 10548 20410 10600
rect 20714 10588 20720 10600
rect 20675 10560 20720 10588
rect 20714 10548 20720 10560
rect 20772 10548 20778 10600
rect 13630 10529 13636 10532
rect 13624 10520 13636 10529
rect 13591 10492 13636 10520
rect 13624 10483 13636 10492
rect 13630 10480 13636 10483
rect 13688 10480 13694 10532
rect 15258 10523 15316 10529
rect 15258 10520 15270 10523
rect 14752 10492 15270 10520
rect 10778 10412 10784 10464
rect 10836 10452 10842 10464
rect 11333 10455 11391 10461
rect 11333 10452 11345 10455
rect 10836 10424 11345 10452
rect 10836 10412 10842 10424
rect 11333 10421 11345 10424
rect 11379 10421 11391 10455
rect 11333 10415 11391 10421
rect 11425 10455 11483 10461
rect 11425 10421 11437 10455
rect 11471 10452 11483 10455
rect 11790 10452 11796 10464
rect 11471 10424 11796 10452
rect 11471 10421 11483 10424
rect 11425 10415 11483 10421
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 14752 10461 14780 10492
rect 15258 10489 15270 10492
rect 15304 10520 15316 10523
rect 15838 10520 15844 10532
rect 15304 10492 15844 10520
rect 15304 10489 15316 10492
rect 15258 10483 15316 10489
rect 15838 10480 15844 10492
rect 15896 10480 15902 10532
rect 15930 10480 15936 10532
rect 15988 10520 15994 10532
rect 17129 10523 17187 10529
rect 17129 10520 17141 10523
rect 15988 10492 17141 10520
rect 15988 10480 15994 10492
rect 17129 10489 17141 10492
rect 17175 10489 17187 10523
rect 17129 10483 17187 10489
rect 18316 10523 18374 10529
rect 18316 10489 18328 10523
rect 18362 10520 18374 10523
rect 18506 10520 18512 10532
rect 18362 10492 18512 10520
rect 18362 10489 18374 10492
rect 18316 10483 18374 10489
rect 18506 10480 18512 10492
rect 18564 10480 18570 10532
rect 14737 10455 14795 10461
rect 14737 10421 14749 10455
rect 14783 10421 14795 10455
rect 17034 10452 17040 10464
rect 16995 10424 17040 10452
rect 14737 10415 14795 10421
rect 17034 10412 17040 10424
rect 17092 10412 17098 10464
rect 19702 10452 19708 10464
rect 19663 10424 19708 10452
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 20162 10412 20168 10464
rect 20220 10452 20226 10464
rect 20220 10424 20265 10452
rect 20220 10412 20226 10424
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 10778 10248 10784 10260
rect 10739 10220 10784 10248
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 12621 10251 12679 10257
rect 12621 10217 12633 10251
rect 12667 10217 12679 10251
rect 12621 10211 12679 10217
rect 11508 10183 11566 10189
rect 11508 10149 11520 10183
rect 11554 10180 11566 10183
rect 11606 10180 11612 10192
rect 11554 10152 11612 10180
rect 11554 10149 11566 10152
rect 11508 10143 11566 10149
rect 11606 10140 11612 10152
rect 11664 10140 11670 10192
rect 12636 10180 12664 10211
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 13688 10220 14289 10248
rect 13688 10208 13694 10220
rect 14277 10217 14289 10220
rect 14323 10217 14335 10251
rect 14277 10211 14335 10217
rect 15289 10251 15347 10257
rect 15289 10217 15301 10251
rect 15335 10248 15347 10251
rect 15930 10248 15936 10260
rect 15335 10220 15936 10248
rect 15335 10217 15347 10220
rect 15289 10211 15347 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16301 10251 16359 10257
rect 16301 10217 16313 10251
rect 16347 10248 16359 10251
rect 17034 10248 17040 10260
rect 16347 10220 17040 10248
rect 16347 10217 16359 10220
rect 16301 10211 16359 10217
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 17586 10208 17592 10260
rect 17644 10248 17650 10260
rect 17865 10251 17923 10257
rect 17865 10248 17877 10251
rect 17644 10220 17877 10248
rect 17644 10208 17650 10220
rect 17865 10217 17877 10220
rect 17911 10217 17923 10251
rect 17865 10211 17923 10217
rect 13142 10183 13200 10189
rect 13142 10180 13154 10183
rect 12636 10152 13154 10180
rect 13142 10149 13154 10152
rect 13188 10180 13200 10183
rect 13262 10180 13268 10192
rect 13188 10152 13268 10180
rect 13188 10149 13200 10152
rect 13142 10143 13200 10149
rect 13262 10140 13268 10152
rect 13320 10140 13326 10192
rect 15749 10183 15807 10189
rect 15749 10149 15761 10183
rect 15795 10180 15807 10183
rect 17126 10180 17132 10192
rect 15795 10152 17132 10180
rect 15795 10149 15807 10152
rect 15749 10143 15807 10149
rect 17126 10140 17132 10152
rect 17184 10140 17190 10192
rect 19052 10183 19110 10189
rect 19052 10149 19064 10183
rect 19098 10180 19110 10183
rect 19426 10180 19432 10192
rect 19098 10152 19432 10180
rect 19098 10149 19110 10152
rect 19052 10143 19110 10149
rect 19426 10140 19432 10152
rect 19484 10140 19490 10192
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10112 12955 10115
rect 13446 10112 13452 10124
rect 12943 10084 13452 10112
rect 12943 10081 12955 10084
rect 12897 10075 12955 10081
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 14366 10072 14372 10124
rect 14424 10112 14430 10124
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 14424 10084 14749 10112
rect 14424 10072 14430 10084
rect 14737 10081 14749 10084
rect 14783 10081 14795 10115
rect 15654 10112 15660 10124
rect 15615 10084 15660 10112
rect 14737 10075 14795 10081
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 16850 10112 16856 10124
rect 16811 10084 16856 10112
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17862 10072 17868 10124
rect 17920 10112 17926 10124
rect 18782 10112 18788 10124
rect 17920 10084 18788 10112
rect 17920 10072 17926 10084
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 10226 10004 10232 10056
rect 10284 10044 10290 10056
rect 11241 10047 11299 10053
rect 11241 10044 11253 10047
rect 10284 10016 11253 10044
rect 10284 10004 10290 10016
rect 11241 10013 11253 10016
rect 11287 10013 11299 10047
rect 15838 10044 15844 10056
rect 15799 10016 15844 10044
rect 11241 10007 11299 10013
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 16758 10004 16764 10056
rect 16816 10044 16822 10056
rect 17037 10047 17095 10053
rect 17037 10044 17049 10047
rect 16816 10016 17049 10044
rect 16816 10004 16822 10016
rect 17037 10013 17049 10016
rect 17083 10013 17095 10047
rect 17037 10007 17095 10013
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10044 18383 10047
rect 18506 10044 18512 10056
rect 18371 10016 18512 10044
rect 18371 10013 18383 10016
rect 18325 10007 18383 10013
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 14553 9911 14611 9917
rect 14553 9877 14565 9911
rect 14599 9908 14611 9911
rect 15010 9908 15016 9920
rect 14599 9880 15016 9908
rect 14599 9877 14611 9880
rect 14553 9871 14611 9877
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 20162 9908 20168 9920
rect 20123 9880 20168 9908
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 11606 9704 11612 9716
rect 11567 9676 11612 9704
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 12434 9704 12440 9716
rect 11756 9676 12440 9704
rect 11756 9664 11762 9676
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 18690 9664 18696 9716
rect 18748 9704 18754 9716
rect 18966 9704 18972 9716
rect 18748 9676 18972 9704
rect 18748 9664 18754 9676
rect 18966 9664 18972 9676
rect 19024 9664 19030 9716
rect 12713 9639 12771 9645
rect 12713 9605 12725 9639
rect 12759 9636 12771 9639
rect 13538 9636 13544 9648
rect 12759 9608 13544 9636
rect 12759 9605 12771 9608
rect 12713 9599 12771 9605
rect 13538 9596 13544 9608
rect 13596 9596 13602 9648
rect 16485 9639 16543 9645
rect 16485 9605 16497 9639
rect 16531 9636 16543 9639
rect 16531 9608 18000 9636
rect 16531 9605 16543 9608
rect 16485 9599 16543 9605
rect 13262 9568 13268 9580
rect 13223 9540 13268 9568
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 17034 9568 17040 9580
rect 16995 9540 17040 9568
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 9858 9500 9864 9512
rect 9732 9472 9864 9500
rect 9732 9460 9738 9472
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 10226 9500 10232 9512
rect 10187 9472 10232 9500
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 13081 9503 13139 9509
rect 13081 9500 13093 9503
rect 10336 9472 13093 9500
rect 7558 9392 7564 9444
rect 7616 9432 7622 9444
rect 10336 9432 10364 9472
rect 13081 9469 13093 9472
rect 13127 9469 13139 9503
rect 13081 9463 13139 9469
rect 7616 9404 10364 9432
rect 10496 9435 10554 9441
rect 7616 9392 7622 9404
rect 10496 9401 10508 9435
rect 10542 9432 10554 9435
rect 11054 9432 11060 9444
rect 10542 9404 11060 9432
rect 10542 9401 10554 9404
rect 10496 9395 10554 9401
rect 11054 9392 11060 9404
rect 11112 9392 11118 9444
rect 16853 9435 16911 9441
rect 16853 9401 16865 9435
rect 16899 9432 16911 9435
rect 17497 9435 17555 9441
rect 17497 9432 17509 9435
rect 16899 9404 17509 9432
rect 16899 9401 16911 9404
rect 16853 9395 16911 9401
rect 17497 9401 17509 9404
rect 17543 9401 17555 9435
rect 17972 9432 18000 9608
rect 18782 9568 18788 9580
rect 18743 9540 18788 9568
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 18233 9503 18291 9509
rect 18233 9469 18245 9503
rect 18279 9500 18291 9503
rect 18598 9500 18604 9512
rect 18279 9472 18604 9500
rect 18279 9469 18291 9472
rect 18233 9463 18291 9469
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 19052 9503 19110 9509
rect 19052 9469 19064 9503
rect 19098 9500 19110 9503
rect 19334 9500 19340 9512
rect 19098 9472 19340 9500
rect 19098 9469 19110 9472
rect 19052 9463 19110 9469
rect 19334 9460 19340 9472
rect 19392 9500 19398 9512
rect 20162 9500 20168 9512
rect 19392 9472 20168 9500
rect 19392 9460 19398 9472
rect 20162 9460 20168 9472
rect 20220 9460 20226 9512
rect 20530 9500 20536 9512
rect 20491 9472 20536 9500
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 19518 9432 19524 9444
rect 17972 9404 19524 9432
rect 17497 9395 17555 9401
rect 19518 9392 19524 9404
rect 19576 9392 19582 9444
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 9585 9367 9643 9373
rect 9585 9364 9597 9367
rect 8996 9336 9597 9364
rect 8996 9324 9002 9336
rect 9585 9333 9597 9336
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 10134 9364 10140 9376
rect 9824 9336 10140 9364
rect 9824 9324 9830 9336
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 13173 9367 13231 9373
rect 13173 9333 13185 9367
rect 13219 9364 13231 9367
rect 13814 9364 13820 9376
rect 13219 9336 13820 9364
rect 13219 9333 13231 9336
rect 13173 9327 13231 9333
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 16945 9367 17003 9373
rect 16945 9364 16957 9367
rect 16724 9336 16957 9364
rect 16724 9324 16730 9336
rect 16945 9333 16957 9336
rect 16991 9333 17003 9367
rect 16945 9327 17003 9333
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18417 9367 18475 9373
rect 18417 9364 18429 9367
rect 18012 9336 18429 9364
rect 18012 9324 18018 9336
rect 18417 9333 18429 9336
rect 18463 9333 18475 9367
rect 18417 9327 18475 9333
rect 19058 9324 19064 9376
rect 19116 9364 19122 9376
rect 19242 9364 19248 9376
rect 19116 9336 19248 9364
rect 19116 9324 19122 9336
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 20162 9364 20168 9376
rect 20123 9336 20168 9364
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 20717 9367 20775 9373
rect 20717 9333 20729 9367
rect 20763 9364 20775 9367
rect 20898 9364 20904 9376
rect 20763 9336 20904 9364
rect 20763 9333 20775 9336
rect 20717 9327 20775 9333
rect 20898 9324 20904 9336
rect 20956 9324 20962 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9129 8631 9163
rect 8938 9160 8944 9172
rect 8899 9132 8944 9160
rect 8573 9123 8631 9129
rect 8588 9092 8616 9123
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9033 9163 9091 9169
rect 9033 9129 9045 9163
rect 9079 9160 9091 9163
rect 11054 9160 11060 9172
rect 9079 9132 10272 9160
rect 11015 9132 11060 9160
rect 9079 9129 9091 9132
rect 9033 9123 9091 9129
rect 10244 9104 10272 9132
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9129 14243 9163
rect 18506 9160 18512 9172
rect 18467 9132 18512 9160
rect 14185 9123 14243 9129
rect 9858 9092 9864 9104
rect 8588 9064 9864 9092
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 10226 9052 10232 9104
rect 10284 9052 10290 9104
rect 14200 9092 14228 9123
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 18601 9163 18659 9169
rect 18601 9129 18613 9163
rect 18647 9160 18659 9163
rect 19702 9160 19708 9172
rect 18647 9132 19708 9160
rect 18647 9129 18659 9132
rect 18601 9123 18659 9129
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 19518 9092 19524 9104
rect 14200 9064 19524 9092
rect 19518 9052 19524 9064
rect 19576 9052 19582 9104
rect 842 8984 848 9036
rect 900 9024 906 9036
rect 7558 9024 7564 9036
rect 900 8996 7564 9024
rect 900 8984 906 8996
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 9950 9033 9956 9036
rect 9944 9024 9956 9033
rect 9232 8996 9956 9024
rect 9232 8965 9260 8996
rect 9944 8987 9956 8996
rect 9950 8984 9956 8987
rect 10008 8984 10014 9036
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 9024 12035 9027
rect 14366 9024 14372 9036
rect 12023 8996 14372 9024
rect 12023 8993 12035 8996
rect 11977 8987 12035 8993
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 14550 9024 14556 9036
rect 14511 8996 14556 9024
rect 14550 8984 14556 8996
rect 14608 8984 14614 9036
rect 15102 8984 15108 9036
rect 15160 9024 15166 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15160 8996 15669 9024
rect 15160 8984 15166 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 15924 9027 15982 9033
rect 15924 8993 15936 9027
rect 15970 9024 15982 9027
rect 16390 9024 16396 9036
rect 15970 8996 16396 9024
rect 15970 8993 15982 8996
rect 15924 8987 15982 8993
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 17405 9027 17463 9033
rect 17405 8993 17417 9027
rect 17451 9024 17463 9027
rect 19420 9027 19478 9033
rect 17451 8996 18184 9024
rect 17451 8993 17463 8996
rect 17405 8987 17463 8993
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 9732 8928 9825 8956
rect 9732 8916 9738 8928
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 14645 8959 14703 8965
rect 14645 8956 14657 8959
rect 13964 8928 14657 8956
rect 13964 8916 13970 8928
rect 14645 8925 14657 8928
rect 14691 8925 14703 8959
rect 14645 8919 14703 8925
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 14792 8928 14837 8956
rect 14792 8916 14798 8928
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17589 8959 17647 8965
rect 17589 8956 17601 8959
rect 17368 8928 17601 8956
rect 17368 8916 17374 8928
rect 17589 8925 17601 8928
rect 17635 8925 17647 8959
rect 17589 8919 17647 8925
rect 8570 8848 8576 8900
rect 8628 8888 8634 8900
rect 9692 8888 9720 8916
rect 18156 8897 18184 8996
rect 19420 8993 19432 9027
rect 19466 9024 19478 9027
rect 20162 9024 20168 9036
rect 19466 8996 20168 9024
rect 19466 8993 19478 8996
rect 19420 8987 19478 8993
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 18785 8959 18843 8965
rect 18785 8925 18797 8959
rect 18831 8956 18843 8959
rect 18831 8928 19012 8956
rect 18831 8925 18843 8928
rect 18785 8919 18843 8925
rect 18141 8891 18199 8897
rect 8628 8860 9720 8888
rect 10612 8860 11928 8888
rect 8628 8848 8634 8860
rect 2958 8780 2964 8832
rect 3016 8820 3022 8832
rect 10612 8820 10640 8860
rect 3016 8792 10640 8820
rect 3016 8780 3022 8792
rect 11606 8780 11612 8832
rect 11664 8820 11670 8832
rect 11793 8823 11851 8829
rect 11793 8820 11805 8823
rect 11664 8792 11805 8820
rect 11664 8780 11670 8792
rect 11793 8789 11805 8792
rect 11839 8789 11851 8823
rect 11900 8820 11928 8860
rect 18141 8857 18153 8891
rect 18187 8857 18199 8891
rect 18141 8851 18199 8857
rect 16850 8820 16856 8832
rect 11900 8792 16856 8820
rect 11793 8783 11851 8789
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 17034 8820 17040 8832
rect 16995 8792 17040 8820
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 18984 8820 19012 8928
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 19153 8959 19211 8965
rect 19153 8956 19165 8959
rect 19116 8928 19165 8956
rect 19116 8916 19122 8928
rect 19153 8925 19165 8928
rect 19199 8925 19211 8959
rect 19153 8919 19211 8925
rect 19334 8820 19340 8832
rect 18984 8792 19340 8820
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 19794 8780 19800 8832
rect 19852 8820 19858 8832
rect 20533 8823 20591 8829
rect 20533 8820 20545 8823
rect 19852 8792 20545 8820
rect 19852 8780 19858 8792
rect 20533 8789 20545 8792
rect 20579 8789 20591 8823
rect 20533 8783 20591 8789
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 1452 8588 10609 8616
rect 1452 8576 1458 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 10597 8579 10655 8585
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8616 10747 8619
rect 11790 8616 11796 8628
rect 10735 8588 11796 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 14734 8616 14740 8628
rect 14695 8588 14740 8616
rect 14734 8576 14740 8588
rect 14792 8576 14798 8628
rect 16390 8616 16396 8628
rect 14844 8588 16068 8616
rect 16351 8588 16396 8616
rect 14844 8548 14872 8588
rect 14384 8520 14872 8548
rect 8570 8480 8576 8492
rect 8531 8452 8576 8480
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 9600 8452 11008 8480
rect 4706 8372 4712 8424
rect 4764 8412 4770 8424
rect 9600 8412 9628 8452
rect 4764 8384 9628 8412
rect 10980 8412 11008 8452
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11241 8483 11299 8489
rect 11241 8480 11253 8483
rect 11112 8452 11253 8480
rect 11112 8440 11118 8452
rect 11241 8449 11253 8452
rect 11287 8449 11299 8483
rect 11241 8443 11299 8449
rect 10980 8384 11192 8412
rect 4764 8372 4770 8384
rect 8840 8347 8898 8353
rect 8840 8313 8852 8347
rect 8886 8344 8898 8347
rect 9582 8344 9588 8356
rect 8886 8316 9588 8344
rect 8886 8313 8898 8316
rect 8840 8307 8898 8313
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 10597 8347 10655 8353
rect 10597 8313 10609 8347
rect 10643 8344 10655 8347
rect 11057 8347 11115 8353
rect 11057 8344 11069 8347
rect 10643 8316 11069 8344
rect 10643 8313 10655 8316
rect 10597 8307 10655 8313
rect 11057 8313 11069 8316
rect 11103 8313 11115 8347
rect 11164 8344 11192 8384
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 13320 8384 13369 8412
rect 13320 8372 13326 8384
rect 13357 8381 13369 8384
rect 13403 8381 13415 8415
rect 14384 8412 14412 8520
rect 14734 8440 14740 8492
rect 14792 8480 14798 8492
rect 14792 8452 15148 8480
rect 14792 8440 14798 8452
rect 13357 8375 13415 8381
rect 13464 8384 14412 8412
rect 15013 8415 15071 8421
rect 13464 8344 13492 8384
rect 15013 8381 15025 8415
rect 15059 8381 15071 8415
rect 15120 8412 15148 8452
rect 15269 8415 15327 8421
rect 15269 8412 15281 8415
rect 15120 8384 15281 8412
rect 15013 8375 15071 8381
rect 15269 8381 15281 8384
rect 15315 8381 15327 8415
rect 16040 8412 16068 8588
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 16666 8616 16672 8628
rect 16627 8588 16672 8616
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 19352 8588 19656 8616
rect 16408 8480 16436 8576
rect 16850 8508 16856 8560
rect 16908 8548 16914 8560
rect 19352 8548 19380 8588
rect 16908 8520 19380 8548
rect 16908 8508 16914 8520
rect 19628 8492 19656 8588
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 16408 8452 17233 8480
rect 17221 8449 17233 8452
rect 17267 8449 17279 8483
rect 19610 8480 19616 8492
rect 19571 8452 19616 8480
rect 17221 8443 17279 8449
rect 19610 8440 19616 8452
rect 19668 8440 19674 8492
rect 20162 8440 20168 8492
rect 20220 8480 20226 8492
rect 20533 8483 20591 8489
rect 20533 8480 20545 8483
rect 20220 8452 20545 8480
rect 20220 8440 20226 8452
rect 20533 8449 20545 8452
rect 20579 8449 20591 8483
rect 20533 8443 20591 8449
rect 17037 8415 17095 8421
rect 17037 8412 17049 8415
rect 16040 8384 17049 8412
rect 15269 8375 15327 8381
rect 17037 8381 17049 8384
rect 17083 8381 17095 8415
rect 20346 8412 20352 8424
rect 20307 8384 20352 8412
rect 17037 8375 17095 8381
rect 11164 8316 13492 8344
rect 13624 8347 13682 8353
rect 11057 8307 11115 8313
rect 13624 8313 13636 8347
rect 13670 8344 13682 8347
rect 13998 8344 14004 8356
rect 13670 8316 14004 8344
rect 13670 8313 13682 8316
rect 13624 8307 13682 8313
rect 13998 8304 14004 8316
rect 14056 8304 14062 8356
rect 9950 8276 9956 8288
rect 9911 8248 9956 8276
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 11149 8279 11207 8285
rect 11149 8245 11161 8279
rect 11195 8276 11207 8279
rect 11790 8276 11796 8288
rect 11195 8248 11796 8276
rect 11195 8245 11207 8248
rect 11149 8239 11207 8245
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 15028 8276 15056 8375
rect 20346 8372 20352 8384
rect 20404 8372 20410 8424
rect 17126 8304 17132 8356
rect 17184 8344 17190 8356
rect 20438 8344 20444 8356
rect 17184 8316 17229 8344
rect 20399 8316 20444 8344
rect 17184 8304 17190 8316
rect 20438 8304 20444 8316
rect 20496 8304 20502 8356
rect 15470 8276 15476 8288
rect 12492 8248 12537 8276
rect 15028 8248 15476 8276
rect 12492 8236 12498 8248
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 18414 8236 18420 8288
rect 18472 8276 18478 8288
rect 18969 8279 19027 8285
rect 18969 8276 18981 8279
rect 18472 8248 18981 8276
rect 18472 8236 18478 8248
rect 18969 8245 18981 8248
rect 19015 8245 19027 8279
rect 19334 8276 19340 8288
rect 19295 8248 19340 8276
rect 18969 8239 19027 8245
rect 19334 8236 19340 8248
rect 19392 8236 19398 8288
rect 19429 8279 19487 8285
rect 19429 8245 19441 8279
rect 19475 8276 19487 8279
rect 19981 8279 20039 8285
rect 19981 8276 19993 8279
rect 19475 8248 19993 8276
rect 19475 8245 19487 8248
rect 19429 8239 19487 8245
rect 19981 8245 19993 8248
rect 20027 8245 20039 8279
rect 19981 8239 20039 8245
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 11606 8032 11612 8084
rect 11664 8032 11670 8084
rect 13998 8072 14004 8084
rect 13959 8044 14004 8072
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14608 8044 14657 8072
rect 14608 8032 14614 8044
rect 14645 8041 14657 8044
rect 14691 8041 14703 8075
rect 15470 8072 15476 8084
rect 15383 8044 15476 8072
rect 14645 8035 14703 8041
rect 15470 8032 15476 8044
rect 15528 8072 15534 8084
rect 19153 8075 19211 8081
rect 15528 8044 16344 8072
rect 15528 8032 15534 8044
rect 8570 8004 8576 8016
rect 7944 7976 8576 8004
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 7944 7945 7972 7976
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 11624 8004 11652 8032
rect 11974 8004 11980 8016
rect 10704 7976 11980 8004
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 7340 7908 7941 7936
rect 7340 7896 7346 7908
rect 7929 7905 7941 7908
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 8196 7939 8254 7945
rect 8196 7905 8208 7939
rect 8242 7936 8254 7939
rect 8662 7936 8668 7948
rect 8242 7908 8668 7936
rect 8242 7905 8254 7908
rect 8196 7899 8254 7905
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 10704 7945 10732 7976
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 12866 8007 12924 8013
rect 12866 8004 12878 8007
rect 12676 7976 12878 8004
rect 12676 7964 12682 7976
rect 12866 7973 12878 7976
rect 12912 7973 12924 8007
rect 12866 7967 12924 7973
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7905 10747 7939
rect 10689 7899 10747 7905
rect 11232 7939 11290 7945
rect 11232 7905 11244 7939
rect 11278 7936 11290 7939
rect 11606 7936 11612 7948
rect 11278 7908 11612 7936
rect 11278 7905 11290 7908
rect 11232 7899 11290 7905
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 13262 7936 13268 7948
rect 12636 7908 13268 7936
rect 12636 7877 12664 7908
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 15010 7896 15016 7948
rect 15068 7936 15074 7948
rect 16316 7945 16344 8044
rect 19153 8041 19165 8075
rect 19199 8072 19211 8075
rect 19334 8072 19340 8084
rect 19199 8044 19340 8072
rect 19199 8041 19211 8044
rect 19153 8035 19211 8041
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 16568 8007 16626 8013
rect 16568 7973 16580 8007
rect 16614 8004 16626 8007
rect 17034 8004 17040 8016
rect 16614 7976 17040 8004
rect 16614 7973 16626 7976
rect 16568 7967 16626 7973
rect 17034 7964 17040 7976
rect 17092 7964 17098 8016
rect 19242 7964 19248 8016
rect 19300 8004 19306 8016
rect 20257 8007 20315 8013
rect 20257 8004 20269 8007
rect 19300 7976 20269 8004
rect 19300 7964 19306 7976
rect 20257 7973 20269 7976
rect 20303 7973 20315 8007
rect 20257 7967 20315 7973
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15068 7908 15669 7936
rect 15068 7896 15074 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 16301 7939 16359 7945
rect 16301 7905 16313 7939
rect 16347 7936 16359 7939
rect 16390 7936 16396 7948
rect 16347 7908 16396 7936
rect 16347 7905 16359 7908
rect 16301 7899 16359 7905
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 18414 7936 18420 7948
rect 18375 7908 18420 7936
rect 18414 7896 18420 7908
rect 18472 7896 18478 7948
rect 20165 7939 20223 7945
rect 20165 7936 20177 7939
rect 18524 7908 20177 7936
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 12621 7871 12679 7877
rect 12621 7837 12633 7871
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 10686 7760 10692 7812
rect 10744 7800 10750 7812
rect 10980 7800 11008 7831
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 18524 7868 18552 7908
rect 20165 7905 20177 7908
rect 20211 7905 20223 7939
rect 20165 7899 20223 7905
rect 18690 7868 18696 7880
rect 17920 7840 18552 7868
rect 18651 7840 18696 7868
rect 17920 7828 17926 7840
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 18966 7828 18972 7880
rect 19024 7868 19030 7880
rect 20349 7871 20407 7877
rect 20349 7868 20361 7871
rect 19024 7840 20361 7868
rect 19024 7828 19030 7840
rect 20349 7837 20361 7840
rect 20395 7837 20407 7871
rect 20349 7831 20407 7837
rect 10744 7772 11008 7800
rect 10744 7760 10750 7772
rect 14550 7760 14556 7812
rect 14608 7800 14614 7812
rect 14608 7772 15608 7800
rect 14608 7760 14614 7772
rect 9309 7735 9367 7741
rect 9309 7701 9321 7735
rect 9355 7732 9367 7735
rect 9582 7732 9588 7744
rect 9355 7704 9588 7732
rect 9355 7701 9367 7704
rect 9309 7695 9367 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 9766 7692 9772 7744
rect 9824 7732 9830 7744
rect 9950 7732 9956 7744
rect 9824 7704 9956 7732
rect 9824 7692 9830 7704
rect 9950 7692 9956 7704
rect 10008 7732 10014 7744
rect 10505 7735 10563 7741
rect 10505 7732 10517 7735
rect 10008 7704 10517 7732
rect 10008 7692 10014 7704
rect 10505 7701 10517 7704
rect 10551 7701 10563 7735
rect 10505 7695 10563 7701
rect 12345 7735 12403 7741
rect 12345 7701 12357 7735
rect 12391 7732 12403 7735
rect 12618 7732 12624 7744
rect 12391 7704 12624 7732
rect 12391 7701 12403 7704
rect 12345 7695 12403 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 15580 7732 15608 7772
rect 17681 7735 17739 7741
rect 17681 7732 17693 7735
rect 15580 7704 17693 7732
rect 17681 7701 17693 7704
rect 17727 7701 17739 7735
rect 17681 7695 17739 7701
rect 19797 7735 19855 7741
rect 19797 7701 19809 7735
rect 19843 7732 19855 7735
rect 20346 7732 20352 7744
rect 19843 7704 20352 7732
rect 19843 7701 19855 7704
rect 19797 7695 19855 7701
rect 20346 7692 20352 7704
rect 20404 7692 20410 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 8846 7488 8852 7540
rect 8904 7528 8910 7540
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 8904 7500 8953 7528
rect 8904 7488 8910 7500
rect 8941 7497 8953 7500
rect 8987 7497 8999 7531
rect 8941 7491 8999 7497
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10226 7528 10232 7540
rect 9999 7500 10232 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 13449 7531 13507 7537
rect 13449 7497 13461 7531
rect 13495 7528 13507 7531
rect 13906 7528 13912 7540
rect 13495 7500 13912 7528
rect 13495 7497 13507 7500
rect 13449 7491 13507 7497
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 14274 7488 14280 7540
rect 14332 7528 14338 7540
rect 14461 7531 14519 7537
rect 14461 7528 14473 7531
rect 14332 7500 14473 7528
rect 14332 7488 14338 7500
rect 14461 7497 14473 7500
rect 14507 7497 14519 7531
rect 14461 7491 14519 7497
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7282 7392 7288 7404
rect 6880 7364 7288 7392
rect 6880 7352 6886 7364
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 8680 7392 8708 7488
rect 11057 7463 11115 7469
rect 11057 7429 11069 7463
rect 11103 7460 11115 7463
rect 12526 7460 12532 7472
rect 11103 7432 12532 7460
rect 11103 7429 11115 7432
rect 11057 7423 11115 7429
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 19610 7460 19616 7472
rect 19523 7432 19616 7460
rect 19610 7420 19616 7432
rect 19668 7460 19674 7472
rect 19668 7432 20484 7460
rect 19668 7420 19674 7432
rect 9493 7395 9551 7401
rect 9493 7392 9505 7395
rect 8680 7364 9505 7392
rect 9493 7361 9505 7364
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 9640 7364 10517 7392
rect 9640 7352 9646 7364
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 11606 7392 11612 7404
rect 11567 7364 11612 7392
rect 10505 7355 10563 7361
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 13998 7392 14004 7404
rect 13959 7364 14004 7392
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 15013 7395 15071 7401
rect 15013 7392 15025 7395
rect 14332 7364 15025 7392
rect 14332 7352 14338 7364
rect 15013 7361 15025 7364
rect 15059 7361 15071 7395
rect 17126 7392 17132 7404
rect 17087 7364 17132 7392
rect 15013 7355 15071 7361
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 20346 7392 20352 7404
rect 20307 7364 20352 7392
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 20456 7401 20484 7432
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 9306 7324 9312 7336
rect 9267 7296 9312 7324
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 13872 7296 13921 7324
rect 13872 7284 13878 7296
rect 13909 7293 13921 7296
rect 13955 7324 13967 7327
rect 15102 7324 15108 7336
rect 13955 7296 15108 7324
rect 13955 7293 13967 7296
rect 13909 7287 13967 7293
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 18233 7327 18291 7333
rect 18233 7293 18245 7327
rect 18279 7293 18291 7327
rect 18233 7287 18291 7293
rect 18500 7327 18558 7333
rect 18500 7293 18512 7327
rect 18546 7324 18558 7327
rect 18782 7324 18788 7336
rect 18546 7296 18788 7324
rect 18546 7293 18558 7296
rect 18500 7287 18558 7293
rect 7552 7259 7610 7265
rect 7552 7225 7564 7259
rect 7598 7256 7610 7259
rect 8386 7256 8392 7268
rect 7598 7228 8392 7256
rect 7598 7225 7610 7228
rect 7552 7219 7610 7225
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 8570 7216 8576 7268
rect 8628 7256 8634 7268
rect 11425 7259 11483 7265
rect 11425 7256 11437 7259
rect 8628 7228 11437 7256
rect 8628 7216 8634 7228
rect 11425 7225 11437 7228
rect 11471 7225 11483 7259
rect 11425 7219 11483 7225
rect 13998 7216 14004 7268
rect 14056 7256 14062 7268
rect 14921 7259 14979 7265
rect 14921 7256 14933 7259
rect 14056 7228 14933 7256
rect 14056 7216 14062 7228
rect 14921 7225 14933 7228
rect 14967 7225 14979 7259
rect 18248 7256 18276 7287
rect 18782 7284 18788 7296
rect 18840 7324 18846 7336
rect 18966 7324 18972 7336
rect 18840 7296 18972 7324
rect 18840 7284 18846 7296
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 18598 7256 18604 7268
rect 18248 7228 18604 7256
rect 14921 7219 14979 7225
rect 18598 7216 18604 7228
rect 18656 7256 18662 7268
rect 19058 7256 19064 7268
rect 18656 7228 19064 7256
rect 18656 7216 18662 7228
rect 19058 7216 19064 7228
rect 19116 7216 19122 7268
rect 9398 7188 9404 7200
rect 9359 7160 9404 7188
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10321 7191 10379 7197
rect 10321 7188 10333 7191
rect 9916 7160 10333 7188
rect 9916 7148 9922 7160
rect 10321 7157 10333 7160
rect 10367 7157 10379 7191
rect 10321 7151 10379 7157
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 11517 7191 11575 7197
rect 10468 7160 10513 7188
rect 10468 7148 10474 7160
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 11790 7188 11796 7200
rect 11563 7160 11796 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 11790 7148 11796 7160
rect 11848 7188 11854 7200
rect 12342 7188 12348 7200
rect 11848 7160 12348 7188
rect 11848 7148 11854 7160
rect 12342 7148 12348 7160
rect 12400 7148 12406 7200
rect 12894 7148 12900 7200
rect 12952 7188 12958 7200
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 12952 7160 13277 7188
rect 12952 7148 12958 7160
rect 13265 7157 13277 7160
rect 13311 7188 13323 7191
rect 13817 7191 13875 7197
rect 13817 7188 13829 7191
rect 13311 7160 13829 7188
rect 13311 7157 13323 7160
rect 13265 7151 13323 7157
rect 13817 7157 13829 7160
rect 13863 7157 13875 7191
rect 13817 7151 13875 7157
rect 14090 7148 14096 7200
rect 14148 7188 14154 7200
rect 14829 7191 14887 7197
rect 14829 7188 14841 7191
rect 14148 7160 14841 7188
rect 14148 7148 14154 7160
rect 14829 7157 14841 7160
rect 14875 7157 14887 7191
rect 14829 7151 14887 7157
rect 16485 7191 16543 7197
rect 16485 7157 16497 7191
rect 16531 7188 16543 7191
rect 16666 7188 16672 7200
rect 16531 7160 16672 7188
rect 16531 7157 16543 7160
rect 16485 7151 16543 7157
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 16850 7188 16856 7200
rect 16811 7160 16856 7188
rect 16850 7148 16856 7160
rect 16908 7148 16914 7200
rect 16942 7148 16948 7200
rect 17000 7188 17006 7200
rect 17000 7160 17045 7188
rect 17000 7148 17006 7160
rect 19702 7148 19708 7200
rect 19760 7188 19766 7200
rect 19889 7191 19947 7197
rect 19889 7188 19901 7191
rect 19760 7160 19901 7188
rect 19760 7148 19766 7160
rect 19889 7157 19901 7160
rect 19935 7157 19947 7191
rect 20254 7188 20260 7200
rect 20215 7160 20260 7188
rect 19889 7151 19947 7157
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 11425 6987 11483 6993
rect 11425 6953 11437 6987
rect 11471 6984 11483 6987
rect 11606 6984 11612 6996
rect 11471 6956 11612 6984
rect 11471 6953 11483 6956
rect 11425 6947 11483 6953
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 12492 6956 12537 6984
rect 12492 6944 12498 6956
rect 16666 6944 16672 6996
rect 16724 6984 16730 6996
rect 17865 6987 17923 6993
rect 17865 6984 17877 6987
rect 16724 6956 17877 6984
rect 16724 6944 16730 6956
rect 17865 6953 17877 6956
rect 17911 6953 17923 6987
rect 17865 6947 17923 6953
rect 12526 6916 12532 6928
rect 12487 6888 12532 6916
rect 12526 6876 12532 6888
rect 12584 6876 12590 6928
rect 13262 6916 13268 6928
rect 12912 6888 13268 6916
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 9306 6848 9312 6860
rect 8251 6820 9312 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 10312 6851 10370 6857
rect 10312 6817 10324 6851
rect 10358 6848 10370 6851
rect 10594 6848 10600 6860
rect 10358 6820 10600 6848
rect 10358 6817 10370 6820
rect 10312 6811 10370 6817
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 11974 6848 11980 6860
rect 11935 6820 11980 6848
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12434 6848 12440 6860
rect 12360 6820 12440 6848
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 12360 6780 12388 6820
rect 12434 6808 12440 6820
rect 12492 6848 12498 6860
rect 12912 6857 12940 6888
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 14550 6876 14556 6928
rect 14608 6876 14614 6928
rect 15746 6876 15752 6928
rect 15804 6916 15810 6928
rect 16390 6916 16396 6928
rect 15804 6888 16396 6916
rect 15804 6876 15810 6888
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 12492 6820 12909 6848
rect 12492 6808 12498 6820
rect 12897 6817 12909 6820
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 13164 6851 13222 6857
rect 13164 6817 13176 6851
rect 13210 6848 13222 6851
rect 14568 6848 14596 6876
rect 16005 6851 16063 6857
rect 16005 6848 16017 6851
rect 13210 6820 14596 6848
rect 15672 6820 16017 6848
rect 13210 6817 13222 6820
rect 13164 6811 13222 6817
rect 12618 6780 12624 6792
rect 10045 6743 10103 6749
rect 11808 6752 12388 6780
rect 12579 6752 12624 6780
rect 10060 6644 10088 6743
rect 11808 6721 11836 6752
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 13964 6752 14565 6780
rect 13964 6740 13970 6752
rect 14553 6749 14565 6752
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 11793 6715 11851 6721
rect 11793 6681 11805 6715
rect 11839 6681 11851 6715
rect 11793 6675 11851 6681
rect 12069 6715 12127 6721
rect 12069 6681 12081 6715
rect 12115 6712 12127 6715
rect 12710 6712 12716 6724
rect 12115 6684 12716 6712
rect 12115 6681 12127 6684
rect 12069 6675 12127 6681
rect 12710 6672 12716 6684
rect 12768 6672 12774 6724
rect 10686 6644 10692 6656
rect 10060 6616 10692 6644
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 14274 6644 14280 6656
rect 14235 6616 14280 6644
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 15672 6644 15700 6820
rect 16005 6817 16017 6820
rect 16051 6817 16063 6851
rect 16005 6811 16063 6817
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 17773 6851 17831 6857
rect 17773 6848 17785 6851
rect 16632 6820 17785 6848
rect 16632 6808 16638 6820
rect 17773 6817 17785 6820
rect 17819 6817 17831 6851
rect 18598 6848 18604 6860
rect 18559 6820 18604 6848
rect 17773 6811 17831 6817
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 18868 6851 18926 6857
rect 18868 6817 18880 6851
rect 18914 6848 18926 6851
rect 19610 6848 19616 6860
rect 18914 6820 19616 6848
rect 18914 6817 18926 6820
rect 18868 6811 18926 6817
rect 19610 6808 19616 6820
rect 19668 6808 19674 6860
rect 15746 6740 15752 6792
rect 15804 6780 15810 6792
rect 15804 6752 15849 6780
rect 15804 6740 15810 6752
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17957 6783 18015 6789
rect 17957 6780 17969 6783
rect 17276 6752 17969 6780
rect 17276 6740 17282 6752
rect 17957 6749 17969 6752
rect 18003 6749 18015 6783
rect 17957 6743 18015 6749
rect 19886 6740 19892 6792
rect 19944 6780 19950 6792
rect 20257 6783 20315 6789
rect 20257 6780 20269 6783
rect 19944 6752 20269 6780
rect 19944 6740 19950 6752
rect 20257 6749 20269 6752
rect 20303 6749 20315 6783
rect 20257 6743 20315 6749
rect 17126 6712 17132 6724
rect 17087 6684 17132 6712
rect 17126 6672 17132 6684
rect 17184 6672 17190 6724
rect 17402 6712 17408 6724
rect 17363 6684 17408 6712
rect 17402 6672 17408 6684
rect 17460 6672 17466 6724
rect 16666 6644 16672 6656
rect 15672 6616 16672 6644
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 19794 6604 19800 6656
rect 19852 6644 19858 6656
rect 19981 6647 20039 6653
rect 19981 6644 19993 6647
rect 19852 6616 19993 6644
rect 19852 6604 19858 6616
rect 19981 6613 19993 6616
rect 20027 6613 20039 6647
rect 19981 6607 20039 6613
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 8386 6440 8392 6452
rect 8347 6412 8392 6440
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 9861 6443 9919 6449
rect 9861 6409 9873 6443
rect 9907 6440 9919 6443
rect 10042 6440 10048 6452
rect 9907 6412 10048 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 13998 6440 14004 6452
rect 13959 6412 14004 6440
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 15746 6440 15752 6452
rect 15028 6412 15752 6440
rect 12989 6375 13047 6381
rect 12989 6341 13001 6375
rect 13035 6372 13047 6375
rect 14090 6372 14096 6384
rect 13035 6344 14096 6372
rect 13035 6341 13047 6344
rect 12989 6335 13047 6341
rect 14090 6332 14096 6344
rect 14148 6332 14154 6384
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 7009 6307 7067 6313
rect 7009 6304 7021 6307
rect 6880 6276 7021 6304
rect 6880 6264 6886 6276
rect 7009 6273 7021 6276
rect 7055 6273 7067 6307
rect 10502 6304 10508 6316
rect 10463 6276 10508 6304
rect 7009 6267 7067 6273
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 13633 6307 13691 6313
rect 13633 6273 13645 6307
rect 13679 6304 13691 6307
rect 14550 6304 14556 6316
rect 13679 6276 14556 6304
rect 13679 6273 13691 6276
rect 13633 6267 13691 6273
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 15028 6313 15056 6412
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 16945 6443 17003 6449
rect 16945 6440 16957 6443
rect 16908 6412 16957 6440
rect 16908 6400 16914 6412
rect 16945 6409 16957 6412
rect 16991 6409 17003 6443
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 16945 6403 17003 6409
rect 17420 6412 19073 6440
rect 16022 6332 16028 6384
rect 16080 6372 16086 6384
rect 17420 6372 17448 6412
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 19061 6403 19119 6409
rect 19150 6400 19156 6452
rect 19208 6440 19214 6452
rect 19245 6443 19303 6449
rect 19245 6440 19257 6443
rect 19208 6412 19257 6440
rect 19208 6400 19214 6412
rect 19245 6409 19257 6412
rect 19291 6409 19303 6443
rect 20254 6440 20260 6452
rect 20215 6412 20260 6440
rect 19245 6403 19303 6409
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 16080 6344 17448 6372
rect 16080 6332 16086 6344
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6236 13415 6239
rect 13906 6236 13912 6248
rect 13403 6208 13912 6236
rect 13403 6205 13415 6208
rect 13357 6199 13415 6205
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 15280 6239 15338 6245
rect 15280 6205 15292 6239
rect 15326 6236 15338 6239
rect 17126 6236 17132 6248
rect 15326 6208 17132 6236
rect 15326 6205 15338 6208
rect 15280 6199 15338 6205
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 17328 6245 17356 6344
rect 18782 6332 18788 6384
rect 18840 6372 18846 6384
rect 18840 6344 20208 6372
rect 18840 6332 18846 6344
rect 17494 6304 17500 6316
rect 17455 6276 17500 6304
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 18892 6313 18920 6344
rect 18877 6307 18935 6313
rect 18877 6273 18889 6307
rect 18923 6304 18935 6307
rect 19702 6304 19708 6316
rect 18923 6276 18957 6304
rect 19663 6276 19708 6304
rect 18923 6273 18935 6276
rect 18877 6267 18935 6273
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 19794 6264 19800 6316
rect 19852 6304 19858 6316
rect 20180 6304 20208 6344
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 19852 6276 19897 6304
rect 20180 6276 20821 6304
rect 19852 6264 19858 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 17402 6196 17408 6248
rect 17460 6236 17466 6248
rect 20717 6239 20775 6245
rect 20717 6236 20729 6239
rect 17460 6208 20729 6236
rect 17460 6196 17466 6208
rect 20717 6205 20729 6208
rect 20763 6236 20775 6239
rect 21082 6236 21088 6248
rect 20763 6208 21088 6236
rect 20763 6205 20775 6208
rect 20717 6199 20775 6205
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 7276 6171 7334 6177
rect 7276 6137 7288 6171
rect 7322 6168 7334 6171
rect 7742 6168 7748 6180
rect 7322 6140 7748 6168
rect 7322 6137 7334 6140
rect 7276 6131 7334 6137
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 10229 6171 10287 6177
rect 10229 6137 10241 6171
rect 10275 6168 10287 6171
rect 10873 6171 10931 6177
rect 10873 6168 10885 6171
rect 10275 6140 10885 6168
rect 10275 6137 10287 6140
rect 10229 6131 10287 6137
rect 10873 6137 10885 6140
rect 10919 6137 10931 6171
rect 10873 6131 10931 6137
rect 15470 6128 15476 6180
rect 15528 6168 15534 6180
rect 18601 6171 18659 6177
rect 18601 6168 18613 6171
rect 15528 6140 18613 6168
rect 15528 6128 15534 6140
rect 18601 6137 18613 6140
rect 18647 6137 18659 6171
rect 18601 6131 18659 6137
rect 19061 6171 19119 6177
rect 19061 6137 19073 6171
rect 19107 6168 19119 6171
rect 20530 6168 20536 6180
rect 19107 6140 20536 6168
rect 19107 6137 19119 6140
rect 19061 6131 19119 6137
rect 20530 6128 20536 6140
rect 20588 6168 20594 6180
rect 20625 6171 20683 6177
rect 20625 6168 20637 6171
rect 20588 6140 20637 6168
rect 20588 6128 20594 6140
rect 20625 6137 20637 6140
rect 20671 6137 20683 6171
rect 20625 6131 20683 6137
rect 10318 6100 10324 6112
rect 10279 6072 10324 6100
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 13449 6103 13507 6109
rect 13449 6100 13461 6103
rect 12308 6072 13461 6100
rect 12308 6060 12314 6072
rect 13449 6069 13461 6072
rect 13495 6069 13507 6103
rect 14366 6100 14372 6112
rect 14327 6072 14372 6100
rect 13449 6063 13507 6069
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 14458 6060 14464 6112
rect 14516 6100 14522 6112
rect 14516 6072 14561 6100
rect 14516 6060 14522 6072
rect 15102 6060 15108 6112
rect 15160 6100 15166 6112
rect 16022 6100 16028 6112
rect 15160 6072 16028 6100
rect 15160 6060 15166 6072
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 16393 6103 16451 6109
rect 16393 6100 16405 6103
rect 16264 6072 16405 6100
rect 16264 6060 16270 6072
rect 16393 6069 16405 6072
rect 16439 6100 16451 6103
rect 17218 6100 17224 6112
rect 16439 6072 17224 6100
rect 16439 6069 16451 6072
rect 16393 6063 16451 6069
rect 17218 6060 17224 6072
rect 17276 6060 17282 6112
rect 17402 6100 17408 6112
rect 17363 6072 17408 6100
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 18230 6100 18236 6112
rect 18191 6072 18236 6100
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 19150 6100 19156 6112
rect 18739 6072 19156 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 19150 6060 19156 6072
rect 19208 6060 19214 6112
rect 19610 6100 19616 6112
rect 19571 6072 19616 6100
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 7742 5896 7748 5908
rect 7703 5868 7748 5896
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8021 5899 8079 5905
rect 8021 5865 8033 5899
rect 8067 5896 8079 5899
rect 8202 5896 8208 5908
rect 8067 5868 8208 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8435 5868 9045 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 10502 5856 10508 5908
rect 10560 5896 10566 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 10560 5868 11069 5896
rect 10560 5856 10566 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 15470 5896 15476 5908
rect 11057 5859 11115 5865
rect 11164 5868 15476 5896
rect 6822 5828 6828 5840
rect 6380 5800 6828 5828
rect 6380 5769 6408 5800
rect 6822 5788 6828 5800
rect 6880 5788 6886 5840
rect 7760 5828 7788 5856
rect 7760 5800 8616 5828
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 6632 5763 6690 5769
rect 6632 5729 6644 5763
rect 6678 5760 6690 5763
rect 8202 5760 8208 5772
rect 6678 5732 8208 5760
rect 6678 5729 6690 5732
rect 6632 5723 6690 5729
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 8478 5692 8484 5704
rect 8439 5664 8484 5692
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 8588 5701 8616 5800
rect 10778 5788 10784 5840
rect 10836 5828 10842 5840
rect 11164 5828 11192 5868
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 15841 5899 15899 5905
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16574 5896 16580 5908
rect 15887 5868 16580 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 16942 5896 16948 5908
rect 16903 5868 16948 5896
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 17218 5856 17224 5908
rect 17276 5896 17282 5908
rect 17313 5899 17371 5905
rect 17313 5896 17325 5899
rect 17276 5868 17325 5896
rect 17276 5856 17282 5868
rect 17313 5865 17325 5868
rect 17359 5896 17371 5899
rect 17862 5896 17868 5908
rect 17359 5868 17868 5896
rect 17359 5865 17371 5868
rect 17313 5859 17371 5865
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 18969 5899 19027 5905
rect 18969 5865 18981 5899
rect 19015 5896 19027 5899
rect 19610 5896 19616 5908
rect 19015 5868 19616 5896
rect 19015 5865 19027 5868
rect 18969 5859 19027 5865
rect 19610 5856 19616 5868
rect 19668 5856 19674 5908
rect 10836 5800 11192 5828
rect 11600 5831 11658 5837
rect 10836 5788 10842 5800
rect 11600 5797 11612 5831
rect 11646 5828 11658 5831
rect 14274 5828 14280 5840
rect 11646 5800 14280 5828
rect 11646 5797 11658 5800
rect 11600 5791 11658 5797
rect 14274 5788 14280 5800
rect 14332 5788 14338 5840
rect 14458 5788 14464 5840
rect 14516 5828 14522 5840
rect 14516 5800 16344 5828
rect 14516 5788 14522 5800
rect 9944 5763 10002 5769
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 10226 5760 10232 5772
rect 9990 5732 10232 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 10226 5720 10232 5732
rect 10284 5720 10290 5772
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 10744 5732 11345 5760
rect 10744 5720 10750 5732
rect 11333 5729 11345 5732
rect 11379 5760 11391 5763
rect 12434 5760 12440 5772
rect 11379 5732 12440 5760
rect 11379 5729 11391 5732
rect 11333 5723 11391 5729
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 15381 5763 15439 5769
rect 15381 5729 15393 5763
rect 15427 5760 15439 5763
rect 16209 5763 16267 5769
rect 16209 5760 16221 5763
rect 15427 5732 16221 5760
rect 15427 5729 15439 5732
rect 15381 5723 15439 5729
rect 16209 5729 16221 5732
rect 16255 5729 16267 5763
rect 16316 5760 16344 5800
rect 18230 5788 18236 5840
rect 18288 5828 18294 5840
rect 19429 5831 19487 5837
rect 19429 5828 19441 5831
rect 18288 5800 19441 5828
rect 18288 5788 18294 5800
rect 19429 5797 19441 5800
rect 19475 5797 19487 5831
rect 19429 5791 19487 5797
rect 19242 5760 19248 5772
rect 16316 5732 17264 5760
rect 16209 5723 16267 5729
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5661 8631 5695
rect 8573 5655 8631 5661
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 16298 5692 16304 5704
rect 16259 5664 16304 5692
rect 9677 5655 9735 5661
rect 9692 5556 9720 5655
rect 16298 5652 16304 5664
rect 16356 5652 16362 5704
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5692 16543 5695
rect 17126 5692 17132 5704
rect 16531 5664 17132 5692
rect 16531 5661 16543 5664
rect 16485 5655 16543 5661
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 17236 5692 17264 5732
rect 17420 5732 19248 5760
rect 17420 5701 17448 5732
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 19337 5763 19395 5769
rect 19337 5729 19349 5763
rect 19383 5760 19395 5763
rect 19886 5760 19892 5772
rect 19383 5732 19892 5760
rect 19383 5729 19395 5732
rect 19337 5723 19395 5729
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 20254 5760 20260 5772
rect 20215 5732 20260 5760
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 17405 5695 17463 5701
rect 17405 5692 17417 5695
rect 17236 5664 17417 5692
rect 17405 5661 17417 5664
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 17494 5652 17500 5704
rect 17552 5692 17558 5704
rect 19518 5692 19524 5704
rect 17552 5664 17645 5692
rect 19479 5664 19524 5692
rect 17552 5652 17558 5664
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 12268 5596 16620 5624
rect 9950 5556 9956 5568
rect 9692 5528 9956 5556
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 12268 5556 12296 5596
rect 12710 5556 12716 5568
rect 10468 5528 12296 5556
rect 12671 5528 12716 5556
rect 10468 5516 10474 5528
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 16592 5556 16620 5596
rect 16666 5584 16672 5636
rect 16724 5624 16730 5636
rect 17512 5624 17540 5652
rect 16724 5596 17540 5624
rect 16724 5584 16730 5596
rect 17402 5556 17408 5568
rect 16592 5528 17408 5556
rect 17402 5516 17408 5528
rect 17460 5516 17466 5568
rect 19058 5516 19064 5568
rect 19116 5556 19122 5568
rect 20441 5559 20499 5565
rect 20441 5556 20453 5559
rect 19116 5528 20453 5556
rect 19116 5516 19122 5528
rect 20441 5525 20453 5528
rect 20487 5525 20499 5559
rect 20441 5519 20499 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 8202 5352 8208 5364
rect 8163 5324 8208 5352
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 8481 5355 8539 5361
rect 8481 5321 8493 5355
rect 8527 5352 8539 5355
rect 9398 5352 9404 5364
rect 8527 5324 9404 5352
rect 8527 5321 8539 5324
rect 8481 5315 8539 5321
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 9585 5355 9643 5361
rect 9585 5321 9597 5355
rect 9631 5352 9643 5355
rect 10318 5352 10324 5364
rect 9631 5324 10324 5352
rect 9631 5321 9643 5324
rect 9585 5315 9643 5321
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 13265 5355 13323 5361
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13354 5352 13360 5364
rect 13311 5324 13360 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 15841 5355 15899 5361
rect 15841 5321 15853 5355
rect 15887 5352 15899 5355
rect 16298 5352 16304 5364
rect 15887 5324 16304 5352
rect 15887 5321 15899 5324
rect 15841 5315 15899 5321
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 18601 5355 18659 5361
rect 18601 5321 18613 5355
rect 18647 5352 18659 5355
rect 20070 5352 20076 5364
rect 18647 5324 20076 5352
rect 18647 5321 18659 5324
rect 18601 5315 18659 5321
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 6822 5216 6828 5228
rect 6783 5188 6828 5216
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 8386 5176 8392 5228
rect 8444 5216 8450 5228
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 8444 5188 9045 5216
rect 8444 5176 8450 5188
rect 9033 5185 9045 5188
rect 9079 5185 9091 5219
rect 10226 5216 10232 5228
rect 10187 5188 10232 5216
rect 9033 5179 9091 5185
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10686 5216 10692 5228
rect 10647 5188 10692 5216
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 13814 5216 13820 5228
rect 13775 5188 13820 5216
rect 13814 5176 13820 5188
rect 13872 5176 13878 5228
rect 14550 5176 14556 5228
rect 14608 5216 14614 5228
rect 14829 5219 14887 5225
rect 14829 5216 14841 5219
rect 14608 5188 14841 5216
rect 14608 5176 14614 5188
rect 14829 5185 14841 5188
rect 14875 5185 14887 5219
rect 14829 5179 14887 5185
rect 16485 5219 16543 5225
rect 16485 5185 16497 5219
rect 16531 5216 16543 5219
rect 16666 5216 16672 5228
rect 16531 5188 16672 5216
rect 16531 5185 16543 5188
rect 16485 5179 16543 5185
rect 16666 5176 16672 5188
rect 16724 5176 16730 5228
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 18598 5216 18604 5228
rect 18012 5188 18604 5216
rect 18012 5176 18018 5188
rect 18598 5176 18604 5188
rect 18656 5216 18662 5228
rect 18969 5219 19027 5225
rect 18969 5216 18981 5219
rect 18656 5188 18981 5216
rect 18656 5176 18662 5188
rect 18969 5185 18981 5188
rect 19015 5185 19027 5219
rect 18969 5179 19027 5185
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 6972 5120 9965 5148
rect 6972 5108 6978 5120
rect 9953 5117 9965 5120
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 10045 5151 10103 5157
rect 10045 5117 10057 5151
rect 10091 5148 10103 5151
rect 10410 5148 10416 5160
rect 10091 5120 10416 5148
rect 10091 5117 10103 5120
rect 10045 5111 10103 5117
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 14458 5108 14464 5160
rect 14516 5148 14522 5160
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 14516 5120 14749 5148
rect 14516 5108 14522 5120
rect 14737 5117 14749 5120
rect 14783 5117 14795 5151
rect 18414 5148 18420 5160
rect 18375 5120 18420 5148
rect 14737 5111 14795 5117
rect 18414 5108 18420 5120
rect 18472 5108 18478 5160
rect 19236 5151 19294 5157
rect 19236 5117 19248 5151
rect 19282 5148 19294 5151
rect 19794 5148 19800 5160
rect 19282 5120 19800 5148
rect 19282 5117 19294 5120
rect 19236 5111 19294 5117
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 20622 5148 20628 5160
rect 20583 5120 20628 5148
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 7092 5083 7150 5089
rect 7092 5049 7104 5083
rect 7138 5080 7150 5083
rect 10956 5083 11014 5089
rect 7138 5052 10456 5080
rect 7138 5049 7150 5052
rect 7092 5043 7150 5049
rect 8846 5012 8852 5024
rect 8807 4984 8852 5012
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 8938 4972 8944 5024
rect 8996 5012 9002 5024
rect 10428 5012 10456 5052
rect 10956 5049 10968 5083
rect 11002 5080 11014 5083
rect 12710 5080 12716 5092
rect 11002 5052 12716 5080
rect 11002 5049 11014 5052
rect 10956 5043 11014 5049
rect 12710 5040 12716 5052
rect 12768 5040 12774 5092
rect 14366 5040 14372 5092
rect 14424 5080 14430 5092
rect 14645 5083 14703 5089
rect 14645 5080 14657 5083
rect 14424 5052 14657 5080
rect 14424 5040 14430 5052
rect 14645 5049 14657 5052
rect 14691 5080 14703 5083
rect 16301 5083 16359 5089
rect 16301 5080 16313 5083
rect 14691 5052 16313 5080
rect 14691 5049 14703 5052
rect 14645 5043 14703 5049
rect 16301 5049 16313 5052
rect 16347 5080 16359 5083
rect 19150 5080 19156 5092
rect 16347 5052 19156 5080
rect 16347 5049 16359 5052
rect 16301 5043 16359 5049
rect 19150 5040 19156 5052
rect 19208 5040 19214 5092
rect 19812 5052 20852 5080
rect 19812 5024 19840 5052
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 8996 4984 9041 5012
rect 10428 4984 12081 5012
rect 8996 4972 9002 4984
rect 12069 4981 12081 4984
rect 12115 5012 12127 5015
rect 12158 5012 12164 5024
rect 12115 4984 12164 5012
rect 12115 4981 12127 4984
rect 12069 4975 12127 4981
rect 12158 4972 12164 4984
rect 12216 4972 12222 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 13630 5012 13636 5024
rect 12492 4984 12537 5012
rect 13591 4984 13636 5012
rect 12492 4972 12498 4984
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13725 5015 13783 5021
rect 13725 4981 13737 5015
rect 13771 5012 13783 5015
rect 14277 5015 14335 5021
rect 14277 5012 14289 5015
rect 13771 4984 14289 5012
rect 13771 4981 13783 4984
rect 13725 4975 13783 4981
rect 14277 4981 14289 4984
rect 14323 4981 14335 5015
rect 14277 4975 14335 4981
rect 15194 4972 15200 5024
rect 15252 5012 15258 5024
rect 16209 5015 16267 5021
rect 16209 5012 16221 5015
rect 15252 4984 16221 5012
rect 15252 4972 15258 4984
rect 16209 4981 16221 4984
rect 16255 4981 16267 5015
rect 16209 4975 16267 4981
rect 19794 4972 19800 5024
rect 19852 4972 19858 5024
rect 20346 5012 20352 5024
rect 20307 4984 20352 5012
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 20824 5021 20852 5052
rect 20809 5015 20867 5021
rect 20809 4981 20821 5015
rect 20855 4981 20867 5015
rect 20809 4975 20867 4981
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 7009 4811 7067 4817
rect 7009 4777 7021 4811
rect 7055 4808 7067 4811
rect 8478 4808 8484 4820
rect 7055 4780 8484 4808
rect 7055 4777 7067 4780
rect 7009 4771 7067 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 10134 4808 10140 4820
rect 8619 4780 10140 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10226 4768 10232 4820
rect 10284 4808 10290 4820
rect 11057 4811 11115 4817
rect 11057 4808 11069 4811
rect 10284 4780 11069 4808
rect 10284 4768 10290 4780
rect 11057 4777 11069 4780
rect 11103 4777 11115 4811
rect 11057 4771 11115 4777
rect 11609 4811 11667 4817
rect 11609 4777 11621 4811
rect 11655 4808 11667 4811
rect 11698 4808 11704 4820
rect 11655 4780 11704 4808
rect 11655 4777 11667 4780
rect 11609 4771 11667 4777
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 11977 4811 12035 4817
rect 11977 4777 11989 4811
rect 12023 4808 12035 4811
rect 12434 4808 12440 4820
rect 12023 4780 12440 4808
rect 12023 4777 12035 4780
rect 11977 4771 12035 4777
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 13630 4768 13636 4820
rect 13688 4808 13694 4820
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 13688 4780 15301 4808
rect 13688 4768 13694 4780
rect 15289 4777 15301 4780
rect 15335 4777 15347 4811
rect 15289 4771 15347 4777
rect 17494 4768 17500 4820
rect 17552 4808 17558 4820
rect 17865 4811 17923 4817
rect 17865 4808 17877 4811
rect 17552 4780 17877 4808
rect 17552 4768 17558 4780
rect 17865 4777 17877 4780
rect 17911 4777 17923 4811
rect 17865 4771 17923 4777
rect 18233 4811 18291 4817
rect 18233 4777 18245 4811
rect 18279 4808 18291 4811
rect 18874 4808 18880 4820
rect 18279 4780 18880 4808
rect 18279 4777 18291 4780
rect 18233 4771 18291 4777
rect 18874 4768 18880 4780
rect 18932 4768 18938 4820
rect 8941 4743 8999 4749
rect 8941 4709 8953 4743
rect 8987 4740 8999 4743
rect 9674 4740 9680 4752
rect 8987 4712 9680 4740
rect 8987 4709 8999 4712
rect 8941 4703 8999 4709
rect 9674 4700 9680 4712
rect 9732 4700 9738 4752
rect 10502 4700 10508 4752
rect 10560 4740 10566 4752
rect 15749 4743 15807 4749
rect 15749 4740 15761 4743
rect 10560 4712 15761 4740
rect 10560 4700 10566 4712
rect 15749 4709 15761 4712
rect 15795 4709 15807 4743
rect 15749 4703 15807 4709
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 5316 4644 7389 4672
rect 5316 4632 5322 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 9766 4672 9772 4684
rect 7377 4635 7435 4641
rect 9232 4644 9772 4672
rect 7466 4604 7472 4616
rect 7427 4576 7472 4604
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 8202 4604 8208 4616
rect 7699 4576 8208 4604
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 9030 4604 9036 4616
rect 8991 4576 9036 4604
rect 9030 4564 9036 4576
rect 9088 4564 9094 4616
rect 9232 4613 9260 4644
rect 9766 4632 9772 4644
rect 9824 4672 9830 4684
rect 9933 4675 9991 4681
rect 9933 4672 9945 4675
rect 9824 4644 9945 4672
rect 9824 4632 9830 4644
rect 9933 4641 9945 4644
rect 9979 4641 9991 4675
rect 12066 4672 12072 4684
rect 12027 4644 12072 4672
rect 9933 4635 9991 4641
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 12526 4632 12532 4684
rect 12584 4672 12590 4684
rect 13078 4672 13084 4684
rect 12584 4644 13084 4672
rect 12584 4632 12590 4644
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13348 4675 13406 4681
rect 13348 4641 13360 4675
rect 13394 4672 13406 4675
rect 14642 4672 14648 4684
rect 13394 4644 14648 4672
rect 13394 4641 13406 4644
rect 13348 4635 13406 4641
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 14783 4644 15669 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 16752 4675 16810 4681
rect 16752 4641 16764 4675
rect 16798 4672 16810 4675
rect 18598 4672 18604 4684
rect 16798 4644 18368 4672
rect 18559 4644 18604 4672
rect 16798 4641 16810 4644
rect 16752 4635 16810 4641
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4573 9735 4607
rect 12158 4604 12164 4616
rect 12119 4576 12164 4604
rect 9677 4567 9735 4573
rect 9692 4468 9720 4567
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 16482 4604 16488 4616
rect 16443 4576 16488 4604
rect 15841 4567 15899 4573
rect 14642 4496 14648 4548
rect 14700 4536 14706 4548
rect 15856 4536 15884 4567
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 18340 4604 18368 4644
rect 18598 4632 18604 4644
rect 18656 4632 18662 4684
rect 18693 4675 18751 4681
rect 18693 4641 18705 4675
rect 18739 4672 18751 4675
rect 19702 4672 19708 4684
rect 18739 4644 19708 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 19702 4632 19708 4644
rect 19760 4632 19766 4684
rect 19886 4672 19892 4684
rect 19847 4644 19892 4672
rect 19886 4632 19892 4644
rect 19944 4632 19950 4684
rect 18782 4604 18788 4616
rect 18340 4576 18788 4604
rect 18782 4564 18788 4576
rect 18840 4564 18846 4616
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19981 4607 20039 4613
rect 19981 4604 19993 4607
rect 19392 4576 19993 4604
rect 19392 4564 19398 4576
rect 19981 4573 19993 4576
rect 20027 4573 20039 4607
rect 20162 4604 20168 4616
rect 20075 4576 20168 4604
rect 19981 4567 20039 4573
rect 20162 4564 20168 4576
rect 20220 4604 20226 4616
rect 20346 4604 20352 4616
rect 20220 4576 20352 4604
rect 20220 4564 20226 4576
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 14700 4508 15884 4536
rect 14700 4496 14706 4508
rect 9950 4468 9956 4480
rect 9692 4440 9956 4468
rect 9950 4428 9956 4440
rect 10008 4468 10014 4480
rect 10318 4468 10324 4480
rect 10008 4440 10324 4468
rect 10008 4428 10014 4440
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 11606 4428 11612 4480
rect 11664 4468 11670 4480
rect 13814 4468 13820 4480
rect 11664 4440 13820 4468
rect 11664 4428 11670 4440
rect 13814 4428 13820 4440
rect 13872 4468 13878 4480
rect 14461 4471 14519 4477
rect 14461 4468 14473 4471
rect 13872 4440 14473 4468
rect 13872 4428 13878 4440
rect 14461 4437 14473 4440
rect 14507 4437 14519 4471
rect 19518 4468 19524 4480
rect 19479 4440 19524 4468
rect 14461 4431 14519 4437
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 7742 4264 7748 4276
rect 7524 4236 7748 4264
rect 7524 4224 7530 4236
rect 7742 4224 7748 4236
rect 7800 4264 7806 4276
rect 7800 4236 9444 4264
rect 7800 4224 7806 4236
rect 9416 4196 9444 4236
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 9861 4267 9919 4273
rect 9861 4264 9873 4267
rect 9824 4236 9873 4264
rect 9824 4224 9830 4236
rect 9861 4233 9873 4236
rect 9907 4233 9919 4267
rect 14642 4264 14648 4276
rect 9861 4227 9919 4233
rect 9968 4236 14504 4264
rect 14603 4236 14648 4264
rect 9968 4196 9996 4236
rect 10962 4196 10968 4208
rect 7944 4168 8340 4196
rect 9416 4168 9996 4196
rect 10923 4168 10968 4196
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 7650 4128 7656 4140
rect 6880 4100 7656 4128
rect 6880 4088 6886 4100
rect 7650 4088 7656 4100
rect 7708 4128 7714 4140
rect 7944 4128 7972 4168
rect 7708 4100 7972 4128
rect 8021 4131 8079 4137
rect 7708 4088 7714 4100
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8202 4128 8208 4140
rect 8067 4100 8208 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8312 4128 8340 4168
rect 10962 4156 10968 4168
rect 11020 4156 11026 4208
rect 14476 4196 14504 4236
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 17218 4264 17224 4276
rect 15488 4236 17224 4264
rect 15488 4196 15516 4236
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 19702 4264 19708 4276
rect 19663 4236 19708 4264
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 11348 4168 11652 4196
rect 14476 4168 15516 4196
rect 20901 4199 20959 4205
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 8312 4100 8493 4128
rect 8481 4097 8493 4100
rect 8527 4097 8539 4131
rect 11348 4128 11376 4168
rect 11514 4128 11520 4140
rect 8481 4091 8539 4097
rect 9508 4100 11376 4128
rect 11475 4100 11520 4128
rect 5350 4020 5356 4072
rect 5408 4060 5414 4072
rect 9508 4060 9536 4100
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 11624 4128 11652 4168
rect 20901 4165 20913 4199
rect 20947 4165 20959 4199
rect 20901 4159 20959 4165
rect 12250 4128 12256 4140
rect 11624 4100 12256 4128
rect 12250 4088 12256 4100
rect 12308 4088 12314 4140
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 13265 4131 13323 4137
rect 13265 4128 13277 4131
rect 13136 4100 13277 4128
rect 13136 4088 13142 4100
rect 13265 4097 13277 4100
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 16482 4088 16488 4140
rect 16540 4128 16546 4140
rect 17862 4128 17868 4140
rect 16540 4100 17868 4128
rect 16540 4088 16546 4100
rect 17862 4088 17868 4100
rect 17920 4128 17926 4140
rect 18046 4128 18052 4140
rect 17920 4100 18052 4128
rect 17920 4088 17926 4100
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 19576 4100 20177 4128
rect 19576 4088 19582 4100
rect 20165 4097 20177 4100
rect 20211 4097 20223 4131
rect 20346 4128 20352 4140
rect 20307 4100 20352 4128
rect 20165 4091 20223 4097
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 20916 4128 20944 4159
rect 20456 4100 20944 4128
rect 12437 4063 12495 4069
rect 5408 4032 9536 4060
rect 10152 4032 11560 4060
rect 5408 4020 5414 4032
rect 7558 3952 7564 4004
rect 7616 3992 7622 4004
rect 7837 3995 7895 4001
rect 7837 3992 7849 3995
rect 7616 3964 7849 3992
rect 7616 3952 7622 3964
rect 7837 3961 7849 3964
rect 7883 3961 7895 3995
rect 7837 3955 7895 3961
rect 8748 3995 8806 4001
rect 8748 3961 8760 3995
rect 8794 3992 8806 3995
rect 9306 3992 9312 4004
rect 8794 3964 9312 3992
rect 8794 3961 8806 3964
rect 8748 3955 8806 3961
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 6362 3884 6368 3936
rect 6420 3924 6426 3936
rect 6914 3924 6920 3936
rect 6420 3896 6920 3924
rect 6420 3884 6426 3896
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 7374 3924 7380 3936
rect 7335 3896 7380 3924
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3924 7803 3927
rect 8294 3924 8300 3936
rect 7791 3896 8300 3924
rect 7791 3893 7803 3896
rect 7745 3887 7803 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 10152 3924 10180 4032
rect 11146 3952 11152 4004
rect 11204 3992 11210 4004
rect 11425 3995 11483 4001
rect 11425 3992 11437 3995
rect 11204 3964 11437 3992
rect 11204 3952 11210 3964
rect 11425 3961 11437 3964
rect 11471 3961 11483 3995
rect 11532 3992 11560 4032
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 12802 4060 12808 4072
rect 12483 4032 12808 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 15378 4060 15384 4072
rect 13464 4032 15384 4060
rect 13464 3992 13492 4032
rect 15378 4020 15384 4032
rect 15436 4020 15442 4072
rect 15473 4063 15531 4069
rect 15473 4029 15485 4063
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 15740 4063 15798 4069
rect 15740 4029 15752 4063
rect 15786 4060 15798 4063
rect 16206 4060 16212 4072
rect 15786 4032 16212 4060
rect 15786 4029 15798 4032
rect 15740 4023 15798 4029
rect 11532 3964 13492 3992
rect 13532 3995 13590 4001
rect 11425 3955 11483 3961
rect 13532 3961 13544 3995
rect 13578 3992 13590 3995
rect 13814 3992 13820 4004
rect 13578 3964 13820 3992
rect 13578 3961 13590 3964
rect 13532 3955 13590 3961
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 15286 3952 15292 4004
rect 15344 3992 15350 4004
rect 15488 3992 15516 4023
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 16500 4060 16528 4088
rect 16316 4032 16528 4060
rect 17405 4063 17463 4069
rect 16316 3992 16344 4032
rect 17405 4029 17417 4063
rect 17451 4060 17463 4063
rect 17954 4060 17960 4072
rect 17451 4032 17960 4060
rect 17451 4029 17463 4032
rect 17405 4023 17463 4029
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 20456 4060 20484 4100
rect 20714 4060 20720 4072
rect 18156 4032 20484 4060
rect 20675 4032 20720 4060
rect 15344 3964 16344 3992
rect 15344 3952 15350 3964
rect 16390 3952 16396 4004
rect 16448 3992 16454 4004
rect 18156 3992 18184 4032
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 18322 4001 18328 4004
rect 18316 3992 18328 4001
rect 16448 3964 18184 3992
rect 18283 3964 18328 3992
rect 16448 3952 16454 3964
rect 18316 3955 18328 3964
rect 18322 3952 18328 3955
rect 18380 3952 18386 4004
rect 20806 3992 20812 4004
rect 18708 3964 20812 3992
rect 8996 3896 10180 3924
rect 11333 3927 11391 3933
rect 8996 3884 9002 3896
rect 11333 3893 11345 3927
rect 11379 3924 11391 3927
rect 11882 3924 11888 3936
rect 11379 3896 11888 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12621 3927 12679 3933
rect 12621 3924 12633 3927
rect 12032 3896 12633 3924
rect 12032 3884 12038 3896
rect 12621 3893 12633 3896
rect 12667 3893 12679 3927
rect 12621 3887 12679 3893
rect 15930 3884 15936 3936
rect 15988 3924 15994 3936
rect 16853 3927 16911 3933
rect 16853 3924 16865 3927
rect 15988 3896 16865 3924
rect 15988 3884 15994 3896
rect 16853 3893 16865 3896
rect 16899 3893 16911 3927
rect 16853 3887 16911 3893
rect 17589 3927 17647 3933
rect 17589 3893 17601 3927
rect 17635 3924 17647 3927
rect 18708 3924 18736 3964
rect 20806 3952 20812 3964
rect 20864 3952 20870 4004
rect 17635 3896 18736 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 18840 3896 19441 3924
rect 18840 3884 18846 3896
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 19429 3887 19487 3893
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 20073 3927 20131 3933
rect 20073 3924 20085 3927
rect 19576 3896 20085 3924
rect 19576 3884 19582 3896
rect 20073 3893 20085 3896
rect 20119 3893 20131 3927
rect 20073 3887 20131 3893
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 9306 3720 9312 3732
rect 9267 3692 9312 3720
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9674 3720 9680 3732
rect 9635 3692 9680 3720
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 11514 3720 11520 3732
rect 10520 3692 11520 3720
rect 3050 3612 3056 3664
rect 3108 3652 3114 3664
rect 5258 3652 5264 3664
rect 3108 3624 5264 3652
rect 3108 3612 3114 3624
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 6822 3652 6828 3664
rect 6288 3624 6828 3652
rect 6288 3593 6316 3624
rect 6822 3612 6828 3624
rect 6880 3612 6886 3664
rect 8202 3661 8208 3664
rect 8196 3652 8208 3661
rect 8163 3624 8208 3652
rect 8196 3615 8208 3624
rect 8202 3612 8208 3615
rect 8260 3612 8266 3664
rect 10520 3652 10548 3692
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 11977 3723 12035 3729
rect 11977 3689 11989 3723
rect 12023 3720 12035 3723
rect 12066 3720 12072 3732
rect 12023 3692 12072 3720
rect 12023 3689 12035 3692
rect 11977 3683 12035 3689
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 13170 3720 13176 3732
rect 12176 3692 13032 3720
rect 13131 3692 13176 3720
rect 9692 3624 10548 3652
rect 10588 3655 10646 3661
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 6540 3587 6598 3593
rect 6540 3553 6552 3587
rect 6586 3584 6598 3587
rect 9692 3584 9720 3624
rect 10588 3621 10600 3655
rect 10634 3652 10646 3655
rect 11606 3652 11612 3664
rect 10634 3624 11612 3652
rect 10634 3621 10646 3624
rect 10588 3615 10646 3621
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 12176 3652 12204 3692
rect 11716 3624 12204 3652
rect 13004 3652 13032 3692
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13633 3723 13691 3729
rect 13633 3689 13645 3723
rect 13679 3720 13691 3723
rect 14185 3723 14243 3729
rect 14185 3720 14197 3723
rect 13679 3692 14197 3720
rect 13679 3689 13691 3692
rect 13633 3683 13691 3689
rect 14185 3689 14197 3692
rect 14231 3689 14243 3723
rect 14185 3683 14243 3689
rect 14645 3723 14703 3729
rect 14645 3689 14657 3723
rect 14691 3720 14703 3723
rect 15289 3723 15347 3729
rect 15289 3720 15301 3723
rect 14691 3692 15301 3720
rect 14691 3689 14703 3692
rect 14645 3683 14703 3689
rect 15289 3689 15301 3692
rect 15335 3689 15347 3723
rect 15289 3683 15347 3689
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15657 3723 15715 3729
rect 15657 3720 15669 3723
rect 15436 3692 15669 3720
rect 15436 3680 15442 3692
rect 15657 3689 15669 3692
rect 15703 3720 15715 3723
rect 17589 3723 17647 3729
rect 17589 3720 17601 3723
rect 15703 3692 17601 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 17589 3689 17601 3692
rect 17635 3689 17647 3723
rect 17589 3683 17647 3689
rect 17681 3723 17739 3729
rect 17681 3689 17693 3723
rect 17727 3720 17739 3723
rect 18598 3720 18604 3732
rect 17727 3692 18604 3720
rect 17727 3689 17739 3692
rect 17681 3683 17739 3689
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 19334 3720 19340 3732
rect 18708 3692 19340 3720
rect 15194 3652 15200 3664
rect 13004 3624 15200 3652
rect 6586 3556 9720 3584
rect 6586 3553 6598 3556
rect 6540 3547 6598 3553
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 11716 3584 11744 3624
rect 15194 3612 15200 3624
rect 15252 3612 15258 3664
rect 17770 3652 17776 3664
rect 15580 3624 17776 3652
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 9824 3556 11744 3584
rect 12176 3556 12357 3584
rect 9824 3544 9830 3556
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 7708 3488 7941 3516
rect 7708 3476 7714 3488
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9858 3516 9864 3528
rect 9272 3488 9864 3516
rect 9272 3476 9278 3488
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 10318 3516 10324 3528
rect 10279 3488 10324 3516
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 12176 3448 12204 3556
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 12492 3556 12537 3584
rect 12492 3544 12498 3556
rect 12986 3544 12992 3596
rect 13044 3584 13050 3596
rect 13541 3587 13599 3593
rect 13541 3584 13553 3587
rect 13044 3556 13553 3584
rect 13044 3544 13050 3556
rect 13541 3553 13553 3556
rect 13587 3553 13599 3587
rect 13541 3547 13599 3553
rect 14553 3587 14611 3593
rect 14553 3553 14565 3587
rect 14599 3584 14611 3587
rect 15470 3584 15476 3596
rect 14599 3556 15476 3584
rect 14599 3553 14611 3556
rect 14553 3547 14611 3553
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3516 12679 3519
rect 12710 3516 12716 3528
rect 12667 3488 12716 3516
rect 12667 3485 12679 3488
rect 12621 3479 12679 3485
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 13814 3516 13820 3528
rect 13775 3488 13820 3516
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 14829 3519 14887 3525
rect 14829 3485 14841 3519
rect 14875 3485 14887 3519
rect 14829 3479 14887 3485
rect 7208 3420 7788 3448
rect 3602 3340 3608 3392
rect 3660 3380 3666 3392
rect 7208 3380 7236 3420
rect 7650 3380 7656 3392
rect 3660 3352 7236 3380
rect 7611 3352 7656 3380
rect 3660 3340 3666 3352
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 7760 3380 7788 3420
rect 11256 3420 12204 3448
rect 11256 3380 11284 3420
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 14844 3448 14872 3479
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 15580 3516 15608 3624
rect 17770 3612 17776 3624
rect 17828 3612 17834 3664
rect 18708 3652 18736 3692
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 20346 3680 20352 3732
rect 20404 3720 20410 3732
rect 20533 3723 20591 3729
rect 20533 3720 20545 3723
rect 20404 3692 20545 3720
rect 20404 3680 20410 3692
rect 20533 3689 20545 3692
rect 20579 3689 20591 3723
rect 20533 3683 20591 3689
rect 20364 3652 20392 3680
rect 17880 3624 18736 3652
rect 19076 3624 20392 3652
rect 15746 3584 15752 3596
rect 15659 3556 15752 3584
rect 15746 3544 15752 3556
rect 15804 3584 15810 3596
rect 17880 3584 17908 3624
rect 15804 3556 17908 3584
rect 18049 3587 18107 3593
rect 15804 3544 15810 3556
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 18693 3587 18751 3593
rect 18693 3584 18705 3587
rect 18095 3556 18705 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 18693 3553 18705 3556
rect 18739 3553 18751 3587
rect 18693 3547 18751 3553
rect 15930 3516 15936 3528
rect 15068 3488 15608 3516
rect 15891 3488 15936 3516
rect 15068 3476 15074 3488
rect 15930 3476 15936 3488
rect 15988 3476 15994 3528
rect 16206 3476 16212 3528
rect 16264 3516 16270 3528
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 16264 3488 18153 3516
rect 16264 3476 16270 3488
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18322 3516 18328 3528
rect 18235 3488 18328 3516
rect 18141 3479 18199 3485
rect 18322 3476 18328 3488
rect 18380 3516 18386 3528
rect 19076 3516 19104 3624
rect 19420 3587 19478 3593
rect 19420 3553 19432 3587
rect 19466 3584 19478 3587
rect 20162 3584 20168 3596
rect 19466 3556 20168 3584
rect 19466 3553 19478 3556
rect 19420 3547 19478 3553
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 18380 3488 19104 3516
rect 19153 3519 19211 3525
rect 18380 3476 18386 3488
rect 19153 3485 19165 3519
rect 19199 3485 19211 3519
rect 19153 3479 19211 3485
rect 16482 3448 16488 3460
rect 13688 3420 16488 3448
rect 13688 3408 13694 3420
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 17589 3451 17647 3457
rect 17589 3417 17601 3451
rect 17635 3448 17647 3451
rect 17635 3420 18184 3448
rect 17635 3417 17647 3420
rect 17589 3411 17647 3417
rect 11698 3380 11704 3392
rect 7760 3352 11284 3380
rect 11659 3352 11704 3380
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 18156 3380 18184 3420
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 19168 3448 19196 3479
rect 18288 3420 19196 3448
rect 18288 3408 18294 3420
rect 19886 3380 19892 3392
rect 18156 3352 19892 3380
rect 19886 3340 19892 3352
rect 19944 3340 19950 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 8202 3176 8208 3188
rect 5868 3148 7788 3176
rect 8163 3148 8208 3176
rect 5868 3136 5874 3148
rect 7760 3108 7788 3148
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8665 3179 8723 3185
rect 8665 3145 8677 3179
rect 8711 3176 8723 3179
rect 9030 3176 9036 3188
rect 8711 3148 9036 3176
rect 8711 3145 8723 3148
rect 8665 3139 8723 3145
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 13136 3148 13676 3176
rect 13136 3136 13142 3148
rect 8478 3108 8484 3120
rect 7760 3080 8484 3108
rect 8478 3068 8484 3080
rect 8536 3068 8542 3120
rect 11606 3068 11612 3120
rect 11664 3108 11670 3120
rect 11793 3111 11851 3117
rect 11793 3108 11805 3111
rect 11664 3080 11805 3108
rect 11664 3068 11670 3080
rect 11793 3077 11805 3080
rect 11839 3077 11851 3111
rect 13648 3108 13676 3148
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14093 3179 14151 3185
rect 14093 3176 14105 3179
rect 13872 3148 14105 3176
rect 13872 3136 13878 3148
rect 14093 3145 14105 3148
rect 14139 3145 14151 3179
rect 16945 3179 17003 3185
rect 16945 3176 16957 3179
rect 14093 3139 14151 3145
rect 14200 3148 16957 3176
rect 14200 3108 14228 3148
rect 16945 3145 16957 3148
rect 16991 3145 17003 3179
rect 16945 3139 17003 3145
rect 17129 3179 17187 3185
rect 17129 3145 17141 3179
rect 17175 3176 17187 3179
rect 19518 3176 19524 3188
rect 17175 3148 18920 3176
rect 19479 3148 19524 3176
rect 17175 3145 17187 3148
rect 17129 3139 17187 3145
rect 16482 3108 16488 3120
rect 13648 3080 14228 3108
rect 16443 3080 16488 3108
rect 11793 3071 11851 3077
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 18785 3111 18843 3117
rect 18785 3108 18797 3111
rect 18012 3080 18797 3108
rect 18012 3068 18018 3080
rect 18785 3077 18797 3080
rect 18831 3077 18843 3111
rect 18892 3108 18920 3148
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 20898 3108 20904 3120
rect 18892 3080 20904 3108
rect 18785 3071 18843 3077
rect 20898 3068 20904 3080
rect 20956 3068 20962 3120
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 8938 3000 8944 3052
rect 8996 3040 9002 3052
rect 9125 3043 9183 3049
rect 9125 3040 9137 3043
rect 8996 3012 9137 3040
rect 8996 3000 9002 3012
rect 9125 3009 9137 3012
rect 9171 3009 9183 3043
rect 9306 3040 9312 3052
rect 9267 3012 9312 3040
rect 9125 3003 9183 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 10376 3012 10425 3040
rect 10376 3000 10382 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 15013 3043 15071 3049
rect 15013 3040 15025 3043
rect 13780 3012 15025 3040
rect 13780 3000 13786 3012
rect 15013 3009 15025 3012
rect 15059 3009 15071 3043
rect 18966 3040 18972 3052
rect 15013 3003 15071 3009
rect 18616 3012 18972 3040
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 6914 2972 6920 2984
rect 4212 2944 6920 2972
rect 4212 2932 4218 2944
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 7092 2975 7150 2981
rect 7092 2941 7104 2975
rect 7138 2972 7150 2975
rect 7650 2972 7656 2984
rect 7138 2944 7656 2972
rect 7138 2941 7150 2944
rect 7092 2935 7150 2941
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 7892 2944 9168 2972
rect 7892 2932 7898 2944
rect 2498 2864 2504 2916
rect 2556 2904 2562 2916
rect 8846 2904 8852 2916
rect 2556 2876 8852 2904
rect 2556 2864 2562 2876
rect 8846 2864 8852 2876
rect 8904 2864 8910 2916
rect 6914 2796 6920 2848
rect 6972 2836 6978 2848
rect 9033 2839 9091 2845
rect 9033 2836 9045 2839
rect 6972 2808 9045 2836
rect 6972 2796 6978 2808
rect 9033 2805 9045 2808
rect 9079 2805 9091 2839
rect 9140 2836 9168 2944
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 10502 2972 10508 2984
rect 9456 2944 10508 2972
rect 9456 2932 9462 2944
rect 10502 2932 10508 2944
rect 10560 2932 10566 2984
rect 10680 2975 10738 2981
rect 10680 2941 10692 2975
rect 10726 2972 10738 2975
rect 11698 2972 11704 2984
rect 10726 2944 11704 2972
rect 10726 2941 10738 2944
rect 10680 2935 10738 2941
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 12713 2975 12771 2981
rect 12713 2972 12725 2975
rect 12584 2944 12725 2972
rect 12584 2932 12590 2944
rect 12713 2941 12725 2944
rect 12759 2941 12771 2975
rect 12713 2935 12771 2941
rect 15105 2975 15163 2981
rect 15105 2941 15117 2975
rect 15151 2972 15163 2975
rect 15194 2972 15200 2984
rect 15151 2944 15200 2972
rect 15151 2941 15163 2944
rect 15105 2935 15163 2941
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 15372 2975 15430 2981
rect 15372 2941 15384 2975
rect 15418 2972 15430 2975
rect 15930 2972 15936 2984
rect 15418 2944 15936 2972
rect 15418 2941 15430 2944
rect 15372 2935 15430 2941
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 16758 2972 16764 2984
rect 16719 2944 16764 2972
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 17310 2972 17316 2984
rect 17271 2944 17316 2972
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2972 18107 2975
rect 18506 2972 18512 2984
rect 18095 2944 18512 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18506 2932 18512 2944
rect 18564 2932 18570 2984
rect 18616 2981 18644 3012
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 20162 3040 20168 3052
rect 20123 3012 20168 3040
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 18601 2975 18659 2981
rect 18601 2941 18613 2975
rect 18647 2941 18659 2975
rect 19889 2975 19947 2981
rect 19889 2972 19901 2975
rect 18601 2935 18659 2941
rect 18708 2944 19901 2972
rect 12980 2907 13038 2913
rect 12980 2873 12992 2907
rect 13026 2904 13038 2907
rect 13630 2904 13636 2916
rect 13026 2876 13636 2904
rect 13026 2873 13038 2876
rect 12980 2867 13038 2873
rect 13630 2864 13636 2876
rect 13688 2864 13694 2916
rect 14182 2864 14188 2916
rect 14240 2904 14246 2916
rect 14240 2876 17540 2904
rect 14240 2864 14246 2876
rect 12158 2836 12164 2848
rect 9140 2808 12164 2836
rect 9033 2799 9091 2805
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 14366 2836 14372 2848
rect 14327 2808 14372 2836
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 17512 2845 17540 2876
rect 17862 2864 17868 2916
rect 17920 2904 17926 2916
rect 18708 2904 18736 2944
rect 19889 2941 19901 2944
rect 19935 2972 19947 2975
rect 19978 2972 19984 2984
rect 19935 2944 19984 2972
rect 19935 2941 19947 2944
rect 19889 2935 19947 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20530 2972 20536 2984
rect 20491 2944 20536 2972
rect 20530 2932 20536 2944
rect 20588 2932 20594 2984
rect 17920 2876 18736 2904
rect 17920 2864 17926 2876
rect 19150 2864 19156 2916
rect 19208 2904 19214 2916
rect 19208 2876 20024 2904
rect 19208 2864 19214 2876
rect 19996 2848 20024 2876
rect 15013 2839 15071 2845
rect 15013 2805 15025 2839
rect 15059 2836 15071 2839
rect 17129 2839 17187 2845
rect 17129 2836 17141 2839
rect 15059 2808 17141 2836
rect 15059 2805 15071 2808
rect 15013 2799 15071 2805
rect 17129 2805 17141 2808
rect 17175 2805 17187 2839
rect 17129 2799 17187 2805
rect 17497 2839 17555 2845
rect 17497 2805 17509 2839
rect 17543 2805 17555 2839
rect 17497 2799 17555 2805
rect 17586 2796 17592 2848
rect 17644 2836 17650 2848
rect 18233 2839 18291 2845
rect 18233 2836 18245 2839
rect 17644 2808 18245 2836
rect 17644 2796 17650 2808
rect 18233 2805 18245 2808
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 20717 2839 20775 2845
rect 20036 2808 20081 2836
rect 20036 2796 20042 2808
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 21910 2836 21916 2848
rect 20763 2808 21916 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 7285 2635 7343 2641
rect 7285 2601 7297 2635
rect 7331 2632 7343 2635
rect 7558 2632 7564 2644
rect 7331 2604 7564 2632
rect 7331 2601 7343 2604
rect 7285 2595 7343 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 7742 2632 7748 2644
rect 7703 2604 7748 2632
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 11057 2635 11115 2641
rect 11057 2601 11069 2635
rect 11103 2632 11115 2635
rect 11146 2632 11152 2644
rect 11103 2604 11152 2632
rect 11103 2601 11115 2604
rect 11057 2595 11115 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11517 2635 11575 2641
rect 11517 2601 11529 2635
rect 11563 2632 11575 2635
rect 11790 2632 11796 2644
rect 11563 2604 11796 2632
rect 11563 2601 11575 2604
rect 11517 2595 11575 2601
rect 11790 2592 11796 2604
rect 11848 2592 11854 2644
rect 11882 2592 11888 2644
rect 11940 2632 11946 2644
rect 12069 2635 12127 2641
rect 12069 2632 12081 2635
rect 11940 2604 12081 2632
rect 11940 2592 11946 2604
rect 12069 2601 12081 2604
rect 12115 2601 12127 2635
rect 12986 2632 12992 2644
rect 12947 2604 12992 2632
rect 12069 2595 12127 2601
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 13357 2635 13415 2641
rect 13357 2601 13369 2635
rect 13403 2632 13415 2635
rect 14366 2632 14372 2644
rect 13403 2604 14372 2632
rect 13403 2601 13415 2604
rect 13357 2595 13415 2601
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 15470 2632 15476 2644
rect 15431 2604 15476 2632
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 15841 2635 15899 2641
rect 15841 2601 15853 2635
rect 15887 2632 15899 2635
rect 17034 2632 17040 2644
rect 15887 2604 17040 2632
rect 15887 2601 15899 2604
rect 15841 2595 15899 2601
rect 17034 2592 17040 2604
rect 17092 2632 17098 2644
rect 17862 2632 17868 2644
rect 17092 2604 17868 2632
rect 17092 2592 17098 2604
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 20717 2635 20775 2641
rect 20717 2601 20729 2635
rect 20763 2601 20775 2635
rect 20717 2595 20775 2601
rect 9122 2524 9128 2576
rect 9180 2564 9186 2576
rect 13449 2567 13507 2573
rect 13449 2564 13461 2567
rect 9180 2536 13461 2564
rect 9180 2524 9186 2536
rect 13449 2533 13461 2536
rect 13495 2533 13507 2567
rect 13449 2527 13507 2533
rect 15286 2524 15292 2576
rect 15344 2564 15350 2576
rect 20732 2564 20760 2595
rect 15344 2536 20760 2564
rect 15344 2524 15350 2536
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 7653 2499 7711 2505
rect 7653 2496 7665 2499
rect 7524 2468 7665 2496
rect 7524 2456 7530 2468
rect 7653 2465 7665 2468
rect 7699 2465 7711 2499
rect 7653 2459 7711 2465
rect 8018 2456 8024 2508
rect 8076 2496 8082 2508
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 8076 2468 11437 2496
rect 8076 2456 8082 2468
rect 11425 2465 11437 2468
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 15654 2496 15660 2508
rect 11664 2468 15660 2496
rect 11664 2456 11670 2468
rect 15654 2456 15660 2468
rect 15712 2456 15718 2508
rect 15933 2499 15991 2505
rect 15933 2496 15945 2499
rect 15764 2468 15945 2496
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2397 7895 2431
rect 11698 2428 11704 2440
rect 11659 2400 11704 2428
rect 7837 2391 7895 2397
rect 7650 2320 7656 2372
rect 7708 2360 7714 2372
rect 7852 2360 7880 2391
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 13630 2428 13636 2440
rect 13591 2400 13636 2428
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 15764 2428 15792 2468
rect 15933 2465 15945 2468
rect 15979 2496 15991 2499
rect 17405 2499 17463 2505
rect 15979 2468 16620 2496
rect 15979 2465 15991 2468
rect 15933 2459 15991 2465
rect 16022 2428 16028 2440
rect 14936 2400 15792 2428
rect 15983 2400 16028 2428
rect 7708 2332 7880 2360
rect 7708 2320 7714 2332
rect 12342 2320 12348 2372
rect 12400 2360 12406 2372
rect 14936 2360 14964 2400
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 16592 2428 16620 2468
rect 17405 2465 17417 2499
rect 17451 2496 17463 2499
rect 17494 2496 17500 2508
rect 17451 2468 17500 2496
rect 17451 2465 17463 2468
rect 17405 2459 17463 2465
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 18690 2496 18696 2508
rect 18651 2468 18696 2496
rect 18690 2456 18696 2468
rect 18748 2456 18754 2508
rect 19242 2456 19248 2508
rect 19300 2496 19306 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 19300 2468 19441 2496
rect 19300 2456 19306 2468
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19429 2459 19487 2465
rect 19981 2499 20039 2505
rect 19981 2465 19993 2499
rect 20027 2465 20039 2499
rect 19981 2459 20039 2465
rect 19150 2428 19156 2440
rect 16592 2400 19156 2428
rect 19150 2388 19156 2400
rect 19208 2388 19214 2440
rect 19996 2428 20024 2459
rect 20438 2456 20444 2508
rect 20496 2496 20502 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20496 2468 20545 2496
rect 20496 2456 20502 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 20990 2428 20996 2440
rect 19996 2400 20996 2428
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 12400 2332 14964 2360
rect 12400 2320 12406 2332
rect 15838 2320 15844 2372
rect 15896 2360 15902 2372
rect 20165 2363 20223 2369
rect 20165 2360 20177 2363
rect 15896 2332 20177 2360
rect 15896 2320 15902 2332
rect 20165 2329 20177 2332
rect 20211 2329 20223 2363
rect 21358 2360 21364 2372
rect 20165 2323 20223 2329
rect 20640 2332 21364 2360
rect 16942 2252 16948 2304
rect 17000 2292 17006 2304
rect 17589 2295 17647 2301
rect 17589 2292 17601 2295
rect 17000 2264 17601 2292
rect 17000 2252 17006 2264
rect 17589 2261 17601 2264
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 18598 2252 18604 2304
rect 18656 2292 18662 2304
rect 18877 2295 18935 2301
rect 18877 2292 18889 2295
rect 18656 2264 18889 2292
rect 18656 2252 18662 2264
rect 18877 2261 18889 2264
rect 18923 2261 18935 2295
rect 18877 2255 18935 2261
rect 19613 2295 19671 2301
rect 19613 2261 19625 2295
rect 19659 2292 19671 2295
rect 20640 2292 20668 2332
rect 21358 2320 21364 2332
rect 21416 2320 21422 2372
rect 19659 2264 20668 2292
rect 19659 2261 19671 2264
rect 19613 2255 19671 2261
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 1946 1776 1952 1828
rect 2004 1816 2010 1828
rect 9214 1816 9220 1828
rect 2004 1788 9220 1816
rect 2004 1776 2010 1788
rect 9214 1776 9220 1788
rect 9272 1776 9278 1828
rect 10226 1640 10232 1692
rect 10284 1680 10290 1692
rect 16206 1680 16212 1692
rect 10284 1652 16212 1680
rect 10284 1640 10290 1652
rect 16206 1640 16212 1652
rect 16264 1640 16270 1692
rect 8570 960 8576 1012
rect 8628 1000 8634 1012
rect 9398 1000 9404 1012
rect 8628 972 9404 1000
rect 8628 960 8634 972
rect 9398 960 9404 972
rect 9456 960 9462 1012
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 20720 20043 20772 20052
rect 20720 20009 20729 20043
rect 20729 20009 20763 20043
rect 20763 20009 20772 20043
rect 20720 20000 20772 20009
rect 20536 19907 20588 19916
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 20168 19499 20220 19508
rect 20168 19465 20177 19499
rect 20177 19465 20211 19499
rect 20211 19465 20220 19499
rect 20168 19456 20220 19465
rect 20720 19499 20772 19508
rect 20720 19465 20729 19499
rect 20729 19465 20763 19499
rect 20763 19465 20772 19499
rect 20720 19456 20772 19465
rect 11704 19252 11756 19304
rect 19984 19295 20036 19304
rect 19984 19261 19993 19295
rect 19993 19261 20027 19295
rect 20027 19261 20036 19295
rect 19984 19252 20036 19261
rect 15200 19184 15252 19236
rect 17960 19116 18012 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 19984 18912 20036 18964
rect 20444 18955 20496 18964
rect 20444 18921 20453 18955
rect 20453 18921 20487 18955
rect 20487 18921 20496 18955
rect 20444 18912 20496 18921
rect 11704 18887 11756 18896
rect 11704 18853 11713 18887
rect 11713 18853 11747 18887
rect 11747 18853 11756 18887
rect 11704 18844 11756 18853
rect 17132 18844 17184 18896
rect 8208 18776 8260 18828
rect 8852 18776 8904 18828
rect 9680 18776 9732 18828
rect 10968 18776 11020 18828
rect 8024 18751 8076 18760
rect 8024 18717 8033 18751
rect 8033 18717 8067 18751
rect 8067 18717 8076 18751
rect 8024 18708 8076 18717
rect 5724 18572 5776 18624
rect 12532 18572 12584 18624
rect 12716 18776 12768 18828
rect 16948 18708 17000 18760
rect 20536 18640 20588 18692
rect 18512 18615 18564 18624
rect 18512 18581 18521 18615
rect 18521 18581 18555 18615
rect 18555 18581 18564 18615
rect 18512 18572 18564 18581
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 8024 18368 8076 18420
rect 15200 18368 15252 18420
rect 17960 18368 18012 18420
rect 20720 18343 20772 18352
rect 20720 18309 20729 18343
rect 20729 18309 20763 18343
rect 20763 18309 20772 18343
rect 20720 18300 20772 18309
rect 12716 18275 12768 18284
rect 12716 18241 12725 18275
rect 12725 18241 12759 18275
rect 12759 18241 12768 18275
rect 12716 18232 12768 18241
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 15108 18207 15160 18216
rect 15108 18173 15117 18207
rect 15117 18173 15151 18207
rect 15151 18173 15160 18207
rect 15108 18164 15160 18173
rect 20076 18164 20128 18216
rect 12532 18096 12584 18148
rect 12716 18096 12768 18148
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 20444 17867 20496 17876
rect 20444 17833 20453 17867
rect 20453 17833 20487 17867
rect 20487 17833 20496 17867
rect 20444 17824 20496 17833
rect 15108 17756 15160 17808
rect 14280 17731 14332 17740
rect 14280 17697 14289 17731
rect 14289 17697 14323 17731
rect 14323 17697 14332 17731
rect 14280 17688 14332 17697
rect 19984 17688 20036 17740
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 20076 17144 20128 17196
rect 19524 17076 19576 17128
rect 16764 17008 16816 17060
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 19984 16711 20036 16720
rect 19984 16677 19993 16711
rect 19993 16677 20027 16711
rect 20027 16677 20036 16711
rect 19984 16668 20036 16677
rect 19432 16600 19484 16652
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 16764 16056 16816 16108
rect 12532 15988 12584 16040
rect 19984 16031 20036 16040
rect 19984 15997 19993 16031
rect 19993 15997 20027 16031
rect 20027 15997 20036 16031
rect 19984 15988 20036 15997
rect 20076 15988 20128 16040
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 10048 15512 10100 15564
rect 19340 15512 19392 15564
rect 19984 15444 20036 15496
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 20168 15147 20220 15156
rect 20168 15113 20177 15147
rect 20177 15113 20211 15147
rect 20211 15113 20220 15147
rect 20168 15104 20220 15113
rect 20720 15079 20772 15088
rect 20720 15045 20729 15079
rect 20729 15045 20763 15079
rect 20763 15045 20772 15079
rect 20720 15036 20772 15045
rect 9772 14900 9824 14952
rect 16212 14900 16264 14952
rect 20352 14900 20404 14952
rect 20076 14832 20128 14884
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 20444 14603 20496 14612
rect 20444 14569 20453 14603
rect 20453 14569 20487 14603
rect 20487 14569 20496 14603
rect 20444 14560 20496 14569
rect 19340 14492 19392 14544
rect 7380 14424 7432 14476
rect 10876 14424 10928 14476
rect 19984 14424 20036 14476
rect 16212 14288 16264 14340
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 20628 13948 20680 14000
rect 20352 13880 20404 13932
rect 13360 13812 13412 13864
rect 19800 13812 19852 13864
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 19340 13515 19392 13524
rect 19340 13481 19349 13515
rect 19349 13481 19383 13515
rect 19383 13481 19392 13515
rect 19340 13472 19392 13481
rect 19984 13447 20036 13456
rect 19984 13413 19993 13447
rect 19993 13413 20027 13447
rect 20027 13413 20036 13447
rect 19984 13404 20036 13413
rect 19156 13379 19208 13388
rect 19156 13345 19165 13379
rect 19165 13345 19199 13379
rect 19199 13345 19208 13379
rect 19156 13336 19208 13345
rect 13268 13268 13320 13320
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 20720 12971 20772 12980
rect 20720 12937 20729 12971
rect 20729 12937 20763 12971
rect 20763 12937 20772 12971
rect 20720 12928 20772 12937
rect 16488 12792 16540 12844
rect 19156 12792 19208 12844
rect 17408 12724 17460 12776
rect 20536 12767 20588 12776
rect 20536 12733 20545 12767
rect 20545 12733 20579 12767
rect 20579 12733 20588 12767
rect 20536 12724 20588 12733
rect 16120 12631 16172 12640
rect 16120 12597 16129 12631
rect 16129 12597 16163 12631
rect 16163 12597 16172 12631
rect 16120 12588 16172 12597
rect 16396 12588 16448 12640
rect 17868 12588 17920 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 16120 12384 16172 12436
rect 19800 12316 19852 12368
rect 20536 12316 20588 12368
rect 15016 12248 15068 12300
rect 16856 12291 16908 12300
rect 16856 12257 16890 12291
rect 16890 12257 16908 12291
rect 16856 12248 16908 12257
rect 18604 12291 18656 12300
rect 18604 12257 18613 12291
rect 18613 12257 18647 12291
rect 18647 12257 18656 12291
rect 18604 12248 18656 12257
rect 18880 12248 18932 12300
rect 19248 12248 19300 12300
rect 11980 12044 12032 12096
rect 16948 12044 17000 12096
rect 17960 12087 18012 12096
rect 17960 12053 17969 12087
rect 17969 12053 18003 12087
rect 18003 12053 18012 12087
rect 17960 12044 18012 12053
rect 22468 12044 22520 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 16856 11883 16908 11892
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 21088 11840 21140 11892
rect 13636 11747 13688 11756
rect 13636 11713 13645 11747
rect 13645 11713 13679 11747
rect 13679 11713 13688 11747
rect 13636 11704 13688 11713
rect 15016 11747 15068 11756
rect 15016 11713 15025 11747
rect 15025 11713 15059 11747
rect 15059 11713 15068 11747
rect 15016 11704 15068 11713
rect 16948 11704 17000 11756
rect 17868 11704 17920 11756
rect 15292 11568 15344 11620
rect 16488 11636 16540 11688
rect 18788 11636 18840 11688
rect 20168 11636 20220 11688
rect 17960 11568 18012 11620
rect 20720 11568 20772 11620
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 13176 11500 13228 11552
rect 13544 11543 13596 11552
rect 13544 11509 13553 11543
rect 13553 11509 13587 11543
rect 13587 11509 13596 11543
rect 13544 11500 13596 11509
rect 18052 11500 18104 11552
rect 18512 11500 18564 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 12992 11296 13044 11348
rect 16304 11296 16356 11348
rect 16488 11296 16540 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 12716 11271 12768 11280
rect 12716 11237 12725 11271
rect 12725 11237 12759 11271
rect 12759 11237 12768 11271
rect 12716 11228 12768 11237
rect 13084 11228 13136 11280
rect 20168 11271 20220 11280
rect 11980 11203 12032 11212
rect 11980 11169 11989 11203
rect 11989 11169 12023 11203
rect 12023 11169 12032 11203
rect 11980 11160 12032 11169
rect 15016 11160 15068 11212
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 16396 11160 16448 11212
rect 17592 11203 17644 11212
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 12808 11092 12860 11144
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 14924 11067 14976 11076
rect 14924 11033 14933 11067
rect 14933 11033 14967 11067
rect 14967 11033 14976 11067
rect 18052 11160 18104 11212
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 19248 11160 19300 11212
rect 20168 11237 20177 11271
rect 20177 11237 20211 11271
rect 20211 11237 20220 11271
rect 20168 11228 20220 11237
rect 17960 11092 18012 11144
rect 14924 11024 14976 11033
rect 16304 11024 16356 11076
rect 16856 10956 16908 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 10968 10795 11020 10804
rect 10968 10761 10977 10795
rect 10977 10761 11011 10795
rect 11011 10761 11020 10795
rect 10968 10752 11020 10761
rect 16396 10795 16448 10804
rect 16396 10761 16405 10795
rect 16405 10761 16439 10795
rect 16439 10761 16448 10795
rect 16396 10752 16448 10761
rect 18788 10752 18840 10804
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 20904 10795 20956 10804
rect 19432 10752 19484 10761
rect 11612 10659 11664 10668
rect 11612 10625 11621 10659
rect 11621 10625 11655 10659
rect 11655 10625 11664 10659
rect 11612 10616 11664 10625
rect 13176 10616 13228 10668
rect 14924 10616 14976 10668
rect 17868 10616 17920 10668
rect 20904 10761 20913 10795
rect 20913 10761 20947 10795
rect 20947 10761 20956 10795
rect 20904 10752 20956 10761
rect 13452 10548 13504 10600
rect 15108 10548 15160 10600
rect 16120 10548 16172 10600
rect 18604 10548 18656 10600
rect 20352 10548 20404 10600
rect 20720 10591 20772 10600
rect 20720 10557 20729 10591
rect 20729 10557 20763 10591
rect 20763 10557 20772 10591
rect 20720 10548 20772 10557
rect 13636 10523 13688 10532
rect 13636 10489 13670 10523
rect 13670 10489 13688 10523
rect 13636 10480 13688 10489
rect 10784 10412 10836 10464
rect 11796 10412 11848 10464
rect 15844 10480 15896 10532
rect 15936 10480 15988 10532
rect 18512 10480 18564 10532
rect 17040 10455 17092 10464
rect 17040 10421 17049 10455
rect 17049 10421 17083 10455
rect 17083 10421 17092 10455
rect 17040 10412 17092 10421
rect 19708 10455 19760 10464
rect 19708 10421 19717 10455
rect 19717 10421 19751 10455
rect 19751 10421 19760 10455
rect 19708 10412 19760 10421
rect 20168 10455 20220 10464
rect 20168 10421 20177 10455
rect 20177 10421 20211 10455
rect 20211 10421 20220 10455
rect 20168 10412 20220 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 10784 10251 10836 10260
rect 10784 10217 10793 10251
rect 10793 10217 10827 10251
rect 10827 10217 10836 10251
rect 10784 10208 10836 10217
rect 11612 10140 11664 10192
rect 13636 10208 13688 10260
rect 15936 10208 15988 10260
rect 17040 10208 17092 10260
rect 17592 10208 17644 10260
rect 13268 10140 13320 10192
rect 17132 10140 17184 10192
rect 19432 10140 19484 10192
rect 13452 10072 13504 10124
rect 14372 10072 14424 10124
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 17868 10072 17920 10124
rect 18788 10115 18840 10124
rect 18788 10081 18797 10115
rect 18797 10081 18831 10115
rect 18831 10081 18840 10115
rect 18788 10072 18840 10081
rect 10232 10004 10284 10056
rect 15844 10047 15896 10056
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 16764 10004 16816 10056
rect 18512 10004 18564 10056
rect 15016 9868 15068 9920
rect 20168 9911 20220 9920
rect 20168 9877 20177 9911
rect 20177 9877 20211 9911
rect 20211 9877 20220 9911
rect 20168 9868 20220 9877
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 11612 9707 11664 9716
rect 11612 9673 11621 9707
rect 11621 9673 11655 9707
rect 11655 9673 11664 9707
rect 11612 9664 11664 9673
rect 11704 9664 11756 9716
rect 12440 9664 12492 9716
rect 18696 9664 18748 9716
rect 18972 9664 19024 9716
rect 13544 9596 13596 9648
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 9680 9460 9732 9512
rect 9864 9460 9916 9512
rect 10232 9503 10284 9512
rect 10232 9469 10241 9503
rect 10241 9469 10275 9503
rect 10275 9469 10284 9503
rect 10232 9460 10284 9469
rect 7564 9392 7616 9444
rect 11060 9392 11112 9444
rect 18788 9571 18840 9580
rect 18788 9537 18797 9571
rect 18797 9537 18831 9571
rect 18831 9537 18840 9571
rect 18788 9528 18840 9537
rect 18604 9460 18656 9512
rect 19340 9460 19392 9512
rect 20168 9460 20220 9512
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 19524 9392 19576 9444
rect 8944 9324 8996 9376
rect 9772 9324 9824 9376
rect 10140 9324 10192 9376
rect 13820 9324 13872 9376
rect 16672 9324 16724 9376
rect 17960 9324 18012 9376
rect 19064 9324 19116 9376
rect 19248 9324 19300 9376
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 20904 9324 20956 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 8944 9163 8996 9172
rect 8944 9129 8953 9163
rect 8953 9129 8987 9163
rect 8987 9129 8996 9163
rect 8944 9120 8996 9129
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 18512 9163 18564 9172
rect 9864 9052 9916 9104
rect 10232 9052 10284 9104
rect 18512 9129 18521 9163
rect 18521 9129 18555 9163
rect 18555 9129 18564 9163
rect 18512 9120 18564 9129
rect 19708 9120 19760 9172
rect 19524 9052 19576 9104
rect 848 8984 900 9036
rect 7564 8984 7616 9036
rect 9956 9027 10008 9036
rect 9956 8993 9990 9027
rect 9990 8993 10008 9027
rect 9956 8984 10008 8993
rect 14372 8984 14424 9036
rect 14556 9027 14608 9036
rect 14556 8993 14565 9027
rect 14565 8993 14599 9027
rect 14599 8993 14608 9027
rect 14556 8984 14608 8993
rect 15108 8984 15160 9036
rect 16396 8984 16448 9036
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 13912 8916 13964 8968
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 17316 8916 17368 8968
rect 8576 8848 8628 8900
rect 20168 8984 20220 9036
rect 2964 8780 3016 8832
rect 11612 8780 11664 8832
rect 16856 8780 16908 8832
rect 17040 8823 17092 8832
rect 17040 8789 17049 8823
rect 17049 8789 17083 8823
rect 17083 8789 17092 8823
rect 17040 8780 17092 8789
rect 19064 8916 19116 8968
rect 19340 8780 19392 8832
rect 19800 8780 19852 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 1400 8576 1452 8628
rect 11796 8576 11848 8628
rect 14740 8619 14792 8628
rect 14740 8585 14749 8619
rect 14749 8585 14783 8619
rect 14783 8585 14792 8619
rect 14740 8576 14792 8585
rect 16396 8619 16448 8628
rect 8576 8483 8628 8492
rect 8576 8449 8585 8483
rect 8585 8449 8619 8483
rect 8619 8449 8628 8483
rect 8576 8440 8628 8449
rect 4712 8372 4764 8424
rect 11060 8440 11112 8492
rect 9588 8304 9640 8356
rect 13268 8372 13320 8424
rect 14740 8440 14792 8492
rect 16396 8585 16405 8619
rect 16405 8585 16439 8619
rect 16439 8585 16448 8619
rect 16396 8576 16448 8585
rect 16672 8619 16724 8628
rect 16672 8585 16681 8619
rect 16681 8585 16715 8619
rect 16715 8585 16724 8619
rect 16672 8576 16724 8585
rect 16856 8508 16908 8560
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 20168 8440 20220 8492
rect 20352 8415 20404 8424
rect 14004 8304 14056 8356
rect 9956 8279 10008 8288
rect 9956 8245 9965 8279
rect 9965 8245 9999 8279
rect 9999 8245 10008 8279
rect 9956 8236 10008 8245
rect 11796 8236 11848 8288
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 20352 8381 20361 8415
rect 20361 8381 20395 8415
rect 20395 8381 20404 8415
rect 20352 8372 20404 8381
rect 17132 8347 17184 8356
rect 17132 8313 17141 8347
rect 17141 8313 17175 8347
rect 17175 8313 17184 8347
rect 20444 8347 20496 8356
rect 17132 8304 17184 8313
rect 20444 8313 20453 8347
rect 20453 8313 20487 8347
rect 20487 8313 20496 8347
rect 20444 8304 20496 8313
rect 12440 8236 12492 8245
rect 15476 8236 15528 8288
rect 18420 8236 18472 8288
rect 19340 8279 19392 8288
rect 19340 8245 19349 8279
rect 19349 8245 19383 8279
rect 19383 8245 19392 8279
rect 19340 8236 19392 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 11612 8032 11664 8084
rect 14004 8075 14056 8084
rect 14004 8041 14013 8075
rect 14013 8041 14047 8075
rect 14047 8041 14056 8075
rect 14004 8032 14056 8041
rect 14556 8032 14608 8084
rect 15476 8075 15528 8084
rect 15476 8041 15485 8075
rect 15485 8041 15519 8075
rect 15519 8041 15528 8075
rect 15476 8032 15528 8041
rect 7288 7896 7340 7948
rect 8576 7964 8628 8016
rect 8668 7896 8720 7948
rect 11980 7964 12032 8016
rect 12624 7964 12676 8016
rect 11612 7896 11664 7948
rect 13268 7896 13320 7948
rect 15016 7896 15068 7948
rect 19340 8032 19392 8084
rect 17040 7964 17092 8016
rect 19248 7964 19300 8016
rect 16396 7896 16448 7948
rect 18420 7939 18472 7948
rect 18420 7905 18429 7939
rect 18429 7905 18463 7939
rect 18463 7905 18472 7939
rect 18420 7896 18472 7905
rect 10692 7760 10744 7812
rect 17868 7828 17920 7880
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 18972 7828 19024 7880
rect 14556 7760 14608 7812
rect 9588 7692 9640 7744
rect 9772 7692 9824 7744
rect 9956 7692 10008 7744
rect 12624 7692 12676 7744
rect 20352 7692 20404 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 8852 7488 8904 7540
rect 10232 7488 10284 7540
rect 13912 7488 13964 7540
rect 14280 7488 14332 7540
rect 6828 7352 6880 7404
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 12532 7420 12584 7472
rect 19616 7463 19668 7472
rect 19616 7429 19625 7463
rect 19625 7429 19659 7463
rect 19659 7429 19668 7463
rect 19616 7420 19668 7429
rect 9588 7352 9640 7404
rect 11612 7395 11664 7404
rect 11612 7361 11621 7395
rect 11621 7361 11655 7395
rect 11655 7361 11664 7395
rect 11612 7352 11664 7361
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 14280 7352 14332 7404
rect 17132 7395 17184 7404
rect 17132 7361 17141 7395
rect 17141 7361 17175 7395
rect 17175 7361 17184 7395
rect 17132 7352 17184 7361
rect 20352 7395 20404 7404
rect 20352 7361 20361 7395
rect 20361 7361 20395 7395
rect 20395 7361 20404 7395
rect 20352 7352 20404 7361
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 13820 7284 13872 7336
rect 15108 7284 15160 7336
rect 8392 7216 8444 7268
rect 8576 7216 8628 7268
rect 14004 7216 14056 7268
rect 18788 7284 18840 7336
rect 18972 7284 19024 7336
rect 18604 7216 18656 7268
rect 19064 7216 19116 7268
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 9864 7148 9916 7200
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 11796 7148 11848 7200
rect 12348 7148 12400 7200
rect 12900 7148 12952 7200
rect 14096 7148 14148 7200
rect 16672 7148 16724 7200
rect 16856 7191 16908 7200
rect 16856 7157 16865 7191
rect 16865 7157 16899 7191
rect 16899 7157 16908 7191
rect 16856 7148 16908 7157
rect 16948 7191 17000 7200
rect 16948 7157 16957 7191
rect 16957 7157 16991 7191
rect 16991 7157 17000 7191
rect 16948 7148 17000 7157
rect 19708 7148 19760 7200
rect 20260 7191 20312 7200
rect 20260 7157 20269 7191
rect 20269 7157 20303 7191
rect 20303 7157 20312 7191
rect 20260 7148 20312 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 11612 6944 11664 6996
rect 12440 6987 12492 6996
rect 12440 6953 12449 6987
rect 12449 6953 12483 6987
rect 12483 6953 12492 6987
rect 12440 6944 12492 6953
rect 16672 6944 16724 6996
rect 12532 6919 12584 6928
rect 12532 6885 12541 6919
rect 12541 6885 12575 6919
rect 12575 6885 12584 6919
rect 12532 6876 12584 6885
rect 9312 6808 9364 6860
rect 10600 6808 10652 6860
rect 11980 6851 12032 6860
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 12440 6808 12492 6860
rect 13268 6876 13320 6928
rect 14556 6876 14608 6928
rect 15752 6876 15804 6928
rect 16396 6876 16448 6928
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 13912 6740 13964 6792
rect 12716 6672 12768 6724
rect 10692 6604 10744 6656
rect 14280 6647 14332 6656
rect 14280 6613 14289 6647
rect 14289 6613 14323 6647
rect 14323 6613 14332 6647
rect 14280 6604 14332 6613
rect 16580 6808 16632 6860
rect 18604 6851 18656 6860
rect 18604 6817 18613 6851
rect 18613 6817 18647 6851
rect 18647 6817 18656 6851
rect 18604 6808 18656 6817
rect 19616 6808 19668 6860
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 17224 6740 17276 6792
rect 19892 6740 19944 6792
rect 17132 6715 17184 6724
rect 17132 6681 17141 6715
rect 17141 6681 17175 6715
rect 17175 6681 17184 6715
rect 17132 6672 17184 6681
rect 17408 6715 17460 6724
rect 17408 6681 17417 6715
rect 17417 6681 17451 6715
rect 17451 6681 17460 6715
rect 17408 6672 17460 6681
rect 16672 6604 16724 6656
rect 19800 6604 19852 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 10048 6400 10100 6452
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 14096 6332 14148 6384
rect 6828 6264 6880 6316
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 14556 6307 14608 6316
rect 14556 6273 14565 6307
rect 14565 6273 14599 6307
rect 14599 6273 14608 6307
rect 14556 6264 14608 6273
rect 15752 6400 15804 6452
rect 16856 6400 16908 6452
rect 16028 6332 16080 6384
rect 19156 6400 19208 6452
rect 20260 6443 20312 6452
rect 20260 6409 20269 6443
rect 20269 6409 20303 6443
rect 20303 6409 20312 6443
rect 20260 6400 20312 6409
rect 13912 6196 13964 6248
rect 17132 6196 17184 6248
rect 18788 6332 18840 6384
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 19708 6307 19760 6316
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 19800 6307 19852 6316
rect 19800 6273 19809 6307
rect 19809 6273 19843 6307
rect 19843 6273 19852 6307
rect 19800 6264 19852 6273
rect 17408 6196 17460 6248
rect 21088 6196 21140 6248
rect 7748 6128 7800 6180
rect 15476 6128 15528 6180
rect 20536 6128 20588 6180
rect 10324 6103 10376 6112
rect 10324 6069 10333 6103
rect 10333 6069 10367 6103
rect 10367 6069 10376 6103
rect 10324 6060 10376 6069
rect 12256 6060 12308 6112
rect 14372 6103 14424 6112
rect 14372 6069 14381 6103
rect 14381 6069 14415 6103
rect 14415 6069 14424 6103
rect 14372 6060 14424 6069
rect 14464 6103 14516 6112
rect 14464 6069 14473 6103
rect 14473 6069 14507 6103
rect 14507 6069 14516 6103
rect 14464 6060 14516 6069
rect 15108 6060 15160 6112
rect 16028 6060 16080 6112
rect 16212 6060 16264 6112
rect 17224 6060 17276 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 18236 6103 18288 6112
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 19156 6060 19208 6112
rect 19616 6103 19668 6112
rect 19616 6069 19625 6103
rect 19625 6069 19659 6103
rect 19659 6069 19668 6103
rect 19616 6060 19668 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 7748 5899 7800 5908
rect 7748 5865 7757 5899
rect 7757 5865 7791 5899
rect 7791 5865 7800 5899
rect 7748 5856 7800 5865
rect 8208 5856 8260 5908
rect 10508 5856 10560 5908
rect 6828 5788 6880 5840
rect 8208 5720 8260 5772
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 10784 5788 10836 5840
rect 15476 5856 15528 5908
rect 16580 5856 16632 5908
rect 16948 5899 17000 5908
rect 16948 5865 16957 5899
rect 16957 5865 16991 5899
rect 16991 5865 17000 5899
rect 16948 5856 17000 5865
rect 17224 5856 17276 5908
rect 17868 5856 17920 5908
rect 19616 5856 19668 5908
rect 14280 5788 14332 5840
rect 14464 5788 14516 5840
rect 10232 5720 10284 5772
rect 10692 5720 10744 5772
rect 12440 5720 12492 5772
rect 18236 5788 18288 5840
rect 16304 5695 16356 5704
rect 16304 5661 16313 5695
rect 16313 5661 16347 5695
rect 16347 5661 16356 5695
rect 16304 5652 16356 5661
rect 17132 5652 17184 5704
rect 19248 5720 19300 5772
rect 19892 5720 19944 5772
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 19524 5695 19576 5704
rect 17500 5652 17552 5661
rect 19524 5661 19533 5695
rect 19533 5661 19567 5695
rect 19567 5661 19576 5695
rect 19524 5652 19576 5661
rect 9956 5516 10008 5568
rect 10416 5516 10468 5568
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 16672 5584 16724 5636
rect 17408 5516 17460 5568
rect 19064 5516 19116 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 9404 5312 9456 5364
rect 10324 5312 10376 5364
rect 13360 5312 13412 5364
rect 16304 5312 16356 5364
rect 20076 5312 20128 5364
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 8392 5176 8444 5228
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 13820 5219 13872 5228
rect 13820 5185 13829 5219
rect 13829 5185 13863 5219
rect 13863 5185 13872 5219
rect 13820 5176 13872 5185
rect 14556 5176 14608 5228
rect 16672 5176 16724 5228
rect 17960 5176 18012 5228
rect 18604 5176 18656 5228
rect 6920 5108 6972 5160
rect 10416 5108 10468 5160
rect 14464 5108 14516 5160
rect 18420 5151 18472 5160
rect 18420 5117 18429 5151
rect 18429 5117 18463 5151
rect 18463 5117 18472 5151
rect 18420 5108 18472 5117
rect 19800 5108 19852 5160
rect 20628 5151 20680 5160
rect 20628 5117 20637 5151
rect 20637 5117 20671 5151
rect 20671 5117 20680 5151
rect 20628 5108 20680 5117
rect 8852 5015 8904 5024
rect 8852 4981 8861 5015
rect 8861 4981 8895 5015
rect 8895 4981 8904 5015
rect 8852 4972 8904 4981
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 12716 5040 12768 5092
rect 14372 5040 14424 5092
rect 19156 5040 19208 5092
rect 8944 4972 8996 4981
rect 12164 4972 12216 5024
rect 12440 5015 12492 5024
rect 12440 4981 12449 5015
rect 12449 4981 12483 5015
rect 12483 4981 12492 5015
rect 13636 5015 13688 5024
rect 12440 4972 12492 4981
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 15200 4972 15252 5024
rect 19800 4972 19852 5024
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 8484 4768 8536 4820
rect 10140 4768 10192 4820
rect 10232 4768 10284 4820
rect 11704 4768 11756 4820
rect 12440 4768 12492 4820
rect 13636 4768 13688 4820
rect 17500 4768 17552 4820
rect 18880 4768 18932 4820
rect 9680 4700 9732 4752
rect 10508 4700 10560 4752
rect 5264 4632 5316 4684
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 8208 4564 8260 4616
rect 9036 4607 9088 4616
rect 9036 4573 9045 4607
rect 9045 4573 9079 4607
rect 9079 4573 9088 4607
rect 9036 4564 9088 4573
rect 9772 4632 9824 4684
rect 12072 4675 12124 4684
rect 12072 4641 12081 4675
rect 12081 4641 12115 4675
rect 12115 4641 12124 4675
rect 12072 4632 12124 4641
rect 12532 4632 12584 4684
rect 13084 4675 13136 4684
rect 13084 4641 13093 4675
rect 13093 4641 13127 4675
rect 13127 4641 13136 4675
rect 13084 4632 13136 4641
rect 14648 4632 14700 4684
rect 18604 4675 18656 4684
rect 12164 4607 12216 4616
rect 12164 4573 12173 4607
rect 12173 4573 12207 4607
rect 12207 4573 12216 4607
rect 12164 4564 12216 4573
rect 16488 4607 16540 4616
rect 14648 4496 14700 4548
rect 16488 4573 16497 4607
rect 16497 4573 16531 4607
rect 16531 4573 16540 4607
rect 16488 4564 16540 4573
rect 18604 4641 18613 4675
rect 18613 4641 18647 4675
rect 18647 4641 18656 4675
rect 18604 4632 18656 4641
rect 19708 4632 19760 4684
rect 19892 4675 19944 4684
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 18788 4607 18840 4616
rect 18788 4573 18797 4607
rect 18797 4573 18831 4607
rect 18831 4573 18840 4607
rect 18788 4564 18840 4573
rect 19340 4564 19392 4616
rect 20168 4607 20220 4616
rect 20168 4573 20177 4607
rect 20177 4573 20211 4607
rect 20211 4573 20220 4607
rect 20168 4564 20220 4573
rect 20352 4564 20404 4616
rect 9956 4428 10008 4480
rect 10324 4428 10376 4480
rect 11612 4428 11664 4480
rect 13820 4428 13872 4480
rect 19524 4471 19576 4480
rect 19524 4437 19533 4471
rect 19533 4437 19567 4471
rect 19567 4437 19576 4471
rect 19524 4428 19576 4437
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 7472 4224 7524 4276
rect 7748 4224 7800 4276
rect 9772 4224 9824 4276
rect 14648 4267 14700 4276
rect 10968 4199 11020 4208
rect 6828 4088 6880 4140
rect 7656 4088 7708 4140
rect 8208 4088 8260 4140
rect 10968 4165 10977 4199
rect 10977 4165 11011 4199
rect 11011 4165 11020 4199
rect 10968 4156 11020 4165
rect 14648 4233 14657 4267
rect 14657 4233 14691 4267
rect 14691 4233 14700 4267
rect 14648 4224 14700 4233
rect 17224 4224 17276 4276
rect 19708 4267 19760 4276
rect 19708 4233 19717 4267
rect 19717 4233 19751 4267
rect 19751 4233 19760 4267
rect 19708 4224 19760 4233
rect 11520 4131 11572 4140
rect 5356 4020 5408 4072
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 12256 4088 12308 4140
rect 13084 4088 13136 4140
rect 16488 4088 16540 4140
rect 17868 4088 17920 4140
rect 18052 4131 18104 4140
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 18052 4088 18104 4097
rect 19524 4088 19576 4140
rect 20352 4131 20404 4140
rect 20352 4097 20361 4131
rect 20361 4097 20395 4131
rect 20395 4097 20404 4131
rect 20352 4088 20404 4097
rect 7564 3952 7616 4004
rect 9312 3952 9364 4004
rect 6368 3884 6420 3936
rect 6920 3884 6972 3936
rect 7380 3927 7432 3936
rect 7380 3893 7389 3927
rect 7389 3893 7423 3927
rect 7423 3893 7432 3927
rect 7380 3884 7432 3893
rect 8300 3884 8352 3936
rect 8944 3884 8996 3936
rect 11152 3952 11204 4004
rect 12808 4020 12860 4072
rect 15384 4020 15436 4072
rect 13820 3952 13872 4004
rect 15292 3952 15344 4004
rect 16212 4020 16264 4072
rect 17960 4020 18012 4072
rect 20720 4063 20772 4072
rect 16396 3952 16448 4004
rect 20720 4029 20729 4063
rect 20729 4029 20763 4063
rect 20763 4029 20772 4063
rect 20720 4020 20772 4029
rect 18328 3995 18380 4004
rect 18328 3961 18362 3995
rect 18362 3961 18380 3995
rect 18328 3952 18380 3961
rect 11888 3884 11940 3936
rect 11980 3884 12032 3936
rect 15936 3884 15988 3936
rect 20812 3952 20864 4004
rect 18788 3884 18840 3936
rect 19524 3884 19576 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 9312 3723 9364 3732
rect 9312 3689 9321 3723
rect 9321 3689 9355 3723
rect 9355 3689 9364 3723
rect 9312 3680 9364 3689
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 3056 3612 3108 3664
rect 5264 3612 5316 3664
rect 6828 3612 6880 3664
rect 8208 3655 8260 3664
rect 8208 3621 8242 3655
rect 8242 3621 8260 3655
rect 8208 3612 8260 3621
rect 11520 3680 11572 3732
rect 12072 3680 12124 3732
rect 13176 3723 13228 3732
rect 11612 3612 11664 3664
rect 13176 3689 13185 3723
rect 13185 3689 13219 3723
rect 13219 3689 13228 3723
rect 13176 3680 13228 3689
rect 15384 3680 15436 3732
rect 18604 3680 18656 3732
rect 9772 3544 9824 3596
rect 15200 3612 15252 3664
rect 7656 3476 7708 3528
rect 9220 3476 9272 3528
rect 9864 3476 9916 3528
rect 10324 3519 10376 3528
rect 10324 3485 10333 3519
rect 10333 3485 10367 3519
rect 10367 3485 10376 3519
rect 10324 3476 10376 3485
rect 12440 3587 12492 3596
rect 12440 3553 12449 3587
rect 12449 3553 12483 3587
rect 12483 3553 12492 3587
rect 12440 3544 12492 3553
rect 12992 3544 13044 3596
rect 15476 3544 15528 3596
rect 12716 3476 12768 3528
rect 13820 3519 13872 3528
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 13820 3476 13872 3485
rect 3608 3340 3660 3392
rect 7656 3383 7708 3392
rect 7656 3349 7665 3383
rect 7665 3349 7699 3383
rect 7699 3349 7708 3383
rect 7656 3340 7708 3349
rect 13636 3408 13688 3460
rect 15016 3476 15068 3528
rect 17776 3612 17828 3664
rect 19340 3680 19392 3732
rect 20352 3680 20404 3732
rect 15752 3587 15804 3596
rect 15752 3553 15761 3587
rect 15761 3553 15795 3587
rect 15795 3553 15804 3587
rect 15752 3544 15804 3553
rect 15936 3519 15988 3528
rect 15936 3485 15945 3519
rect 15945 3485 15979 3519
rect 15979 3485 15988 3519
rect 15936 3476 15988 3485
rect 16212 3476 16264 3528
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 20168 3544 20220 3596
rect 18328 3476 18380 3485
rect 16488 3408 16540 3460
rect 11704 3383 11756 3392
rect 11704 3349 11713 3383
rect 11713 3349 11747 3383
rect 11747 3349 11756 3383
rect 11704 3340 11756 3349
rect 18236 3408 18288 3460
rect 19892 3340 19944 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 5816 3136 5868 3188
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 9036 3136 9088 3188
rect 13084 3136 13136 3188
rect 8484 3068 8536 3120
rect 11612 3068 11664 3120
rect 13820 3136 13872 3188
rect 19524 3179 19576 3188
rect 16488 3111 16540 3120
rect 16488 3077 16497 3111
rect 16497 3077 16531 3111
rect 16531 3077 16540 3111
rect 16488 3068 16540 3077
rect 17960 3068 18012 3120
rect 19524 3145 19533 3179
rect 19533 3145 19567 3179
rect 19567 3145 19576 3179
rect 19524 3136 19576 3145
rect 20904 3068 20956 3120
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 8944 3000 8996 3052
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 10324 3000 10376 3052
rect 13728 3000 13780 3052
rect 4160 2932 4212 2984
rect 6920 2932 6972 2984
rect 7656 2932 7708 2984
rect 7840 2932 7892 2984
rect 2504 2864 2556 2916
rect 8852 2864 8904 2916
rect 6920 2796 6972 2848
rect 9404 2932 9456 2984
rect 10508 2932 10560 2984
rect 11704 2932 11756 2984
rect 12532 2932 12584 2984
rect 15200 2932 15252 2984
rect 15936 2932 15988 2984
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 17316 2975 17368 2984
rect 17316 2941 17325 2975
rect 17325 2941 17359 2975
rect 17359 2941 17368 2975
rect 17316 2932 17368 2941
rect 18512 2932 18564 2984
rect 18972 3000 19024 3052
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 13636 2864 13688 2916
rect 14188 2864 14240 2916
rect 12164 2796 12216 2848
rect 14372 2839 14424 2848
rect 14372 2805 14381 2839
rect 14381 2805 14415 2839
rect 14415 2805 14424 2839
rect 14372 2796 14424 2805
rect 17868 2864 17920 2916
rect 19984 2932 20036 2984
rect 20536 2975 20588 2984
rect 20536 2941 20545 2975
rect 20545 2941 20579 2975
rect 20579 2941 20588 2975
rect 20536 2932 20588 2941
rect 19156 2864 19208 2916
rect 17592 2796 17644 2848
rect 19984 2839 20036 2848
rect 19984 2805 19993 2839
rect 19993 2805 20027 2839
rect 20027 2805 20036 2839
rect 19984 2796 20036 2805
rect 21916 2796 21968 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 7564 2592 7616 2644
rect 7748 2635 7800 2644
rect 7748 2601 7757 2635
rect 7757 2601 7791 2635
rect 7791 2601 7800 2635
rect 7748 2592 7800 2601
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 11152 2592 11204 2644
rect 11796 2592 11848 2644
rect 11888 2592 11940 2644
rect 12992 2635 13044 2644
rect 12992 2601 13001 2635
rect 13001 2601 13035 2635
rect 13035 2601 13044 2635
rect 12992 2592 13044 2601
rect 14372 2592 14424 2644
rect 15476 2635 15528 2644
rect 15476 2601 15485 2635
rect 15485 2601 15519 2635
rect 15519 2601 15528 2635
rect 15476 2592 15528 2601
rect 17040 2592 17092 2644
rect 17868 2592 17920 2644
rect 9128 2524 9180 2576
rect 15292 2524 15344 2576
rect 7472 2456 7524 2508
rect 8024 2456 8076 2508
rect 11612 2456 11664 2508
rect 15660 2456 15712 2508
rect 11704 2431 11756 2440
rect 7656 2320 7708 2372
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 16028 2431 16080 2440
rect 12348 2320 12400 2372
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 17500 2456 17552 2508
rect 18696 2499 18748 2508
rect 18696 2465 18705 2499
rect 18705 2465 18739 2499
rect 18739 2465 18748 2499
rect 18696 2456 18748 2465
rect 19248 2456 19300 2508
rect 19156 2388 19208 2440
rect 20444 2456 20496 2508
rect 20996 2388 21048 2440
rect 15844 2320 15896 2372
rect 16948 2252 17000 2304
rect 18604 2252 18656 2304
rect 21364 2320 21416 2372
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 1952 1776 2004 1828
rect 9220 1776 9272 1828
rect 10232 1640 10284 1692
rect 16212 1640 16264 1692
rect 8576 960 8628 1012
rect 9404 960 9456 1012
<< metal2 >>
rect 5722 22320 5778 22800
rect 17130 22320 17186 22800
rect 19062 22536 19118 22545
rect 19062 22471 19118 22480
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 5736 18630 5764 22320
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 11716 18902 11744 19246
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 8036 18426 8064 18702
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 2962 11520 3018 11529
rect 2962 11455 3018 11464
rect 848 9036 900 9042
rect 848 8978 900 8984
rect 294 3496 350 3505
rect 294 3431 350 3440
rect 308 480 336 3431
rect 860 480 888 8978
rect 2976 8838 3004 11455
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1412 480 1440 8570
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 1952 1828 2004 1834
rect 1952 1770 2004 1776
rect 1964 480 1992 1770
rect 2516 480 2544 2858
rect 3068 480 3096 3606
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3620 480 3648 3334
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4172 480 4200 2926
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 480 4752 8366
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7300 7410 7328 7890
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 6840 6322 6868 7346
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6840 5846 6868 6258
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6840 5234 6868 5782
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5276 3670 5304 4626
rect 6840 4146 6868 5170
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5368 3346 5396 4014
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 5276 3318 5396 3346
rect 5276 480 5304 3318
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5828 480 5856 3130
rect 6380 480 6408 3878
rect 6840 3670 6868 4082
rect 6932 3942 6960 5102
rect 7392 3942 7420 14418
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7576 9042 7604 9386
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7760 5914 7788 6122
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8220 5914 8248 18770
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8588 8498 8616 8842
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8588 8022 8616 8434
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8680 7546 8708 7890
rect 8864 7546 8892 18770
rect 9692 9518 9720 18770
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9784 9382 9812 14894
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 8956 9178 8984 9318
rect 9770 9208 9826 9217
rect 8944 9172 8996 9178
rect 9770 9143 9826 9152
rect 8944 9114 8996 9120
rect 9680 8968 9732 8974
rect 9784 8956 9812 9143
rect 9876 9110 9904 9454
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9732 8928 9812 8956
rect 9680 8910 9732 8916
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9600 7750 9628 8298
rect 9784 7750 9812 8928
rect 9968 8294 9996 8978
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 9600 7410 9628 7686
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8404 6458 8432 7210
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8220 5370 8248 5714
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8220 4622 8248 5306
rect 8404 5234 8432 6394
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8496 4826 8524 5646
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7484 4282 7512 4558
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6840 3058 6868 3606
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6920 2984 6972 2990
rect 6918 2952 6920 2961
rect 6972 2952 6974 2961
rect 6918 2887 6974 2896
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6932 480 6960 2790
rect 7576 2650 7604 3946
rect 7668 3534 7696 4082
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7668 2990 7696 3334
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7484 480 7512 2450
rect 7668 2378 7696 2926
rect 7760 2650 7788 4218
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8220 3670 8248 4082
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8220 3194 8248 3606
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 7840 2984 7892 2990
rect 7838 2952 7840 2961
rect 7892 2952 7894 2961
rect 7838 2887 7894 2896
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8312 2650 8340 3878
rect 8588 3210 8616 7210
rect 9324 6866 9352 7278
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9416 5370 9444 7142
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8496 3182 8616 3210
rect 8496 3126 8524 3182
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 8864 2922 8892 4966
rect 8956 3942 8984 4966
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 3058 8984 3878
rect 9048 3194 9076 4558
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9324 3738 9352 3946
rect 9692 3738 9720 4694
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9784 4282 9812 4626
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 8036 480 8064 2450
rect 8576 1012 8628 1018
rect 8576 954 8628 960
rect 8588 480 8616 954
rect 9140 480 9168 2518
rect 9232 1834 9260 3470
rect 9324 3058 9352 3674
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9220 1828 9272 1834
rect 9220 1770 9272 1776
rect 9416 1018 9444 2926
rect 9784 2530 9812 3538
rect 9876 3534 9904 7142
rect 9968 5574 9996 7686
rect 10060 6458 10088 15506
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10888 10690 10916 14418
rect 10980 10810 11008 18770
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11992 11218 12020 12038
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10888 10662 11100 10690
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10796 10266 10824 10406
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10244 9518 10272 9998
rect 11072 9568 11100 10662
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11624 10198 11652 10610
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11624 9722 11652 10134
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 10980 9540 11100 9568
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9968 4486 9996 5510
rect 10152 4826 10180 9318
rect 10244 9217 10272 9454
rect 10230 9208 10286 9217
rect 10230 9143 10286 9152
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10244 7546 10272 9046
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10244 5234 10272 5714
rect 10336 5370 10364 6054
rect 10428 5574 10456 7142
rect 10600 6860 10652 6866
rect 10520 6820 10600 6848
rect 10520 6322 10548 6820
rect 10600 6802 10652 6808
rect 10704 6662 10732 7754
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10520 5914 10548 6258
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10704 5778 10732 6598
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10244 4826 10272 5170
rect 10428 5166 10456 5510
rect 10704 5234 10732 5714
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10336 3534 10364 4422
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10336 3058 10364 3470
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10520 2990 10548 4694
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 9692 2502 9812 2530
rect 9404 1012 9456 1018
rect 9404 954 9456 960
rect 9692 480 9720 2502
rect 10232 1692 10284 1698
rect 10232 1634 10284 1640
rect 10244 480 10272 1634
rect 10796 480 10824 5782
rect 10980 4214 11008 9540
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11072 9178 11100 9386
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11072 8498 11100 9114
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11624 8090 11652 8774
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11624 7410 11652 7890
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11624 7002 11652 7346
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11716 4826 11744 9658
rect 11808 8634 11836 10406
rect 12452 9722 12480 18158
rect 12544 18154 12572 18566
rect 12728 18290 12756 18770
rect 15212 18426 15240 19178
rect 17144 18902 17172 22320
rect 17958 21176 18014 21185
rect 17958 21111 18014 21120
rect 17972 19174 18000 21111
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17958 18864 18014 18873
rect 17958 18799 18014 18808
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 11808 7206 11836 8230
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11992 6866 12020 7958
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 10968 4208 11020 4214
rect 10968 4150 11020 4156
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 11164 2650 11192 3946
rect 11532 3738 11560 4082
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11532 3482 11560 3674
rect 11624 3670 11652 4422
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11794 3632 11850 3641
rect 11794 3567 11850 3576
rect 11532 3454 11652 3482
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11624 3126 11652 3454
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 11716 2990 11744 3334
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11624 1986 11652 2450
rect 11716 2446 11744 2926
rect 11808 2650 11836 3567
rect 11900 2650 11928 3878
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11348 1958 11652 1986
rect 11348 480 11376 1958
rect 11992 480 12020 3878
rect 12084 3738 12112 4626
rect 12176 4622 12204 4966
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12268 4298 12296 6054
rect 12176 4270 12296 4298
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12176 2854 12204 4270
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12268 4049 12296 4082
rect 12254 4040 12310 4049
rect 12254 3975 12310 3984
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 12360 2378 12388 7142
rect 12452 7002 12480 8230
rect 12544 8106 12572 15982
rect 12728 11286 12756 18090
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 15120 17814 15148 18158
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12544 8078 12756 8106
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12636 7750 12664 7958
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12544 6934 12572 7414
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12452 5778 12480 6802
rect 12636 6798 12664 7686
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12728 6730 12756 8078
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12452 5114 12480 5714
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12452 5086 12572 5114
rect 12728 5098 12756 5510
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12452 4826 12480 4966
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12544 4690 12572 5086
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12438 3632 12494 3641
rect 12438 3567 12440 3576
rect 12492 3567 12494 3576
rect 12440 3538 12492 3544
rect 12544 2990 12572 4626
rect 12728 3534 12756 5034
rect 12820 4078 12848 11086
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12808 4072 12860 4078
rect 12912 4049 12940 7142
rect 12808 4014 12860 4020
rect 12898 4040 12954 4049
rect 12898 3975 12954 3984
rect 13004 3754 13032 11290
rect 13096 11286 13124 11494
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13188 10674 13216 11494
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13280 10282 13308 13262
rect 13188 10254 13308 10282
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13096 4146 13124 4626
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12912 3726 13032 3754
rect 13188 3738 13216 10254
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13280 9586 13308 10134
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 7954 13308 8366
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13280 6934 13308 7890
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13372 5370 13400 13806
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 10130 13492 10542
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13556 9654 13584 11494
rect 13648 10538 13676 11698
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13648 10266 13676 10474
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13832 7342 13860 9318
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13924 7546 13952 8910
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 14016 8090 14044 8298
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14016 7410 14044 8026
rect 14292 7546 14320 17682
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 16776 16114 16804 17002
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 16224 14346 16252 14894
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 16132 12442 16160 12582
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15028 11762 15056 12242
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15304 11218 15332 11562
rect 16408 11506 16436 12582
rect 16500 11694 16528 12786
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16868 11898 16896 12242
rect 16960 12102 16988 18702
rect 17972 18426 18000 18799
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16960 11762 16988 12038
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16132 11478 16436 11506
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14384 10130 14412 11086
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14936 10674 14964 11018
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14384 9042 14412 10066
rect 15028 9926 15056 11154
rect 16132 10606 16160 11478
rect 16500 11354 16528 11630
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16316 11082 16344 11290
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16408 10810 16436 11154
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14568 8090 14596 8978
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14752 8634 14780 8910
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14752 8498 14780 8570
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 15028 7954 15056 9862
rect 15120 9042 15148 10542
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15488 8090 15516 8230
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13924 6254 13952 6734
rect 14016 6458 14044 7210
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14108 6390 14136 7142
rect 14292 6662 14320 7346
rect 14568 6934 14596 7754
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14556 6928 14608 6934
rect 14556 6870 14608 6876
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 14292 5846 14320 6598
rect 14568 6322 14596 6870
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 15120 6118 15148 7278
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 14280 5840 14332 5846
rect 14280 5782 14332 5788
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4826 13676 4966
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13832 4486 13860 5170
rect 14384 5098 14412 6054
rect 14476 5846 14504 6054
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 15488 5914 15516 6122
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14476 5166 14504 5782
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14568 4672 14596 5170
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14648 4684 14700 4690
rect 14568 4644 14648 4672
rect 14648 4626 14700 4632
rect 14660 4554 14688 4626
rect 14648 4548 14700 4554
rect 14648 4490 14700 4496
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 14660 4282 14688 4490
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13176 3732 13228 3738
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12912 2802 12940 3726
rect 13176 3674 13228 3680
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 12544 2774 12940 2802
rect 12348 2372 12400 2378
rect 12348 2314 12400 2320
rect 12544 480 12572 2774
rect 13004 2650 13032 3538
rect 13832 3534 13860 3946
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 15212 3670 15240 4966
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13096 480 13124 3130
rect 13648 2922 13676 3402
rect 13832 3194 13860 3470
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13636 2916 13688 2922
rect 13636 2858 13688 2864
rect 13648 2446 13676 2858
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13740 1986 13768 2994
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 13648 1958 13768 1986
rect 13648 480 13676 1958
rect 14200 480 14228 2858
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14384 2650 14412 2790
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 15028 1850 15056 3470
rect 15304 3074 15332 3946
rect 15396 3738 15424 4014
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15212 3046 15332 3074
rect 15212 2990 15240 3046
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15488 2650 15516 3538
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 14752 1822 15056 1850
rect 14752 480 14780 1822
rect 15304 480 15332 2518
rect 15672 2514 15700 10066
rect 15856 10062 15884 10474
rect 15948 10266 15976 10474
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15764 6798 15792 6870
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15764 6458 15792 6734
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16040 6118 16068 6326
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15750 3632 15806 3641
rect 15750 3567 15752 3576
rect 15804 3567 15806 3576
rect 15752 3538 15804 3544
rect 15948 3534 15976 3878
rect 15936 3528 15988 3534
rect 16132 3505 16160 10542
rect 16868 10130 16896 10950
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 17052 10266 17080 10406
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16408 8634 16436 8978
rect 16684 8634 16712 9318
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16408 6934 16436 7890
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16684 7002 16712 7142
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 4078 16252 6054
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16316 5370 16344 5646
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16408 4604 16436 6870
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16592 5914 16620 6802
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16684 5642 16712 6598
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16684 5234 16712 5578
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16488 4616 16540 4622
rect 16408 4576 16488 4604
rect 16488 4558 16540 4564
rect 16500 4146 16528 4558
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16212 3528 16264 3534
rect 15936 3470 15988 3476
rect 16118 3496 16174 3505
rect 15948 2990 15976 3470
rect 16212 3470 16264 3476
rect 16118 3431 16174 3440
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15948 2802 15976 2926
rect 15948 2774 16048 2802
rect 16020 2666 16048 2774
rect 16020 2638 16068 2666
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 16040 2446 16068 2638
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15844 2372 15896 2378
rect 15844 2314 15896 2320
rect 15856 480 15884 2314
rect 16224 1698 16252 3470
rect 16212 1692 16264 1698
rect 16212 1634 16264 1640
rect 16408 480 16436 3946
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16500 3126 16528 3402
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16776 2990 16804 9998
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 17052 8838 17080 9522
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16868 8566 16896 8774
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 17052 8022 17080 8774
rect 17144 8362 17172 10134
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17144 7562 17172 8298
rect 17052 7534 17172 7562
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16868 6458 16896 7142
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16960 5914 16988 7142
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 17052 2650 17080 7534
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17144 6730 17172 7346
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 17144 6254 17172 6666
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17144 5710 17172 6190
rect 17236 6118 17264 6734
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17236 4282 17264 5850
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17236 2825 17264 4218
rect 17328 2990 17356 8910
rect 17420 6730 17448 12718
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17880 12345 17908 12582
rect 17866 12336 17922 12345
rect 17866 12271 17922 12280
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17604 10266 17632 11154
rect 17880 10674 17908 11698
rect 17972 11626 18000 12038
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18524 11642 18552 18566
rect 18602 12744 18658 12753
rect 18602 12679 18658 12688
rect 18616 12306 18644 12679
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 18432 11614 18552 11642
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 17972 11150 18000 11562
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 11218 18092 11494
rect 18432 11257 18460 11614
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18418 11248 18474 11257
rect 18052 11212 18104 11218
rect 18418 11183 18474 11192
rect 18052 11154 18104 11160
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17880 10130 17908 10610
rect 18524 10538 18552 11494
rect 18694 11384 18750 11393
rect 18694 11319 18696 11328
rect 18748 11319 18750 11328
rect 18696 11290 18748 11296
rect 18694 11248 18750 11257
rect 18604 11212 18656 11218
rect 18694 11183 18750 11192
rect 18604 11154 18656 11160
rect 18616 10606 18644 11154
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18602 10024 18658 10033
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17590 8120 17646 8129
rect 17590 8055 17646 8064
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17420 6118 17448 6190
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17420 5574 17448 6054
rect 17512 5710 17540 6258
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17408 5568 17460 5574
rect 17408 5510 17460 5516
rect 17512 4826 17540 5646
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17604 4706 17632 8055
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 5914 17908 7822
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17972 5794 18000 9318
rect 18524 9178 18552 9998
rect 18602 9959 18658 9968
rect 18616 9518 18644 9959
rect 18708 9722 18736 11183
rect 18800 10810 18828 11630
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18800 9586 18828 10066
rect 18892 9602 18920 12242
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18883 9574 18920 9602
rect 18604 9512 18656 9518
rect 18883 9500 18911 9574
rect 18883 9472 18920 9500
rect 18604 9454 18656 9460
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18432 7954 18460 8230
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18510 7576 18566 7585
rect 18510 7511 18566 7520
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18248 5846 18276 6054
rect 17512 4678 17632 4706
rect 17788 5766 18000 5794
rect 18236 5840 18288 5846
rect 18236 5782 18288 5788
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17222 2816 17278 2825
rect 17222 2751 17278 2760
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 17512 2514 17540 4678
rect 17788 3670 17816 5766
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18418 5264 18474 5273
rect 17960 5228 18012 5234
rect 18418 5199 18474 5208
rect 17960 5170 18012 5176
rect 17972 4978 18000 5170
rect 18432 5166 18460 5199
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 17880 4950 18000 4978
rect 17880 4146 17908 4950
rect 17958 4856 18014 4865
rect 17958 4791 18014 4800
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17972 4078 18000 4791
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 18064 3448 18092 4082
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 18340 3534 18368 3946
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18236 3460 18288 3466
rect 18064 3420 18236 3448
rect 18236 3402 18288 3408
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 17592 2848 17644 2854
rect 17592 2790 17644 2796
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 16960 480 16988 2246
rect 17604 1442 17632 2790
rect 17880 2650 17908 2858
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 17512 1414 17632 1442
rect 17972 1442 18000 3062
rect 18524 2990 18552 7511
rect 18604 7268 18656 7274
rect 18604 7210 18656 7216
rect 18616 6866 18644 7210
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18616 5234 18644 6802
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18616 3738 18644 4626
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18708 2514 18736 7822
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18800 6390 18828 7278
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18892 4826 18920 9472
rect 18984 7886 19012 9658
rect 19076 9382 19104 22471
rect 20902 22128 20958 22137
rect 20902 22063 20958 22072
rect 20166 20632 20222 20641
rect 20166 20567 20222 20576
rect 20180 19514 20208 20567
rect 20718 20224 20774 20233
rect 20718 20159 20774 20168
rect 20732 20058 20760 20159
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 20442 19272 20498 19281
rect 19996 18970 20024 19246
rect 20442 19207 20498 19216
rect 20456 18970 20484 19207
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20548 18698 20576 19858
rect 20718 19816 20774 19825
rect 20718 19751 20774 19760
rect 20732 19514 20760 19751
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 20720 18352 20772 18358
rect 20718 18320 20720 18329
rect 20772 18320 20774 18329
rect 20718 18255 20774 18264
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19352 14550 19380 15506
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19338 14104 19394 14113
rect 19338 14039 19394 14048
rect 19352 13530 19380 14039
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19168 12850 19196 13330
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19260 11914 19288 12242
rect 19168 11886 19288 11914
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18984 7342 19012 7822
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 19076 7274 19104 8910
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 18970 7168 19026 7177
rect 18970 7103 19026 7112
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18800 3942 18828 4558
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18984 3058 19012 7103
rect 19168 6458 19196 11886
rect 19246 11792 19302 11801
rect 19246 11727 19302 11736
rect 19260 11218 19288 11727
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19444 10962 19472 16594
rect 19352 10934 19472 10962
rect 19352 10010 19380 10934
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19444 10198 19472 10746
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19352 9982 19472 10010
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19260 8022 19288 9318
rect 19352 8838 19380 9454
rect 19444 9092 19472 9982
rect 19536 9450 19564 17070
rect 19996 16726 20024 17682
rect 20088 17202 20116 18158
rect 20442 17912 20498 17921
rect 20442 17847 20444 17856
rect 20496 17847 20498 17856
rect 20444 17818 20496 17824
rect 20718 17368 20774 17377
rect 20718 17303 20720 17312
rect 20772 17303 20774 17312
rect 20720 17274 20772 17280
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20166 16960 20222 16969
rect 20166 16895 20222 16904
rect 19984 16720 20036 16726
rect 19984 16662 20036 16668
rect 20180 16250 20208 16895
rect 20718 16552 20774 16561
rect 20718 16487 20774 16496
rect 20732 16250 20760 16487
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 20442 16008 20498 16017
rect 19996 15502 20024 15982
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 20088 14890 20116 15982
rect 20442 15943 20498 15952
rect 20456 15706 20484 15943
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20166 15600 20222 15609
rect 20166 15535 20222 15544
rect 20180 15162 20208 15535
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20720 15088 20772 15094
rect 20718 15056 20720 15065
rect 20772 15056 20774 15065
rect 20718 14991 20774 15000
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19812 12374 19840 13806
rect 19996 13462 20024 14418
rect 20364 13938 20392 14894
rect 20442 14648 20498 14657
rect 20442 14583 20444 14592
rect 20496 14583 20498 14592
rect 20444 14554 20496 14560
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20640 13705 20668 13942
rect 20626 13696 20682 13705
rect 20626 13631 20682 13640
rect 19984 13456 20036 13462
rect 19984 13398 20036 13404
rect 20718 13288 20774 13297
rect 20718 13223 20774 13232
rect 20732 12986 20760 13223
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20548 12374 20576 12718
rect 19800 12368 19852 12374
rect 19800 12310 19852 12316
rect 20536 12368 20588 12374
rect 20536 12310 20588 12316
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20180 11286 20208 11630
rect 20720 11620 20772 11626
rect 20720 11562 20772 11568
rect 20168 11280 20220 11286
rect 20168 11222 20220 11228
rect 20534 10840 20590 10849
rect 20534 10775 20590 10784
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 19708 10464 19760 10470
rect 20168 10464 20220 10470
rect 19708 10406 19760 10412
rect 20166 10432 20168 10441
rect 20220 10432 20222 10441
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19720 9178 19748 10406
rect 20166 10367 20222 10376
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20180 9518 20208 9862
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19524 9104 19576 9110
rect 19444 9064 19524 9092
rect 19524 9046 19576 9052
rect 20180 9042 20208 9318
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19616 8492 19668 8498
rect 19812 8480 19840 8774
rect 20180 8498 20208 8978
rect 19668 8452 19840 8480
rect 20168 8492 20220 8498
rect 19616 8434 19668 8440
rect 20168 8434 20220 8440
rect 20364 8430 20392 10542
rect 20548 9518 20576 10775
rect 20732 10606 20760 11562
rect 20916 10810 20944 22063
rect 21086 21584 21142 21593
rect 21086 21519 21142 21528
rect 21100 11898 21128 21519
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20626 9480 20682 9489
rect 20626 9415 20682 9424
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19352 8090 19380 8230
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1414 18092 1442
rect 17512 480 17540 1414
rect 18064 480 18092 1414
rect 18616 480 18644 2246
rect 19076 1850 19104 5510
rect 19168 5098 19196 6054
rect 19260 5778 19288 7958
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 19616 7472 19668 7478
rect 19616 7414 19668 7420
rect 19628 6866 19656 7414
rect 20364 7410 20392 7686
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19628 6746 19656 6802
rect 19536 6718 19656 6746
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19536 5710 19564 6718
rect 19720 6322 19748 7142
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 19812 6322 19840 6598
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19628 5914 19656 6054
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19812 5166 19840 6258
rect 19904 5778 19932 6734
rect 20272 6458 20300 7142
rect 20456 6769 20484 8298
rect 20442 6760 20498 6769
rect 20442 6695 20498 6704
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20640 6338 20668 9415
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20718 8528 20774 8537
rect 20718 8463 20774 8472
rect 20456 6310 20668 6338
rect 20258 6216 20314 6225
rect 20258 6151 20314 6160
rect 20272 5778 20300 6151
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 19168 3505 19196 5034
rect 19800 5024 19852 5030
rect 19800 4966 19852 4972
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19246 4312 19302 4321
rect 19246 4247 19302 4256
rect 19154 3496 19210 3505
rect 19154 3431 19210 3440
rect 19156 2916 19208 2922
rect 19156 2858 19208 2864
rect 19168 2446 19196 2858
rect 19260 2514 19288 4247
rect 19352 3738 19380 4558
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19536 4146 19564 4422
rect 19720 4282 19748 4626
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19156 2440 19208 2446
rect 19352 2394 19380 3674
rect 19536 3194 19564 3878
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19812 2530 19840 4966
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19904 3398 19932 4626
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19156 2382 19208 2388
rect 19260 2366 19380 2394
rect 19720 2502 19840 2530
rect 19076 1822 19196 1850
rect 19168 480 19196 1822
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3054 0 3110 480
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4710 0 4766 480
rect 5262 0 5318 480
rect 5814 0 5870 480
rect 6366 0 6422 480
rect 6918 0 6974 480
rect 7470 0 7526 480
rect 8022 0 8078 480
rect 8574 0 8630 480
rect 9126 0 9182 480
rect 9678 0 9734 480
rect 10230 0 10286 480
rect 10782 0 10838 480
rect 11334 0 11390 480
rect 11978 0 12034 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14186 0 14242 480
rect 14738 0 14794 480
rect 15290 0 15346 480
rect 15842 0 15898 480
rect 16394 0 16450 480
rect 16946 0 17002 480
rect 17498 0 17554 480
rect 18050 0 18106 480
rect 18602 0 18658 480
rect 19154 0 19210 480
rect 19260 241 19288 2366
rect 19720 480 19748 2502
rect 19904 1057 19932 3334
rect 19984 2984 20036 2990
rect 19982 2952 19984 2961
rect 20036 2952 20038 2961
rect 19982 2887 20038 2896
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19996 2009 20024 2790
rect 20088 2530 20116 5306
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20364 4622 20392 4966
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20180 3602 20208 4558
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20364 3738 20392 4082
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 20180 3058 20208 3538
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20088 2502 20300 2530
rect 20456 2514 20484 6310
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20548 5012 20576 6122
rect 20626 5808 20682 5817
rect 20626 5743 20682 5752
rect 20640 5166 20668 5743
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20548 4984 20668 5012
rect 20534 3904 20590 3913
rect 20534 3839 20590 3848
rect 20548 2990 20576 3839
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20640 2553 20668 4984
rect 20732 4078 20760 8463
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20626 2544 20682 2553
rect 19982 2000 20038 2009
rect 19982 1935 20038 1944
rect 19890 1048 19946 1057
rect 19890 983 19946 992
rect 20272 480 20300 2502
rect 20444 2508 20496 2514
rect 20626 2479 20682 2488
rect 20444 2450 20496 2456
rect 20824 480 20852 3946
rect 20916 3126 20944 9318
rect 20994 9072 21050 9081
rect 20994 9007 21050 9016
rect 20904 3120 20956 3126
rect 20904 3062 20956 3068
rect 20902 2816 20958 2825
rect 20902 2751 20958 2760
rect 20916 649 20944 2751
rect 21008 2446 21036 9007
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 21100 1601 21128 6190
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 21086 1592 21142 1601
rect 21086 1527 21142 1536
rect 20902 640 20958 649
rect 20902 575 20958 584
rect 21376 480 21404 2314
rect 21928 480 21956 2790
rect 22480 480 22508 12038
rect 19246 232 19302 241
rect 19246 167 19302 176
rect 19706 0 19762 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
<< via2 >>
rect 19062 22480 19118 22536
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 2962 11464 3018 11520
rect 294 3440 350 3496
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 9770 9152 9826 9208
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 6918 2932 6920 2952
rect 6920 2932 6972 2952
rect 6972 2932 6974 2952
rect 6918 2896 6974 2932
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7838 2932 7840 2952
rect 7840 2932 7892 2952
rect 7892 2932 7894 2952
rect 7838 2896 7894 2932
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 10230 9152 10286 9208
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 17958 21120 18014 21176
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 17958 18808 18014 18864
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11794 3576 11850 3632
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12254 3984 12310 4040
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 12438 3596 12494 3632
rect 12438 3576 12440 3596
rect 12440 3576 12492 3596
rect 12492 3576 12494 3596
rect 12898 3984 12954 4040
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15750 3596 15806 3632
rect 15750 3576 15752 3596
rect 15752 3576 15804 3596
rect 15804 3576 15806 3596
rect 16118 3440 16174 3496
rect 17866 12280 17922 12336
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18602 12688 18658 12744
rect 18418 11192 18474 11248
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18694 11348 18750 11384
rect 18694 11328 18696 11348
rect 18696 11328 18748 11348
rect 18748 11328 18750 11348
rect 18694 11192 18750 11248
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 17590 8064 17646 8120
rect 18602 9968 18658 10024
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18510 7520 18566 7576
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 17222 2760 17278 2816
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18418 5208 18474 5264
rect 17958 4800 18014 4856
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 20902 22072 20958 22128
rect 20166 20576 20222 20632
rect 20718 20168 20774 20224
rect 20442 19216 20498 19272
rect 20718 19760 20774 19816
rect 20718 18300 20720 18320
rect 20720 18300 20772 18320
rect 20772 18300 20774 18320
rect 20718 18264 20774 18300
rect 19338 14048 19394 14104
rect 18970 7112 19026 7168
rect 19246 11736 19302 11792
rect 20442 17876 20498 17912
rect 20442 17856 20444 17876
rect 20444 17856 20496 17876
rect 20496 17856 20498 17876
rect 20718 17332 20774 17368
rect 20718 17312 20720 17332
rect 20720 17312 20772 17332
rect 20772 17312 20774 17332
rect 20166 16904 20222 16960
rect 20718 16496 20774 16552
rect 20442 15952 20498 16008
rect 20166 15544 20222 15600
rect 20718 15036 20720 15056
rect 20720 15036 20772 15056
rect 20772 15036 20774 15056
rect 20718 15000 20774 15036
rect 20442 14612 20498 14648
rect 20442 14592 20444 14612
rect 20444 14592 20496 14612
rect 20496 14592 20498 14612
rect 20626 13640 20682 13696
rect 20718 13232 20774 13288
rect 20534 10784 20590 10840
rect 20166 10412 20168 10432
rect 20168 10412 20220 10432
rect 20220 10412 20222 10432
rect 20166 10376 20222 10412
rect 21086 21528 21142 21584
rect 20626 9424 20682 9480
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 20442 6704 20498 6760
rect 20718 8472 20774 8528
rect 20258 6160 20314 6216
rect 19246 4256 19302 4312
rect 19154 3440 19210 3496
rect 19982 2932 19984 2952
rect 19984 2932 20036 2952
rect 20036 2932 20038 2952
rect 19982 2896 20038 2932
rect 20626 5752 20682 5808
rect 20534 3848 20590 3904
rect 19982 1944 20038 2000
rect 19890 992 19946 1048
rect 20626 2488 20682 2544
rect 20994 9016 21050 9072
rect 20902 2760 20958 2816
rect 21086 1536 21142 1592
rect 20902 584 20958 640
rect 19246 176 19302 232
<< metal3 >>
rect 19057 22538 19123 22541
rect 22320 22538 22800 22568
rect 19057 22536 22800 22538
rect 19057 22480 19062 22536
rect 19118 22480 22800 22536
rect 19057 22478 22800 22480
rect 19057 22475 19123 22478
rect 22320 22448 22800 22478
rect 20897 22130 20963 22133
rect 22320 22130 22800 22160
rect 20897 22128 22800 22130
rect 20897 22072 20902 22128
rect 20958 22072 22800 22128
rect 20897 22070 22800 22072
rect 20897 22067 20963 22070
rect 22320 22040 22800 22070
rect 21081 21586 21147 21589
rect 22320 21586 22800 21616
rect 21081 21584 22800 21586
rect 21081 21528 21086 21584
rect 21142 21528 22800 21584
rect 21081 21526 22800 21528
rect 21081 21523 21147 21526
rect 22320 21496 22800 21526
rect 17953 21178 18019 21181
rect 22320 21178 22800 21208
rect 17953 21176 22800 21178
rect 17953 21120 17958 21176
rect 18014 21120 22800 21176
rect 17953 21118 22800 21120
rect 17953 21115 18019 21118
rect 22320 21088 22800 21118
rect 20161 20634 20227 20637
rect 22320 20634 22800 20664
rect 20161 20632 22800 20634
rect 20161 20576 20166 20632
rect 20222 20576 22800 20632
rect 20161 20574 22800 20576
rect 20161 20571 20227 20574
rect 22320 20544 22800 20574
rect 20713 20226 20779 20229
rect 22320 20226 22800 20256
rect 20713 20224 22800 20226
rect 20713 20168 20718 20224
rect 20774 20168 22800 20224
rect 20713 20166 22800 20168
rect 20713 20163 20779 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 20713 19818 20779 19821
rect 22320 19818 22800 19848
rect 20713 19816 22800 19818
rect 20713 19760 20718 19816
rect 20774 19760 22800 19816
rect 20713 19758 22800 19760
rect 20713 19755 20779 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 20437 19274 20503 19277
rect 22320 19274 22800 19304
rect 20437 19272 22800 19274
rect 20437 19216 20442 19272
rect 20498 19216 22800 19272
rect 20437 19214 22800 19216
rect 20437 19211 20503 19214
rect 22320 19184 22800 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 17953 18866 18019 18869
rect 22320 18866 22800 18896
rect 17953 18864 22800 18866
rect 17953 18808 17958 18864
rect 18014 18808 22800 18864
rect 17953 18806 22800 18808
rect 17953 18803 18019 18806
rect 22320 18776 22800 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 20713 18322 20779 18325
rect 22320 18322 22800 18352
rect 20713 18320 22800 18322
rect 20713 18264 20718 18320
rect 20774 18264 22800 18320
rect 20713 18262 22800 18264
rect 20713 18259 20779 18262
rect 22320 18232 22800 18262
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 20437 17914 20503 17917
rect 22320 17914 22800 17944
rect 20437 17912 22800 17914
rect 20437 17856 20442 17912
rect 20498 17856 22800 17912
rect 20437 17854 22800 17856
rect 20437 17851 20503 17854
rect 22320 17824 22800 17854
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 20713 17370 20779 17373
rect 22320 17370 22800 17400
rect 20713 17368 22800 17370
rect 20713 17312 20718 17368
rect 20774 17312 22800 17368
rect 20713 17310 22800 17312
rect 20713 17307 20779 17310
rect 22320 17280 22800 17310
rect 20161 16962 20227 16965
rect 22320 16962 22800 16992
rect 20161 16960 22800 16962
rect 20161 16904 20166 16960
rect 20222 16904 22800 16960
rect 20161 16902 22800 16904
rect 20161 16899 20227 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22320 16872 22800 16902
rect 14672 16831 14992 16832
rect 20713 16554 20779 16557
rect 22320 16554 22800 16584
rect 20713 16552 22800 16554
rect 20713 16496 20718 16552
rect 20774 16496 22800 16552
rect 20713 16494 22800 16496
rect 20713 16491 20779 16494
rect 22320 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 20437 16010 20503 16013
rect 22320 16010 22800 16040
rect 20437 16008 22800 16010
rect 20437 15952 20442 16008
rect 20498 15952 22800 16008
rect 20437 15950 22800 15952
rect 20437 15947 20503 15950
rect 22320 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 20161 15602 20227 15605
rect 22320 15602 22800 15632
rect 20161 15600 22800 15602
rect 20161 15544 20166 15600
rect 20222 15544 22800 15600
rect 20161 15542 22800 15544
rect 20161 15539 20227 15542
rect 22320 15512 22800 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 20713 15058 20779 15061
rect 22320 15058 22800 15088
rect 20713 15056 22800 15058
rect 20713 15000 20718 15056
rect 20774 15000 22800 15056
rect 20713 14998 22800 15000
rect 20713 14995 20779 14998
rect 22320 14968 22800 14998
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 20437 14650 20503 14653
rect 22320 14650 22800 14680
rect 20437 14648 22800 14650
rect 20437 14592 20442 14648
rect 20498 14592 22800 14648
rect 20437 14590 22800 14592
rect 20437 14587 20503 14590
rect 22320 14560 22800 14590
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 19333 14106 19399 14109
rect 22320 14106 22800 14136
rect 19333 14104 22800 14106
rect 19333 14048 19338 14104
rect 19394 14048 22800 14104
rect 19333 14046 22800 14048
rect 19333 14043 19399 14046
rect 22320 14016 22800 14046
rect 20621 13698 20687 13701
rect 22320 13698 22800 13728
rect 20621 13696 22800 13698
rect 20621 13640 20626 13696
rect 20682 13640 22800 13696
rect 20621 13638 22800 13640
rect 20621 13635 20687 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22320 13608 22800 13638
rect 14672 13567 14992 13568
rect 20713 13290 20779 13293
rect 22320 13290 22800 13320
rect 20713 13288 22800 13290
rect 20713 13232 20718 13288
rect 20774 13232 22800 13288
rect 20713 13230 22800 13232
rect 20713 13227 20779 13230
rect 22320 13200 22800 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 18597 12746 18663 12749
rect 22320 12746 22800 12776
rect 18597 12744 22800 12746
rect 18597 12688 18602 12744
rect 18658 12688 22800 12744
rect 18597 12686 22800 12688
rect 18597 12683 18663 12686
rect 22320 12656 22800 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 17861 12338 17927 12341
rect 22320 12338 22800 12368
rect 17861 12336 22800 12338
rect 17861 12280 17866 12336
rect 17922 12280 22800 12336
rect 17861 12278 22800 12280
rect 17861 12275 17927 12278
rect 22320 12248 22800 12278
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 19241 11794 19307 11797
rect 22320 11794 22800 11824
rect 19241 11792 22800 11794
rect 19241 11736 19246 11792
rect 19302 11736 22800 11792
rect 19241 11734 22800 11736
rect 19241 11731 19307 11734
rect 22320 11704 22800 11734
rect 0 11522 480 11552
rect 2957 11522 3023 11525
rect 0 11520 3023 11522
rect 0 11464 2962 11520
rect 3018 11464 3023 11520
rect 0 11462 3023 11464
rect 0 11432 480 11462
rect 2957 11459 3023 11462
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 18689 11386 18755 11389
rect 22320 11386 22800 11416
rect 18689 11384 22800 11386
rect 18689 11328 18694 11384
rect 18750 11328 22800 11384
rect 18689 11326 22800 11328
rect 18689 11323 18755 11326
rect 22320 11296 22800 11326
rect 18413 11250 18479 11253
rect 18689 11250 18755 11253
rect 18413 11248 18755 11250
rect 18413 11192 18418 11248
rect 18474 11192 18694 11248
rect 18750 11192 18755 11248
rect 18413 11190 18755 11192
rect 18413 11187 18479 11190
rect 18689 11187 18755 11190
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 20529 10842 20595 10845
rect 22320 10842 22800 10872
rect 20529 10840 22800 10842
rect 20529 10784 20534 10840
rect 20590 10784 22800 10840
rect 20529 10782 22800 10784
rect 20529 10779 20595 10782
rect 22320 10752 22800 10782
rect 20161 10434 20227 10437
rect 22320 10434 22800 10464
rect 20161 10432 22800 10434
rect 20161 10376 20166 10432
rect 20222 10376 22800 10432
rect 20161 10374 22800 10376
rect 20161 10371 20227 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22320 10344 22800 10374
rect 14672 10303 14992 10304
rect 18597 10026 18663 10029
rect 22320 10026 22800 10056
rect 18597 10024 22800 10026
rect 18597 9968 18602 10024
rect 18658 9968 22800 10024
rect 18597 9966 22800 9968
rect 18597 9963 18663 9966
rect 22320 9936 22800 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 20621 9482 20687 9485
rect 22320 9482 22800 9512
rect 20621 9480 22800 9482
rect 20621 9424 20626 9480
rect 20682 9424 22800 9480
rect 20621 9422 22800 9424
rect 20621 9419 20687 9422
rect 22320 9392 22800 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 9765 9210 9831 9213
rect 10225 9210 10291 9213
rect 9765 9208 10291 9210
rect 9765 9152 9770 9208
rect 9826 9152 10230 9208
rect 10286 9152 10291 9208
rect 9765 9150 10291 9152
rect 9765 9147 9831 9150
rect 10225 9147 10291 9150
rect 20989 9074 21055 9077
rect 22320 9074 22800 9104
rect 20989 9072 22800 9074
rect 20989 9016 20994 9072
rect 21050 9016 22800 9072
rect 20989 9014 22800 9016
rect 20989 9011 21055 9014
rect 22320 8984 22800 9014
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 20713 8530 20779 8533
rect 22320 8530 22800 8560
rect 20713 8528 22800 8530
rect 20713 8472 20718 8528
rect 20774 8472 22800 8528
rect 20713 8470 22800 8472
rect 20713 8467 20779 8470
rect 22320 8440 22800 8470
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 17585 8122 17651 8125
rect 22320 8122 22800 8152
rect 17585 8120 22800 8122
rect 17585 8064 17590 8120
rect 17646 8064 22800 8120
rect 17585 8062 22800 8064
rect 17585 8059 17651 8062
rect 22320 8032 22800 8062
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 18505 7578 18571 7581
rect 22320 7578 22800 7608
rect 18505 7576 22800 7578
rect 18505 7520 18510 7576
rect 18566 7520 22800 7576
rect 18505 7518 22800 7520
rect 18505 7515 18571 7518
rect 22320 7488 22800 7518
rect 18965 7170 19031 7173
rect 22320 7170 22800 7200
rect 18965 7168 22800 7170
rect 18965 7112 18970 7168
rect 19026 7112 22800 7168
rect 18965 7110 22800 7112
rect 18965 7107 19031 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22320 7080 22800 7110
rect 14672 7039 14992 7040
rect 20437 6762 20503 6765
rect 22320 6762 22800 6792
rect 20437 6760 22800 6762
rect 20437 6704 20442 6760
rect 20498 6704 22800 6760
rect 20437 6702 22800 6704
rect 20437 6699 20503 6702
rect 22320 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 20253 6218 20319 6221
rect 22320 6218 22800 6248
rect 20253 6216 22800 6218
rect 20253 6160 20258 6216
rect 20314 6160 22800 6216
rect 20253 6158 22800 6160
rect 20253 6155 20319 6158
rect 22320 6128 22800 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 20621 5810 20687 5813
rect 22320 5810 22800 5840
rect 20621 5808 22800 5810
rect 20621 5752 20626 5808
rect 20682 5752 22800 5808
rect 20621 5750 22800 5752
rect 20621 5747 20687 5750
rect 22320 5720 22800 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 18413 5266 18479 5269
rect 22320 5266 22800 5296
rect 18413 5264 22800 5266
rect 18413 5208 18418 5264
rect 18474 5208 22800 5264
rect 18413 5206 22800 5208
rect 18413 5203 18479 5206
rect 22320 5176 22800 5206
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 17953 4858 18019 4861
rect 22320 4858 22800 4888
rect 17953 4856 22800 4858
rect 17953 4800 17958 4856
rect 18014 4800 22800 4856
rect 17953 4798 22800 4800
rect 17953 4795 18019 4798
rect 22320 4768 22800 4798
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 19241 4314 19307 4317
rect 22320 4314 22800 4344
rect 19241 4312 22800 4314
rect 19241 4256 19246 4312
rect 19302 4256 22800 4312
rect 19241 4254 22800 4256
rect 19241 4251 19307 4254
rect 22320 4224 22800 4254
rect 12249 4042 12315 4045
rect 12893 4042 12959 4045
rect 12249 4040 12959 4042
rect 12249 3984 12254 4040
rect 12310 3984 12898 4040
rect 12954 3984 12959 4040
rect 12249 3982 12959 3984
rect 12249 3979 12315 3982
rect 12893 3979 12959 3982
rect 20529 3906 20595 3909
rect 22320 3906 22800 3936
rect 20529 3904 22800 3906
rect 20529 3848 20534 3904
rect 20590 3848 22800 3904
rect 20529 3846 22800 3848
rect 20529 3843 20595 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22320 3816 22800 3846
rect 14672 3775 14992 3776
rect 11789 3634 11855 3637
rect 12433 3634 12499 3637
rect 15745 3634 15811 3637
rect 11789 3632 15811 3634
rect 11789 3576 11794 3632
rect 11850 3576 12438 3632
rect 12494 3576 15750 3632
rect 15806 3576 15811 3632
rect 11789 3574 15811 3576
rect 11789 3571 11855 3574
rect 12433 3571 12499 3574
rect 15745 3571 15811 3574
rect 289 3498 355 3501
rect 16113 3498 16179 3501
rect 289 3496 16179 3498
rect 289 3440 294 3496
rect 350 3440 16118 3496
rect 16174 3440 16179 3496
rect 289 3438 16179 3440
rect 289 3435 355 3438
rect 16113 3435 16179 3438
rect 19149 3498 19215 3501
rect 22320 3498 22800 3528
rect 19149 3496 22800 3498
rect 19149 3440 19154 3496
rect 19210 3440 22800 3496
rect 19149 3438 22800 3440
rect 19149 3435 19215 3438
rect 22320 3408 22800 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 6913 2954 6979 2957
rect 7833 2954 7899 2957
rect 6913 2952 7899 2954
rect 6913 2896 6918 2952
rect 6974 2896 7838 2952
rect 7894 2896 7899 2952
rect 6913 2894 7899 2896
rect 6913 2891 6979 2894
rect 7833 2891 7899 2894
rect 19977 2954 20043 2957
rect 22320 2954 22800 2984
rect 19977 2952 22800 2954
rect 19977 2896 19982 2952
rect 20038 2896 22800 2952
rect 19977 2894 22800 2896
rect 19977 2891 20043 2894
rect 22320 2864 22800 2894
rect 17217 2818 17283 2821
rect 20897 2818 20963 2821
rect 17217 2816 20963 2818
rect 17217 2760 17222 2816
rect 17278 2760 20902 2816
rect 20958 2760 20963 2816
rect 17217 2758 20963 2760
rect 17217 2755 17283 2758
rect 20897 2755 20963 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 20621 2546 20687 2549
rect 22320 2546 22800 2576
rect 20621 2544 22800 2546
rect 20621 2488 20626 2544
rect 20682 2488 22800 2544
rect 20621 2486 22800 2488
rect 20621 2483 20687 2486
rect 22320 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 19977 2002 20043 2005
rect 22320 2002 22800 2032
rect 19977 2000 22800 2002
rect 19977 1944 19982 2000
rect 20038 1944 22800 2000
rect 19977 1942 22800 1944
rect 19977 1939 20043 1942
rect 22320 1912 22800 1942
rect 21081 1594 21147 1597
rect 22320 1594 22800 1624
rect 21081 1592 22800 1594
rect 21081 1536 21086 1592
rect 21142 1536 22800 1592
rect 21081 1534 22800 1536
rect 21081 1531 21147 1534
rect 22320 1504 22800 1534
rect 19885 1050 19951 1053
rect 22320 1050 22800 1080
rect 19885 1048 22800 1050
rect 19885 992 19890 1048
rect 19946 992 22800 1048
rect 19885 990 22800 992
rect 19885 987 19951 990
rect 22320 960 22800 990
rect 20897 642 20963 645
rect 22320 642 22800 672
rect 20897 640 22800 642
rect 20897 584 20902 640
rect 20958 584 22800 640
rect 20897 582 22800 584
rect 20897 579 20963 582
rect 22320 552 22800 582
rect 19241 234 19307 237
rect 22320 234 22800 264
rect 19241 232 22800 234
rect 19241 176 19246 232
rect 19302 176 22800 232
rect 19241 174 22800 176
rect 19241 171 19307 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1605641404
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1605641404
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _41_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 8280 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7268 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8648 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1605641404
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_81
timestamp 1605641404
transform 1 0 8556 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1605641404
transform 1 0 8280 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10396 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_91
timestamp 1605641404
transform 1 0 9476 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_99
timestamp 1605641404
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106
timestamp 1605641404
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11040 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1605641404
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1605641404
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1605641404
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1605641404
transform 1 0 12052 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1605641404
transform 1 0 14352 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12696 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12972 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_0_138
timestamp 1605641404
transform 1 0 13800 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1605641404
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15088 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1605641404
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1605641404
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_165
timestamp 1605641404
transform 1 0 16284 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_147
timestamp 1605641404
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_151
timestamp 1605641404
transform 1 0 14996 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_168
timestamp 1605641404
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _85_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 16744 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_174
timestamp 1605641404
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1605641404
transform 1 0 17296 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_180
timestamp 1605641404
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1605641404
transform 1 0 17756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1605641404
transform 1 0 17388 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1605641404
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1605641404
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1605641404
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1605641404
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1605641404
transform 1 0 18676 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1605641404
transform 1 0 18584 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1605641404
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 19504 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_195
timestamp 1605641404
transform 1 0 19044 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1605641404
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1605641404
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_194
timestamp 1605641404
transform 1 0 18952 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1605641404
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1605641404
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1605641404
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1605641404
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1605641404
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1605641404
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1605641404
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1605641404
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1605641404
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1605641404
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6256 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1605641404
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7912 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_72
timestamp 1605641404
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10304 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1605641404
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1605641404
transform 1 0 9936 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11960 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1605641404
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_127
timestamp 1605641404
transform 1 0 12788 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1605641404
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1605641404
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_163
timestamp 1605641404
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 17664 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1605641404
transform 1 0 17204 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_179
timestamp 1605641404
transform 1 0 17572 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1605641404
transform 1 0 18676 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 19136 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_189
timestamp 1605641404
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1605641404
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1605641404
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1605641404
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1605641404
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1605641404
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1605641404
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1605641404
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1605641404
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1605641404
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_62
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8464 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7360 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_77
timestamp 1605641404
transform 1 0 8188 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_96
timestamp 1605641404
transform 1 0 9936 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_104
timestamp 1605641404
transform 1 0 10672 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10948 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_116
timestamp 1605641404
transform 1 0 11776 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13248 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1605641404
transform 1 0 12788 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_131
timestamp 1605641404
transform 1 0 13156 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15456 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_3_148
timestamp 1605641404
transform 1 0 14720 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1605641404
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1605641404
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_176
timestamp 1605641404
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1605641404
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19688 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1605641404
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1605641404
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1605641404
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1605641404
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1605641404
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1605641404
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_56
timestamp 1605641404
transform 1 0 6256 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6992 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_73
timestamp 1605641404
transform 1 0 7820 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1605641404
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11592 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp 1605641404
transform 1 0 11132 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_113
timestamp 1605641404
transform 1 0 11500 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_123
timestamp 1605641404
transform 1 0 12420 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13064 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_129
timestamp 1605641404
transform 1 0 12972 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1605641404
transform 1 0 14720 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_146
timestamp 1605641404
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1605641404
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1605641404
transform 1 0 16100 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16468 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 18216 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_183
timestamp 1605641404
transform 1 0 17940 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19504 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_195
timestamp 1605641404
transform 1 0 19044 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_199
timestamp 1605641404
transform 1 0 19412 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1605641404
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1605641404
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1605641404
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1605641404
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1605641404
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1605641404
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1605641404
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1605641404
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8464 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1605641404
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10672 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9568 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_89
timestamp 1605641404
transform 1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_101
timestamp 1605641404
transform 1 0 10396 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1605641404
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14260 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13248 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_126
timestamp 1605641404
transform 1 0 12696 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_141
timestamp 1605641404
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 15824 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_152
timestamp 1605641404
transform 1 0 15088 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1605641404
transform 1 0 16652 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1605641404
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1605641404
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1605641404
transform 1 0 18400 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18952 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_192
timestamp 1605641404
transform 1 0 18768 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1605641404
transform 1 0 20608 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1605641404
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_216
timestamp 1605641404
transform 1 0 20976 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1605641404
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1605641404
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1605641404
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1605641404
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6348 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1605641404
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_56
timestamp 1605641404
transform 1 0 6256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1605641404
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1605641404
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6992 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_73
timestamp 1605641404
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1605641404
transform 1 0 8464 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1605641404
transform 1 0 9016 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1605641404
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1605641404
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_92
timestamp 1605641404
transform 1 0 9568 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1605641404
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1605641404
transform 1 0 10856 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11316 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1605641404
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_109
timestamp 1605641404
transform 1 0 11132 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1605641404
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_123
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13984 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12972 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_127
timestamp 1605641404
transform 1 0 12788 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1605641404
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_138
timestamp 1605641404
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1605641404
transform 1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14996 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15824 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_158
timestamp 1605641404
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 1605641404
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_171
timestamp 1605641404
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_167
timestamp 1605641404
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_169
timestamp 1605641404
transform 1 0 16652 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16928 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16928 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1605641404
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1605641404
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 18216 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_181
timestamp 1605641404
transform 1 0 17756 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1605641404
transform 1 0 20240 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 20240 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 18952 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 19228 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_193
timestamp 1605641404
transform 1 0 18860 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_203
timestamp 1605641404
transform 1 0 19780 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_207
timestamp 1605641404
transform 1 0 20148 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp 1605641404
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_206
timestamp 1605641404
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1605641404
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1605641404
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1605641404
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp 1605641404
transform 1 0 21068 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1605641404
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1605641404
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1605641404
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1605641404
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1605641404
transform 1 0 8188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_68
timestamp 1605641404
transform 1 0 7360 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_76
timestamp 1605641404
transform 1 0 8096 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1605641404
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10028 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11776 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_113
timestamp 1605641404
transform 1 0 11500 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12880 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1605641404
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1605641404
transform 1 0 14536 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15732 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1605641404
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_158
timestamp 1605641404
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 17388 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_175
timestamp 1605641404
transform 1 0 17204 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1605641404
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1605641404
transform 1 0 20240 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 18584 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1605641404
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1605641404
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1605641404
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1605641404
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1605641404
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1605641404
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1605641404
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1605641404
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1605641404
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7268 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1605641404
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1605641404
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8924 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9936 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_94
timestamp 1605641404
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11040 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_105
timestamp 1605641404
transform 1 0 10764 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1605641404
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1605641404
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_123
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_131
timestamp 1605641404
transform 1 0 13156 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_143
timestamp 1605641404
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1605641404
transform 1 0 15272 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_166
timestamp 1605641404
transform 1 0 16376 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18216 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16468 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_176
timestamp 1605641404
transform 1 0 17296 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1605641404
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1605641404
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19872 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_202
timestamp 1605641404
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_213
timestamp 1605641404
transform 1 0 20700 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1605641404
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1605641404
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1605641404
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1605641404
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1605641404
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7912 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_10_68
timestamp 1605641404
transform 1 0 7360 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 10488 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1605641404
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_101
timestamp 1605641404
transform 1 0 10396 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10948 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12604 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_105
timestamp 1605641404
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_123
timestamp 1605641404
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1605641404
transform 1 0 14076 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1605641404
transform 1 0 14628 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16284 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1605641404
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_159
timestamp 1605641404
transform 1 0 15732 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_181
timestamp 1605641404
transform 1 0 17756 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_187
timestamp 1605641404
transform 1 0 18308 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1605641404
transform 1 0 19136 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 18400 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19780 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1605641404
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_199
timestamp 1605641404
transform 1 0 19412 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1605641404
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1605641404
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1605641404
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1605641404
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1605641404
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1605641404
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1605641404
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1605641404
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8556 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_11_74
timestamp 1605641404
transform 1 0 7912 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_80
timestamp 1605641404
transform 1 0 8464 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10672 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_97
timestamp 1605641404
transform 1 0 10028 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1605641404
transform 1 0 10580 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1605641404
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1605641404
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13340 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_11_126
timestamp 1605641404
transform 1 0 12696 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_132
timestamp 1605641404
transform 1 0 13248 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14996 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_149
timestamp 1605641404
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16652 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_167
timestamp 1605641404
transform 1 0 16468 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1605641404
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1605641404
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_184
timestamp 1605641404
transform 1 0 18032 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19964 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18952 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_192
timestamp 1605641404
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp 1605641404
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_214
timestamp 1605641404
transform 1 0 20792 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1605641404
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1605641404
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1605641404
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1605641404
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1605641404
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_80
timestamp 1605641404
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1605641404
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 11776 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_109
timestamp 1605641404
transform 1 0 11132 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_115
timestamp 1605641404
transform 1 0 11684 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_119
timestamp 1605641404
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_131
timestamp 1605641404
transform 1 0 13156 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_139
timestamp 1605641404
transform 1 0 13892 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15640 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1605641404
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18124 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17388 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_174
timestamp 1605641404
transform 1 0 17112 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1605641404
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 19136 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1605641404
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1605641404
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1605641404
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1605641404
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1605641404
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1605641404
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1605641404
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1605641404
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1605641404
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1605641404
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1605641404
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1605641404
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1605641404
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1605641404
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1605641404
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1605641404
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1605641404
transform 1 0 9568 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10212 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_86
timestamp 1605641404
transform 1 0 9016 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_95
timestamp 1605641404
transform 1 0 9844 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1605641404
transform 1 0 10764 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11224 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_115
timestamp 1605641404
transform 1 0 11684 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1605641404
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_123
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_108
timestamp 1605641404
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12880 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12696 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1605641404
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_126
timestamp 1605641404
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1605641404
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1605641404
transform 1 0 16284 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 14536 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1605641404
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_159
timestamp 1605641404
transform 1 0 15732 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1605641404
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1605641404
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_168
timestamp 1605641404
transform 1 0 16560 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_176
timestamp 1605641404
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16468 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16836 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_185
timestamp 1605641404
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_181
timestamp 1605641404
transform 1 0 17756 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_177
timestamp 1605641404
transform 1 0 17388 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1605641404
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1605641404
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1605641404
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1605641404
transform 1 0 18216 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1605641404
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1605641404
transform 1 0 17848 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1605641404
transform 1 0 18308 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18768 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18768 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_13_190
timestamp 1605641404
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_208
timestamp 1605641404
transform 1 0 20240 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1605641404
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_208
timestamp 1605641404
transform 1 0 20240 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1605641404
transform 1 0 20516 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1605641404
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1605641404
transform 1 0 20884 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1605641404
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1605641404
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1605641404
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1605641404
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1605641404
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1605641404
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1605641404
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1605641404
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1605641404
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1605641404
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_98
timestamp 1605641404
transform 1 0 10120 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10948 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1605641404
transform 1 0 10856 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_116
timestamp 1605641404
transform 1 0 11776 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1605641404
transform 1 0 12880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13340 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_127
timestamp 1605641404
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_131
timestamp 1605641404
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14996 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1605641404
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16652 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1605641404
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_167
timestamp 1605641404
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1605641404
transform 1 0 17480 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1605641404
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19688 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1605641404
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1605641404
transform 1 0 20700 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_211
timestamp 1605641404
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_217
timestamp 1605641404
transform 1 0 21068 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1605641404
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1605641404
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1605641404
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1605641404
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1605641404
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1605641404
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11960 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1605641404
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_117
timestamp 1605641404
transform 1 0 11868 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_124
timestamp 1605641404
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 12696 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp 1605641404
transform 1 0 14536 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18216 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 17204 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1605641404
transform 1 0 16744 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_174
timestamp 1605641404
transform 1 0 17112 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_184
timestamp 1605641404
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1605641404
transform 1 0 19320 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19872 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_195
timestamp 1605641404
transform 1 0 19044 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_202
timestamp 1605641404
transform 1 0 19688 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1605641404
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1605641404
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1605641404
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1605641404
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1605641404
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1605641404
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1605641404
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1605641404
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1605641404
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1605641404
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1605641404
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1605641404
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1605641404
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13064 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1605641404
transform 1 0 12972 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1605641404
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1605641404
transform 1 0 14996 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15456 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_154
timestamp 1605641404
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18032 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1605641404
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_172
timestamp 1605641404
transform 1 0 16928 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1605641404
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19780 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_200
timestamp 1605641404
transform 1 0 19504 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1605641404
transform 1 0 20516 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_209
timestamp 1605641404
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_215
timestamp 1605641404
transform 1 0 20884 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_219
timestamp 1605641404
transform 1 0 21252 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1605641404
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1605641404
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1605641404
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1605641404
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1605641404
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1605641404
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1605641404
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1605641404
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1605641404
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1605641404
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15548 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_166
timestamp 1605641404
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16560 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_184
timestamp 1605641404
transform 1 0 18032 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1605641404
transform 1 0 18584 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19872 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19136 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1605641404
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_202
timestamp 1605641404
transform 1 0 19688 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1605641404
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1605641404
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1605641404
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1605641404
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1605641404
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1605641404
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1605641404
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1605641404
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1605641404
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1605641404
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1605641404
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1605641404
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1605641404
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1605641404
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1605641404
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1605641404
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1605641404
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1605641404
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1605641404
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1605641404
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1605641404
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1605641404
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1605641404
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16100 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1605641404
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_159
timestamp 1605641404
transform 1 0 15732 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1605641404
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1605641404
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_172
timestamp 1605641404
transform 1 0 16928 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1605641404
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1605641404
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1605641404
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1605641404
transform 1 0 19136 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19596 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19688 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_196
timestamp 1605641404
transform 1 0 19136 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_200
timestamp 1605641404
transform 1 0 19504 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_207
timestamp 1605641404
transform 1 0 20148 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1605641404
transform 1 0 18584 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_200
timestamp 1605641404
transform 1 0 19504 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1605641404
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1605641404
transform 1 0 20516 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1605641404
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_215
timestamp 1605641404
transform 1 0 20884 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_219
timestamp 1605641404
transform 1 0 21252 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1605641404
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1605641404
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1605641404
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1605641404
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1605641404
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1605641404
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1605641404
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1605641404
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1605641404
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1605641404
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1605641404
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1605641404
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1605641404
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1605641404
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1605641404
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1605641404
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19688 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_196
timestamp 1605641404
transform 1 0 19136 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_208
timestamp 1605641404
transform 1 0 20240 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1605641404
transform 1 0 20516 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp 1605641404
transform 1 0 20884 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_219
timestamp 1605641404
transform 1 0 21252 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1605641404
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1605641404
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1605641404
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1605641404
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 7912 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_68
timestamp 1605641404
transform 1 0 7360 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1605641404
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11592 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_105
timestamp 1605641404
transform 1 0 10764 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_113
timestamp 1605641404
transform 1 0 11500 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_120
timestamp 1605641404
transform 1 0 12144 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_132
timestamp 1605641404
transform 1 0 13248 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_144
timestamp 1605641404
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1605641404
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1605641404
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1605641404
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1605641404
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1605641404
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_202
timestamp 1605641404
transform 1 0 19688 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1605641404
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1605641404
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1605641404
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1605641404
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1605641404
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1605641404
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1605641404
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1605641404
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1605641404
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1605641404
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 9844 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_86
timestamp 1605641404
transform 1 0 9016 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_94
timestamp 1605641404
transform 1 0 9752 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_101
timestamp 1605641404
transform 1 0 10396 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1605641404
transform 1 0 11500 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1605641404
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1605641404
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1605641404
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1605641404
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1605641404
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1605641404
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1605641404
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1605641404
transform 1 0 19964 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_196
timestamp 1605641404
transform 1 0 19136 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_204
timestamp 1605641404
transform 1 0 19872 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1605641404
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1605641404
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1605641404
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1605641404
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1605641404
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1605641404
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1605641404
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1605641404
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1605641404
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1605641404
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 10488 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1605641404
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_93
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1605641404
transform 1 0 10396 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_108
timestamp 1605641404
transform 1 0 11040 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_120
timestamp 1605641404
transform 1 0 12144 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_132
timestamp 1605641404
transform 1 0 13248 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1605641404
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1605641404
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1605641404
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1605641404
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1605641404
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1605641404
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1605641404
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1605641404
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_202
timestamp 1605641404
transform 1 0 19688 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1605641404
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1605641404
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1605641404
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1605641404
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1605641404
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1605641404
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1605641404
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1605641404
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1605641404
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1605641404
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1605641404
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1605641404
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1605641404
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1605641404
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1605641404
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1605641404
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12420 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1605641404
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1605641404
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_129
timestamp 1605641404
transform 1 0 12972 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_141
timestamp 1605641404
transform 1 0 14076 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_153
timestamp 1605641404
transform 1 0 15180 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_165
timestamp 1605641404
transform 1 0 16284 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1605641404
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_177
timestamp 1605641404
transform 1 0 17388 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1605641404
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1605641404
transform 1 0 19964 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_196
timestamp 1605641404
transform 1 0 19136 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_204
timestamp 1605641404
transform 1 0 19872 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1605641404
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1605641404
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1605641404
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1605641404
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1605641404
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1605641404
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1605641404
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1605641404
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1605641404
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1605641404
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1605641404
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1605641404
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1605641404
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1605641404
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1605641404
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1605641404
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1605641404
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1605641404
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1605641404
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1605641404
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1605641404
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1605641404
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1605641404
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1605641404
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1605641404
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1605641404
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1605641404
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1605641404
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1605641404
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1605641404
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1605641404
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1605641404
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1605641404
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1605641404
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1605641404
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1605641404
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1605641404
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1605641404
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1605641404
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1605641404
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1605641404
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1605641404
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1605641404
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1605641404
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1605641404
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1605641404
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19688 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19688 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1605641404
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1605641404
transform 1 0 20240 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_196
timestamp 1605641404
transform 1 0 19136 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_208
timestamp 1605641404
transform 1 0 20240 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1605641404
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1605641404
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1605641404
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1605641404
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1605641404
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1605641404
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1605641404
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1605641404
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1605641404
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1605641404
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1605641404
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1605641404
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1605641404
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1605641404
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1605641404
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1605641404
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1605641404
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1605641404
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1605641404
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1605641404
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1605641404
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1605641404
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14260 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1605641404
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1605641404
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1605641404
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1605641404
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1605641404
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1605641404
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1605641404
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1605641404
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1605641404
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_202
timestamp 1605641404
transform 1 0 19688 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1605641404
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1605641404
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1605641404
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1605641404
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1605641404
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1605641404
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1605641404
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1605641404
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1605641404
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1605641404
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1605641404
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1605641404
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1605641404
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1605641404
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1605641404
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1605641404
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1605641404
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12420 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1605641404
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1605641404
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_129
timestamp 1605641404
transform 1 0 12972 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_141
timestamp 1605641404
transform 1 0 14076 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1605641404
transform 1 0 15088 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_149
timestamp 1605641404
transform 1 0 14812 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_156
timestamp 1605641404
transform 1 0 15456 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1605641404
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_168
timestamp 1605641404
transform 1 0 16560 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1605641404
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1605641404
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1605641404
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_208
timestamp 1605641404
transform 1 0 20240 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1605641404
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1605641404
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1605641404
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1605641404
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1605641404
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1605641404
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1605641404
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1605641404
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1605641404
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1605641404
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1605641404
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1605641404
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 7728 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 8648 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_68
timestamp 1605641404
transform 1 0 7360 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_78
timestamp 1605641404
transform 1 0 8280 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 9844 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1605641404
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1605641404
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1605641404
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_101
timestamp 1605641404
transform 1 0 10396 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11408 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_109
timestamp 1605641404
transform 1 0 11132 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_118
timestamp 1605641404
transform 1 0 11960 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_130
timestamp 1605641404
transform 1 0 13064 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_142
timestamp 1605641404
transform 1 0 14168 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1605641404
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1605641404
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1605641404
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_166
timestamp 1605641404
transform 1 0 16376 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17112 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1605641404
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1605641404
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_202
timestamp 1605641404
transform 1 0 19688 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1605641404
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1605641404
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1605641404
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1605641404
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1605641404
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1605641404
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1605641404
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1605641404
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1605641404
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1605641404
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1605641404
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1605641404
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1605641404
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1605641404
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1605641404
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1605641404
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1605641404
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1605641404
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1605641404
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1605641404
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1605641404
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1605641404
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1605641404
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_163
timestamp 1605641404
transform 1 0 16100 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1605641404
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_175
timestamp 1605641404
transform 1 0 17204 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1605641404
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1605641404
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_196
timestamp 1605641404
transform 1 0 19136 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_204
timestamp 1605641404
transform 1 0 19872 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1605641404
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1605641404
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1605641404
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1605641404
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1605641404
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1605641404
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1605641404
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1605641404
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1605641404
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1605641404
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1605641404
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1605641404
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1605641404
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1605641404
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1605641404
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1605641404
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1605641404
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1605641404
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1605641404
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1605641404
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1605641404
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1605641404
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1605641404
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1605641404
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1605641404
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1605641404
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1605641404
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1605641404
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1605641404
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1605641404
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1605641404
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1605641404
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1605641404
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1605641404
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1605641404
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1605641404
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1605641404
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal2 s 17130 22320 17186 22800 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 11432 480 11552 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 22320 3816 22800 3936 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 22320 8440 22800 8560 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 22320 8984 22800 9104 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 22320 9392 22800 9512 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 22320 11296 22800 11416 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 22320 11704 22800 11824 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 22320 6128 22800 6248 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 22320 6672 22800 6792 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 22320 7080 22800 7200 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 22320 7488 22800 7608 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 22320 8032 22800 8152 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 22320 13200 22800 13320 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 22320 13608 22800 13728 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 22320 14016 22800 14136 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 22320 14560 22800 14680 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 22320 14968 22800 15088 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 22320 15512 22800 15632 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 22320 15920 22800 16040 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 22320 16872 22800 16992 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 846 0 902 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 7470 0 7526 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 9678 0 9734 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 10230 0 10286 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 1950 0 2006 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2502 0 2558 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3054 0 3110 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 17498 0 17554 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 16394 0 16450 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 5722 22320 5778 22800 6 prog_clk
port 83 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 84 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_35_
port 85 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_36_
port 86 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_37_
port 87 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_38_
port 88 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_39_
port 89 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_40_
port 90 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_41_
port 91 nsew default input
rlabel metal3 s 22320 22448 22800 22568 6 right_top_grid_pin_1_
port 92 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 93 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 94 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
