* NGSPICE file created from grid_io_top.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_1 abstract view
.subckt scs8hd_ebufn_1 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_and4_4 abstract view
.subckt scs8hd_and4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

.subckt grid_io_top address[0] address[1] address[2] address[3] bottom_width_0_height_0__pin_0_
+ bottom_width_0_height_0__pin_10_ bottom_width_0_height_0__pin_11_ bottom_width_0_height_0__pin_12_
+ bottom_width_0_height_0__pin_13_ bottom_width_0_height_0__pin_14_ bottom_width_0_height_0__pin_15_
+ bottom_width_0_height_0__pin_1_ bottom_width_0_height_0__pin_2_ bottom_width_0_height_0__pin_3_
+ bottom_width_0_height_0__pin_4_ bottom_width_0_height_0__pin_5_ bottom_width_0_height_0__pin_6_
+ bottom_width_0_height_0__pin_7_ bottom_width_0_height_0__pin_8_ bottom_width_0_height_0__pin_9_
+ data_in enable gfpga_pad_GPIO_PAD[0] gfpga_pad_GPIO_PAD[1] gfpga_pad_GPIO_PAD[2]
+ gfpga_pad_GPIO_PAD[3] gfpga_pad_GPIO_PAD[4] gfpga_pad_GPIO_PAD[5] gfpga_pad_GPIO_PAD[6]
+ gfpga_pad_GPIO_PAD[7] vpwr vgnd
XFILLER_11_818 vgnd vpwr scs8hd_decap_12
XFILLER_11_1086 vgnd vpwr scs8hd_decap_12
XFILLER_14_678 vgnd vpwr scs8hd_decap_12
XFILLER_6_800 vgnd vpwr scs8hd_decap_12
XFILLER_6_855 vgnd vpwr scs8hd_decap_12
XFILLER_9_159 vgnd vpwr scs8hd_decap_12
XFILLER_10_873 vgnd vpwr scs8hd_decap_12
XFILLER_3_23 vgnd vpwr scs8hd_decap_12
XFILLER_5_354 vgnd vpwr scs8hd_decap_12
XFILLER_7_1143 vgnd vpwr scs8hd_decap_3
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_11_659 vgnd vpwr scs8hd_decap_12
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_2_379 vgnd vpwr scs8hd_fill_1
XFILLER_2_324 vgnd vpwr scs8hd_decap_12
XFILLER_3_847 vpwr vgnd scs8hd_fill_2
XFILLER_6_663 vgnd vpwr scs8hd_decap_8
XFILLER_2_880 vgnd vpwr scs8hd_decap_4
XFILLER_5_195 vgnd vpwr scs8hd_decap_12
XFILLER_16_707 vgnd vpwr scs8hd_decap_6
XFILLER_11_489 vgnd vpwr scs8hd_decap_12
XFILLER_3_611 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XFILLER_6_471 vgnd vpwr scs8hd_decap_12
XFILLER_9_1013 vgnd vpwr scs8hd_decap_12
XFILLER_0_614 vgnd vpwr scs8hd_decap_6
XFILLER_16_559 vgnd vpwr scs8hd_decap_12
XFILLER_12_776 vgnd vpwr scs8hd_decap_12
XFILLER_8_703 vgnd vpwr scs8hd_decap_12
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
XFILLER_3_452 vgnd vpwr scs8hd_decap_12
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_728 vgnd vpwr scs8hd_decap_4
XFILLER_1_989 vgnd vpwr scs8hd_decap_12
XFILLER_0_466 vgnd vpwr scs8hd_decap_12
XFILLER_16_323 vgnd vpwr scs8hd_decap_12
XPHY_373 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_362 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_351 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_340 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_544 vgnd vpwr scs8hd_decap_12
XFILLER_3_293 vgnd vpwr scs8hd_decap_12
XFILLER_4_750 vgnd vpwr scs8hd_decap_12
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_14_849 vgnd vpwr scs8hd_decap_12
XFILLER_15_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_5_525 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_385 vgnd vpwr scs8hd_decap_12
XFILLER_9_842 vgnd vpwr scs8hd_decap_12
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_6_812 vgnd vpwr scs8hd_decap_12
XFILLER_6_867 vgnd vpwr scs8hd_decap_12
XFILLER_1_550 vgnd vpwr scs8hd_decap_6
XFILLER_3_35 vgnd vpwr scs8hd_decap_12
XFILLER_5_388 vpwr vgnd scs8hd_fill_2
XFILLER_7_1111 vgnd vpwr scs8hd_decap_12
XFILLER_9_672 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_15_977 vgnd vpwr scs8hd_decap_12
XFILLER_14_410 vgnd vpwr scs8hd_decap_12
XFILLER_0_807 vgnd vpwr scs8hd_decap_12
XFILLER_12_947 vgnd vpwr scs8hd_decap_12
XFILLER_7_428 vgnd vpwr scs8hd_decap_12
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XFILLER_7_940 vgnd vpwr scs8hd_decap_12
XFILLER_6_483 vgnd vpwr scs8hd_decap_12
XFILLER_9_1025 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _10_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_788 vgnd vpwr scs8hd_decap_12
XFILLER_8_715 vgnd vpwr scs8hd_decap_12
XFILLER_11_232 vgnd vpwr scs8hd_decap_12
XFILLER_3_420 vgnd vpwr scs8hd_decap_6
XFILLER_3_464 vgnd vpwr scs8hd_decap_12
XFILLER_4_910 vgnd vpwr scs8hd_decap_12
XFILLER_7_269 vgnd vpwr scs8hd_decap_12
XFILLER_7_781 vgnd vpwr scs8hd_decap_12
XFILLER_1_902 vgnd vpwr scs8hd_decap_12
XFILLER_0_412 vgnd vpwr scs8hd_decap_3
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_1_957 vgnd vpwr scs8hd_decap_12
XFILLER_0_478 vgnd vpwr scs8hd_decap_12
XFILLER_0_423 vgnd vpwr scs8hd_decap_8
XFILLER_16_335 vgnd vpwr scs8hd_decap_6
XPHY_352 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_341 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_330 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_374 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_363 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_556 vgnd vpwr scs8hd_decap_12
XFILLER_4_762 vgnd vpwr scs8hd_fill_1
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XFILLER_5_537 vgnd vpwr scs8hd_decap_6
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XFILLER_5_1050 vgnd vpwr scs8hd_decap_12
XFILLER_16_187 vgnd vpwr scs8hd_decap_12
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_581 vgnd vpwr scs8hd_decap_12
XFILLER_11_1099 vgnd vpwr scs8hd_decap_12
XFILLER_2_507 vgnd vpwr scs8hd_decap_12
XFILLER_13_135 vgnd vpwr scs8hd_decap_12
XFILLER_5_367 vgnd vpwr scs8hd_decap_12
XFILLER_6_879 vgnd vpwr scs8hd_decap_6
XFILLER_10_886 vgnd vpwr scs8hd_decap_12
XFILLER_3_47 vgnd vpwr scs8hd_decap_12
XFILLER_7_1123 vgnd vpwr scs8hd_decap_12
XFILLER_12_190 vgnd vpwr scs8hd_decap_12
XFILLER_9_684 vgnd vpwr scs8hd_decap_12
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_337 vgnd vpwr scs8hd_decap_12
XFILLER_14_422 vgnd vpwr scs8hd_decap_12
XFILLER_2_1020 vgnd vpwr scs8hd_decap_12
XFILLER_15_989 vgnd vpwr scs8hd_decap_12
XFILLER_0_819 vgnd vpwr scs8hd_decap_12
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_12_959 vgnd vpwr scs8hd_decap_12
XFILLER_11_403 vgnd vpwr scs8hd_decap_12
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_720 vgnd vpwr scs8hd_decap_12
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XFILLER_6_451 vgnd vpwr scs8hd_decap_6
XFILLER_7_952 vgnd vpwr scs8hd_decap_12
XFILLER_6_495 vgnd vpwr scs8hd_decap_12
XFILLER_16_528 vgnd vpwr scs8hd_decap_12
XFILLER_8_727 vgnd vpwr scs8hd_decap_12
XFILLER_3_476 vgnd vpwr scs8hd_decap_12
XFILLER_4_922 vgnd vpwr scs8hd_decap_12
XFILLER_4_944 vpwr vgnd scs8hd_fill_2
XFILLER_8_1081 vgnd vpwr scs8hd_decap_12
XFILLER_15_550 vgnd vpwr scs8hd_decap_12
XFILLER_14_1020 vgnd vpwr scs8hd_decap_12
XFILLER_1_969 vgnd vpwr scs8hd_decap_6
XFILLER_1_914 vgnd vpwr scs8hd_fill_1
XFILLER_0_435 vgnd vpwr scs8hd_decap_12
XPHY_375 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_364 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_353 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_342 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_331 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_320 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_520 vgnd vpwr scs8hd_decap_12
XFILLER_8_568 vgnd vpwr scs8hd_decap_12
XFILLER_16_881 vgnd vpwr scs8hd_decap_12
XFILLER_15_391 vgnd vpwr scs8hd_decap_12
XFILLER_13_306 vgnd vpwr scs8hd_decap_12
XANTENNA__04__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_1_733 vgnd vpwr scs8hd_decap_12
XFILLER_5_1062 vgnd vpwr scs8hd_decap_12
XFILLER_16_199 vgnd vpwr scs8hd_decap_12
XFILLER_12_361 vgnd vpwr scs8hd_decap_12
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_855 vgnd vpwr scs8hd_decap_12
XFILLER_4_593 vgnd vpwr scs8hd_decap_12
XFILLER_8_398 vpwr vgnd scs8hd_fill_2
XFILLER_11_1001 vgnd vpwr scs8hd_decap_12
XFILLER_13_147 vgnd vpwr scs8hd_decap_12
XFILLER_5_379 vgnd vpwr scs8hd_decap_6
XFILLER_6_825 vgnd vpwr scs8hd_decap_4
XFILLER_10_898 vgnd vpwr scs8hd_decap_12
XFILLER_1_563 vgnd vpwr scs8hd_decap_12
XFILLER_7_1135 vgnd vpwr scs8hd_decap_8
XFILLER_9_696 vgnd vpwr scs8hd_decap_12
XFILLER_4_390 vgnd vpwr scs8hd_fill_1
XFILLER_5_891 vgnd vpwr scs8hd_decap_12
XFILLER_10_117 vgnd vpwr scs8hd_decap_12
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_3_806 vgnd vpwr scs8hd_decap_12
XFILLER_2_349 vgnd vpwr scs8hd_decap_12
XFILLER_14_434 vgnd vpwr scs8hd_decap_12
XFILLER_2_1032 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_382 vpwr vgnd scs8hd_fill_2
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_8_ logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[4] vgnd vpwr scs8hd_ebufn_1
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XFILLER_11_415 vgnd vpwr scs8hd_decap_12
XANTENNA__12__A _06_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_4_1105 vgnd vpwr scs8hd_decap_12
XFILLER_7_964 vgnd vpwr scs8hd_decap_12
XFILLER_9_1038 vgnd vpwr scs8hd_decap_12
XANTENNA__07__A _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_400 vpwr vgnd scs8hd_fill_2
XFILLER_4_934 vgnd vpwr scs8hd_decap_8
XFILLER_8_739 vgnd vpwr scs8hd_decap_12
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XFILLER_8_1093 vgnd vpwr scs8hd_decap_12
XFILLER_15_562 vgnd vpwr scs8hd_decap_12
XFILLER_7_794 vgnd vpwr scs8hd_decap_12
XFILLER_14_1032 vgnd vpwr scs8hd_decap_12
XFILLER_0_447 vgnd vpwr scs8hd_decap_12
XFILLER_16_304 vgnd vpwr scs8hd_decap_6
XPHY_376 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_365 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_354 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_343 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_332 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_321 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_310 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_532 vgnd vpwr scs8hd_decap_12
XFILLER_3_241 vgnd vpwr scs8hd_decap_3
XFILLER_4_764 vgnd vpwr scs8hd_decap_12
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_6_1008 vgnd vpwr scs8hd_decap_12
XFILLER_16_893 vgnd vpwr scs8hd_decap_6
XFILLER_13_318 vgnd vpwr scs8hd_decap_12
XFILLER_0_1141 vgnd vpwr scs8hd_decap_4
XANTENNA__20__A gfpga_pad_GPIO_PAD[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_745 vgnd vpwr scs8hd_decap_12
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_16_156 vgnd vpwr scs8hd_decap_12
XFILLER_5_1074 vgnd vpwr scs8hd_decap_12
XFILLER_13_830 vgnd vpwr scs8hd_decap_12
XFILLER_12_373 vgnd vpwr scs8hd_decap_12
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_300 vgnd vpwr scs8hd_decap_12
XFILLER_9_867 vgnd vpwr scs8hd_decap_12
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_11_1013 vgnd vpwr scs8hd_decap_12
XFILLER_14_605 vgnd vpwr scs8hd_decap_12
XFILLER_13_159 vgnd vpwr scs8hd_decap_12
XANTENNA__15__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_10_800 vgnd vpwr scs8hd_decap_12
XFILLER_1_575 vgnd vpwr scs8hd_decap_12
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_3_818 vgnd vpwr scs8hd_decap_12
XFILLER_15_903 vgnd vpwr scs8hd_decap_12
XFILLER_14_446 vgnd vpwr scs8hd_decap_12
XFILLER_2_1044 vgnd vpwr scs8hd_decap_12
XFILLER_2_884 vgnd vpwr scs8hd_fill_1
XFILLER_12_1130 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _12_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__12__B _14_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_615 vgnd vpwr scs8hd_decap_12
XFILLER_4_1117 vgnd vpwr scs8hd_decap_12
XFILLER_15_733 vgnd vpwr scs8hd_decap_12
XFILLER_14_276 vgnd vpwr scs8hd_decap_12
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_10_471 vgnd vpwr scs8hd_decap_12
XFILLER_12_703 vgnd vpwr scs8hd_decap_12
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
XANTENNA__07__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__23__A gfpga_pad_GPIO_PAD[4] vgnd vpwr scs8hd_diode_2
XFILLER_3_489 vgnd vpwr scs8hd_decap_12
XFILLER_15_574 vgnd vpwr scs8hd_decap_12
XFILLER_14_1044 vgnd vpwr scs8hd_decap_12
XFILLER_1_949 vpwr vgnd scs8hd_fill_2
XFILLER_1_916 vgnd vpwr scs8hd_decap_12
XFILLER_0_459 vgnd vpwr scs8hd_decap_6
XFILLER_0_404 vgnd vpwr scs8hd_decap_8
XPHY_300 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__18__A gfpga_pad_GPIO_PAD[7] vgnd vpwr scs8hd_diode_2
XPHY_377 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_366 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_355 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_344 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_333 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_322 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_311 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_544 vgnd vpwr scs8hd_decap_12
XFILLER_4_776 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_0_993 vgnd vpwr scs8hd_decap_12
XFILLER_16_850 vgnd vpwr scs8hd_decap_12
XFILLER_16_1117 vgnd vpwr scs8hd_decap_12
XFILLER_1_757 vgnd vpwr scs8hd_decap_12
XFILLER_16_168 vgnd vpwr scs8hd_decap_12
XFILLER_13_842 vgnd vpwr scs8hd_decap_12
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_5_1086 vgnd vpwr scs8hd_decap_12
XFILLER_12_385 vgnd vpwr scs8hd_decap_12
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_312 vgnd vpwr scs8hd_decap_12
XFILLER_9_879 vgnd vpwr scs8hd_decap_12
XFILLER_4_551 vgnd vpwr scs8hd_decap_12
XFILLER_11_1025 vgnd vpwr scs8hd_decap_12
XFILLER_14_617 vgnd vpwr scs8hd_decap_12
XANTENNA__15__B _14_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_812 vgnd vpwr scs8hd_decap_12
XFILLER_1_587 vgnd vpwr scs8hd_decap_12
XFILLER_13_672 vgnd vpwr scs8hd_decap_12
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_9 vgnd vpwr scs8hd_fill_1
XFILLER_2_1056 vgnd vpwr scs8hd_decap_12
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XFILLER_10_642 vgnd vpwr scs8hd_decap_12
XFILLER_9_440 vgnd vpwr scs8hd_decap_12
XFILLER_12_1142 vgnd vpwr scs8hd_decap_4
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_11_428 vgnd vpwr scs8hd_decap_12
XFILLER_3_627 vgnd vpwr scs8hd_decap_12
XANTENNA__12__C _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_745 vgnd vpwr scs8hd_decap_12
XFILLER_14_288 vgnd vpwr scs8hd_decap_12
XFILLER_11_940 vgnd vpwr scs8hd_decap_12
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
XFILLER_7_977 vgnd vpwr scs8hd_decap_12
XFILLER_10_483 vgnd vpwr scs8hd_decap_12
XFILLER_9_281 vgnd vpwr scs8hd_decap_12
XFILLER_16_509 vgnd vpwr scs8hd_decap_12
XANTENNA__07__C _06_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_715 vgnd vpwr scs8hd_decap_12
XFILLER_11_269 vgnd vpwr scs8hd_decap_12
XFILLER_4_958 vgnd vpwr scs8hd_decap_12
XFILLER_15_586 vgnd vpwr scs8hd_decap_12
XFILLER_11_781 vgnd vpwr scs8hd_decap_12
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
XFILLER_14_1056 vgnd vpwr scs8hd_decap_12
XFILLER_1_928 vgnd vpwr scs8hd_decap_12
XPHY_334 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_323 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_301 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_312 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_378 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_367 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_356 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_345 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_556 vgnd vpwr scs8hd_decap_12
XFILLER_3_221 vgnd vpwr scs8hd_decap_12
XFILLER_4_788 vgnd vpwr scs8hd_decap_12
XFILLER_16_862 vgnd vpwr scs8hd_decap_6
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_1110 vgnd vpwr scs8hd_decap_6
XFILLER_16_1129 vgnd vpwr scs8hd_decap_12
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_1_769 vgnd vpwr scs8hd_decap_12
XFILLER_16_125 vgnd vpwr scs8hd_decap_12
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_324 vgnd vpwr scs8hd_decap_12
XFILLER_4_563 vgnd vpwr scs8hd_decap_12
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_14_629 vgnd vpwr scs8hd_decap_12
XANTENNA__15__C _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_599 vgnd vpwr scs8hd_decap_8
XFILLER_13_684 vgnd vpwr scs8hd_decap_12
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XFILLER_9_611 vgnd vpwr scs8hd_decap_12
XFILLER_4_382 vgnd vpwr scs8hd_decap_8
XFILLER_4_393 vpwr vgnd scs8hd_fill_2
XFILLER_5_850 vgnd vpwr scs8hd_decap_4
XFILLER_10_1081 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XFILLER_15_916 vgnd vpwr scs8hd_decap_12
XFILLER_14_459 vgnd vpwr scs8hd_decap_12
XFILLER_10_654 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_1_330 vgnd vpwr scs8hd_decap_12
XFILLER_2_886 vgnd vpwr scs8hd_decap_12
XFILLER_14_971 vgnd vpwr scs8hd_decap_12
XFILLER_9_452 vgnd vpwr scs8hd_decap_12
XFILLER_5_680 vgnd vpwr scs8hd_decap_12
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XFILLER_3_639 vgnd vpwr scs8hd_decap_12
XANTENNA__12__D _09_/D vgnd vpwr scs8hd_diode_2
XFILLER_15_757 vgnd vpwr scs8hd_decap_12
XFILLER_11_952 vgnd vpwr scs8hd_decap_12
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_495 vgnd vpwr scs8hd_decap_12
XFILLER_2_694 vgnd vpwr scs8hd_decap_8
XFILLER_7_989 vgnd vpwr scs8hd_decap_12
XFILLER_9_293 vgnd vpwr scs8hd_decap_12
XANTENNA__07__D enable vgnd vpwr scs8hd_diode_2
XFILLER_12_727 vgnd vpwr scs8hd_decap_12
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
XFILLER_15_598 vgnd vpwr scs8hd_decap_12
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
XFILLER_7_720 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XPHY_368 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_357 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_346 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_335 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_324 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_302 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_313 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_379 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_568 vgnd vpwr scs8hd_decap_12
XFILLER_4_701 vgnd vpwr scs8hd_fill_1
XFILLER_0_962 vgnd vpwr scs8hd_decap_12
XFILLER_3_233 vgnd vpwr scs8hd_decap_8
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_550 vgnd vpwr scs8hd_decap_12
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
X_09_ address[1] enable address[3] _09_/D _09_/X vgnd vpwr scs8hd_and4_4
XFILLER_1_704 vgnd vpwr scs8hd_decap_12
XFILLER_16_137 vgnd vpwr scs8hd_decap_12
XFILLER_5_1099 vgnd vpwr scs8hd_decap_12
XFILLER_13_855 vgnd vpwr scs8hd_decap_12
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_398 vgnd vpwr scs8hd_decap_12
XFILLER_4_520 vgnd vpwr scs8hd_decap_8
XFILLER_4_575 vgnd vpwr scs8hd_decap_4
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_11_1038 vgnd vpwr scs8hd_decap_12
XANTENNA__15__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_10_825 vgnd vpwr scs8hd_decap_12
XFILLER_1_501 vgnd vpwr scs8hd_decap_12
XFILLER_5_306 vgnd vpwr scs8hd_decap_12
XFILLER_1_556 vgnd vpwr scs8hd_fill_1
XFILLER_13_696 vgnd vpwr scs8hd_decap_12
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XFILLER_9_623 vgnd vpwr scs8hd_decap_12
XFILLER_4_361 vgnd vpwr scs8hd_decap_8
XFILLER_10_1093 vgnd vpwr scs8hd_decap_12
XFILLER_16_490 vgnd vpwr scs8hd_decap_6
XFILLER_15_928 vgnd vpwr scs8hd_decap_12
XFILLER_2_1003 vgnd vpwr scs8hd_decap_4
XFILLER_2_1069 vgnd vpwr scs8hd_decap_12
XFILLER_10_666 vgnd vpwr scs8hd_decap_12
XFILLER_1_342 vgnd vpwr scs8hd_decap_12
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_386 vgnd vpwr scs8hd_decap_12
XFILLER_2_898 vgnd vpwr scs8hd_decap_12
XFILLER_14_983 vgnd vpwr scs8hd_decap_12
XFILLER_9_464 vgnd vpwr scs8hd_decap_12
XFILLER_4_51 vgnd vpwr scs8hd_decap_12
XFILLER_5_692 vgnd vpwr scs8hd_decap_12
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_769 vgnd vpwr scs8hd_decap_12
XFILLER_14_202 vgnd vpwr scs8hd_decap_12
XFILLER_11_964 vgnd vpwr scs8hd_decap_12
XFILLER_12_739 vgnd vpwr scs8hd_decap_12
XFILLER_3_404 vpwr vgnd scs8hd_fill_2
XFILLER_3_426 vgnd vpwr scs8hd_fill_1
XFILLER_8_1020 vgnd vpwr scs8hd_decap_12
XFILLER_11_794 vgnd vpwr scs8hd_decap_12
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XFILLER_14_1069 vgnd vpwr scs8hd_decap_12
XPHY_369 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_358 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_347 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_336 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_325 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_303 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_314 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_507 vgnd vpwr scs8hd_decap_12
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_974 vgnd vpwr scs8hd_decap_12
XFILLER_16_831 vgnd vpwr scs8hd_decap_6
XFILLER_15_330 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_10_ logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[5] vgnd vpwr scs8hd_ebufn_1
XFILLER_7_562 vgnd vpwr scs8hd_decap_12
X_08_ address[2] _09_/D vgnd vpwr scs8hd_inv_8
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_0_1145 vgnd vpwr scs8hd_fill_1
XFILLER_1_716 vgnd vpwr scs8hd_decap_12
XFILLER_5_1001 vgnd vpwr scs8hd_decap_12
XFILLER_16_149 vgnd vpwr scs8hd_decap_6
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_14_ vgnd vpwr scs8hd_diode_2
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_867 vgnd vpwr scs8hd_decap_12
XFILLER_12_300 vgnd vpwr scs8hd_decap_12
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_337 vgnd vpwr scs8hd_decap_12
XFILLER_16_683 vgnd vpwr scs8hd_decap_12
XFILLER_15_171 vgnd vpwr scs8hd_decap_12
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_7_392 vpwr vgnd scs8hd_fill_2
XFILLER_10_837 vgnd vpwr scs8hd_decap_12
XFILLER_1_513 vgnd vpwr scs8hd_decap_12
XFILLER_5_318 vgnd vpwr scs8hd_decap_12
XFILLER_12_141 vgnd vpwr scs8hd_decap_12
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XFILLER_9_635 vgnd vpwr scs8hd_decap_12
XFILLER_0_590 vgnd vpwr scs8hd_decap_12
XFILLER_8_690 vgnd vpwr scs8hd_decap_12
XFILLER_6_605 vgnd vpwr scs8hd_decap_12
XFILLER_10_678 vgnd vpwr scs8hd_decap_12
XFILLER_1_354 vgnd vpwr scs8hd_decap_12
XFILLER_2_800 vgnd vpwr scs8hd_decap_12
XFILLER_2_833 vgnd vpwr scs8hd_decap_3
XFILLER_2_844 vgnd vpwr scs8hd_decap_12
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XFILLER_1_398 vgnd vpwr scs8hd_decap_12
XFILLER_14_995 vgnd vpwr scs8hd_decap_12
XFILLER_9_476 vgnd vpwr scs8hd_decap_12
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XFILLER_4_63 vgnd vpwr scs8hd_decap_12
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XFILLER_3_608 vpwr vgnd scs8hd_fill_2
XFILLER_6_457 vgnd vpwr scs8hd_fill_1
XFILLER_7_903 vgnd vpwr scs8hd_decap_12
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_10_ vgnd vpwr scs8hd_diode_2
XFILLER_3_1143 vgnd vpwr scs8hd_decap_3
XFILLER_8_1032 vgnd vpwr scs8hd_decap_12
XFILLER_15_501 vgnd vpwr scs8hd_decap_12
XFILLER_7_733 vgnd vpwr scs8hd_decap_12
XFILLER_6_276 vgnd vpwr scs8hd_decap_12
XFILLER_2_471 vgnd vpwr scs8hd_decap_12
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XFILLER_0_419 vpwr vgnd scs8hd_fill_2
XPHY_359 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_348 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_337 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_326 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_304 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_315 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_714 vgnd vpwr scs8hd_decap_12
XFILLER_0_986 vgnd vpwr scs8hd_decap_6
XFILLER_0_931 vgnd vpwr scs8hd_decap_12
XFILLER_15_342 vgnd vpwr scs8hd_decap_12
XFILLER_7_574 vgnd vpwr scs8hd_decap_12
X_07_ _04_/X address[2] _06_/Y enable _07_/X vgnd vpwr scs8hd_and4_4
XFILLER_1_728 vgnd vpwr scs8hd_decap_4
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
XFILLER_5_1013 vgnd vpwr scs8hd_decap_12
XFILLER_16_106 vgnd vpwr scs8hd_decap_12
XFILLER_12_312 vgnd vpwr scs8hd_decap_12
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_879 vgnd vpwr scs8hd_decap_12
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_349 vgnd vpwr scs8hd_decap_12
XFILLER_9_806 vgnd vpwr scs8hd_decap_12
XFILLER_16_695 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_1143 vgnd vpwr scs8hd_decap_3
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_8_861 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_6_ vgnd vpwr scs8hd_diode_2
XFILLER_10_849 vgnd vpwr scs8hd_decap_12
XFILLER_1_525 vgnd vpwr scs8hd_decap_12
XFILLER_16_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_647 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_1130 vgnd vpwr scs8hd_decap_12
XFILLER_6_617 vgnd vpwr scs8hd_decap_12
XFILLER_2_812 vgnd vpwr scs8hd_decap_12
XFILLER_2_856 vgnd vpwr scs8hd_decap_12
XFILLER_13_440 vgnd vpwr scs8hd_decap_12
XFILLER_5_672 vpwr vgnd scs8hd_fill_2
XFILLER_4_75 vgnd vpwr scs8hd_decap_12
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_977 vgnd vpwr scs8hd_decap_12
XFILLER_10_410 vgnd vpwr scs8hd_decap_12
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_2_642 vgnd vpwr scs8hd_decap_12
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XFILLER_13_281 vgnd vpwr scs8hd_decap_12
XFILLER_3_1111 vgnd vpwr scs8hd_decap_12
XFILLER_3_428 vgnd vpwr scs8hd_decap_12
XFILLER_1_7 vpwr vgnd scs8hd_fill_2
XFILLER_8_1044 vgnd vpwr scs8hd_decap_12
XFILLER_15_513 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_2_ vgnd vpwr scs8hd_diode_2
XFILLER_7_745 vgnd vpwr scs8hd_decap_12
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
XFILLER_2_483 vgnd vpwr scs8hd_decap_12
XFILLER_3_940 vgnd vpwr scs8hd_decap_6
XFILLER_3_973 vgnd vpwr scs8hd_decap_3
XFILLER_6_288 vgnd vpwr scs8hd_decap_12
X_23_ gfpga_pad_GPIO_PAD[4] bottom_width_0_height_0__pin_9_ vgnd vpwr scs8hd_buf_2
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _12_/Y vgnd vpwr scs8hd_diode_2
XPHY_305 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_316 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_349 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_338 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_327 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_269 vgnd vpwr scs8hd_decap_12
XFILLER_4_726 vgnd vpwr scs8hd_decap_12
XFILLER_16_800 vgnd vpwr scs8hd_decap_6
XFILLER_0_943 vgnd vpwr scs8hd_decap_12
XFILLER_15_354 vgnd vpwr scs8hd_decap_12
XFILLER_7_586 vgnd vpwr scs8hd_decap_12
XFILLER_3_781 vgnd vpwr scs8hd_decap_12
X_06_ address[1] _06_/Y vgnd vpwr scs8hd_inv_8
XFILLER_5_1025 vgnd vpwr scs8hd_decap_12
XFILLER_16_118 vgnd vpwr scs8hd_decap_6
XFILLER_12_324 vgnd vpwr scs8hd_decap_12
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_818 vgnd vpwr scs8hd_decap_12
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_652 vgnd vpwr scs8hd_decap_12
XFILLER_15_1111 vgnd vpwr scs8hd_decap_12
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_8_873 vgnd vpwr scs8hd_decap_12
XFILLER_1_559 vpwr vgnd scs8hd_fill_2
XFILLER_1_537 vgnd vpwr scs8hd_decap_12
XFILLER_13_611 vgnd vpwr scs8hd_decap_12
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XFILLER_9_659 vgnd vpwr scs8hd_decap_12
XFILLER_6_1142 vgnd vpwr scs8hd_decap_4
XFILLER_6_629 vgnd vpwr scs8hd_decap_12
XFILLER_1_367 vgnd vpwr scs8hd_decap_12
XFILLER_2_868 vgnd vpwr scs8hd_decap_12
XFILLER_13_452 vgnd vpwr scs8hd_decap_12
XFILLER_9_489 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_4
XFILLER_5_640 vpwr vgnd scs8hd_fill_2
XFILLER_1_890 vgnd vpwr scs8hd_decap_12
XFILLER_4_87 vgnd vpwr scs8hd_decap_4
XFILLER_1_1050 vgnd vpwr scs8hd_decap_12
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
XFILLER_11_989 vgnd vpwr scs8hd_decap_12
XFILLER_6_415 vgnd vpwr scs8hd_decap_12
XFILLER_7_916 vgnd vpwr scs8hd_decap_12
XFILLER_10_422 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_131 vgnd vpwr scs8hd_decap_12
XFILLER_2_654 vgnd vpwr scs8hd_decap_12
XFILLER_6_459 vgnd vpwr scs8hd_decap_12
XFILLER_13_293 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _05_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_971 vgnd vpwr scs8hd_decap_12
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XFILLER_3_1123 vgnd vpwr scs8hd_decap_12
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XFILLER_8_1056 vgnd vpwr scs8hd_decap_12
XFILLER_15_525 vgnd vpwr scs8hd_decap_12
XFILLER_11_720 vgnd vpwr scs8hd_decap_12
XFILLER_7_757 vgnd vpwr scs8hd_decap_12
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
XFILLER_2_495 vgnd vpwr scs8hd_decap_12
X_22_ gfpga_pad_GPIO_PAD[3] bottom_width_0_height_0__pin_7_ vgnd vpwr scs8hd_buf_2
XFILLER_1_11 vgnd vpwr scs8hd_decap_12
XPHY_339 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_328 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_306 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_317 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_955 vgnd vpwr scs8hd_decap_6
XFILLER_0_900 vgnd vpwr scs8hd_decap_12
XFILLER_3_204 vgnd vpwr scs8hd_decap_3
XFILLER_4_738 vgnd vpwr scs8hd_decap_12
XFILLER_11_550 vgnd vpwr scs8hd_decap_12
XFILLER_13_1050 vgnd vpwr scs8hd_decap_12
XFILLER_7_598 vgnd vpwr scs8hd_decap_12
X_05_ _04_/X address[2] address[1] enable _05_/X vgnd vpwr scs8hd_and4_4
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_579 vgnd vpwr scs8hd_fill_1
XFILLER_16_664 vgnd vpwr scs8hd_decap_12
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_1123 vgnd vpwr scs8hd_decap_12
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XFILLER_11_391 vgnd vpwr scs8hd_decap_12
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XFILLER_4_1081 vgnd vpwr scs8hd_decap_12
XFILLER_16_63 vgnd vpwr scs8hd_decap_12
XFILLER_13_623 vgnd vpwr scs8hd_decap_12
XFILLER_12_166 vgnd vpwr scs8hd_decap_12
XFILLER_5_822 vgnd vpwr scs8hd_fill_1
XFILLER_5_855 vgnd vpwr scs8hd_decap_12
XFILLER_10_1020 vgnd vpwr scs8hd_decap_12
XFILLER_0_571 vpwr vgnd scs8hd_fill_2
XFILLER_2_825 vgnd vpwr scs8hd_decap_8
XFILLER_1_379 vgnd vpwr scs8hd_fill_1
XFILLER_14_910 vgnd vpwr scs8hd_decap_12
XFILLER_13_464 vgnd vpwr scs8hd_decap_12
XFILLER_4_11 vgnd vpwr scs8hd_fill_1
XFILLER_5_652 vgnd vpwr scs8hd_decap_12
XFILLER_16_280 vgnd vpwr scs8hd_decap_12
XFILLER_1_1062 vgnd vpwr scs8hd_decap_12
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
XFILLER_13_86 vgnd vpwr scs8hd_decap_12
XFILLER_6_427 vgnd vpwr scs8hd_decap_12
XFILLER_7_928 vgnd vpwr scs8hd_decap_12
XFILLER_10_434 vgnd vpwr scs8hd_decap_12
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_143 vgnd vpwr scs8hd_decap_12
XFILLER_2_666 vgnd vpwr scs8hd_decap_12
XFILLER_14_751 vgnd vpwr scs8hd_decap_12
XFILLER_9_232 vgnd vpwr scs8hd_decap_12
XFILLER_6_983 vgnd vpwr scs8hd_decap_12
XFILLER_3_1135 vgnd vpwr scs8hd_decap_8
XFILLER_3_408 vgnd vpwr scs8hd_decap_12
XFILLER_15_537 vgnd vpwr scs8hd_decap_12
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
XFILLER_7_769 vgnd vpwr scs8hd_decap_12
XFILLER_1_23 vgnd vpwr scs8hd_decap_12
X_21_ gfpga_pad_GPIO_PAD[2] bottom_width_0_height_0__pin_5_ vgnd vpwr scs8hd_buf_2
XFILLER_3_953 vgnd vpwr scs8hd_decap_12
XFILLER_14_581 vgnd vpwr scs8hd_decap_12
XPHY_329 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_307 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_318 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_507 vgnd vpwr scs8hd_decap_12
XFILLER_0_912 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_15_367 vgnd vpwr scs8hd_decap_12
XFILLER_11_562 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _13_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_1062 vgnd vpwr scs8hd_decap_12
XFILLER_3_794 vgnd vpwr scs8hd_decap_12
X_04_ address[3] _04_/X vgnd vpwr scs8hd_buf_1
XFILLER_5_1038 vgnd vpwr scs8hd_decap_12
XFILLER_12_337 vgnd vpwr scs8hd_decap_12
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_742 vpwr vgnd scs8hd_fill_2
XFILLER_16_676 vgnd vpwr scs8hd_decap_6
XFILLER_16_621 vgnd vpwr scs8hd_decap_12
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_1135 vgnd vpwr scs8hd_decap_8
XFILLER_7_330 vgnd vpwr scs8hd_decap_12
XFILLER_8_886 vgnd vpwr scs8hd_decap_12
XFILLER_7_385 vgnd vpwr scs8hd_fill_1
XFILLER_4_1093 vgnd vpwr scs8hd_decap_12
XFILLER_16_75 vgnd vpwr scs8hd_decap_12
XFILLER_13_635 vgnd vpwr scs8hd_decap_12
XFILLER_12_178 vgnd vpwr scs8hd_decap_12
XFILLER_4_300 vgnd vpwr scs8hd_decap_12
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_5_867 vgnd vpwr scs8hd_decap_12
XFILLER_10_1032 vgnd vpwr scs8hd_decap_12
XFILLER_12_690 vgnd vpwr scs8hd_decap_12
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XFILLER_2_1008 vgnd vpwr scs8hd_decap_12
XFILLER_10_605 vgnd vpwr scs8hd_decap_12
XFILLER_14_922 vgnd vpwr scs8hd_decap_12
XFILLER_13_476 vgnd vpwr scs8hd_decap_12
XFILLER_9_403 vgnd vpwr scs8hd_decap_12
XFILLER_12_1105 vgnd vpwr scs8hd_decap_12
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_5_664 vgnd vpwr scs8hd_decap_4
XFILLER_1_1074 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_12_ logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[6] vgnd vpwr scs8hd_ebufn_1
XFILLER_16_292 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_708 vgnd vpwr scs8hd_decap_12
XFILLER_11_903 vgnd vpwr scs8hd_decap_12
XFILLER_13_98 vgnd vpwr scs8hd_decap_12
XFILLER_6_439 vgnd vpwr scs8hd_decap_12
XFILLER_10_446 vgnd vpwr scs8hd_decap_12
XFILLER_1_155 vgnd vpwr scs8hd_decap_12
XFILLER_2_678 vgnd vpwr scs8hd_decap_8
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_995 vgnd vpwr scs8hd_decap_12
XFILLER_8_1069 vgnd vpwr scs8hd_decap_12
XFILLER_11_733 vgnd vpwr scs8hd_decap_12
XFILLER_3_965 vgnd vpwr scs8hd_decap_8
XFILLER_10_276 vgnd vpwr scs8hd_decap_12
XFILLER_1_35 vgnd vpwr scs8hd_decap_12
X_20_ gfpga_pad_GPIO_PAD[1] bottom_width_0_height_0__pin_3_ vgnd vpwr scs8hd_buf_2
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_1008 vgnd vpwr scs8hd_decap_12
XFILLER_14_593 vgnd vpwr scs8hd_decap_12
XPHY_308 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_319 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_0_924 vgnd vpwr scs8hd_decap_6
XFILLER_16_869 vgnd vpwr scs8hd_decap_12
XFILLER_15_379 vgnd vpwr scs8hd_decap_12
XFILLER_11_574 vgnd vpwr scs8hd_decap_12
XFILLER_7_501 vgnd vpwr scs8hd_decap_12
XFILLER_13_1074 vgnd vpwr scs8hd_decap_12
XFILLER_0_1117 vgnd vpwr scs8hd_decap_12
XFILLER_15_891 vgnd vpwr scs8hd_decap_12
XFILLER_13_806 vgnd vpwr scs8hd_decap_12
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_349 vgnd vpwr scs8hd_decap_12
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_776 vgnd vpwr scs8hd_decap_12
XFILLER_16_633 vgnd vpwr scs8hd_decap_12
XFILLER_15_110 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_12_861 vgnd vpwr scs8hd_decap_12
XFILLER_7_342 vgnd vpwr scs8hd_decap_12
XFILLER_8_898 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _05_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_87 vgnd vpwr scs8hd_decap_6
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_647 vgnd vpwr scs8hd_decap_12
XFILLER_4_312 vgnd vpwr scs8hd_decap_12
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XFILLER_0_540 vgnd vpwr scs8hd_decap_12
XFILLER_5_879 vgnd vpwr scs8hd_decap_12
XFILLER_10_1044 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_617 vgnd vpwr scs8hd_decap_12
XFILLER_14_934 vgnd vpwr scs8hd_decap_12
XFILLER_9_415 vgnd vpwr scs8hd_decap_12
XFILLER_12_1117 vgnd vpwr scs8hd_decap_12
XFILLER_5_676 vpwr vgnd scs8hd_fill_2
XFILLER_4_186 vgnd vpwr scs8hd_decap_12
XFILLER_1_1086 vgnd vpwr scs8hd_decap_12
XFILLER_1_167 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_764 vgnd vpwr scs8hd_decap_12
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_440 vgnd vpwr scs8hd_decap_12
XFILLER_11_745 vgnd vpwr scs8hd_decap_12
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_2_410 vgnd vpwr scs8hd_decap_12
XFILLER_3_977 vgnd vpwr scs8hd_decap_12
XFILLER_10_288 vgnd vpwr scs8hd_decap_12
XFILLER_1_47 vgnd vpwr scs8hd_decap_12
XFILLER_5_281 vgnd vpwr scs8hd_decap_12
XPHY_309 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_1086 vgnd vpwr scs8hd_decap_12
XFILLER_11_586 vgnd vpwr scs8hd_decap_12
XFILLER_7_513 vgnd vpwr scs8hd_decap_12
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_0_1129 vgnd vpwr scs8hd_decap_12
XFILLER_9_1143 vgnd vpwr scs8hd_decap_3
XFILLER_13_818 vgnd vpwr scs8hd_decap_12
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_722 vgnd vpwr scs8hd_decap_12
XFILLER_0_788 vgnd vpwr scs8hd_decap_12
XFILLER_16_645 vgnd vpwr scs8hd_decap_6
XFILLER_12_873 vgnd vpwr scs8hd_decap_12
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_8_800 vgnd vpwr scs8hd_decap_12
XFILLER_7_354 vgnd vpwr scs8hd_decap_12
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_659 vgnd vpwr scs8hd_decap_12
XFILLER_4_324 vgnd vpwr scs8hd_decap_12
XFILLER_5_825 vpwr vgnd scs8hd_fill_2
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XFILLER_10_1056 vgnd vpwr scs8hd_decap_12
XFILLER_0_552 vgnd vpwr scs8hd_decap_6
XFILLER_16_497 vgnd vpwr scs8hd_decap_12
XFILLER_4_880 vgnd vpwr scs8hd_decap_4
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
XFILLER_10_629 vgnd vpwr scs8hd_decap_12
XFILLER_13_489 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_14 vgnd vpwr scs8hd_decap_12
XFILLER_4_36 vgnd vpwr scs8hd_fill_1
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_4_198 vgnd vpwr scs8hd_decap_12
XFILLER_5_611 vgnd vpwr scs8hd_decap_12
XFILLER_5_644 vpwr vgnd scs8hd_fill_2
XFILLER_16_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_471 vgnd vpwr scs8hd_decap_12
XFILLER_11_916 vgnd vpwr scs8hd_decap_12
XFILLER_10_459 vgnd vpwr scs8hd_decap_12
XFILLER_1_179 vgnd vpwr scs8hd_decap_4
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XFILLER_14_776 vgnd vpwr scs8hd_decap_12
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_971 vgnd vpwr scs8hd_decap_12
XFILLER_5_452 vgnd vpwr scs8hd_decap_12
XFILLER_11_757 vgnd vpwr scs8hd_decap_12
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XFILLER_2_422 vgnd vpwr scs8hd_decap_12
XFILLER_3_989 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XFILLER_5_293 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_16_838 vgnd vpwr scs8hd_decap_12
XFILLER_11_598 vgnd vpwr scs8hd_decap_12
XFILLER_7_525 vgnd vpwr scs8hd_decap_12
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_9_1111 vgnd vpwr scs8hd_decap_12
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_528 vpwr vgnd scs8hd_fill_2
XFILLER_4_539 vgnd vpwr scs8hd_decap_12
XFILLER_0_745 vgnd vpwr scs8hd_decap_12
XFILLER_0_734 vgnd vpwr scs8hd_decap_8
XANTENNA__10__A _06_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_602 vgnd vpwr scs8hd_decap_12
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_8_812 vgnd vpwr scs8hd_decap_12
XFILLER_3_550 vgnd vpwr scs8hd_decap_12
XFILLER_7_388 vpwr vgnd scs8hd_fill_2
XFILLER_16_56 vgnd vpwr scs8hd_decap_6
XANTENNA__05__A _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_369 vpwr vgnd scs8hd_fill_2
XFILLER_0_575 vgnd vpwr scs8hd_decap_12
XFILLER_8_642 vgnd vpwr scs8hd_decap_12
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XFILLER_1_306 vgnd vpwr scs8hd_decap_12
XFILLER_14_947 vgnd vpwr scs8hd_decap_12
XFILLER_5_623 vgnd vpwr scs8hd_decap_12
XFILLER_9_428 vgnd vpwr scs8hd_decap_12
XFILLER_1_862 vpwr vgnd scs8hd_fill_2
XFILLER_4_26 vgnd vpwr scs8hd_decap_4
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_16_273 vgnd vpwr scs8hd_decap_6
XFILLER_1_1099 vgnd vpwr scs8hd_decap_12
XPHY_290 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_450 vgnd vpwr scs8hd_decap_8
XFILLER_8_483 vgnd vpwr scs8hd_decap_12
XFILLER_9_940 vgnd vpwr scs8hd_decap_12
XFILLER_11_928 vgnd vpwr scs8hd_decap_12
XFILLER_14_788 vgnd vpwr scs8hd_decap_12
XFILLER_13_232 vgnd vpwr scs8hd_decap_12
XFILLER_5_464 vgnd vpwr scs8hd_decap_12
XFILLER_6_910 vgnd vpwr scs8hd_decap_12
XFILLER_9_269 vgnd vpwr scs8hd_decap_12
XFILLER_10_983 vgnd vpwr scs8hd_decap_12
XFILLER_1_692 vgnd vpwr scs8hd_decap_12
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_9_781 vgnd vpwr scs8hd_decap_12
XFILLER_11_769 vgnd vpwr scs8hd_decap_12
XANTENNA__13__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_10_202 vgnd vpwr scs8hd_decap_12
XFILLER_2_434 vgnd vpwr scs8hd_decap_12
XFILLER_3_946 vgnd vpwr scs8hd_fill_1
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_762 vgnd vpwr scs8hd_fill_1
XFILLER_7_1050 vgnd vpwr scs8hd_decap_12
XFILLER_3_209 vpwr vgnd scs8hd_fill_2
XANTENNA__08__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_13_1099 vgnd vpwr scs8hd_decap_12
XFILLER_3_721 vgnd vpwr scs8hd_decap_8
XFILLER_7_537 vgnd vpwr scs8hd_decap_12
XFILLER_6_581 vgnd vpwr scs8hd_decap_12
XFILLER_9_1123 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_507 vgnd vpwr scs8hd_decap_12
XFILLER_0_757 vgnd vpwr scs8hd_decap_12
XANTENNA__10__B enable vgnd vpwr scs8hd_diode_2
XFILLER_16_614 vgnd vpwr scs8hd_decap_6
XFILLER_15_135 vgnd vpwr scs8hd_decap_12
XFILLER_12_886 vgnd vpwr scs8hd_decap_12
XFILLER_11_330 vgnd vpwr scs8hd_decap_12
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_562 vgnd vpwr scs8hd_decap_12
XFILLER_7_367 vgnd vpwr scs8hd_decap_12
XFILLER_4_1020 vgnd vpwr scs8hd_decap_12
XFILLER_14_190 vgnd vpwr scs8hd_decap_12
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XANTENNA__05__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_521 vgnd vpwr scs8hd_decap_6
XANTENNA__21__A gfpga_pad_GPIO_PAD[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_337 vgnd vpwr scs8hd_decap_12
XFILLER_5_838 vgnd vpwr scs8hd_decap_12
XFILLER_10_1069 vgnd vpwr scs8hd_decap_12
XFILLER_0_587 vpwr vgnd scs8hd_fill_2
XFILLER_16_466 vgnd vpwr scs8hd_decap_12
XFILLER_8_654 vgnd vpwr scs8hd_decap_12
XFILLER_11_171 vgnd vpwr scs8hd_decap_12
XFILLER_1_318 vgnd vpwr scs8hd_decap_12
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XFILLER_14_959 vgnd vpwr scs8hd_decap_12
XFILLER_13_403 vgnd vpwr scs8hd_decap_12
XANTENNA__16__A gfpga_pad_GPIO_PAD[5] vgnd vpwr scs8hd_diode_2
XFILLER_5_635 vgnd vpwr scs8hd_decap_3
XFILLER_1_830 vgnd vpwr scs8hd_decap_6
XFILLER_0_373 vgnd vpwr scs8hd_decap_12
XFILLER_4_178 vgnd vpwr scs8hd_decap_6
XFILLER_5_668 vgnd vpwr scs8hd_fill_1
XFILLER_16_230 vgnd vpwr scs8hd_decap_12
XFILLER_1_1001 vgnd vpwr scs8hd_decap_12
XPHY_291 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_952 vgnd vpwr scs8hd_decap_12
XFILLER_8_495 vgnd vpwr scs8hd_decap_12
XFILLER_2_605 vgnd vpwr scs8hd_decap_12
XFILLER_16_1086 vgnd vpwr scs8hd_decap_12
XFILLER_5_421 vgnd vpwr scs8hd_decap_6
XFILLER_5_476 vgnd vpwr scs8hd_decap_12
XFILLER_6_922 vgnd vpwr scs8hd_decap_12
XFILLER_6_944 vpwr vgnd scs8hd_fill_2
XFILLER_10_995 vgnd vpwr scs8hd_decap_12
XFILLER_3_903 vgnd vpwr scs8hd_decap_12
XANTENNA__13__B _14_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_708 vgnd vpwr scs8hd_decap_12
XFILLER_2_446 vgnd vpwr scs8hd_decap_12
XFILLER_14_520 vgnd vpwr scs8hd_decap_12
XFILLER_2_991 vgnd vpwr scs8hd_decap_12
XFILLER_7_1062 vgnd vpwr scs8hd_decap_12
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_807 vgnd vpwr scs8hd_decap_12
XFILLER_15_306 vgnd vpwr scs8hd_decap_12
XFILLER_13_1001 vgnd vpwr scs8hd_decap_12
XFILLER_11_501 vgnd vpwr scs8hd_decap_12
XFILLER_3_733 vgnd vpwr scs8hd_decap_12
XFILLER_2_276 vgnd vpwr scs8hd_decap_12
XFILLER_14_361 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_14_ logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[7] vgnd vpwr scs8hd_ebufn_1
XFILLER_6_593 vgnd vpwr scs8hd_decap_12
XFILLER_9_1135 vgnd vpwr scs8hd_decap_8
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__10__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_0_769 vgnd vpwr scs8hd_decap_6
XANTENNA__19__A gfpga_pad_GPIO_PAD[0] vgnd vpwr scs8hd_diode_2
XFILLER_15_147 vgnd vpwr scs8hd_decap_12
XFILLER_12_898 vgnd vpwr scs8hd_decap_12
XFILLER_11_342 vgnd vpwr scs8hd_decap_12
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XFILLER_7_379 vgnd vpwr scs8hd_decap_6
XFILLER_8_825 vgnd vpwr scs8hd_decap_12
XFILLER_3_574 vgnd vpwr scs8hd_decap_12
XFILLER_4_1032 vgnd vpwr scs8hd_decap_12
XFILLER_7_891 vgnd vpwr scs8hd_decap_12
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XFILLER_5_806 vgnd vpwr scs8hd_decap_12
XANTENNA__05__C address[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_349 vgnd vpwr scs8hd_decap_12
XFILLER_16_478 vgnd vpwr scs8hd_decap_12
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
XFILLER_8_666 vgnd vpwr scs8hd_decap_12
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_393 vgnd vpwr scs8hd_fill_1
XFILLER_6_1105 vgnd vpwr scs8hd_decap_12
XFILLER_13_415 vgnd vpwr scs8hd_decap_12
XFILLER_1_842 vgnd vpwr scs8hd_decap_12
XFILLER_0_385 vgnd vpwr scs8hd_decap_12
XFILLER_4_39 vgnd vpwr scs8hd_decap_12
XFILLER_16_242 vgnd vpwr scs8hd_decap_6
XFILLER_1_1013 vgnd vpwr scs8hd_decap_12
XPHY_292 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_964 vgnd vpwr scs8hd_decap_12
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XFILLER_11_1143 vgnd vpwr scs8hd_decap_3
XFILLER_2_617 vgnd vpwr scs8hd_decap_12
XFILLER_1_127 vpwr vgnd scs8hd_fill_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_16_1098 vgnd vpwr scs8hd_decap_12
XFILLER_6_934 vgnd vpwr scs8hd_decap_8
XFILLER_1_672 vgnd vpwr scs8hd_decap_12
XFILLER_9_794 vgnd vpwr scs8hd_decap_12
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XFILLER_8_1008 vgnd vpwr scs8hd_decap_12
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XANTENNA__13__C _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_532 vgnd vpwr scs8hd_decap_12
XFILLER_2_1130 vgnd vpwr scs8hd_decap_12
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_764 vgnd vpwr scs8hd_decap_12
XFILLER_7_1074 vgnd vpwr scs8hd_decap_12
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_819 vgnd vpwr scs8hd_decap_12
XFILLER_15_318 vgnd vpwr scs8hd_decap_12
XFILLER_13_1013 vgnd vpwr scs8hd_decap_12
XFILLER_11_513 vgnd vpwr scs8hd_decap_12
XFILLER_2_288 vgnd vpwr scs8hd_decap_12
XFILLER_3_745 vgnd vpwr scs8hd_decap_12
XFILLER_15_830 vgnd vpwr scs8hd_decap_12
XFILLER_14_373 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _13_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__10__D _09_/D vgnd vpwr scs8hd_diode_2
XFILLER_15_159 vgnd vpwr scs8hd_decap_12
XFILLER_12_800 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _07_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_354 vgnd vpwr scs8hd_decap_12
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XFILLER_8_837 vgnd vpwr scs8hd_decap_12
XFILLER_3_586 vgnd vpwr scs8hd_decap_12
XFILLER_4_1044 vgnd vpwr scs8hd_decap_12
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_129 vgnd vpwr scs8hd_decap_12
XANTENNA__05__D enable vgnd vpwr scs8hd_diode_2
XFILLER_14_1130 vgnd vpwr scs8hd_decap_12
XFILLER_5_818 vgnd vpwr scs8hd_decap_4
XFILLER_16_435 vgnd vpwr scs8hd_decap_12
XFILLER_4_884 vgnd vpwr scs8hd_fill_1
XFILLER_8_678 vgnd vpwr scs8hd_decap_12
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XFILLER_6_1117 vgnd vpwr scs8hd_decap_12
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_648 vpwr vgnd scs8hd_fill_2
XFILLER_0_397 vgnd vpwr scs8hd_decap_6
XFILLER_0_342 vgnd vpwr scs8hd_decap_12
XFILLER_1_1025 vgnd vpwr scs8hd_decap_12
XPHY_293 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_471 vgnd vpwr scs8hd_decap_12
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_670 vgnd vpwr scs8hd_fill_1
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_11_1111 vgnd vpwr scs8hd_decap_12
XFILLER_2_629 vgnd vpwr scs8hd_decap_12
XFILLER_14_703 vgnd vpwr scs8hd_decap_12
XFILLER_16_1055 vgnd vpwr scs8hd_decap_12
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_489 vgnd vpwr scs8hd_decap_12
XFILLER_1_684 vpwr vgnd scs8hd_fill_2
XANTENNA__13__D _09_/D vgnd vpwr scs8hd_diode_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XFILLER_2_459 vgnd vpwr scs8hd_decap_12
XFILLER_3_916 vgnd vpwr scs8hd_decap_12
XFILLER_3_949 vpwr vgnd scs8hd_fill_2
XFILLER_14_544 vgnd vpwr scs8hd_decap_12
XFILLER_2_1142 vgnd vpwr scs8hd_decap_4
XFILLER_5_231 vgnd vpwr scs8hd_decap_12
XFILLER_6_776 vgnd vpwr scs8hd_decap_12
XFILLER_7_1086 vgnd vpwr scs8hd_decap_12
XFILLER_13_1025 vgnd vpwr scs8hd_decap_12
XFILLER_11_525 vgnd vpwr scs8hd_decap_12
XFILLER_3_702 vgnd vpwr scs8hd_fill_1
XFILLER_3_757 vgnd vpwr scs8hd_decap_12
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XFILLER_15_842 vgnd vpwr scs8hd_decap_12
XFILLER_14_385 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_540 vgnd vpwr scs8hd_decap_3
XFILLER_12_812 vgnd vpwr scs8hd_decap_12
XFILLER_3_532 vgnd vpwr scs8hd_decap_12
XFILLER_8_849 vgnd vpwr scs8hd_decap_12
XFILLER_3_598 vgnd vpwr scs8hd_decap_8
XFILLER_15_672 vgnd vpwr scs8hd_decap_12
XFILLER_4_1056 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_14_1142 vgnd vpwr scs8hd_decap_4
XFILLER_16_447 vgnd vpwr scs8hd_decap_12
XFILLER_12_642 vgnd vpwr scs8hd_decap_12
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_373 vpwr vgnd scs8hd_fill_2
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _14_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_428 vgnd vpwr scs8hd_decap_12
XFILLER_1_866 vgnd vpwr scs8hd_decap_12
XFILLER_1_855 vgnd vpwr scs8hd_decap_3
XFILLER_0_354 vgnd vpwr scs8hd_decap_12
XFILLER_16_211 vgnd vpwr scs8hd_decap_6
XFILLER_13_940 vgnd vpwr scs8hd_decap_12
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_294 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_483 vgnd vpwr scs8hd_decap_12
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_977 vgnd vpwr scs8hd_decap_12
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_11_1123 vgnd vpwr scs8hd_decap_12
XFILLER_14_715 vgnd vpwr scs8hd_decap_12
XFILLER_16_1067 vgnd vpwr scs8hd_decap_12
XFILLER_13_269 vgnd vpwr scs8hd_decap_12
XFILLER_6_947 vgnd vpwr scs8hd_decap_12
XFILLER_10_910 vgnd vpwr scs8hd_decap_12
XFILLER_13_781 vgnd vpwr scs8hd_decap_12
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
XFILLER_3_928 vgnd vpwr scs8hd_decap_12
XFILLER_14_556 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_243 vgnd vpwr scs8hd_fill_1
XFILLER_6_700 vpwr vgnd scs8hd_fill_2
XFILLER_6_744 vgnd vpwr scs8hd_decap_12
XFILLER_6_788 vgnd vpwr scs8hd_decap_12
XFILLER_10_751 vgnd vpwr scs8hd_decap_12
XFILLER_11_537 vgnd vpwr scs8hd_decap_12
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_769 vgnd vpwr scs8hd_decap_12
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_10_581 vgnd vpwr scs8hd_decap_12
XFILLER_6_552 vgnd vpwr scs8hd_decap_12
XFILLER_12_1081 vgnd vpwr scs8hd_decap_12
XFILLER_11_367 vgnd vpwr scs8hd_decap_12
XFILLER_3_544 vgnd vpwr scs8hd_decap_4
XFILLER_15_684 vgnd vpwr scs8hd_decap_12
XFILLER_6_393 vpwr vgnd scs8hd_fill_2
XFILLER_16_459 vgnd vpwr scs8hd_decap_6
XFILLER_16_404 vgnd vpwr scs8hd_decap_12
XFILLER_12_654 vgnd vpwr scs8hd_decap_12
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XFILLER_3_330 vgnd vpwr scs8hd_decap_12
XFILLER_3_396 vpwr vgnd scs8hd_fill_2
XFILLER_4_831 vgnd vpwr scs8hd_decap_12
XFILLER_4_886 vgnd vpwr scs8hd_decap_12
XFILLER_16_993 vgnd vpwr scs8hd_decap_12
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XFILLER_1_878 vgnd vpwr scs8hd_decap_12
XFILLER_0_311 vgnd vpwr scs8hd_decap_12
XFILLER_1_1038 vgnd vpwr scs8hd_decap_12
XFILLER_0_366 vgnd vpwr scs8hd_decap_6
XFILLER_13_952 vgnd vpwr scs8hd_decap_12
XPHY_295 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_495 vgnd vpwr scs8hd_decap_12
XFILLER_9_989 vgnd vpwr scs8hd_decap_12
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_11_1135 vgnd vpwr scs8hd_decap_8
XFILLER_16_1024 vgnd vpwr scs8hd_decap_12
XFILLER_14_727 vgnd vpwr scs8hd_decap_12
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
XFILLER_16_1079 vgnd vpwr scs8hd_decap_6
XFILLER_6_959 vgnd vpwr scs8hd_decap_12
XFILLER_10_922 vgnd vpwr scs8hd_decap_12
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_9_720 vgnd vpwr scs8hd_decap_12
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_11_708 vgnd vpwr scs8hd_decap_12
XFILLER_14_568 vgnd vpwr scs8hd_decap_12
XFILLER_6_756 vgnd vpwr scs8hd_decap_6
XFILLER_7_1099 vgnd vpwr scs8hd_decap_12
XFILLER_9_550 vgnd vpwr scs8hd_decap_12
XFILLER_13_1038 vgnd vpwr scs8hd_decap_12
XFILLER_15_855 vgnd vpwr scs8hd_decap_12
XPHY_60 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_14_398 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_520 vgnd vpwr scs8hd_decap_12
XFILLER_10_593 vgnd vpwr scs8hd_decap_12
XFILLER_6_564 vgnd vpwr scs8hd_decap_12
XFILLER_2_64 vgnd vpwr scs8hd_decap_12
XFILLER_12_1093 vgnd vpwr scs8hd_decap_12
XFILLER_9_391 vgnd vpwr scs8hd_decap_12
XFILLER_0_718 vpwr vgnd scs8hd_fill_2
XFILLER_0_707 vgnd vpwr scs8hd_decap_6
XFILLER_12_825 vgnd vpwr scs8hd_decap_12
XFILLER_11_379 vgnd vpwr scs8hd_decap_12
XFILLER_7_306 vgnd vpwr scs8hd_decap_12
XFILLER_3_501 vgnd vpwr scs8hd_decap_12
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XFILLER_4_1069 vgnd vpwr scs8hd_decap_12
XFILLER_15_696 vgnd vpwr scs8hd_decap_12
XFILLER_11_891 vgnd vpwr scs8hd_decap_12
XFILLER_6_361 vgnd vpwr scs8hd_decap_12
XFILLER_10_1008 vgnd vpwr scs8hd_decap_12
XFILLER_0_559 vgnd vpwr scs8hd_decap_8
XFILLER_16_416 vgnd vpwr scs8hd_decap_12
XFILLER_11_110 vgnd vpwr scs8hd_decap_12
XFILLER_12_666 vgnd vpwr scs8hd_decap_12
XFILLER_4_843 vpwr vgnd scs8hd_fill_2
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
XFILLER_3_342 vgnd vpwr scs8hd_decap_12
XFILLER_4_898 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_0_ logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[0] vgnd vpwr scs8hd_ebufn_1
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _07_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XFILLER_0_323 vgnd vpwr scs8hd_decap_12
XFILLER_13_964 vgnd vpwr scs8hd_decap_12
XPHY_296 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_673 vgnd vpwr scs8hd_decap_12
XFILLER_16_1036 vgnd vpwr scs8hd_decap_12
XFILLER_14_739 vgnd vpwr scs8hd_decap_12
XFILLER_10_934 vgnd vpwr scs8hd_decap_12
XFILLER_13_794 vgnd vpwr scs8hd_decap_12
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_10_764 vgnd vpwr scs8hd_decap_12
XFILLER_1_440 vgnd vpwr scs8hd_decap_12
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_7_1001 vgnd vpwr scs8hd_decap_12
XFILLER_9_562 vgnd vpwr scs8hd_decap_12
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_3_705 vpwr vgnd scs8hd_fill_2
XFILLER_15_867 vgnd vpwr scs8hd_decap_12
XFILLER_14_300 vgnd vpwr scs8hd_decap_12
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_61 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_532 vgnd vpwr scs8hd_decap_8
XFILLER_6_576 vgnd vpwr scs8hd_decap_4
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_2_76 vgnd vpwr scs8hd_decap_12
XFILLER_12_837 vgnd vpwr scs8hd_decap_12
XFILLER_7_318 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vpwr vgnd scs8hd_fill_2
XFILLER_3_513 vgnd vpwr scs8hd_decap_12
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_14_141 vgnd vpwr scs8hd_decap_12
XFILLER_6_373 vgnd vpwr scs8hd_decap_12
XFILLER_16_428 vgnd vpwr scs8hd_decap_6
XFILLER_12_678 vgnd vpwr scs8hd_decap_12
XFILLER_8_605 vgnd vpwr scs8hd_decap_12
XFILLER_3_354 vgnd vpwr scs8hd_decap_12
XFILLER_4_800 vgnd vpwr scs8hd_decap_12
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
XFILLER_16_962 vgnd vpwr scs8hd_decap_12
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_0_335 vgnd vpwr scs8hd_decap_6
XFILLER_5_1143 vgnd vpwr scs8hd_decap_3
XPHY_297 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_286 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_402 vgnd vpwr scs8hd_decap_12
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_903 vgnd vpwr scs8hd_decap_12
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XFILLER_4_685 vgnd vpwr scs8hd_decap_12
XFILLER_16_1048 vgnd vpwr scs8hd_decap_6
XFILLER_1_611 vgnd vpwr scs8hd_decap_12
XFILLER_1_688 vpwr vgnd scs8hd_fill_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_8_276 vgnd vpwr scs8hd_decap_12
XFILLER_9_733 vgnd vpwr scs8hd_decap_12
XFILLER_4_471 vgnd vpwr scs8hd_decap_12
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_6_703 vgnd vpwr scs8hd_decap_12
XFILLER_10_776 vgnd vpwr scs8hd_decap_12
XFILLER_1_452 vgnd vpwr scs8hd_decap_12
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_7_1013 vgnd vpwr scs8hd_decap_12
XFILLER_9_574 vgnd vpwr scs8hd_decap_12
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XFILLER_4_7 vgnd vpwr scs8hd_decap_4
XFILLER_15_879 vgnd vpwr scs8hd_decap_12
XFILLER_14_312 vgnd vpwr scs8hd_decap_12
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_62 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_51 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_2_88 vgnd vpwr scs8hd_decap_4
XFILLER_12_849 vgnd vpwr scs8hd_decap_12
XFILLER_3_525 vgnd vpwr scs8hd_decap_4
XFILLER_8_1130 vgnd vpwr scs8hd_decap_12
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
XFILLER_7_831 vpwr vgnd scs8hd_fill_2
XFILLER_6_385 vgnd vpwr scs8hd_decap_8
XFILLER_7_853 vgnd vpwr scs8hd_fill_1
XFILLER_0_528 vgnd vpwr scs8hd_decap_12
XFILLER_8_617 vgnd vpwr scs8hd_decap_12
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
XFILLER_3_377 vgnd vpwr scs8hd_decap_12
XFILLER_4_812 vgnd vpwr scs8hd_decap_12
XFILLER_4_856 vgnd vpwr scs8hd_decap_12
XFILLER_16_974 vgnd vpwr scs8hd_decap_12
XFILLER_15_440 vgnd vpwr scs8hd_decap_12
XFILLER_7_672 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
X_19_ gfpga_pad_GPIO_PAD[0] bottom_width_0_height_0__pin_1_ vgnd vpwr scs8hd_buf_2
XFILLER_5_1111 vgnd vpwr scs8hd_decap_12
XFILLER_12_410 vgnd vpwr scs8hd_decap_12
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_977 vgnd vpwr scs8hd_decap_12
XPHY_298 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_287 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_414 vgnd vpwr scs8hd_decap_12
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_196 vgnd vpwr scs8hd_decap_8
XFILLER_4_642 vgnd vpwr scs8hd_decap_12
XFILLER_4_697 vgnd vpwr scs8hd_decap_4
XFILLER_0_881 vgnd vpwr scs8hd_decap_12
XFILLER_15_281 vgnd vpwr scs8hd_decap_12
XFILLER_16_1005 vgnd vpwr scs8hd_decap_12
XFILLER_5_417 vpwr vgnd scs8hd_fill_2
XFILLER_5_428 vgnd vpwr scs8hd_decap_12
XFILLER_10_947 vgnd vpwr scs8hd_decap_12
XFILLER_1_623 vgnd vpwr scs8hd_decap_12
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XFILLER_9_745 vgnd vpwr scs8hd_decap_12
XFILLER_5_951 vgnd vpwr scs8hd_decap_12
XFILLER_8_288 vgnd vpwr scs8hd_decap_12
XFILLER_4_483 vgnd vpwr scs8hd_decap_12
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_16_590 vgnd vpwr scs8hd_decap_12
XFILLER_5_269 vgnd vpwr scs8hd_decap_12
XFILLER_6_715 vgnd vpwr scs8hd_decap_12
XFILLER_10_788 vgnd vpwr scs8hd_decap_12
XFILLER_1_464 vgnd vpwr scs8hd_decap_12
XFILLER_2_910 vgnd vpwr scs8hd_decap_12
XFILLER_7_1025 vgnd vpwr scs8hd_decap_12
XFILLER_9_586 vgnd vpwr scs8hd_decap_12
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XFILLER_3_729 vgnd vpwr scs8hd_decap_3
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_14_324 vgnd vpwr scs8hd_decap_12
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_63 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_52 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_751 vgnd vpwr scs8hd_decap_12
XFILLER_2_56 vgnd vpwr scs8hd_decap_6
XFILLER_3_548 vgnd vpwr scs8hd_fill_1
XFILLER_11_98 vgnd vpwr scs8hd_decap_12
XFILLER_4_1006 vgnd vpwr scs8hd_fill_1
XFILLER_8_1142 vgnd vpwr scs8hd_decap_4
XFILLER_15_611 vgnd vpwr scs8hd_decap_12
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
XFILLER_2_581 vgnd vpwr scs8hd_decap_12
XFILLER_3_1050 vgnd vpwr scs8hd_decap_12
XFILLER_8_629 vgnd vpwr scs8hd_decap_12
XFILLER_11_135 vgnd vpwr scs8hd_decap_12
XFILLER_3_367 vgnd vpwr scs8hd_decap_4
XFILLER_3_389 vgnd vpwr scs8hd_decap_4
XFILLER_4_868 vgnd vpwr scs8hd_decap_12
XFILLER_16_986 vgnd vpwr scs8hd_decap_6
XFILLER_16_931 vgnd vpwr scs8hd_decap_12
XFILLER_15_452 vgnd vpwr scs8hd_decap_12
XFILLER_7_684 vgnd vpwr scs8hd_decap_12
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_190 vgnd vpwr scs8hd_decap_12
X_18_ gfpga_pad_GPIO_PAD[7] bottom_width_0_height_0__pin_15_ vgnd vpwr scs8hd_buf_2
XFILLER_1_838 vpwr vgnd scs8hd_fill_2
XFILLER_0_304 vgnd vpwr scs8hd_decap_6
XFILLER_5_1123 vgnd vpwr scs8hd_decap_12
XFILLER_16_249 vgnd vpwr scs8hd_decap_12
XFILLER_12_422 vgnd vpwr scs8hd_decap_12
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_916 vgnd vpwr scs8hd_decap_12
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_989 vgnd vpwr scs8hd_decap_12
XPHY_299 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_288 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_426 vgnd vpwr scs8hd_decap_12
XFILLER_8_459 vgnd vpwr scs8hd_decap_12
XFILLER_0_893 vgnd vpwr scs8hd_decap_6
XFILLER_4_654 vgnd vpwr scs8hd_decap_12
XFILLER_15_293 vgnd vpwr scs8hd_decap_12
XFILLER_8_971 vgnd vpwr scs8hd_decap_12
XFILLER_16_1017 vgnd vpwr scs8hd_decap_6
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_1086 vgnd vpwr scs8hd_decap_12
XFILLER_10_959 vgnd vpwr scs8hd_decap_12
XFILLER_1_635 vgnd vpwr scs8hd_decap_12
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_13_720 vgnd vpwr scs8hd_decap_12
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XFILLER_9_757 vgnd vpwr scs8hd_decap_12
XFILLER_4_451 vgnd vpwr scs8hd_decap_6
XFILLER_4_495 vgnd vpwr scs8hd_decap_12
XFILLER_5_23 vgnd vpwr scs8hd_decap_12
XFILLER_5_963 vgnd vpwr scs8hd_decap_12
XFILLER_15_1050 vgnd vpwr scs8hd_decap_12
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_1_410 vgnd vpwr scs8hd_decap_12
XFILLER_2_922 vgnd vpwr scs8hd_decap_12
XFILLER_6_727 vgnd vpwr scs8hd_decap_8
XFILLER_1_476 vgnd vpwr scs8hd_decap_12
XFILLER_2_955 vgnd vpwr scs8hd_decap_12
XFILLER_13_550 vgnd vpwr scs8hd_decap_12
XFILLER_9_598 vgnd vpwr scs8hd_decap_12
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_53 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_42 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_1081 vgnd vpwr scs8hd_decap_12
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_10_520 vgnd vpwr scs8hd_decap_12
XFILLER_1_273 vgnd vpwr scs8hd_decap_12
XFILLER_13_391 vgnd vpwr scs8hd_decap_12
XFILLER_12_1020 vgnd vpwr scs8hd_decap_12
XFILLER_11_306 vgnd vpwr scs8hd_decap_12
XFILLER_15_623 vgnd vpwr scs8hd_decap_12
XFILLER_14_166 vgnd vpwr scs8hd_decap_12
XFILLER_7_855 vgnd vpwr scs8hd_decap_12
XFILLER_10_361 vgnd vpwr scs8hd_decap_12
XFILLER_2_593 vgnd vpwr scs8hd_decap_12
XFILLER_3_1062 vgnd vpwr scs8hd_decap_12
XFILLER_4_825 vgnd vpwr scs8hd_decap_4
XFILLER_11_147 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_16_943 vgnd vpwr scs8hd_decap_12
XFILLER_15_464 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
XFILLER_7_696 vgnd vpwr scs8hd_decap_12
XFILLER_3_891 vgnd vpwr scs8hd_decap_12
X_17_ gfpga_pad_GPIO_PAD[6] bottom_width_0_height_0__pin_13_ vgnd vpwr scs8hd_buf_2
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_806 vgnd vpwr scs8hd_decap_12
XFILLER_5_1135 vgnd vpwr scs8hd_decap_8
XPHY_289 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_434 vgnd vpwr scs8hd_decap_12
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_928 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_666 vgnd vpwr scs8hd_decap_4
XFILLER_8_438 vgnd vpwr scs8hd_decap_12
XFILLER_0_850 vgnd vpwr scs8hd_decap_12
XFILLER_8_983 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _09_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_1098 vgnd vpwr scs8hd_decap_12
XFILLER_1_647 vgnd vpwr scs8hd_decap_12
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XFILLER_9_769 vgnd vpwr scs8hd_decap_12
XFILLER_5_975 vgnd vpwr scs8hd_fill_1
XFILLER_15_1062 vgnd vpwr scs8hd_decap_12
XFILLER_14_507 vgnd vpwr scs8hd_decap_12
XFILLER_2_1105 vgnd vpwr scs8hd_decap_12
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_422 vgnd vpwr scs8hd_decap_4
XFILLER_2_934 vgnd vpwr scs8hd_decap_12
XFILLER_2_967 vgnd vpwr scs8hd_decap_12
XFILLER_7_1038 vgnd vpwr scs8hd_decap_12
XFILLER_13_562 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_2_ logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[1] vgnd vpwr scs8hd_ebufn_1
XFILLER_5_761 vgnd vpwr scs8hd_decap_12
XFILLER_5_794 vgnd vpwr scs8hd_decap_12
XFILLER_3_709 vgnd vpwr scs8hd_decap_12
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_14_337 vgnd vpwr scs8hd_decap_12
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_54 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_43 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XFILLER_6_1093 vgnd vpwr scs8hd_decap_12
XPHY_21 vgnd vpwr scs8hd_decap_3
XFILLER_10_532 vgnd vpwr scs8hd_decap_12
XFILLER_1_285 vgnd vpwr scs8hd_decap_12
XFILLER_2_764 vgnd vpwr scs8hd_decap_12
XFILLER_9_330 vgnd vpwr scs8hd_decap_12
XFILLER_12_1032 vgnd vpwr scs8hd_decap_12
XFILLER_11_318 vgnd vpwr scs8hd_decap_12
XFILLER_2_7 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _14_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_1008 vgnd vpwr scs8hd_decap_12
XFILLER_15_635 vgnd vpwr scs8hd_decap_12
XFILLER_14_178 vgnd vpwr scs8hd_decap_12
XFILLER_11_830 vgnd vpwr scs8hd_decap_12
XFILLER_6_300 vgnd vpwr scs8hd_decap_12
XFILLER_7_867 vgnd vpwr scs8hd_decap_12
XFILLER_10_373 vgnd vpwr scs8hd_decap_12
XFILLER_14_1105 vgnd vpwr scs8hd_decap_12
XFILLER_14_690 vgnd vpwr scs8hd_decap_12
XFILLER_9_171 vgnd vpwr scs8hd_decap_12
XFILLER_0_509 vgnd vpwr scs8hd_decap_12
XFILLER_12_605 vgnd vpwr scs8hd_decap_12
XFILLER_3_1074 vgnd vpwr scs8hd_decap_12
XFILLER_11_159 vgnd vpwr scs8hd_decap_12
XFILLER_16_955 vgnd vpwr scs8hd_decap_6
XFILLER_16_900 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_12_ vgnd vpwr scs8hd_diode_2
XFILLER_15_476 vgnd vpwr scs8hd_decap_12
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
X_16_ gfpga_pad_GPIO_PAD[5] bottom_width_0_height_0__pin_11_ vgnd vpwr scs8hd_buf_2
XFILLER_1_818 vgnd vpwr scs8hd_decap_12
XFILLER_16_218 vgnd vpwr scs8hd_decap_12
XFILLER_13_903 vgnd vpwr scs8hd_decap_12
XFILLER_12_446 vgnd vpwr scs8hd_decap_12
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_862 vgnd vpwr scs8hd_decap_6
XFILLER_8_995 vgnd vpwr scs8hd_decap_12
XFILLER_0_1055 vgnd vpwr scs8hd_decap_12
XFILLER_1_659 vgnd vpwr scs8hd_decap_12
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_13_733 vgnd vpwr scs8hd_decap_12
XFILLER_12_276 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_1130 vgnd vpwr scs8hd_decap_12
XFILLER_16_571 vgnd vpwr scs8hd_decap_12
XFILLER_15_1074 vgnd vpwr scs8hd_decap_12
XFILLER_2_1117 vgnd vpwr scs8hd_decap_12
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_703 vgnd vpwr scs8hd_decap_12
XFILLER_2_979 vgnd vpwr scs8hd_decap_12
XFILLER_1_489 vgnd vpwr scs8hd_decap_12
XFILLER_13_574 vgnd vpwr scs8hd_decap_12
XFILLER_9_501 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _15_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_773 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_8_ vgnd vpwr scs8hd_diode_2
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_15_806 vgnd vpwr scs8hd_decap_12
XFILLER_14_349 vgnd vpwr scs8hd_decap_12
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_55 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_44 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XFILLER_10_544 vgnd vpwr scs8hd_decap_12
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_1_297 vgnd vpwr scs8hd_decap_8
XFILLER_2_776 vgnd vpwr scs8hd_decap_12
XFILLER_14_861 vgnd vpwr scs8hd_decap_12
XFILLER_9_342 vgnd vpwr scs8hd_decap_12
XFILLER_12_1044 vgnd vpwr scs8hd_decap_12
XFILLER_3_529 vgnd vpwr scs8hd_fill_1
XFILLER_15_647 vgnd vpwr scs8hd_decap_12
XFILLER_11_842 vgnd vpwr scs8hd_decap_12
XFILLER_6_312 vgnd vpwr scs8hd_decap_12
XFILLER_7_835 vgnd vpwr scs8hd_decap_12
XFILLER_7_879 vgnd vpwr scs8hd_decap_12
XFILLER_10_385 vgnd vpwr scs8hd_decap_12
XFILLER_14_1117 vgnd vpwr scs8hd_decap_12
XFILLER_3_1086 vgnd vpwr scs8hd_decap_12
XFILLER_12_617 vgnd vpwr scs8hd_decap_12
XANTENNA__11__A enable vgnd vpwr scs8hd_diode_2
XFILLER_16_912 vgnd vpwr scs8hd_decap_12
XFILLER_11_672 vgnd vpwr scs8hd_decap_12
X_15_ address[1] _14_/B _04_/X address[2] _15_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_4_ vgnd vpwr scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__06__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_7_440 vgnd vpwr scs8hd_decap_12
XFILLER_0_1067 vgnd vpwr scs8hd_decap_12
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_13_745 vgnd vpwr scs8hd_decap_12
XFILLER_12_288 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_1142 vgnd vpwr scs8hd_decap_4
XFILLER_5_48 vgnd vpwr scs8hd_decap_12
XFILLER_5_977 vgnd vpwr scs8hd_decap_12
XFILLER_16_583 vgnd vpwr scs8hd_decap_6
XFILLER_15_1086 vgnd vpwr scs8hd_decap_12
XFILLER_7_281 vgnd vpwr scs8hd_decap_12
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_5_207 vgnd vpwr scs8hd_decap_12
XFILLER_10_715 vgnd vpwr scs8hd_decap_12
XFILLER_13_586 vgnd vpwr scs8hd_decap_12
XFILLER_9_513 vgnd vpwr scs8hd_decap_12
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_785 vgnd vpwr scs8hd_decap_8
XFILLER_0_490 vgnd vpwr scs8hd_decap_6
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XFILLER_15_818 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_56 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_34 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_45 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__14__A _06_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_556 vgnd vpwr scs8hd_decap_12
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_2_788 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_0_ vgnd vpwr scs8hd_diode_2
XFILLER_14_873 vgnd vpwr scs8hd_decap_12
XFILLER_9_354 vgnd vpwr scs8hd_decap_12
XFILLER_12_1056 vgnd vpwr scs8hd_decap_12
XFILLER_15_659 vgnd vpwr scs8hd_decap_12
XANTENNA__09__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_6_324 vgnd vpwr scs8hd_decap_12
XFILLER_7_847 vgnd vpwr scs8hd_decap_6
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_70 vgnd vpwr scs8hd_decap_12
XFILLER_12_629 vgnd vpwr scs8hd_decap_12
XFILLER_16_924 vgnd vpwr scs8hd_decap_6
XFILLER_15_489 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_684 vgnd vpwr scs8hd_decap_12
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XFILLER_7_611 vgnd vpwr scs8hd_decap_12
X_14_ _06_/Y _14_/B _04_/X address[2] _14_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_916 vgnd vpwr scs8hd_decap_12
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_459 vgnd vpwr scs8hd_decap_12
XANTENNA__22__A gfpga_pad_GPIO_PAD[3] vgnd vpwr scs8hd_diode_2
XFILLER_0_831 vgnd vpwr scs8hd_decap_6
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
XFILLER_16_776 vgnd vpwr scs8hd_decap_12
XFILLER_12_971 vgnd vpwr scs8hd_decap_12
XFILLER_7_452 vgnd vpwr scs8hd_decap_12
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XFILLER_0_1079 vgnd vpwr scs8hd_decap_6
XFILLER_0_1024 vgnd vpwr scs8hd_decap_12
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XANTENNA__17__A gfpga_pad_GPIO_PAD[6] vgnd vpwr scs8hd_diode_2
XFILLER_13_757 vgnd vpwr scs8hd_decap_12
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_989 vgnd vpwr scs8hd_decap_12
XFILLER_0_683 vgnd vpwr scs8hd_decap_12
XFILLER_16_540 vgnd vpwr scs8hd_decap_12
XFILLER_7_293 vgnd vpwr scs8hd_decap_12
XFILLER_10_727 vgnd vpwr scs8hd_decap_12
XFILLER_5_219 vgnd vpwr scs8hd_decap_12
XFILLER_13_598 vgnd vpwr scs8hd_decap_12
XFILLER_9_525 vgnd vpwr scs8hd_decap_12
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_35 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_57 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__14__B _14_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_568 vgnd vpwr scs8hd_decap_12
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_550 vgnd vpwr scs8hd_decap_12
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XANTENNA__09__B enable vgnd vpwr scs8hd_diode_2
XFILLER_11_855 vgnd vpwr scs8hd_decap_12
XFILLER_7_826 vpwr vgnd scs8hd_fill_2
XFILLER_10_398 vgnd vpwr scs8hd_decap_12
XFILLER_2_520 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_82 vgnd vpwr scs8hd_decap_12
XFILLER_3_1099 vgnd vpwr scs8hd_decap_12
XFILLER_3_306 vgnd vpwr scs8hd_decap_12
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XFILLER_11_696 vgnd vpwr scs8hd_decap_12
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_7_623 vgnd vpwr scs8hd_decap_12
XFILLER_2_361 vgnd vpwr scs8hd_decap_12
XFILLER_3_851 vgnd vpwr scs8hd_decap_3
X_13_ address[1] _14_/B _04_/X _09_/D _13_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_928 vgnd vpwr scs8hd_decap_12
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _09_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_788 vgnd vpwr scs8hd_decap_12
XFILLER_12_983 vgnd vpwr scs8hd_decap_12
XFILLER_8_910 vgnd vpwr scs8hd_decap_12
XFILLER_7_464 vgnd vpwr scs8hd_decap_12
XFILLER_0_1036 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_1_607 vgnd vpwr scs8hd_decap_3
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_9_1050 vgnd vpwr scs8hd_decap_12
XFILLER_13_769 vgnd vpwr scs8hd_decap_12
XFILLER_12_202 vgnd vpwr scs8hd_decap_12
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XFILLER_0_695 vgnd vpwr scs8hd_decap_12
XFILLER_16_552 vgnd vpwr scs8hd_decap_6
XFILLER_15_1099 vgnd vpwr scs8hd_decap_12
XFILLER_8_751 vgnd vpwr scs8hd_decap_12
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_739 vgnd vpwr scs8hd_decap_12
XFILLER_1_426 vgnd vpwr scs8hd_fill_1
XFILLER_9_537 vgnd vpwr scs8hd_decap_12
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_581 vgnd vpwr scs8hd_decap_12
XFILLER_6_1020 vgnd vpwr scs8hd_decap_12
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_58 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_47 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_36 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XANTENNA__14__C _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_507 vgnd vpwr scs8hd_decap_12
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_14_886 vgnd vpwr scs8hd_decap_12
XFILLER_13_330 vgnd vpwr scs8hd_decap_12
XFILLER_12_1069 vgnd vpwr scs8hd_decap_12
XFILLER_5_562 vgnd vpwr scs8hd_decap_12
XFILLER_9_367 vgnd vpwr scs8hd_decap_12
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XANTENNA__09__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_300 vgnd vpwr scs8hd_decap_12
XFILLER_11_867 vgnd vpwr scs8hd_decap_12
XFILLER_6_337 vgnd vpwr scs8hd_decap_12
XFILLER_2_565 vgnd vpwr scs8hd_decap_12
XFILLER_2_532 vgnd vpwr scs8hd_decap_12
XFILLER_13_171 vgnd vpwr scs8hd_decap_12
XFILLER_5_392 vpwr vgnd scs8hd_fill_2
XFILLER_3_94 vgnd vpwr scs8hd_decap_12
XFILLER_3_1001 vgnd vpwr scs8hd_decap_12
XFILLER_3_318 vgnd vpwr scs8hd_decap_12
XFILLER_15_403 vgnd vpwr scs8hd_decap_12
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
XFILLER_3_830 vgnd vpwr scs8hd_decap_12
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_635 vgnd vpwr scs8hd_decap_12
XFILLER_2_373 vgnd vpwr scs8hd_decap_6
X_12_ _06_/Y _14_/B _04_/X _09_/D _12_/Y vgnd vpwr scs8hd_nor4_4
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_4_ logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[2] vgnd vpwr scs8hd_ebufn_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
XFILLER_4_605 vgnd vpwr scs8hd_fill_1
XFILLER_0_800 vgnd vpwr scs8hd_decap_6
XFILLER_16_745 vgnd vpwr scs8hd_decap_12
XFILLER_12_995 vgnd vpwr scs8hd_decap_12
XFILLER_7_476 vgnd vpwr scs8hd_decap_12
XFILLER_8_922 vgnd vpwr scs8hd_decap_12
XFILLER_0_1048 vgnd vpwr scs8hd_decap_6
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XFILLER_9_1062 vgnd vpwr scs8hd_decap_12
XFILLER_5_903 vgnd vpwr scs8hd_decap_12
XFILLER_9_708 vgnd vpwr scs8hd_decap_12
XFILLER_4_457 vgnd vpwr scs8hd_fill_1
XFILLER_0_652 vgnd vpwr scs8hd_decap_12
XFILLER_15_1001 vgnd vpwr scs8hd_decap_12
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_501 vgnd vpwr scs8hd_decap_12
XFILLER_4_210 vgnd vpwr scs8hd_decap_4
XFILLER_5_733 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_decap_12
XFILLER_1_1143 vgnd vpwr scs8hd_decap_3
XFILLER_8_593 vgnd vpwr scs8hd_decap_12
XFILLER_6_1032 vgnd vpwr scs8hd_decap_12
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_48 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_37 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_15 vgnd vpwr scs8hd_decap_3
XANTENNA__14__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_19 vgnd vpwr scs8hd_decap_12
XFILLER_1_257 vgnd vpwr scs8hd_decap_8
XFILLER_2_703 vgnd vpwr scs8hd_decap_12
XFILLER_14_898 vgnd vpwr scs8hd_decap_12
XFILLER_13_342 vgnd vpwr scs8hd_decap_12
XFILLER_5_574 vgnd vpwr scs8hd_decap_12
XFILLER_9_379 vgnd vpwr scs8hd_decap_12
XFILLER_16_180 vgnd vpwr scs8hd_decap_6
XFILLER_9_891 vgnd vpwr scs8hd_decap_12
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XFILLER_8_1105 vgnd vpwr scs8hd_decap_12
XANTENNA__09__D _09_/D vgnd vpwr scs8hd_diode_2
XFILLER_14_117 vgnd vpwr scs8hd_decap_12
XFILLER_7_806 vgnd vpwr scs8hd_decap_12
XFILLER_10_312 vgnd vpwr scs8hd_decap_12
XFILLER_11_879 vgnd vpwr scs8hd_decap_12
XFILLER_6_349 vgnd vpwr scs8hd_decap_12
XFILLER_2_577 vgnd vpwr scs8hd_decap_3
XFILLER_2_544 vgnd vpwr scs8hd_decap_12
XFILLER_9_110 vgnd vpwr scs8hd_decap_12
XFILLER_3_1013 vgnd vpwr scs8hd_decap_12
XFILLER_15_415 vgnd vpwr scs8hd_decap_12
XFILLER_13_1143 vgnd vpwr scs8hd_decap_3
XFILLER_7_647 vgnd vpwr scs8hd_decap_12
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
XFILLER_3_842 vgnd vpwr scs8hd_decap_3
XFILLER_2_396 vgnd vpwr scs8hd_fill_1
X_11_ enable _14_/B vgnd vpwr scs8hd_inv_8
XFILLER_6_680 vgnd vpwr scs8hd_decap_12
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_4_617 vgnd vpwr scs8hd_decap_12
XFILLER_16_757 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
XFILLER_11_440 vgnd vpwr scs8hd_decap_12
XFILLER_8_934 vgnd vpwr scs8hd_decap_12
XFILLER_3_672 vgnd vpwr scs8hd_decap_12
XFILLER_0_1005 vgnd vpwr scs8hd_decap_12
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_4_1130 vgnd vpwr scs8hd_decap_12
XFILLER_9_1074 vgnd vpwr scs8hd_decap_12
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_0_664 vgnd vpwr scs8hd_decap_12
XFILLER_16_521 vgnd vpwr scs8hd_decap_6
XFILLER_15_1013 vgnd vpwr scs8hd_decap_12
XFILLER_11_281 vgnd vpwr scs8hd_decap_12
XFILLER_4_970 vgnd vpwr scs8hd_decap_12
XFILLER_8_764 vgnd vpwr scs8hd_decap_12
XFILLER_1_428 vgnd vpwr scs8hd_decap_12
XFILLER_13_513 vgnd vpwr scs8hd_decap_12
XFILLER_1_940 vgnd vpwr scs8hd_decap_3
XFILLER_4_288 vgnd vpwr scs8hd_decap_12
XFILLER_16_373 vgnd vpwr scs8hd_decap_12
XFILLER_1_1111 vgnd vpwr scs8hd_decap_12
XFILLER_6_1044 vgnd vpwr scs8hd_decap_12
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_38 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_16 vgnd vpwr scs8hd_decap_3
XFILLER_2_715 vgnd vpwr scs8hd_decap_12
XFILLER_1_269 vpwr vgnd scs8hd_fill_2
XFILLER_14_800 vgnd vpwr scs8hd_decap_12
XFILLER_16_1141 vgnd vpwr scs8hd_decap_4
XFILLER_13_354 vgnd vpwr scs8hd_decap_12
XFILLER_5_586 vgnd vpwr scs8hd_decap_12
XFILLER_1_781 vgnd vpwr scs8hd_decap_12
XFILLER_0_280 vgnd vpwr scs8hd_decap_12
XFILLER_8_1117 vgnd vpwr scs8hd_decap_12
XFILLER_14_129 vgnd vpwr scs8hd_decap_12
XFILLER_7_818 vgnd vpwr scs8hd_decap_8
XFILLER_10_324 vgnd vpwr scs8hd_decap_12
XFILLER_2_556 vgnd vpwr scs8hd_fill_1
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_1025 vgnd vpwr scs8hd_decap_12
XFILLER_13_1111 vgnd vpwr scs8hd_decap_12
XFILLER_11_611 vgnd vpwr scs8hd_decap_12
XFILLER_7_659 vgnd vpwr scs8hd_decap_12
XFILLER_10_154 vgnd vpwr scs8hd_decap_12
X_10_ _06_/Y enable address[3] _09_/D _10_/X vgnd vpwr scs8hd_and4_4
XFILLER_14_471 vgnd vpwr scs8hd_decap_12
XFILLER_6_692 vgnd vpwr scs8hd_decap_8
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_106 vgnd vpwr scs8hd_decap_12
XFILLER_4_629 vgnd vpwr scs8hd_decap_12
XFILLER_16_714 vgnd vpwr scs8hd_decap_12
XFILLER_16_769 vgnd vpwr scs8hd_decap_6
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
XFILLER_11_452 vgnd vpwr scs8hd_decap_12
XFILLER_7_489 vgnd vpwr scs8hd_decap_12
XFILLER_3_651 vgnd vpwr scs8hd_decap_12
XFILLER_3_684 vgnd vpwr scs8hd_decap_12
XFILLER_0_1017 vgnd vpwr scs8hd_decap_6
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_4_1142 vgnd vpwr scs8hd_decap_4
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_9_1086 vgnd vpwr scs8hd_decap_12
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XFILLER_4_415 vgnd vpwr scs8hd_decap_12
XFILLER_5_916 vgnd vpwr scs8hd_decap_12
XFILLER_5_938 vpwr vgnd scs8hd_fill_2
XFILLER_0_676 vgnd vpwr scs8hd_decap_6
XFILLER_0_621 vgnd vpwr scs8hd_decap_12
XFILLER_4_459 vgnd vpwr scs8hd_decap_12
XFILLER_15_1025 vgnd vpwr scs8hd_decap_12
XFILLER_11_293 vgnd vpwr scs8hd_decap_12
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
XFILLER_4_982 vgnd vpwr scs8hd_decap_12
XFILLER_8_776 vgnd vpwr scs8hd_decap_12
XFILLER_13_525 vgnd vpwr scs8hd_decap_12
XFILLER_16_385 vgnd vpwr scs8hd_decap_12
XFILLER_1_1123 vgnd vpwr scs8hd_decap_12
XPHY_380 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_6_1056 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_727 vgnd vpwr scs8hd_decap_12
XFILLER_14_812 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _10_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_598 vgnd vpwr scs8hd_decap_12
XFILLER_0_292 vgnd vpwr scs8hd_decap_12
XFILLER_11_1050 vgnd vpwr scs8hd_decap_12
XFILLER_14_642 vgnd vpwr scs8hd_decap_12
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XFILLER_15_428 vgnd vpwr scs8hd_decap_12
XFILLER_11_623 vgnd vpwr scs8hd_decap_12
XFILLER_13_1123 vgnd vpwr scs8hd_decap_12
XFILLER_10_166 vgnd vpwr scs8hd_decap_12
XFILLER_2_398 vgnd vpwr scs8hd_decap_12
XFILLER_3_855 vgnd vpwr scs8hd_decap_12
XFILLER_15_940 vgnd vpwr scs8hd_decap_12
XFILLER_2_1081 vgnd vpwr scs8hd_decap_12
XFILLER_14_483 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_869 vgnd vpwr scs8hd_decap_12
XFILLER_3_118 vgnd vpwr scs8hd_decap_4
XFILLER_16_726 vgnd vpwr scs8hd_decap_12
XFILLER_15_269 vgnd vpwr scs8hd_decap_12
XFILLER_12_910 vgnd vpwr scs8hd_decap_12
XFILLER_11_464 vgnd vpwr scs8hd_decap_12
XFILLER_7_413 vgnd vpwr scs8hd_decap_12
XFILLER_8_947 vgnd vpwr scs8hd_decap_12
XFILLER_3_663 vgnd vpwr scs8hd_decap_8
XFILLER_3_696 vgnd vpwr scs8hd_decap_6
XFILLER_15_781 vgnd vpwr scs8hd_decap_12
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XFILLER_4_427 vgnd vpwr scs8hd_decap_12
XFILLER_5_928 vgnd vpwr scs8hd_decap_8
XFILLER_0_633 vgnd vpwr scs8hd_decap_12
XFILLER_12_751 vgnd vpwr scs8hd_decap_12
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_788 vgnd vpwr scs8hd_decap_12
XFILLER_4_994 vgnd vpwr scs8hd_decap_12
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XFILLER_13_537 vgnd vpwr scs8hd_decap_12
XFILLER_14_1081 vgnd vpwr scs8hd_decap_12
XFILLER_1_953 vpwr vgnd scs8hd_fill_2
XFILLER_1_975 vgnd vpwr scs8hd_fill_1
XPHY_370 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_397 vgnd vpwr scs8hd_decap_6
XFILLER_16_342 vgnd vpwr scs8hd_decap_12
XFILLER_1_1135 vgnd vpwr scs8hd_decap_8
XPHY_381 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_581 vgnd vpwr scs8hd_decap_12
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_10_507 vgnd vpwr scs8hd_decap_12
XFILLER_2_739 vgnd vpwr scs8hd_decap_12
XFILLER_16_1110 vgnd vpwr scs8hd_decap_6
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_367 vgnd vpwr scs8hd_decap_12
XFILLER_1_794 vgnd vpwr scs8hd_decap_12
XFILLER_10_337 vgnd vpwr scs8hd_decap_12
XFILLER_11_1062 vgnd vpwr scs8hd_decap_12
XFILLER_14_654 vgnd vpwr scs8hd_decap_12
XFILLER_9_135 vgnd vpwr scs8hd_decap_12
XFILLER_5_330 vgnd vpwr scs8hd_decap_12
XFILLER_5_385 vgnd vpwr scs8hd_fill_1
XFILLER_5_396 vpwr vgnd scs8hd_fill_2
XFILLER_6_831 vgnd vpwr scs8hd_decap_12
XFILLER_6_886 vgnd vpwr scs8hd_decap_12
XFILLER_3_1038 vgnd vpwr scs8hd_decap_12
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _15_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_635 vgnd vpwr scs8hd_decap_12
XFILLER_13_1135 vgnd vpwr scs8hd_decap_8
XFILLER_2_300 vgnd vpwr scs8hd_decap_12
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_178 vgnd vpwr scs8hd_decap_12
XFILLER_2_388 vgnd vpwr scs8hd_decap_8
XFILLER_3_867 vgnd vpwr scs8hd_decap_12
XFILLER_15_952 vgnd vpwr scs8hd_decap_12
XFILLER_2_1093 vgnd vpwr scs8hd_decap_12
XFILLER_14_495 vgnd vpwr scs8hd_decap_12
XFILLER_10_690 vgnd vpwr scs8hd_decap_12
XFILLER_5_171 vgnd vpwr scs8hd_decap_8
XFILLER_16_738 vgnd vpwr scs8hd_decap_6
XFILLER_12_922 vgnd vpwr scs8hd_decap_12
XFILLER_11_476 vgnd vpwr scs8hd_decap_12
XFILLER_7_425 vpwr vgnd scs8hd_fill_2
XFILLER_8_959 vgnd vpwr scs8hd_decap_12
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
XFILLER_13_708 vgnd vpwr scs8hd_decap_12
XFILLER_9_1099 vgnd vpwr scs8hd_decap_12
XFILLER_4_439 vgnd vpwr scs8hd_decap_12
XFILLER_10_1105 vgnd vpwr scs8hd_decap_12
XFILLER_0_645 vgnd vpwr scs8hd_decap_6
XFILLER_15_1038 vgnd vpwr scs8hd_decap_12
XFILLER_14_1093 vgnd vpwr scs8hd_decap_12
XFILLER_5_704 vgnd vpwr scs8hd_decap_12
XFILLER_5_737 vgnd vpwr scs8hd_decap_12
XFILLER_0_431 vgnd vpwr scs8hd_decap_3
XFILLER_0_497 vgnd vpwr scs8hd_decap_12
XPHY_382 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_371 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_360 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_354 vgnd vpwr scs8hd_decap_12
XFILLER_8_520 vgnd vpwr scs8hd_decap_12
XFILLER_12_593 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_6_ logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[3] vgnd vpwr scs8hd_ebufn_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_1069 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_14_825 vgnd vpwr scs8hd_decap_12
XFILLER_13_379 vgnd vpwr scs8hd_decap_12
XFILLER_9_306 vgnd vpwr scs8hd_decap_12
XFILLER_12_1008 vgnd vpwr scs8hd_decap_12
XFILLER_5_501 vgnd vpwr scs8hd_decap_12
XFILLER_5_545 vgnd vpwr scs8hd_decap_4
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
XFILLER_13_891 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_361 vgnd vpwr scs8hd_decap_12
XFILLER_11_806 vgnd vpwr scs8hd_decap_12
XFILLER_11_1074 vgnd vpwr scs8hd_decap_12
XFILLER_10_349 vgnd vpwr scs8hd_decap_12
XFILLER_14_666 vgnd vpwr scs8hd_decap_12
XFILLER_13_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_147 vgnd vpwr scs8hd_decap_12
XFILLER_10_861 vgnd vpwr scs8hd_decap_12
XFILLER_3_11 vgnd vpwr scs8hd_decap_12
XFILLER_5_342 vgnd vpwr scs8hd_decap_12
XFILLER_6_843 vgnd vpwr scs8hd_decap_12
XFILLER_6_898 vgnd vpwr scs8hd_decap_12
XFILLER_11_647 vgnd vpwr scs8hd_decap_12
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XFILLER_2_312 vgnd vpwr scs8hd_decap_12
XFILLER_3_879 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_6
XFILLER_15_964 vgnd vpwr scs8hd_decap_12
XFILLER_6_651 vgnd vpwr scs8hd_decap_12
XFILLER_0_838 vgnd vpwr scs8hd_decap_12
XFILLER_12_934 vgnd vpwr scs8hd_decap_12
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_15_794 vgnd vpwr scs8hd_decap_12
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
XFILLER_9_1001 vgnd vpwr scs8hd_decap_12
XFILLER_0_602 vgnd vpwr scs8hd_decap_12
XFILLER_10_1117 vgnd vpwr scs8hd_decap_12
XFILLER_12_764 vgnd vpwr scs8hd_decap_12
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XFILLER_3_440 vgnd vpwr scs8hd_decap_12
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_716 vgnd vpwr scs8hd_decap_12
XFILLER_5_749 vgnd vpwr scs8hd_decap_12
XFILLER_1_977 vgnd vpwr scs8hd_decap_12
XFILLER_16_366 vgnd vpwr scs8hd_decap_6
XFILLER_16_311 vgnd vpwr scs8hd_decap_12
XPHY_372 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_361 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_350 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_532 vgnd vpwr scs8hd_decap_12
XFILLER_3_281 vgnd vpwr scs8hd_decap_12
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_1145 vgnd vpwr scs8hd_fill_1
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XFILLER_14_837 vgnd vpwr scs8hd_decap_12
XFILLER_9_318 vgnd vpwr scs8hd_decap_12
XFILLER_5_513 vgnd vpwr scs8hd_decap_12
XFILLER_0_273 vgnd vpwr scs8hd_decap_6
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_373 vgnd vpwr scs8hd_decap_12
XFILLER_9_830 vgnd vpwr scs8hd_decap_12
.ends

