magic
tech sky130A
magscale 1 2
timestamp 1608157227
<< obsli1 >>
rect 1104 2159 21620 20145
<< obsm1 >>
rect 198 1164 22618 20176
<< metal2 >>
rect 5722 22000 5778 22800
rect 17130 22000 17186 22800
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2410 0 2466 800
rect 2870 0 2926 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7746 0 7802 800
rect 8206 0 8262 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12254 0 12310 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 14922 0 14978 800
rect 15382 0 15438 800
rect 15842 0 15898 800
rect 16302 0 16358 800
rect 16670 0 16726 800
rect 17130 0 17186 800
rect 17590 0 17646 800
rect 18050 0 18106 800
rect 18510 0 18566 800
rect 18970 0 19026 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20258 0 20314 800
rect 20718 0 20774 800
rect 21178 0 21234 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
<< obsm2 >>
rect 204 21944 5666 22545
rect 5834 21944 17074 22545
rect 17242 21944 22612 22545
rect 204 856 22612 21944
rect 314 167 514 856
rect 682 167 974 856
rect 1142 167 1434 856
rect 1602 167 1894 856
rect 2062 167 2354 856
rect 2522 167 2814 856
rect 2982 167 3274 856
rect 3442 167 3642 856
rect 3810 167 4102 856
rect 4270 167 4562 856
rect 4730 167 5022 856
rect 5190 167 5482 856
rect 5650 167 5942 856
rect 6110 167 6402 856
rect 6570 167 6770 856
rect 6938 167 7230 856
rect 7398 167 7690 856
rect 7858 167 8150 856
rect 8318 167 8610 856
rect 8778 167 9070 856
rect 9238 167 9530 856
rect 9698 167 9898 856
rect 10066 167 10358 856
rect 10526 167 10818 856
rect 10986 167 11278 856
rect 11446 167 11738 856
rect 11906 167 12198 856
rect 12366 167 12658 856
rect 12826 167 13118 856
rect 13286 167 13486 856
rect 13654 167 13946 856
rect 14114 167 14406 856
rect 14574 167 14866 856
rect 15034 167 15326 856
rect 15494 167 15786 856
rect 15954 167 16246 856
rect 16414 167 16614 856
rect 16782 167 17074 856
rect 17242 167 17534 856
rect 17702 167 17994 856
rect 18162 167 18454 856
rect 18622 167 18914 856
rect 19082 167 19374 856
rect 19542 167 19742 856
rect 19910 167 20202 856
rect 20370 167 20662 856
rect 20830 167 21122 856
rect 21290 167 21582 856
rect 21750 167 22042 856
rect 22210 167 22502 856
<< metal3 >>
rect 0 22448 800 22568
rect 22000 22448 22800 22568
rect 0 22040 800 22160
rect 22000 22040 22800 22160
rect 0 21496 800 21616
rect 22000 21496 22800 21616
rect 0 21088 800 21208
rect 22000 21088 22800 21208
rect 0 20544 800 20664
rect 22000 20544 22800 20664
rect 0 20136 800 20256
rect 22000 20136 22800 20256
rect 0 19728 800 19848
rect 22000 19728 22800 19848
rect 0 19184 800 19304
rect 22000 19184 22800 19304
rect 0 18776 800 18896
rect 22000 18776 22800 18896
rect 0 18232 800 18352
rect 22000 18232 22800 18352
rect 0 17824 800 17944
rect 22000 17824 22800 17944
rect 0 17280 800 17400
rect 22000 17280 22800 17400
rect 0 16872 800 16992
rect 22000 16872 22800 16992
rect 0 16464 800 16584
rect 22000 16464 22800 16584
rect 0 15920 800 16040
rect 22000 15920 22800 16040
rect 0 15512 800 15632
rect 22000 15512 22800 15632
rect 0 14968 800 15088
rect 22000 14968 22800 15088
rect 0 14560 800 14680
rect 22000 14560 22800 14680
rect 0 14016 800 14136
rect 22000 14016 22800 14136
rect 0 13608 800 13728
rect 22000 13608 22800 13728
rect 0 13200 800 13320
rect 22000 13200 22800 13320
rect 0 12656 800 12776
rect 22000 12656 22800 12776
rect 0 12248 800 12368
rect 22000 12248 22800 12368
rect 0 11704 800 11824
rect 22000 11704 22800 11824
rect 0 11296 800 11416
rect 22000 11296 22800 11416
rect 0 10752 800 10872
rect 22000 10752 22800 10872
rect 0 10344 800 10464
rect 22000 10344 22800 10464
rect 0 9936 800 10056
rect 22000 9936 22800 10056
rect 0 9392 800 9512
rect 22000 9392 22800 9512
rect 0 8984 800 9104
rect 22000 8984 22800 9104
rect 0 8440 800 8560
rect 22000 8440 22800 8560
rect 0 8032 800 8152
rect 22000 8032 22800 8152
rect 0 7488 800 7608
rect 22000 7488 22800 7608
rect 0 7080 800 7200
rect 22000 7080 22800 7200
rect 0 6672 800 6792
rect 22000 6672 22800 6792
rect 0 6128 800 6248
rect 22000 6128 22800 6248
rect 0 5720 800 5840
rect 22000 5720 22800 5840
rect 0 5176 800 5296
rect 22000 5176 22800 5296
rect 0 4768 800 4888
rect 22000 4768 22800 4888
rect 0 4224 800 4344
rect 22000 4224 22800 4344
rect 0 3816 800 3936
rect 22000 3816 22800 3936
rect 0 3408 800 3528
rect 22000 3408 22800 3528
rect 0 2864 800 2984
rect 22000 2864 22800 2984
rect 0 2456 800 2576
rect 22000 2456 22800 2576
rect 0 1912 800 2032
rect 22000 1912 22800 2032
rect 0 1504 800 1624
rect 22000 1504 22800 1624
rect 0 960 800 1080
rect 22000 960 22800 1080
rect 0 552 800 672
rect 22000 552 22800 672
rect 0 144 800 264
rect 22000 144 22800 264
<< obsm3 >>
rect 880 22368 21920 22541
rect 800 22240 22000 22368
rect 880 21960 21920 22240
rect 800 21696 22000 21960
rect 880 21416 21920 21696
rect 800 21288 22000 21416
rect 880 21008 21920 21288
rect 800 20744 22000 21008
rect 880 20464 21920 20744
rect 800 20336 22000 20464
rect 880 20056 21920 20336
rect 800 19928 22000 20056
rect 880 19648 21920 19928
rect 800 19384 22000 19648
rect 880 19104 21920 19384
rect 800 18976 22000 19104
rect 880 18696 21920 18976
rect 800 18432 22000 18696
rect 880 18152 21920 18432
rect 800 18024 22000 18152
rect 880 17744 21920 18024
rect 800 17480 22000 17744
rect 880 17200 21920 17480
rect 800 17072 22000 17200
rect 880 16792 21920 17072
rect 800 16664 22000 16792
rect 880 16384 21920 16664
rect 800 16120 22000 16384
rect 880 15840 21920 16120
rect 800 15712 22000 15840
rect 880 15432 21920 15712
rect 800 15168 22000 15432
rect 880 14888 21920 15168
rect 800 14760 22000 14888
rect 880 14480 21920 14760
rect 800 14216 22000 14480
rect 880 13936 21920 14216
rect 800 13808 22000 13936
rect 880 13528 21920 13808
rect 800 13400 22000 13528
rect 880 13120 21920 13400
rect 800 12856 22000 13120
rect 880 12576 21920 12856
rect 800 12448 22000 12576
rect 880 12168 21920 12448
rect 800 11904 22000 12168
rect 880 11624 21920 11904
rect 800 11496 22000 11624
rect 880 11216 21920 11496
rect 800 10952 22000 11216
rect 880 10672 21920 10952
rect 800 10544 22000 10672
rect 880 10264 21920 10544
rect 800 10136 22000 10264
rect 880 9856 21920 10136
rect 800 9592 22000 9856
rect 880 9312 21920 9592
rect 800 9184 22000 9312
rect 880 8904 21920 9184
rect 800 8640 22000 8904
rect 880 8360 21920 8640
rect 800 8232 22000 8360
rect 880 7952 21920 8232
rect 800 7688 22000 7952
rect 880 7408 21920 7688
rect 800 7280 22000 7408
rect 880 7000 21920 7280
rect 800 6872 22000 7000
rect 880 6592 21920 6872
rect 800 6328 22000 6592
rect 880 6048 21920 6328
rect 800 5920 22000 6048
rect 880 5640 21920 5920
rect 800 5376 22000 5640
rect 880 5096 21920 5376
rect 800 4968 22000 5096
rect 880 4688 21920 4968
rect 800 4424 22000 4688
rect 880 4144 21920 4424
rect 800 4016 22000 4144
rect 880 3736 21920 4016
rect 800 3608 22000 3736
rect 880 3328 21920 3608
rect 800 3064 22000 3328
rect 880 2784 21920 3064
rect 800 2656 22000 2784
rect 880 2376 21920 2656
rect 800 2112 22000 2376
rect 880 1832 21920 2112
rect 800 1704 22000 1832
rect 880 1424 21920 1704
rect 800 1160 22000 1424
rect 880 880 21920 1160
rect 800 752 22000 880
rect 880 472 21920 752
rect 800 344 22000 472
rect 880 171 21920 344
<< metal4 >>
rect 4376 2128 4696 20176
rect 7808 2128 8128 20176
<< obsm4 >>
rect 5211 2048 7728 20176
rect 8208 2048 19445 20176
rect 5211 1939 19445 2048
<< labels >>
rlabel metal2 s 21638 0 21694 800 6 SC_IN_BOT
port 1 nsew default input
rlabel metal2 s 22098 0 22154 800 6 SC_OUT_BOT
port 2 nsew default output
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 3 nsew default input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 4 nsew default input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 5 nsew default input
rlabel metal2 s 1490 0 1546 800 6 bottom_left_grid_pin_45_
port 6 nsew default input
rlabel metal2 s 1950 0 2006 800 6 bottom_left_grid_pin_46_
port 7 nsew default input
rlabel metal2 s 2410 0 2466 800 6 bottom_left_grid_pin_47_
port 8 nsew default input
rlabel metal2 s 2870 0 2926 800 6 bottom_left_grid_pin_48_
port 9 nsew default input
rlabel metal2 s 3330 0 3386 800 6 bottom_left_grid_pin_49_
port 10 nsew default input
rlabel metal2 s 5722 22000 5778 22800 6 ccff_head
port 11 nsew default input
rlabel metal2 s 17130 22000 17186 22800 6 ccff_tail
port 12 nsew default output
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[0]
port 13 nsew default input
rlabel metal3 s 0 8440 800 8560 6 chanx_left_in[10]
port 14 nsew default input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[11]
port 15 nsew default input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[12]
port 16 nsew default input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[13]
port 17 nsew default input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[14]
port 18 nsew default input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[15]
port 19 nsew default input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[16]
port 20 nsew default input
rlabel metal3 s 0 11704 800 11824 6 chanx_left_in[17]
port 21 nsew default input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 22 nsew default input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[19]
port 23 nsew default input
rlabel metal3 s 0 4224 800 4344 6 chanx_left_in[1]
port 24 nsew default input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[2]
port 25 nsew default input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[3]
port 26 nsew default input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[4]
port 27 nsew default input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[5]
port 28 nsew default input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[6]
port 29 nsew default input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[7]
port 30 nsew default input
rlabel metal3 s 0 7488 800 7608 6 chanx_left_in[8]
port 31 nsew default input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[9]
port 32 nsew default input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[0]
port 33 nsew default output
rlabel metal3 s 0 17824 800 17944 6 chanx_left_out[10]
port 34 nsew default output
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[11]
port 35 nsew default output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[12]
port 36 nsew default output
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[13]
port 37 nsew default output
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[14]
port 38 nsew default output
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[15]
port 39 nsew default output
rlabel metal3 s 0 20544 800 20664 6 chanx_left_out[16]
port 40 nsew default output
rlabel metal3 s 0 21088 800 21208 6 chanx_left_out[17]
port 41 nsew default output
rlabel metal3 s 0 21496 800 21616 6 chanx_left_out[18]
port 42 nsew default output
rlabel metal3 s 0 22040 800 22160 6 chanx_left_out[19]
port 43 nsew default output
rlabel metal3 s 0 13608 800 13728 6 chanx_left_out[1]
port 44 nsew default output
rlabel metal3 s 0 14016 800 14136 6 chanx_left_out[2]
port 45 nsew default output
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[3]
port 46 nsew default output
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[4]
port 47 nsew default output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 48 nsew default output
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[6]
port 49 nsew default output
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[7]
port 50 nsew default output
rlabel metal3 s 0 16872 800 16992 6 chanx_left_out[8]
port 51 nsew default output
rlabel metal3 s 0 17280 800 17400 6 chanx_left_out[9]
port 52 nsew default output
rlabel metal3 s 22000 3816 22800 3936 6 chanx_right_in[0]
port 53 nsew default input
rlabel metal3 s 22000 8440 22800 8560 6 chanx_right_in[10]
port 54 nsew default input
rlabel metal3 s 22000 8984 22800 9104 6 chanx_right_in[11]
port 55 nsew default input
rlabel metal3 s 22000 9392 22800 9512 6 chanx_right_in[12]
port 56 nsew default input
rlabel metal3 s 22000 9936 22800 10056 6 chanx_right_in[13]
port 57 nsew default input
rlabel metal3 s 22000 10344 22800 10464 6 chanx_right_in[14]
port 58 nsew default input
rlabel metal3 s 22000 10752 22800 10872 6 chanx_right_in[15]
port 59 nsew default input
rlabel metal3 s 22000 11296 22800 11416 6 chanx_right_in[16]
port 60 nsew default input
rlabel metal3 s 22000 11704 22800 11824 6 chanx_right_in[17]
port 61 nsew default input
rlabel metal3 s 22000 12248 22800 12368 6 chanx_right_in[18]
port 62 nsew default input
rlabel metal3 s 22000 12656 22800 12776 6 chanx_right_in[19]
port 63 nsew default input
rlabel metal3 s 22000 4224 22800 4344 6 chanx_right_in[1]
port 64 nsew default input
rlabel metal3 s 22000 4768 22800 4888 6 chanx_right_in[2]
port 65 nsew default input
rlabel metal3 s 22000 5176 22800 5296 6 chanx_right_in[3]
port 66 nsew default input
rlabel metal3 s 22000 5720 22800 5840 6 chanx_right_in[4]
port 67 nsew default input
rlabel metal3 s 22000 6128 22800 6248 6 chanx_right_in[5]
port 68 nsew default input
rlabel metal3 s 22000 6672 22800 6792 6 chanx_right_in[6]
port 69 nsew default input
rlabel metal3 s 22000 7080 22800 7200 6 chanx_right_in[7]
port 70 nsew default input
rlabel metal3 s 22000 7488 22800 7608 6 chanx_right_in[8]
port 71 nsew default input
rlabel metal3 s 22000 8032 22800 8152 6 chanx_right_in[9]
port 72 nsew default input
rlabel metal3 s 22000 13200 22800 13320 6 chanx_right_out[0]
port 73 nsew default output
rlabel metal3 s 22000 17824 22800 17944 6 chanx_right_out[10]
port 74 nsew default output
rlabel metal3 s 22000 18232 22800 18352 6 chanx_right_out[11]
port 75 nsew default output
rlabel metal3 s 22000 18776 22800 18896 6 chanx_right_out[12]
port 76 nsew default output
rlabel metal3 s 22000 19184 22800 19304 6 chanx_right_out[13]
port 77 nsew default output
rlabel metal3 s 22000 19728 22800 19848 6 chanx_right_out[14]
port 78 nsew default output
rlabel metal3 s 22000 20136 22800 20256 6 chanx_right_out[15]
port 79 nsew default output
rlabel metal3 s 22000 20544 22800 20664 6 chanx_right_out[16]
port 80 nsew default output
rlabel metal3 s 22000 21088 22800 21208 6 chanx_right_out[17]
port 81 nsew default output
rlabel metal3 s 22000 21496 22800 21616 6 chanx_right_out[18]
port 82 nsew default output
rlabel metal3 s 22000 22040 22800 22160 6 chanx_right_out[19]
port 83 nsew default output
rlabel metal3 s 22000 13608 22800 13728 6 chanx_right_out[1]
port 84 nsew default output
rlabel metal3 s 22000 14016 22800 14136 6 chanx_right_out[2]
port 85 nsew default output
rlabel metal3 s 22000 14560 22800 14680 6 chanx_right_out[3]
port 86 nsew default output
rlabel metal3 s 22000 14968 22800 15088 6 chanx_right_out[4]
port 87 nsew default output
rlabel metal3 s 22000 15512 22800 15632 6 chanx_right_out[5]
port 88 nsew default output
rlabel metal3 s 22000 15920 22800 16040 6 chanx_right_out[6]
port 89 nsew default output
rlabel metal3 s 22000 16464 22800 16584 6 chanx_right_out[7]
port 90 nsew default output
rlabel metal3 s 22000 16872 22800 16992 6 chanx_right_out[8]
port 91 nsew default output
rlabel metal3 s 22000 17280 22800 17400 6 chanx_right_out[9]
port 92 nsew default output
rlabel metal2 s 3698 0 3754 800 6 chany_bottom_in[0]
port 93 nsew default input
rlabel metal2 s 8206 0 8262 800 6 chany_bottom_in[10]
port 94 nsew default input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[11]
port 95 nsew default input
rlabel metal2 s 9126 0 9182 800 6 chany_bottom_in[12]
port 96 nsew default input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[13]
port 97 nsew default input
rlabel metal2 s 9954 0 10010 800 6 chany_bottom_in[14]
port 98 nsew default input
rlabel metal2 s 10414 0 10470 800 6 chany_bottom_in[15]
port 99 nsew default input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[16]
port 100 nsew default input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_in[17]
port 101 nsew default input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[18]
port 102 nsew default input
rlabel metal2 s 12254 0 12310 800 6 chany_bottom_in[19]
port 103 nsew default input
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_in[1]
port 104 nsew default input
rlabel metal2 s 4618 0 4674 800 6 chany_bottom_in[2]
port 105 nsew default input
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_in[3]
port 106 nsew default input
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_in[4]
port 107 nsew default input
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_in[5]
port 108 nsew default input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[6]
port 109 nsew default input
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_in[7]
port 110 nsew default input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[8]
port 111 nsew default input
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_in[9]
port 112 nsew default input
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_out[0]
port 113 nsew default output
rlabel metal2 s 17130 0 17186 800 6 chany_bottom_out[10]
port 114 nsew default output
rlabel metal2 s 17590 0 17646 800 6 chany_bottom_out[11]
port 115 nsew default output
rlabel metal2 s 18050 0 18106 800 6 chany_bottom_out[12]
port 116 nsew default output
rlabel metal2 s 18510 0 18566 800 6 chany_bottom_out[13]
port 117 nsew default output
rlabel metal2 s 18970 0 19026 800 6 chany_bottom_out[14]
port 118 nsew default output
rlabel metal2 s 19430 0 19486 800 6 chany_bottom_out[15]
port 119 nsew default output
rlabel metal2 s 19798 0 19854 800 6 chany_bottom_out[16]
port 120 nsew default output
rlabel metal2 s 20258 0 20314 800 6 chany_bottom_out[17]
port 121 nsew default output
rlabel metal2 s 20718 0 20774 800 6 chany_bottom_out[18]
port 122 nsew default output
rlabel metal2 s 21178 0 21234 800 6 chany_bottom_out[19]
port 123 nsew default output
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_out[1]
port 124 nsew default output
rlabel metal2 s 13542 0 13598 800 6 chany_bottom_out[2]
port 125 nsew default output
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_out[3]
port 126 nsew default output
rlabel metal2 s 14462 0 14518 800 6 chany_bottom_out[4]
port 127 nsew default output
rlabel metal2 s 14922 0 14978 800 6 chany_bottom_out[5]
port 128 nsew default output
rlabel metal2 s 15382 0 15438 800 6 chany_bottom_out[6]
port 129 nsew default output
rlabel metal2 s 15842 0 15898 800 6 chany_bottom_out[7]
port 130 nsew default output
rlabel metal2 s 16302 0 16358 800 6 chany_bottom_out[8]
port 131 nsew default output
rlabel metal2 s 16670 0 16726 800 6 chany_bottom_out[9]
port 132 nsew default output
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 133 nsew default input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 134 nsew default input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 135 nsew default input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 136 nsew default input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_38_
port 137 nsew default input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 138 nsew default input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_40_
port 139 nsew default input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 140 nsew default input
rlabel metal3 s 0 22448 800 22568 6 left_top_grid_pin_1_
port 141 nsew default input
rlabel metal2 s 22558 0 22614 800 6 prog_clk_0_S_in
port 142 nsew default input
rlabel metal3 s 22000 144 22800 264 6 right_bottom_grid_pin_34_
port 143 nsew default input
rlabel metal3 s 22000 552 22800 672 6 right_bottom_grid_pin_35_
port 144 nsew default input
rlabel metal3 s 22000 960 22800 1080 6 right_bottom_grid_pin_36_
port 145 nsew default input
rlabel metal3 s 22000 1504 22800 1624 6 right_bottom_grid_pin_37_
port 146 nsew default input
rlabel metal3 s 22000 1912 22800 2032 6 right_bottom_grid_pin_38_
port 147 nsew default input
rlabel metal3 s 22000 2456 22800 2576 6 right_bottom_grid_pin_39_
port 148 nsew default input
rlabel metal3 s 22000 2864 22800 2984 6 right_bottom_grid_pin_40_
port 149 nsew default input
rlabel metal3 s 22000 3408 22800 3528 6 right_bottom_grid_pin_41_
port 150 nsew default input
rlabel metal3 s 22000 22448 22800 22568 6 right_top_grid_pin_1_
port 151 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 152 nsew power input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 153 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22800 22800
string LEFview TRUE
<< end >>
