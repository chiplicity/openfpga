VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__1_
  CLASS BLOCK ;
  FOREIGN sb_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 2.400 ;
    END
  END bottom_left_grid_pin_11_
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 2.400 ;
    END
  END bottom_left_grid_pin_15_
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN bottom_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.400 ;
    END
  END bottom_left_grid_pin_3_
  PIN bottom_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 2.400 ;
    END
  END bottom_left_grid_pin_5_
  PIN bottom_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 2.400 ;
    END
  END bottom_left_grid_pin_7_
  PIN bottom_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 2.400 ;
    END
  END bottom_left_grid_pin_9_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 2.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 8.880 140.000 9.480 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 15.680 140.000 16.280 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 22.480 140.000 23.080 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 29.280 140.000 29.880 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 36.080 140.000 36.680 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 42.200 140.000 42.800 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 49.000 140.000 49.600 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 55.800 140.000 56.400 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 62.600 140.000 63.200 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 82.320 140.000 82.920 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 89.120 140.000 89.720 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.920 140.000 96.520 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 102.720 140.000 103.320 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 108.840 140.000 109.440 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 115.640 140.000 116.240 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 122.440 140.000 123.040 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.240 140.000 129.840 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.040 140.000 136.640 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 137.600 4.050 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 137.600 11.410 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 137.600 19.230 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 137.600 27.050 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 137.600 34.870 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 137.600 42.690 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 137.600 50.510 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 137.600 58.330 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 137.600 66.150 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 137.600 73.970 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 137.600 81.330 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 137.600 89.150 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 137.600 96.970 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.510 137.600 104.790 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 137.600 112.610 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.150 137.600 120.430 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.970 137.600 128.250 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.790 137.600 136.070 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 2.400 ;
    END
  END enable
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 75.520 140.000 76.120 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END top_left_grid_pin_11_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.400 113.520 ;
    END
  END top_left_grid_pin_13_
  PIN top_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.400 131.200 ;
    END
  END top_left_grid_pin_15_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END top_left_grid_pin_1_
  PIN top_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END top_left_grid_pin_3_
  PIN top_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END top_left_grid_pin_5_
  PIN top_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 2.400 61.160 ;
    END
  END top_left_grid_pin_7_
  PIN top_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.400 78.840 ;
    END
  END top_left_grid_pin_9_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 2.760 140.000 3.360 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    USE POWER ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.530 0.040 138.390 137.660 ;
      LAYER met2 ;
        RECT 0.550 137.320 3.490 137.770 ;
        RECT 4.330 137.320 10.850 137.770 ;
        RECT 11.690 137.320 18.670 137.770 ;
        RECT 19.510 137.320 26.490 137.770 ;
        RECT 27.330 137.320 34.310 137.770 ;
        RECT 35.150 137.320 42.130 137.770 ;
        RECT 42.970 137.320 49.950 137.770 ;
        RECT 50.790 137.320 57.770 137.770 ;
        RECT 58.610 137.320 65.590 137.770 ;
        RECT 66.430 137.320 73.410 137.770 ;
        RECT 74.250 137.320 80.770 137.770 ;
        RECT 81.610 137.320 88.590 137.770 ;
        RECT 89.430 137.320 96.410 137.770 ;
        RECT 97.250 137.320 104.230 137.770 ;
        RECT 105.070 137.320 112.050 137.770 ;
        RECT 112.890 137.320 119.870 137.770 ;
        RECT 120.710 137.320 127.690 137.770 ;
        RECT 128.530 137.320 135.510 137.770 ;
        RECT 136.350 137.320 138.370 137.770 ;
        RECT 0.550 2.680 138.370 137.320 ;
        RECT 0.550 0.010 1.650 2.680 ;
        RECT 2.490 0.010 5.330 2.680 ;
        RECT 6.170 0.010 9.010 2.680 ;
        RECT 9.850 0.010 13.150 2.680 ;
        RECT 13.990 0.010 16.830 2.680 ;
        RECT 17.670 0.010 20.970 2.680 ;
        RECT 21.810 0.010 24.650 2.680 ;
        RECT 25.490 0.010 28.790 2.680 ;
        RECT 29.630 0.010 32.470 2.680 ;
        RECT 33.310 0.010 36.610 2.680 ;
        RECT 37.450 0.010 40.290 2.680 ;
        RECT 41.130 0.010 43.970 2.680 ;
        RECT 44.810 0.010 48.110 2.680 ;
        RECT 48.950 0.010 51.790 2.680 ;
        RECT 52.630 0.010 55.930 2.680 ;
        RECT 56.770 0.010 59.610 2.680 ;
        RECT 60.450 0.010 63.750 2.680 ;
        RECT 64.590 0.010 67.430 2.680 ;
        RECT 68.270 0.010 71.570 2.680 ;
        RECT 72.410 0.010 75.250 2.680 ;
        RECT 76.090 0.010 78.930 2.680 ;
        RECT 79.770 0.010 83.070 2.680 ;
        RECT 83.910 0.010 86.750 2.680 ;
        RECT 87.590 0.010 90.890 2.680 ;
        RECT 91.730 0.010 94.570 2.680 ;
        RECT 95.410 0.010 98.710 2.680 ;
        RECT 99.550 0.010 102.390 2.680 ;
        RECT 103.230 0.010 106.530 2.680 ;
        RECT 107.370 0.010 110.210 2.680 ;
        RECT 111.050 0.010 113.890 2.680 ;
        RECT 114.730 0.010 118.030 2.680 ;
        RECT 118.870 0.010 121.710 2.680 ;
        RECT 122.550 0.010 125.850 2.680 ;
        RECT 126.690 0.010 129.530 2.680 ;
        RECT 130.370 0.010 133.670 2.680 ;
        RECT 134.510 0.010 137.350 2.680 ;
        RECT 138.190 0.010 138.370 2.680 ;
      LAYER met3 ;
        RECT 0.310 137.040 138.650 137.865 ;
        RECT 0.310 135.640 137.200 137.040 ;
        RECT 0.310 131.600 138.650 135.640 ;
        RECT 2.800 130.240 138.650 131.600 ;
        RECT 2.800 130.200 137.200 130.240 ;
        RECT 0.310 128.840 137.200 130.200 ;
        RECT 0.310 123.440 138.650 128.840 ;
        RECT 0.310 122.040 137.200 123.440 ;
        RECT 0.310 116.640 138.650 122.040 ;
        RECT 0.310 115.240 137.200 116.640 ;
        RECT 0.310 113.920 138.650 115.240 ;
        RECT 2.800 112.520 138.650 113.920 ;
        RECT 0.310 109.840 138.650 112.520 ;
        RECT 0.310 108.440 137.200 109.840 ;
        RECT 0.310 103.720 138.650 108.440 ;
        RECT 0.310 102.320 137.200 103.720 ;
        RECT 0.310 96.920 138.650 102.320 ;
        RECT 0.310 96.240 137.200 96.920 ;
        RECT 2.800 95.520 137.200 96.240 ;
        RECT 2.800 94.840 138.650 95.520 ;
        RECT 0.310 90.120 138.650 94.840 ;
        RECT 0.310 88.720 137.200 90.120 ;
        RECT 0.310 83.320 138.650 88.720 ;
        RECT 0.310 81.920 137.200 83.320 ;
        RECT 0.310 79.240 138.650 81.920 ;
        RECT 2.800 77.840 138.650 79.240 ;
        RECT 0.310 76.520 138.650 77.840 ;
        RECT 0.310 75.120 137.200 76.520 ;
        RECT 0.310 70.400 138.650 75.120 ;
        RECT 0.310 69.000 137.200 70.400 ;
        RECT 0.310 63.600 138.650 69.000 ;
        RECT 0.310 62.200 137.200 63.600 ;
        RECT 0.310 61.560 138.650 62.200 ;
        RECT 2.800 60.160 138.650 61.560 ;
        RECT 0.310 56.800 138.650 60.160 ;
        RECT 0.310 55.400 137.200 56.800 ;
        RECT 0.310 50.000 138.650 55.400 ;
        RECT 0.310 48.600 137.200 50.000 ;
        RECT 0.310 43.880 138.650 48.600 ;
        RECT 2.800 43.200 138.650 43.880 ;
        RECT 2.800 42.480 137.200 43.200 ;
        RECT 0.310 41.800 137.200 42.480 ;
        RECT 0.310 37.080 138.650 41.800 ;
        RECT 0.310 35.680 137.200 37.080 ;
        RECT 0.310 30.280 138.650 35.680 ;
        RECT 0.310 28.880 137.200 30.280 ;
        RECT 0.310 26.200 138.650 28.880 ;
        RECT 2.800 24.800 138.650 26.200 ;
        RECT 0.310 23.480 138.650 24.800 ;
        RECT 0.310 22.080 137.200 23.480 ;
        RECT 0.310 16.680 138.650 22.080 ;
        RECT 0.310 15.280 137.200 16.680 ;
        RECT 0.310 9.880 138.650 15.280 ;
        RECT 0.310 9.200 137.200 9.880 ;
        RECT 2.800 8.480 137.200 9.200 ;
        RECT 2.800 7.800 138.650 8.480 ;
        RECT 0.310 3.760 138.650 7.800 ;
        RECT 0.310 3.360 137.200 3.760 ;
      LAYER met4 ;
        RECT 20.110 128.480 138.625 137.865 ;
        RECT 20.110 10.240 27.655 128.480 ;
        RECT 30.055 10.240 50.985 128.480 ;
        RECT 53.385 10.240 138.625 128.480 ;
        RECT 20.110 4.510 138.625 10.240 ;
      LAYER met5 ;
        RECT 19.900 4.300 96.940 19.500 ;
  END
END sb_0__1_
END LIBRARY

