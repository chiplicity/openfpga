magic
tech sky130A
magscale 1 2
timestamp 1605205362
<< locali >>
rect 12633 19159 12667 19465
rect 7113 18615 7147 18921
rect 10517 18615 10551 18921
rect 21005 18343 21039 19125
rect 9689 9979 9723 10081
rect 12265 9503 12299 9673
rect 12265 9469 12357 9503
rect 10057 8415 10091 8585
rect 15393 8279 15427 8517
rect 9689 7735 9723 8041
rect 12081 7871 12115 8041
rect 8677 6647 8711 6817
rect 15117 6783 15151 6953
rect 21005 6919 21039 8041
rect 21005 5695 21039 6681
<< viali >>
rect 7665 19465 7699 19499
rect 12633 19465 12667 19499
rect 2329 19329 2363 19363
rect 3157 19329 3191 19363
rect 4721 19329 4755 19363
rect 5457 19329 5491 19363
rect 6653 19329 6687 19363
rect 8217 19329 8251 19363
rect 9505 19329 9539 19363
rect 10977 19329 11011 19363
rect 11805 19329 11839 19363
rect 2053 19261 2087 19295
rect 3341 19261 3375 19295
rect 6377 19261 6411 19295
rect 6929 19261 6963 19295
rect 7297 19261 7331 19295
rect 8493 19261 8527 19295
rect 9229 19261 9263 19295
rect 9787 19261 9821 19295
rect 12173 19261 12207 19295
rect 4537 19193 4571 19227
rect 5365 19193 5399 19227
rect 14197 19397 14231 19431
rect 14841 19329 14875 19363
rect 17693 19329 17727 19363
rect 18797 19329 18831 19363
rect 18981 19329 19015 19363
rect 19717 19329 19751 19363
rect 12725 19261 12759 19295
rect 15025 19261 15059 19295
rect 15676 19261 15710 19295
rect 19625 19261 19659 19295
rect 19993 19261 20027 19295
rect 12992 19193 13026 19227
rect 15914 19193 15948 19227
rect 19533 19193 19567 19227
rect 1685 19125 1719 19159
rect 2145 19125 2179 19159
rect 2513 19125 2547 19159
rect 2881 19125 2915 19159
rect 2973 19125 3007 19159
rect 3525 19125 3559 19159
rect 4077 19125 4111 19159
rect 4445 19125 4479 19159
rect 4905 19125 4939 19159
rect 5273 19125 5307 19159
rect 6009 19125 6043 19159
rect 6469 19125 6503 19159
rect 7113 19125 7147 19159
rect 7481 19125 7515 19159
rect 8033 19125 8067 19159
rect 8125 19125 8159 19159
rect 8677 19125 8711 19159
rect 8861 19125 8895 19159
rect 9321 19125 9355 19159
rect 9965 19125 9999 19159
rect 10333 19125 10367 19159
rect 10701 19125 10735 19159
rect 10793 19125 10827 19159
rect 11161 19125 11195 19159
rect 11529 19125 11563 19159
rect 11621 19125 11655 19159
rect 12357 19125 12391 19159
rect 12633 19125 12667 19159
rect 14105 19125 14139 19159
rect 14565 19125 14599 19159
rect 14657 19125 14691 19159
rect 15209 19125 15243 19159
rect 17049 19125 17083 19159
rect 17141 19125 17175 19159
rect 17509 19125 17543 19159
rect 17601 19125 17635 19159
rect 18337 19125 18371 19159
rect 18705 19125 18739 19159
rect 19165 19125 19199 19159
rect 20177 19125 20211 19159
rect 21005 19125 21039 19159
rect 1593 18921 1627 18955
rect 3525 18921 3559 18955
rect 3801 18921 3835 18955
rect 7113 18921 7147 18955
rect 9229 18921 9263 18955
rect 9689 18921 9723 18955
rect 10517 18921 10551 18955
rect 14013 18921 14047 18955
rect 14105 18921 14139 18955
rect 17141 18921 17175 18955
rect 19809 18921 19843 18955
rect 20085 18921 20119 18955
rect 1409 18785 1443 18819
rect 1777 18785 1811 18819
rect 2145 18785 2179 18819
rect 2412 18785 2446 18819
rect 3617 18785 3651 18819
rect 4344 18785 4378 18819
rect 5816 18785 5850 18819
rect 4077 18717 4111 18751
rect 5549 18717 5583 18751
rect 5457 18649 5491 18683
rect 7472 18785 7506 18819
rect 9137 18785 9171 18819
rect 10057 18785 10091 18819
rect 7205 18717 7239 18751
rect 9321 18717 9355 18751
rect 10149 18717 10183 18751
rect 10241 18717 10275 18751
rect 8769 18649 8803 18683
rect 10968 18853 11002 18887
rect 14933 18853 14967 18887
rect 16028 18853 16062 18887
rect 17969 18853 18003 18887
rect 10701 18785 10735 18819
rect 12173 18785 12207 18819
rect 12633 18785 12667 18819
rect 12900 18785 12934 18819
rect 14473 18785 14507 18819
rect 15301 18785 15335 18819
rect 15485 18785 15519 18819
rect 17233 18785 17267 18819
rect 18061 18785 18095 18819
rect 18696 18785 18730 18819
rect 19901 18785 19935 18819
rect 20269 18785 20303 18819
rect 14565 18717 14599 18751
rect 14657 18717 14691 18751
rect 15761 18717 15795 18751
rect 18153 18717 18187 18751
rect 18429 18717 18463 18751
rect 17601 18649 17635 18683
rect 20453 18649 20487 18683
rect 1961 18581 1995 18615
rect 6929 18581 6963 18615
rect 7113 18581 7147 18615
rect 8585 18581 8619 18615
rect 10517 18581 10551 18615
rect 12081 18581 12115 18615
rect 12357 18581 12391 18615
rect 15669 18581 15703 18615
rect 17417 18581 17451 18615
rect 2789 18377 2823 18411
rect 4353 18377 4387 18411
rect 9229 18377 9263 18411
rect 12173 18377 12207 18411
rect 14933 18377 14967 18411
rect 19533 18377 19567 18411
rect 6653 18309 6687 18343
rect 6837 18309 6871 18343
rect 17325 18309 17359 18343
rect 17785 18309 17819 18343
rect 19441 18309 19475 18343
rect 21005 18309 21039 18343
rect 5089 18241 5123 18275
rect 5273 18241 5307 18275
rect 7389 18241 7423 18275
rect 14473 18241 14507 18275
rect 15577 18241 15611 18275
rect 15669 18241 15703 18275
rect 15945 18241 15979 18275
rect 20085 18241 20119 18275
rect 1409 18173 1443 18207
rect 2973 18173 3007 18207
rect 3240 18173 3274 18207
rect 4905 18173 4939 18207
rect 5540 18173 5574 18207
rect 7849 18173 7883 18207
rect 9321 18173 9355 18207
rect 9577 18173 9611 18207
rect 10793 18173 10827 18207
rect 12449 18173 12483 18207
rect 12716 18173 12750 18207
rect 14381 18173 14415 18207
rect 14749 18173 14783 18207
rect 15485 18173 15519 18207
rect 16212 18173 16246 18207
rect 17601 18173 17635 18207
rect 18061 18173 18095 18207
rect 1676 18105 1710 18139
rect 7297 18105 7331 18139
rect 8116 18105 8150 18139
rect 11060 18105 11094 18139
rect 14289 18105 14323 18139
rect 18328 18105 18362 18139
rect 19993 18105 20027 18139
rect 4445 18037 4479 18071
rect 4813 18037 4847 18071
rect 7205 18037 7239 18071
rect 10701 18037 10735 18071
rect 13829 18037 13863 18071
rect 13921 18037 13955 18071
rect 15117 18037 15151 18071
rect 19901 18037 19935 18071
rect 2789 17833 2823 17867
rect 3525 17833 3559 17867
rect 5733 17833 5767 17867
rect 9321 17833 9355 17867
rect 11253 17833 11287 17867
rect 12817 17833 12851 17867
rect 13921 17833 13955 17867
rect 15853 17833 15887 17867
rect 16405 17833 16439 17867
rect 16497 17833 16531 17867
rect 19349 17833 19383 17867
rect 6101 17765 6135 17799
rect 6285 17765 6319 17799
rect 6469 17765 6503 17799
rect 6920 17765 6954 17799
rect 10140 17765 10174 17799
rect 11612 17765 11646 17799
rect 17601 17765 17635 17799
rect 19809 17765 19843 17799
rect 1409 17697 1443 17731
rect 1676 17697 1710 17731
rect 3617 17697 3651 17731
rect 4077 17697 4111 17731
rect 4721 17697 4755 17731
rect 5641 17697 5675 17731
rect 8493 17697 8527 17731
rect 8585 17697 8619 17731
rect 8953 17697 8987 17731
rect 13185 17697 13219 17731
rect 13737 17697 13771 17731
rect 14749 17697 14783 17731
rect 15301 17697 15335 17731
rect 15669 17697 15703 17731
rect 17509 17697 17543 17731
rect 18236 17697 18270 17731
rect 20269 17697 20303 17731
rect 3801 17629 3835 17663
rect 4813 17629 4847 17663
rect 4997 17629 5031 17663
rect 5825 17629 5859 17663
rect 6653 17629 6687 17663
rect 8677 17629 8711 17663
rect 9873 17629 9907 17663
rect 11345 17629 11379 17663
rect 13277 17629 13311 17663
rect 13369 17629 13403 17663
rect 14105 17629 14139 17663
rect 14841 17629 14875 17663
rect 15025 17629 15059 17663
rect 16589 17629 16623 17663
rect 17693 17629 17727 17663
rect 17969 17629 18003 17663
rect 19901 17629 19935 17663
rect 20085 17629 20119 17663
rect 8033 17561 8067 17595
rect 8125 17561 8159 17595
rect 12725 17561 12759 17595
rect 15485 17561 15519 17595
rect 16037 17561 16071 17595
rect 19441 17561 19475 17595
rect 3157 17493 3191 17527
rect 4353 17493 4387 17527
rect 5273 17493 5307 17527
rect 9137 17493 9171 17527
rect 14381 17493 14415 17527
rect 17141 17493 17175 17527
rect 20453 17493 20487 17527
rect 5733 17289 5767 17323
rect 8585 17289 8619 17323
rect 13277 17289 13311 17323
rect 17785 17289 17819 17323
rect 19441 17289 19475 17323
rect 19533 17289 19567 17323
rect 1593 17221 1627 17255
rect 15761 17221 15795 17255
rect 3893 17153 3927 17187
rect 4721 17153 4755 17187
rect 5457 17153 5491 17187
rect 6377 17153 6411 17187
rect 10609 17153 10643 17187
rect 10885 17153 10919 17187
rect 13093 17153 13127 17187
rect 13829 17153 13863 17187
rect 14197 17153 14231 17187
rect 16313 17153 16347 17187
rect 17141 17153 17175 17187
rect 20085 17153 20119 17187
rect 1409 17085 1443 17119
rect 1777 17085 1811 17119
rect 3617 17085 3651 17119
rect 3709 17085 3743 17119
rect 4445 17085 4479 17119
rect 6929 17085 6963 17119
rect 8401 17085 8435 17119
rect 8769 17085 8803 17119
rect 9036 17085 9070 17119
rect 10241 17085 10275 17119
rect 12817 17085 12851 17119
rect 13645 17085 13679 17119
rect 13737 17085 13771 17119
rect 16129 17085 16163 17119
rect 17601 17085 17635 17119
rect 18061 17085 18095 17119
rect 18328 17085 18362 17119
rect 19901 17085 19935 17119
rect 2044 17017 2078 17051
rect 5273 17017 5307 17051
rect 7196 17017 7230 17051
rect 11152 17017 11186 17051
rect 14464 17017 14498 17051
rect 19993 17017 20027 17051
rect 3157 16949 3191 16983
rect 3249 16949 3283 16983
rect 4077 16949 4111 16983
rect 4537 16949 4571 16983
rect 4905 16949 4939 16983
rect 5365 16949 5399 16983
rect 6101 16949 6135 16983
rect 6193 16949 6227 16983
rect 8309 16949 8343 16983
rect 10149 16949 10183 16983
rect 10425 16949 10459 16983
rect 12265 16949 12299 16983
rect 12449 16949 12483 16983
rect 12909 16949 12943 16983
rect 15577 16949 15611 16983
rect 16221 16949 16255 16983
rect 16589 16949 16623 16983
rect 16957 16949 16991 16983
rect 17049 16949 17083 16983
rect 1593 16745 1627 16779
rect 3157 16745 3191 16779
rect 3433 16745 3467 16779
rect 4353 16745 4387 16779
rect 4537 16745 4571 16779
rect 5365 16745 5399 16779
rect 6377 16745 6411 16779
rect 7297 16745 7331 16779
rect 8131 16745 8165 16779
rect 9505 16745 9539 16779
rect 11621 16745 11655 16779
rect 11989 16745 12023 16779
rect 14013 16745 14047 16779
rect 15301 16745 15335 16779
rect 17785 16745 17819 16779
rect 19257 16745 19291 16779
rect 20361 16745 20395 16779
rect 2044 16677 2078 16711
rect 4905 16677 4939 16711
rect 12808 16677 12842 16711
rect 14381 16677 14415 16711
rect 18122 16677 18156 16711
rect 1409 16609 1443 16643
rect 1777 16609 1811 16643
rect 3249 16609 3283 16643
rect 3617 16609 3651 16643
rect 4169 16609 4203 16643
rect 4997 16609 5031 16643
rect 5733 16609 5767 16643
rect 5825 16609 5859 16643
rect 6193 16609 6227 16643
rect 6561 16609 6595 16643
rect 7205 16609 7239 16643
rect 8401 16609 8435 16643
rect 10425 16609 10459 16643
rect 12541 16609 12575 16643
rect 14841 16609 14875 16643
rect 15669 16609 15703 16643
rect 15761 16609 15795 16643
rect 16405 16609 16439 16643
rect 16672 16609 16706 16643
rect 17877 16609 17911 16643
rect 19717 16609 19751 16643
rect 20177 16609 20211 16643
rect 5089 16541 5123 16575
rect 6009 16541 6043 16575
rect 7481 16541 7515 16575
rect 7665 16541 7699 16575
rect 8128 16541 8162 16575
rect 9689 16541 9723 16575
rect 10012 16541 10046 16575
rect 10152 16541 10186 16575
rect 12081 16541 12115 16575
rect 12173 16541 12207 16575
rect 14473 16541 14507 16575
rect 14565 16541 14599 16575
rect 15853 16541 15887 16575
rect 19809 16541 19843 16575
rect 19993 16541 20027 16575
rect 3801 16473 3835 16507
rect 13921 16473 13955 16507
rect 6837 16405 6871 16439
rect 11529 16405 11563 16439
rect 15025 16405 15059 16439
rect 19349 16405 19383 16439
rect 3617 16201 3651 16235
rect 6469 16201 6503 16235
rect 7297 16201 7331 16235
rect 9965 16201 9999 16235
rect 12173 16201 12207 16235
rect 14197 16201 14231 16235
rect 15945 16201 15979 16235
rect 17417 16201 17451 16235
rect 19441 16201 19475 16235
rect 3249 16133 3283 16167
rect 17693 16133 17727 16167
rect 1869 16065 1903 16099
rect 4077 16065 4111 16099
rect 4169 16065 4203 16099
rect 4813 16065 4847 16099
rect 7757 16065 7791 16099
rect 7849 16065 7883 16099
rect 8588 16065 8622 16099
rect 8861 16065 8895 16099
rect 10057 16065 10091 16099
rect 10796 16065 10830 16099
rect 11069 16065 11103 16099
rect 16037 16065 16071 16099
rect 20085 16065 20119 16099
rect 1501 15997 1535 16031
rect 2136 15997 2170 16031
rect 3525 15997 3559 16031
rect 4445 15997 4479 16031
rect 6285 15997 6319 16031
rect 6929 15997 6963 16031
rect 7665 15997 7699 16031
rect 8125 15997 8159 16031
rect 8448 15997 8482 16031
rect 10333 15997 10367 16031
rect 12449 15997 12483 16031
rect 12817 15997 12851 16031
rect 13084 15997 13118 16031
rect 14565 15997 14599 16031
rect 14832 15997 14866 16031
rect 16304 15997 16338 16031
rect 17509 15997 17543 16031
rect 18061 15997 18095 16031
rect 3985 15929 4019 15963
rect 5080 15929 5114 15963
rect 14289 15929 14323 15963
rect 18306 15929 18340 15963
rect 19901 15929 19935 15963
rect 1685 15861 1719 15895
rect 3341 15861 3375 15895
rect 4629 15861 4663 15895
rect 6193 15861 6227 15895
rect 7113 15861 7147 15895
rect 10799 15861 10833 15895
rect 12633 15861 12667 15895
rect 19533 15861 19567 15895
rect 19993 15861 20027 15895
rect 3433 15657 3467 15691
rect 8401 15657 8435 15691
rect 8493 15657 8527 15691
rect 11069 15657 11103 15691
rect 14381 15657 14415 15691
rect 14657 15657 14691 15691
rect 16865 15657 16899 15691
rect 18521 15657 18555 15691
rect 19993 15657 20027 15691
rect 2044 15589 2078 15623
rect 4344 15589 4378 15623
rect 5816 15589 5850 15623
rect 15730 15589 15764 15623
rect 17386 15589 17420 15623
rect 1777 15521 1811 15555
rect 3249 15521 3283 15555
rect 3617 15521 3651 15555
rect 5549 15521 5583 15555
rect 7277 15521 7311 15555
rect 8861 15521 8895 15555
rect 9321 15521 9355 15555
rect 9945 15521 9979 15555
rect 11529 15521 11563 15555
rect 11796 15521 11830 15555
rect 13268 15521 13302 15555
rect 14473 15521 14507 15555
rect 14841 15521 14875 15555
rect 17141 15521 17175 15555
rect 18613 15521 18647 15555
rect 18880 15521 18914 15555
rect 20085 15521 20119 15555
rect 4077 15453 4111 15487
rect 7021 15453 7055 15487
rect 8953 15453 8987 15487
rect 9137 15453 9171 15487
rect 9689 15453 9723 15487
rect 11253 15453 11287 15487
rect 13001 15453 13035 15487
rect 15485 15453 15519 15487
rect 3157 15385 3191 15419
rect 12909 15385 12943 15419
rect 3801 15317 3835 15351
rect 5457 15317 5491 15351
rect 6929 15317 6963 15351
rect 15025 15317 15059 15351
rect 20269 15317 20303 15351
rect 2881 15113 2915 15147
rect 4813 15113 4847 15147
rect 5733 15113 5767 15147
rect 8217 15113 8251 15147
rect 9689 15113 9723 15147
rect 12449 15113 12483 15147
rect 13001 15113 13035 15147
rect 15209 15113 15243 15147
rect 15393 15113 15427 15147
rect 17693 15113 17727 15147
rect 10885 15045 10919 15079
rect 1501 14977 1535 15011
rect 3433 14977 3467 15011
rect 5457 14977 5491 15011
rect 6193 14977 6227 15011
rect 6285 14977 6319 15011
rect 10425 14977 10459 15011
rect 11437 14977 11471 15011
rect 13185 14977 13219 15011
rect 16037 14977 16071 15011
rect 18981 14977 19015 15011
rect 19165 14977 19199 15011
rect 1768 14909 1802 14943
rect 3065 14909 3099 14943
rect 5365 14909 5399 14943
rect 6837 14909 6871 14943
rect 8309 14909 8343 14943
rect 10149 14909 10183 14943
rect 11253 14909 11287 14943
rect 11897 14909 11931 14943
rect 12265 14909 12299 14943
rect 12633 14909 12667 14943
rect 12817 14909 12851 14943
rect 13452 14909 13486 14943
rect 14657 14909 14691 14943
rect 15025 14909 15059 14943
rect 16221 14909 16255 14943
rect 17877 14909 17911 14943
rect 18705 14909 18739 14943
rect 19432 14909 19466 14943
rect 3700 14841 3734 14875
rect 5273 14841 5307 14875
rect 6101 14841 6135 14875
rect 7104 14841 7138 14875
rect 8576 14841 8610 14875
rect 10241 14841 10275 14875
rect 11345 14841 11379 14875
rect 15853 14841 15887 14875
rect 16488 14841 16522 14875
rect 18797 14841 18831 14875
rect 3249 14773 3283 14807
rect 4905 14773 4939 14807
rect 9781 14773 9815 14807
rect 10609 14773 10643 14807
rect 11713 14773 11747 14807
rect 12081 14773 12115 14807
rect 14565 14773 14599 14807
rect 14841 14773 14875 14807
rect 15761 14773 15795 14807
rect 17601 14773 17635 14807
rect 18337 14773 18371 14807
rect 20545 14773 20579 14807
rect 2789 14569 2823 14603
rect 2881 14569 2915 14603
rect 4445 14569 4479 14603
rect 4905 14569 4939 14603
rect 7205 14569 7239 14603
rect 9229 14569 9263 14603
rect 13185 14569 13219 14603
rect 13277 14569 13311 14603
rect 20085 14569 20119 14603
rect 3249 14501 3283 14535
rect 5365 14501 5399 14535
rect 7542 14501 7576 14535
rect 9137 14501 9171 14535
rect 10057 14501 10091 14535
rect 10589 14501 10623 14535
rect 18972 14501 19006 14535
rect 20177 14501 20211 14535
rect 1409 14433 1443 14467
rect 1676 14433 1710 14467
rect 3893 14433 3927 14467
rect 5273 14433 5307 14467
rect 5825 14433 5859 14467
rect 6092 14433 6126 14467
rect 7297 14433 7331 14467
rect 9689 14433 9723 14467
rect 10333 14433 10367 14467
rect 11805 14433 11839 14467
rect 12072 14433 12106 14467
rect 13820 14433 13854 14467
rect 15393 14433 15427 14467
rect 15761 14433 15795 14467
rect 16028 14433 16062 14467
rect 17233 14433 17267 14467
rect 17500 14433 17534 14467
rect 18705 14433 18739 14467
rect 20361 14433 20395 14467
rect 3341 14365 3375 14399
rect 3433 14365 3467 14399
rect 4537 14365 4571 14399
rect 4629 14365 4663 14399
rect 5549 14365 5583 14399
rect 9413 14365 9447 14399
rect 13553 14365 13587 14399
rect 4077 14297 4111 14331
rect 14933 14297 14967 14331
rect 3709 14229 3743 14263
rect 8677 14229 8711 14263
rect 8769 14229 8803 14263
rect 9873 14229 9907 14263
rect 11713 14229 11747 14263
rect 15577 14229 15611 14263
rect 17141 14229 17175 14263
rect 18613 14229 18647 14263
rect 20545 14229 20579 14263
rect 3065 14025 3099 14059
rect 3341 14025 3375 14059
rect 4997 14025 5031 14059
rect 5825 14025 5859 14059
rect 7481 14025 7515 14059
rect 10609 14025 10643 14059
rect 12817 14025 12851 14059
rect 15025 14025 15059 14059
rect 15301 14025 15335 14059
rect 16865 13957 16899 13991
rect 1685 13889 1719 13923
rect 3525 13889 3559 13923
rect 5549 13889 5583 13923
rect 6377 13889 6411 13923
rect 7941 13889 7975 13923
rect 8125 13889 8159 13923
rect 9232 13889 9266 13923
rect 9505 13889 9539 13923
rect 13185 13889 13219 13923
rect 13691 13889 13725 13923
rect 15485 13889 15519 13923
rect 17417 13889 17451 13923
rect 17601 13889 17635 13923
rect 18705 13889 18739 13923
rect 18889 13889 18923 13923
rect 3157 13821 3191 13855
rect 3792 13821 3826 13855
rect 5457 13821 5491 13855
rect 6193 13821 6227 13855
rect 6929 13821 6963 13855
rect 7113 13821 7147 13855
rect 7297 13821 7331 13855
rect 8309 13821 8343 13855
rect 8769 13821 8803 13855
rect 10701 13821 10735 13855
rect 10968 13821 11002 13855
rect 13001 13821 13035 13855
rect 13921 13821 13955 13855
rect 15117 13821 15151 13855
rect 15752 13821 15786 13855
rect 19073 13821 19107 13855
rect 19340 13821 19374 13855
rect 1952 13753 1986 13787
rect 7849 13753 7883 13787
rect 17325 13753 17359 13787
rect 4905 13685 4939 13719
rect 5365 13685 5399 13719
rect 6285 13685 6319 13719
rect 8493 13685 8527 13719
rect 9235 13685 9269 13719
rect 12081 13685 12115 13719
rect 12449 13685 12483 13719
rect 13651 13685 13685 13719
rect 16957 13685 16991 13719
rect 18245 13685 18279 13719
rect 18613 13685 18647 13719
rect 20453 13685 20487 13719
rect 3709 13481 3743 13515
rect 6469 13481 6503 13515
rect 8217 13481 8251 13515
rect 9229 13481 9263 13515
rect 12633 13481 12667 13515
rect 14933 13481 14967 13515
rect 16037 13481 16071 13515
rect 16773 13481 16807 13515
rect 18061 13481 18095 13515
rect 4721 13413 4755 13447
rect 5356 13413 5390 13447
rect 7757 13413 7791 13447
rect 8585 13413 8619 13447
rect 11520 13413 11554 13447
rect 17141 13413 17175 13447
rect 1676 13345 1710 13379
rect 3249 13345 3283 13379
rect 3893 13345 3927 13379
rect 4629 13345 4663 13379
rect 6929 13345 6963 13379
rect 9045 13345 9079 13379
rect 9945 13345 9979 13379
rect 11253 13345 11287 13379
rect 12725 13345 12759 13379
rect 13093 13345 13127 13379
rect 13461 13345 13495 13379
rect 13728 13345 13762 13379
rect 15117 13345 15151 13379
rect 15301 13345 15335 13379
rect 16681 13345 16715 13379
rect 17969 13345 18003 13379
rect 18797 13345 18831 13379
rect 19625 13345 19659 13379
rect 20085 13345 20119 13379
rect 1409 13277 1443 13311
rect 3341 13277 3375 13311
rect 3525 13277 3559 13311
rect 4813 13277 4847 13311
rect 5089 13277 5123 13311
rect 7021 13277 7055 13311
rect 7205 13277 7239 13311
rect 7849 13277 7883 13311
rect 8033 13277 8067 13311
rect 8677 13277 8711 13311
rect 8769 13277 8803 13311
rect 9689 13277 9723 13311
rect 16129 13277 16163 13311
rect 16313 13277 16347 13311
rect 17233 13277 17267 13311
rect 17417 13277 17451 13311
rect 18245 13277 18279 13311
rect 18889 13277 18923 13311
rect 18981 13277 19015 13311
rect 19717 13277 19751 13311
rect 19809 13277 19843 13311
rect 2881 13209 2915 13243
rect 6561 13209 6595 13243
rect 14841 13209 14875 13243
rect 15485 13209 15519 13243
rect 17601 13209 17635 13243
rect 20269 13209 20303 13243
rect 2789 13141 2823 13175
rect 4261 13141 4295 13175
rect 7389 13141 7423 13175
rect 11069 13141 11103 13175
rect 12909 13141 12943 13175
rect 13277 13141 13311 13175
rect 15669 13141 15703 13175
rect 16497 13141 16531 13175
rect 18429 13141 18463 13175
rect 19257 13141 19291 13175
rect 2881 12937 2915 12971
rect 4353 12937 4387 12971
rect 5825 12937 5859 12971
rect 5917 12937 5951 12971
rect 10793 12937 10827 12971
rect 14473 12937 14507 12971
rect 16773 12937 16807 12971
rect 17785 12937 17819 12971
rect 9965 12869 9999 12903
rect 14289 12869 14323 12903
rect 16681 12869 16715 12903
rect 4445 12801 4479 12835
rect 6377 12801 6411 12835
rect 6469 12801 6503 12835
rect 6837 12801 6871 12835
rect 8309 12801 8343 12835
rect 10517 12801 10551 12835
rect 12081 12801 12115 12835
rect 12909 12801 12943 12835
rect 15117 12801 15151 12835
rect 17325 12801 17359 12835
rect 18797 12801 18831 12835
rect 19073 12801 19107 12835
rect 1501 12733 1535 12767
rect 2973 12733 3007 12767
rect 3240 12733 3274 12767
rect 4712 12733 4746 12767
rect 7104 12733 7138 12767
rect 10977 12733 11011 12767
rect 11897 12733 11931 12767
rect 15301 12733 15335 12767
rect 17601 12733 17635 12767
rect 18521 12733 18555 12767
rect 19340 12733 19374 12767
rect 1768 12665 1802 12699
rect 6285 12665 6319 12699
rect 8576 12665 8610 12699
rect 10425 12665 10459 12699
rect 11069 12665 11103 12699
rect 11253 12665 11287 12699
rect 13176 12665 13210 12699
rect 14841 12665 14875 12699
rect 15568 12665 15602 12699
rect 8217 12597 8251 12631
rect 9689 12597 9723 12631
rect 10333 12597 10367 12631
rect 11437 12597 11471 12631
rect 11529 12597 11563 12631
rect 11989 12597 12023 12631
rect 12449 12597 12483 12631
rect 12817 12597 12851 12631
rect 14933 12597 14967 12631
rect 17141 12597 17175 12631
rect 17233 12597 17267 12631
rect 18153 12597 18187 12631
rect 18613 12597 18647 12631
rect 20453 12597 20487 12631
rect 2789 12393 2823 12427
rect 3157 12393 3191 12427
rect 5549 12393 5583 12427
rect 5825 12393 5859 12427
rect 7665 12393 7699 12427
rect 9413 12393 9447 12427
rect 9689 12393 9723 12427
rect 14381 12393 14415 12427
rect 15025 12393 15059 12427
rect 18613 12393 18647 12427
rect 1676 12325 1710 12359
rect 3525 12325 3559 12359
rect 6552 12325 6586 12359
rect 17969 12325 18003 12359
rect 19156 12325 19190 12359
rect 1409 12257 1443 12291
rect 3065 12257 3099 12291
rect 3617 12257 3651 12291
rect 4436 12257 4470 12291
rect 5641 12257 5675 12291
rect 6193 12257 6227 12291
rect 7941 12257 7975 12291
rect 8033 12257 8067 12291
rect 8289 12257 8323 12291
rect 10057 12257 10091 12291
rect 10609 12257 10643 12291
rect 10932 12257 10966 12291
rect 12864 12257 12898 12291
rect 13277 12257 13311 12291
rect 14473 12257 14507 12291
rect 14841 12257 14875 12291
rect 15568 12257 15602 12291
rect 17141 12257 17175 12291
rect 18429 12257 18463 12291
rect 3709 12189 3743 12223
rect 4169 12189 4203 12223
rect 6285 12189 6319 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 11072 12189 11106 12223
rect 11345 12189 11379 12223
rect 12541 12189 12575 12223
rect 13004 12189 13038 12223
rect 15301 12189 15335 12223
rect 17233 12189 17267 12223
rect 17417 12189 17451 12223
rect 18061 12189 18095 12223
rect 18153 12189 18187 12223
rect 18889 12189 18923 12223
rect 20361 12189 20395 12223
rect 2881 12121 2915 12155
rect 7757 12121 7791 12155
rect 16773 12121 16807 12155
rect 6009 12053 6043 12087
rect 12449 12053 12483 12087
rect 14657 12053 14691 12087
rect 16681 12053 16715 12087
rect 17601 12053 17635 12087
rect 20269 12053 20303 12087
rect 3709 11849 3743 11883
rect 5365 11849 5399 11883
rect 5917 11849 5951 11883
rect 10517 11849 10551 11883
rect 14013 11849 14047 11883
rect 17877 11849 17911 11883
rect 1869 11781 1903 11815
rect 5733 11781 5767 11815
rect 8309 11781 8343 11815
rect 16313 11781 16347 11815
rect 2513 11713 2547 11747
rect 3341 11713 3375 11747
rect 6561 11713 6595 11747
rect 8861 11713 8895 11747
rect 9965 11713 9999 11747
rect 10701 11713 10735 11747
rect 12541 11713 12575 11747
rect 14565 11713 14599 11747
rect 20269 11713 20303 11747
rect 20361 11713 20395 11747
rect 3525 11645 3559 11679
rect 3985 11645 4019 11679
rect 5549 11645 5583 11679
rect 6844 11645 6878 11679
rect 8677 11645 8711 11679
rect 8769 11645 8803 11679
rect 10333 11645 10367 11679
rect 10968 11645 11002 11679
rect 14381 11645 14415 11679
rect 14933 11645 14967 11679
rect 15200 11645 15234 11679
rect 16497 11645 16531 11679
rect 18061 11645 18095 11679
rect 18317 11645 18351 11679
rect 20177 11645 20211 11679
rect 2237 11577 2271 11611
rect 3065 11577 3099 11611
rect 4252 11577 4286 11611
rect 6285 11577 6319 11611
rect 7104 11577 7138 11611
rect 12808 11577 12842 11611
rect 16764 11577 16798 11611
rect 2329 11509 2363 11543
rect 2697 11509 2731 11543
rect 3157 11509 3191 11543
rect 6377 11509 6411 11543
rect 8217 11509 8251 11543
rect 9321 11509 9355 11543
rect 9689 11509 9723 11543
rect 9781 11509 9815 11543
rect 12081 11509 12115 11543
rect 13921 11509 13955 11543
rect 14473 11509 14507 11543
rect 19441 11509 19475 11543
rect 19809 11509 19843 11543
rect 2881 11305 2915 11339
rect 3709 11305 3743 11339
rect 5457 11305 5491 11339
rect 5917 11305 5951 11339
rect 7941 11305 7975 11339
rect 8309 11305 8343 11339
rect 8401 11305 8435 11339
rect 8769 11305 8803 11339
rect 11345 11305 11379 11339
rect 12265 11305 12299 11339
rect 14749 11305 14783 11339
rect 16681 11305 16715 11339
rect 17233 11305 17267 11339
rect 20545 11305 20579 11339
rect 12633 11237 12667 11271
rect 13360 11237 13394 11271
rect 17684 11237 17718 11271
rect 19432 11237 19466 11271
rect 1665 11169 1699 11203
rect 3249 11169 3283 11203
rect 3893 11169 3927 11203
rect 4344 11169 4378 11203
rect 5733 11169 5767 11203
rect 6368 11169 6402 11203
rect 7573 11169 7607 11203
rect 9137 11169 9171 11203
rect 9965 11169 9999 11203
rect 10232 11169 10266 11203
rect 11805 11169 11839 11203
rect 12725 11169 12759 11203
rect 14565 11169 14599 11203
rect 15117 11169 15151 11203
rect 15568 11169 15602 11203
rect 16957 11169 16991 11203
rect 17049 11169 17083 11203
rect 1409 11101 1443 11135
rect 3341 11101 3375 11135
rect 3433 11101 3467 11135
rect 4077 11101 4111 11135
rect 6101 11101 6135 11135
rect 8493 11101 8527 11135
rect 9229 11101 9263 11135
rect 9413 11101 9447 11135
rect 9689 11101 9723 11135
rect 11897 11101 11931 11135
rect 12081 11101 12115 11135
rect 12817 11101 12851 11135
rect 13093 11101 13127 11135
rect 15301 11101 15335 11135
rect 17417 11101 17451 11135
rect 18889 11101 18923 11135
rect 19165 11101 19199 11135
rect 2789 11033 2823 11067
rect 7757 11033 7791 11067
rect 14473 11033 14507 11067
rect 16773 11033 16807 11067
rect 7481 10965 7515 10999
rect 11437 10965 11471 10999
rect 14933 10965 14967 10999
rect 18797 10965 18831 10999
rect 2789 10761 2823 10795
rect 4261 10761 4295 10795
rect 5733 10761 5767 10795
rect 6837 10761 6871 10795
rect 7665 10761 7699 10795
rect 10057 10761 10091 10795
rect 11621 10761 11655 10795
rect 13829 10761 13863 10795
rect 16773 10761 16807 10795
rect 19441 10693 19475 10727
rect 6285 10625 6319 10659
rect 6469 10625 6503 10659
rect 7481 10625 7515 10659
rect 8309 10625 8343 10659
rect 12449 10625 12483 10659
rect 13921 10625 13955 10659
rect 17325 10625 17359 10659
rect 17417 10625 17451 10659
rect 20085 10625 20119 10659
rect 1409 10557 1443 10591
rect 1676 10557 1710 10591
rect 2881 10557 2915 10591
rect 3148 10557 3182 10591
rect 4353 10557 4387 10591
rect 4609 10557 4643 10591
rect 7205 10557 7239 10591
rect 8677 10557 8711 10591
rect 12705 10557 12739 10591
rect 14188 10557 14222 10591
rect 15393 10557 15427 10591
rect 17233 10557 17267 10591
rect 17877 10557 17911 10591
rect 18061 10557 18095 10591
rect 20361 10557 20395 10591
rect 8125 10489 8159 10523
rect 8922 10489 8956 10523
rect 10333 10489 10367 10523
rect 15660 10489 15694 10523
rect 18328 10489 18362 10523
rect 5825 10421 5859 10455
rect 6193 10421 6227 10455
rect 7297 10421 7331 10455
rect 8033 10421 8067 10455
rect 15301 10421 15335 10455
rect 16865 10421 16899 10455
rect 17693 10421 17727 10455
rect 19533 10421 19567 10455
rect 19901 10421 19935 10455
rect 19993 10421 20027 10455
rect 3157 10217 3191 10251
rect 5549 10217 5583 10251
rect 6745 10217 6779 10251
rect 7021 10217 7055 10251
rect 7849 10217 7883 10251
rect 8769 10217 8803 10251
rect 11989 10217 12023 10251
rect 17417 10217 17451 10251
rect 20269 10217 20303 10251
rect 2044 10149 2078 10183
rect 4344 10149 4378 10183
rect 10394 10149 10428 10183
rect 12081 10149 12115 10183
rect 15761 10149 15795 10183
rect 15945 10149 15979 10183
rect 1777 10081 1811 10115
rect 3893 10081 3927 10115
rect 5917 10081 5951 10115
rect 6561 10081 6595 10115
rect 7389 10081 7423 10115
rect 8217 10081 8251 10115
rect 8309 10081 8343 10115
rect 9137 10081 9171 10115
rect 9229 10081 9263 10115
rect 9689 10081 9723 10115
rect 9781 10081 9815 10115
rect 12449 10081 12483 10115
rect 12909 10081 12943 10115
rect 14749 10081 14783 10115
rect 15577 10081 15611 10115
rect 16304 10081 16338 10115
rect 17509 10081 17543 10115
rect 17877 10081 17911 10115
rect 20177 10081 20211 10115
rect 4077 10013 4111 10047
rect 6009 10013 6043 10047
rect 6193 10013 6227 10047
rect 7481 10013 7515 10047
rect 7665 10013 7699 10047
rect 8493 10013 8527 10047
rect 9413 10013 9447 10047
rect 10149 10013 10183 10047
rect 12173 10013 12207 10047
rect 15301 10013 15335 10047
rect 16037 10013 16071 10047
rect 18200 10013 18234 10047
rect 18383 10013 18417 10047
rect 18613 10013 18647 10047
rect 20361 10013 20395 10047
rect 9689 9945 9723 9979
rect 9965 9945 9999 9979
rect 11529 9945 11563 9979
rect 12633 9945 12667 9979
rect 14933 9945 14967 9979
rect 3709 9877 3743 9911
rect 5457 9877 5491 9911
rect 11621 9877 11655 9911
rect 14197 9877 14231 9911
rect 17693 9877 17727 9911
rect 19717 9877 19751 9911
rect 19809 9877 19843 9911
rect 6837 9673 6871 9707
rect 10701 9673 10735 9707
rect 12265 9673 12299 9707
rect 15117 9673 15151 9707
rect 1777 9605 1811 9639
rect 2973 9605 3007 9639
rect 6653 9605 6687 9639
rect 9229 9605 9263 9639
rect 2421 9537 2455 9571
rect 3617 9537 3651 9571
rect 5273 9537 5307 9571
rect 7389 9537 7423 9571
rect 7849 9537 7883 9571
rect 13461 9605 13495 9639
rect 18429 9605 18463 9639
rect 13093 9537 13127 9571
rect 15393 9537 15427 9571
rect 17509 9537 17543 9571
rect 18613 9537 18647 9571
rect 2145 9469 2179 9503
rect 3801 9469 3835 9503
rect 4068 9469 4102 9503
rect 9321 9469 9355 9503
rect 9577 9469 9611 9503
rect 10793 9469 10827 9503
rect 12357 9469 12391 9503
rect 13277 9469 13311 9503
rect 13737 9469 13771 9503
rect 14004 9469 14038 9503
rect 15660 9469 15694 9503
rect 17877 9469 17911 9503
rect 18245 9469 18279 9503
rect 20085 9469 20119 9503
rect 2237 9401 2271 9435
rect 5540 9401 5574 9435
rect 7205 9401 7239 9435
rect 8116 9401 8150 9435
rect 11060 9401 11094 9435
rect 12909 9401 12943 9435
rect 18858 9401 18892 9435
rect 2881 9333 2915 9367
rect 3341 9333 3375 9367
rect 3433 9333 3467 9367
rect 5181 9333 5215 9367
rect 7297 9333 7331 9367
rect 12173 9333 12207 9367
rect 12449 9333 12483 9367
rect 12817 9333 12851 9367
rect 16773 9333 16807 9367
rect 16865 9333 16899 9367
rect 17233 9333 17267 9367
rect 17325 9333 17359 9367
rect 17693 9333 17727 9367
rect 19993 9333 20027 9367
rect 20269 9333 20303 9367
rect 2697 9129 2731 9163
rect 4077 9129 4111 9163
rect 5733 9129 5767 9163
rect 7205 9129 7239 9163
rect 8677 9129 8711 9163
rect 12449 9129 12483 9163
rect 13921 9129 13955 9163
rect 14197 9129 14231 9163
rect 17969 9129 18003 9163
rect 18061 9129 18095 9163
rect 18613 9129 18647 9163
rect 3617 9061 3651 9095
rect 4620 9061 4654 9095
rect 6092 9061 6126 9095
rect 7564 9061 7598 9095
rect 10701 9061 10735 9095
rect 12786 9061 12820 9095
rect 15568 9061 15602 9095
rect 2789 8993 2823 9027
rect 3525 8993 3559 9027
rect 4261 8993 4295 9027
rect 4353 8993 4387 9027
rect 5825 8993 5859 9027
rect 7297 8993 7331 9027
rect 9137 8993 9171 9027
rect 9689 8993 9723 9027
rect 10609 8993 10643 9027
rect 11069 8993 11103 9027
rect 11336 8993 11370 9027
rect 14013 8993 14047 9027
rect 14749 8993 14783 9027
rect 14841 8993 14875 9027
rect 17141 8993 17175 9027
rect 18429 8993 18463 9027
rect 18797 8993 18831 9027
rect 19432 8993 19466 9027
rect 2881 8925 2915 8959
rect 3801 8925 3835 8959
rect 9229 8925 9263 8959
rect 9321 8925 9355 8959
rect 10885 8925 10919 8959
rect 12541 8925 12575 8959
rect 15025 8925 15059 8959
rect 15301 8925 15335 8959
rect 17233 8925 17267 8959
rect 17325 8925 17359 8959
rect 18153 8925 18187 8959
rect 19165 8925 19199 8959
rect 16773 8857 16807 8891
rect 2329 8789 2363 8823
rect 3157 8789 3191 8823
rect 8769 8789 8803 8823
rect 9873 8789 9907 8823
rect 10241 8789 10275 8823
rect 14381 8789 14415 8823
rect 16681 8789 16715 8823
rect 17601 8789 17635 8823
rect 18981 8789 19015 8823
rect 20545 8789 20579 8823
rect 2421 8585 2455 8619
rect 4077 8585 4111 8619
rect 6285 8585 6319 8619
rect 8309 8585 8343 8619
rect 10057 8585 10091 8619
rect 13277 8585 13311 8619
rect 15117 8585 15151 8619
rect 16957 8585 16991 8619
rect 19901 8585 19935 8619
rect 3249 8517 3283 8551
rect 6469 8517 6503 8551
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 3893 8449 3927 8483
rect 4537 8449 4571 8483
rect 4721 8449 4755 8483
rect 6929 8449 6963 8483
rect 8493 8449 8527 8483
rect 11529 8517 11563 8551
rect 12173 8517 12207 8551
rect 12449 8517 12483 8551
rect 14105 8517 14139 8551
rect 15393 8517 15427 8551
rect 10149 8449 10183 8483
rect 13093 8449 13127 8483
rect 13829 8449 13863 8483
rect 14657 8449 14691 8483
rect 2789 8381 2823 8415
rect 3709 8381 3743 8415
rect 4445 8381 4479 8415
rect 4905 8381 4939 8415
rect 5172 8381 5206 8415
rect 6653 8381 6687 8415
rect 10057 8381 10091 8415
rect 11621 8381 11655 8415
rect 11989 8381 12023 8415
rect 14473 8381 14507 8415
rect 14933 8381 14967 8415
rect 3617 8313 3651 8347
rect 7196 8313 7230 8347
rect 8760 8313 8794 8347
rect 10416 8313 10450 8347
rect 12817 8313 12851 8347
rect 15485 8449 15519 8483
rect 17509 8449 17543 8483
rect 18061 8449 18095 8483
rect 18524 8449 18558 8483
rect 15752 8381 15786 8415
rect 17417 8381 17451 8415
rect 18384 8381 18418 8415
rect 18797 8381 18831 8415
rect 20177 8313 20211 8347
rect 20361 8313 20395 8347
rect 9873 8245 9907 8279
rect 11805 8245 11839 8279
rect 12909 8245 12943 8279
rect 13645 8245 13679 8279
rect 13737 8245 13771 8279
rect 14565 8245 14599 8279
rect 15393 8245 15427 8279
rect 16865 8245 16899 8279
rect 17325 8245 17359 8279
rect 5089 8041 5123 8075
rect 5457 8041 5491 8075
rect 6745 8041 6779 8075
rect 9689 8041 9723 8075
rect 11161 8041 11195 8075
rect 11253 8041 11287 8075
rect 12081 8041 12115 8075
rect 13645 8041 13679 8075
rect 15117 8041 15151 8075
rect 15669 8041 15703 8075
rect 15761 8041 15795 8075
rect 16129 8041 16163 8075
rect 20545 8041 20579 8075
rect 21005 8041 21039 8075
rect 3525 7973 3559 8007
rect 5825 7973 5859 8007
rect 7665 7973 7699 8007
rect 3617 7905 3651 7939
rect 4997 7905 5031 7939
rect 6653 7905 6687 7939
rect 7757 7905 7791 7939
rect 8125 7905 8159 7939
rect 8392 7905 8426 7939
rect 3801 7837 3835 7871
rect 5273 7837 5307 7871
rect 5917 7837 5951 7871
rect 6101 7837 6135 7871
rect 6837 7837 6871 7871
rect 7941 7837 7975 7871
rect 11621 7973 11655 8007
rect 10048 7905 10082 7939
rect 12532 7973 12566 8007
rect 14004 7905 14038 7939
rect 16405 7905 16439 7939
rect 16728 7905 16762 7939
rect 17141 7905 17175 7939
rect 18705 7905 18739 7939
rect 19165 7905 19199 7939
rect 19432 7905 19466 7939
rect 9781 7837 9815 7871
rect 11713 7837 11747 7871
rect 11897 7837 11931 7871
rect 12081 7837 12115 7871
rect 12265 7837 12299 7871
rect 13737 7837 13771 7871
rect 15945 7837 15979 7871
rect 16911 7837 16945 7871
rect 18797 7837 18831 7871
rect 18889 7837 18923 7871
rect 3157 7701 3191 7735
rect 4629 7701 4663 7735
rect 6285 7701 6319 7735
rect 7297 7701 7331 7735
rect 9505 7701 9539 7735
rect 9689 7701 9723 7735
rect 15301 7701 15335 7735
rect 18245 7701 18279 7735
rect 18337 7701 18371 7735
rect 4445 7497 4479 7531
rect 8585 7497 8619 7531
rect 12265 7497 12299 7531
rect 13829 7497 13863 7531
rect 17785 7497 17819 7531
rect 3617 7429 3651 7463
rect 19533 7429 19567 7463
rect 4077 7361 4111 7395
rect 4261 7361 4295 7395
rect 5089 7361 5123 7395
rect 5273 7361 5307 7395
rect 6837 7361 6871 7395
rect 9229 7361 9263 7395
rect 9413 7361 9447 7395
rect 14013 7361 14047 7395
rect 14519 7361 14553 7395
rect 16129 7361 16163 7395
rect 19993 7361 20027 7395
rect 20085 7361 20119 7395
rect 4905 7293 4939 7327
rect 8493 7293 8527 7327
rect 9669 7293 9703 7327
rect 10885 7293 10919 7327
rect 12449 7293 12483 7327
rect 14749 7293 14783 7327
rect 16396 7293 16430 7327
rect 17601 7293 17635 7327
rect 18061 7293 18095 7327
rect 18328 7293 18362 7327
rect 3525 7225 3559 7259
rect 3985 7225 4019 7259
rect 5540 7225 5574 7259
rect 7082 7225 7116 7259
rect 8953 7225 8987 7259
rect 11152 7225 11186 7259
rect 12716 7225 12750 7259
rect 19901 7225 19935 7259
rect 20361 7225 20395 7259
rect 4813 7157 4847 7191
rect 6653 7157 6687 7191
rect 8217 7157 8251 7191
rect 8309 7157 8343 7191
rect 9045 7157 9079 7191
rect 10793 7157 10827 7191
rect 14479 7157 14513 7191
rect 15853 7157 15887 7191
rect 17509 7157 17543 7191
rect 19441 7157 19475 7191
rect 6285 6953 6319 6987
rect 8493 6953 8527 6987
rect 9873 6953 9907 6987
rect 11437 6953 11471 6987
rect 13369 6953 13403 6987
rect 15025 6953 15059 6987
rect 15117 6953 15151 6987
rect 15761 6953 15795 6987
rect 16589 6953 16623 6987
rect 16681 6953 16715 6987
rect 18429 6953 18463 6987
rect 7380 6885 7414 6919
rect 9137 6885 9171 6919
rect 5172 6817 5206 6851
rect 6561 6817 6595 6851
rect 6653 6817 6687 6851
rect 6837 6817 6871 6851
rect 8677 6817 8711 6851
rect 9689 6817 9723 6851
rect 10324 6817 10358 6851
rect 11529 6817 11563 6851
rect 11785 6817 11819 6851
rect 13001 6817 13035 6851
rect 13553 6817 13587 6851
rect 13912 6817 13946 6851
rect 4905 6749 4939 6783
rect 7113 6749 7147 6783
rect 17316 6885 17350 6919
rect 19533 6885 19567 6919
rect 21005 6885 21039 6919
rect 15669 6817 15703 6851
rect 18705 6817 18739 6851
rect 18797 6817 18831 6851
rect 19993 6817 20027 6851
rect 9229 6749 9263 6783
rect 9413 6749 9447 6783
rect 10057 6749 10091 6783
rect 13645 6749 13679 6783
rect 15117 6749 15151 6783
rect 15853 6749 15887 6783
rect 16865 6749 16899 6783
rect 17049 6749 17083 6783
rect 19625 6749 19659 6783
rect 19717 6749 19751 6783
rect 12909 6681 12943 6715
rect 15301 6681 15335 6715
rect 20177 6681 20211 6715
rect 21005 6681 21039 6715
rect 6377 6613 6411 6647
rect 7021 6613 7055 6647
rect 8677 6613 8711 6647
rect 8769 6613 8803 6647
rect 13185 6613 13219 6647
rect 16221 6613 16255 6647
rect 18521 6613 18555 6647
rect 18981 6613 19015 6647
rect 19165 6613 19199 6647
rect 5917 6409 5951 6443
rect 6837 6409 6871 6443
rect 12633 6409 12667 6443
rect 20545 6409 20579 6443
rect 6561 6341 6595 6375
rect 11989 6341 12023 6375
rect 18429 6341 18463 6375
rect 7481 6273 7515 6307
rect 13461 6273 13495 6307
rect 15761 6273 15795 6307
rect 16589 6273 16623 6307
rect 17417 6273 17451 6307
rect 18705 6273 18739 6307
rect 4537 6205 4571 6239
rect 6009 6205 6043 6239
rect 6377 6205 6411 6239
rect 7665 6205 7699 6239
rect 9137 6205 9171 6239
rect 10609 6205 10643 6239
rect 12081 6205 12115 6239
rect 12449 6205 12483 6239
rect 13645 6205 13679 6239
rect 16405 6205 16439 6239
rect 18061 6205 18095 6239
rect 18613 6205 18647 6239
rect 20177 6205 20211 6239
rect 4804 6137 4838 6171
rect 7932 6137 7966 6171
rect 9404 6137 9438 6171
rect 10876 6137 10910 6171
rect 13912 6137 13946 6171
rect 16497 6137 16531 6171
rect 17233 6137 17267 6171
rect 17693 6137 17727 6171
rect 18972 6137 19006 6171
rect 20361 6137 20395 6171
rect 6193 6069 6227 6103
rect 7205 6069 7239 6103
rect 7297 6069 7331 6103
rect 9045 6069 9079 6103
rect 10517 6069 10551 6103
rect 12817 6069 12851 6103
rect 13185 6069 13219 6103
rect 13277 6069 13311 6103
rect 15025 6069 15059 6103
rect 15209 6069 15243 6103
rect 15577 6069 15611 6103
rect 15669 6069 15703 6103
rect 16037 6069 16071 6103
rect 16865 6069 16899 6103
rect 17325 6069 17359 6103
rect 18245 6069 18279 6103
rect 20085 6069 20119 6103
rect 3617 5865 3651 5899
rect 4261 5865 4295 5899
rect 5917 5865 5951 5899
rect 6745 5865 6779 5899
rect 9505 5865 9539 5899
rect 17141 5865 17175 5899
rect 19533 5865 19567 5899
rect 19993 5865 20027 5899
rect 3525 5797 3559 5831
rect 7665 5797 7699 5831
rect 17233 5797 17267 5831
rect 4445 5729 4479 5763
rect 4537 5729 4571 5763
rect 4804 5729 4838 5763
rect 6009 5729 6043 5763
rect 7573 5729 7607 5763
rect 8125 5729 8159 5763
rect 8392 5729 8426 5763
rect 10149 5729 10183 5763
rect 10977 5729 11011 5763
rect 13268 5729 13302 5763
rect 14657 5729 14691 5763
rect 14841 5729 14875 5763
rect 15568 5729 15602 5763
rect 17601 5729 17635 5763
rect 18420 5729 18454 5763
rect 20085 5729 20119 5763
rect 3801 5661 3835 5695
rect 6837 5661 6871 5695
rect 6929 5661 6963 5695
rect 7849 5661 7883 5695
rect 10241 5661 10275 5695
rect 10333 5661 10367 5695
rect 11069 5661 11103 5695
rect 11392 5661 11426 5695
rect 11575 5661 11609 5695
rect 11805 5661 11839 5695
rect 13001 5661 13035 5695
rect 15301 5661 15335 5695
rect 17417 5661 17451 5695
rect 18153 5661 18187 5695
rect 20269 5661 20303 5695
rect 21005 5661 21039 5695
rect 3157 5593 3191 5627
rect 6193 5593 6227 5627
rect 16773 5593 16807 5627
rect 6377 5525 6411 5559
rect 7205 5525 7239 5559
rect 9781 5525 9815 5559
rect 10793 5525 10827 5559
rect 12909 5525 12943 5559
rect 14381 5525 14415 5559
rect 14473 5525 14507 5559
rect 15025 5525 15059 5559
rect 16681 5525 16715 5559
rect 17785 5525 17819 5559
rect 19625 5525 19659 5559
rect 6009 5321 6043 5355
rect 6469 5321 6503 5355
rect 7297 5321 7331 5355
rect 8125 5321 8159 5355
rect 10701 5321 10735 5355
rect 12449 5321 12483 5355
rect 19441 5321 19475 5355
rect 19533 5321 19567 5355
rect 7849 5185 7883 5219
rect 8677 5185 8711 5219
rect 9321 5185 9355 5219
rect 10793 5185 10827 5219
rect 11989 5185 12023 5219
rect 13001 5185 13035 5219
rect 13277 5185 13311 5219
rect 17693 5185 17727 5219
rect 19993 5185 20027 5219
rect 20085 5185 20119 5219
rect 4629 5117 4663 5151
rect 6285 5117 6319 5151
rect 6929 5117 6963 5151
rect 8953 5117 8987 5151
rect 9588 5117 9622 5151
rect 12909 5117 12943 5151
rect 13645 5117 13679 5151
rect 13912 5117 13946 5151
rect 15117 5117 15151 5151
rect 15669 5117 15703 5151
rect 15936 5117 15970 5151
rect 17601 5117 17635 5151
rect 18061 5117 18095 5151
rect 19901 5117 19935 5151
rect 4896 5049 4930 5083
rect 8585 5049 8619 5083
rect 11897 5049 11931 5083
rect 18328 5049 18362 5083
rect 7113 4981 7147 5015
rect 7665 4981 7699 5015
rect 7757 4981 7791 5015
rect 8493 4981 8527 5015
rect 9137 4981 9171 5015
rect 11437 4981 11471 5015
rect 11805 4981 11839 5015
rect 12817 4981 12851 5015
rect 15025 4981 15059 5015
rect 15301 4981 15335 5015
rect 17049 4981 17083 5015
rect 17141 4981 17175 5015
rect 17509 4981 17543 5015
rect 6009 4777 6043 4811
rect 6469 4777 6503 4811
rect 6837 4777 6871 4811
rect 7205 4777 7239 4811
rect 7849 4777 7883 4811
rect 8401 4777 8435 4811
rect 12081 4777 12115 4811
rect 12633 4777 12667 4811
rect 13001 4777 13035 4811
rect 15669 4777 15703 4811
rect 17509 4777 17543 4811
rect 20545 4777 20579 4811
rect 4804 4709 4838 4743
rect 7297 4709 7331 4743
rect 8493 4709 8527 4743
rect 13093 4709 13127 4743
rect 15761 4709 15795 4743
rect 19432 4709 19466 4743
rect 4537 4641 4571 4675
rect 6377 4641 6411 4675
rect 7665 4641 7699 4675
rect 8861 4641 8895 4675
rect 9321 4641 9355 4675
rect 10012 4641 10046 4675
rect 10425 4641 10459 4675
rect 11989 4641 12023 4675
rect 13461 4641 13495 4675
rect 13728 4641 13762 4675
rect 15117 4641 15151 4675
rect 16385 4641 16419 4675
rect 17857 4641 17891 4675
rect 6653 4573 6687 4607
rect 7389 4573 7423 4607
rect 8677 4573 8711 4607
rect 9689 4573 9723 4607
rect 10152 4573 10186 4607
rect 12173 4573 12207 4607
rect 13185 4573 13219 4607
rect 15853 4573 15887 4607
rect 16129 4573 16163 4607
rect 17601 4573 17635 4607
rect 19165 4573 19199 4607
rect 5917 4505 5951 4539
rect 9137 4505 9171 4539
rect 11621 4505 11655 4539
rect 14933 4505 14967 4539
rect 8033 4437 8067 4471
rect 11529 4437 11563 4471
rect 14841 4437 14875 4471
rect 15301 4437 15335 4471
rect 18981 4437 19015 4471
rect 5825 4233 5859 4267
rect 5917 4233 5951 4267
rect 6837 4233 6871 4267
rect 7849 4233 7883 4267
rect 11345 4233 11379 4267
rect 14197 4233 14231 4267
rect 15025 4233 15059 4267
rect 16129 4233 16163 4267
rect 20545 4233 20579 4267
rect 9781 4165 9815 4199
rect 18061 4165 18095 4199
rect 6377 4097 6411 4131
rect 6561 4097 6595 4131
rect 7389 4097 7423 4131
rect 11989 4097 12023 4131
rect 14749 4097 14783 4131
rect 15485 4097 15519 4131
rect 15577 4097 15611 4131
rect 16957 4097 16991 4131
rect 17785 4097 17819 4131
rect 18613 4097 18647 4131
rect 4445 4029 4479 4063
rect 4712 4029 4746 4063
rect 6285 4029 6319 4063
rect 7665 4029 7699 4063
rect 8401 4029 8435 4063
rect 9873 4029 9907 4063
rect 11713 4029 11747 4063
rect 12449 4029 12483 4063
rect 12716 4029 12750 4063
rect 15945 4029 15979 4063
rect 18429 4029 18463 4063
rect 19165 4029 19199 4063
rect 8668 3961 8702 3995
rect 10140 3961 10174 3995
rect 11805 3961 11839 3995
rect 13921 3961 13955 3995
rect 15393 3961 15427 3995
rect 17509 3961 17543 3995
rect 19432 3961 19466 3995
rect 7205 3893 7239 3927
rect 7297 3893 7331 3927
rect 11253 3893 11287 3927
rect 13829 3893 13863 3927
rect 14565 3893 14599 3927
rect 14657 3893 14691 3927
rect 16313 3893 16347 3927
rect 16681 3893 16715 3927
rect 16773 3893 16807 3927
rect 17141 3893 17175 3927
rect 17601 3893 17635 3927
rect 18521 3893 18555 3927
rect 15025 3689 15059 3723
rect 16957 3689 16991 3723
rect 18705 3689 18739 3723
rect 20545 3689 20579 3723
rect 4712 3621 4746 3655
rect 8392 3621 8426 3655
rect 10149 3621 10183 3655
rect 4445 3553 4479 3587
rect 6193 3553 6227 3587
rect 6460 3553 6494 3587
rect 8125 3553 8159 3587
rect 10057 3553 10091 3587
rect 12725 3553 12759 3587
rect 13415 3553 13449 3587
rect 14841 3553 14875 3587
rect 15301 3553 15335 3587
rect 15844 3553 15878 3587
rect 17316 3553 17350 3587
rect 18521 3553 18555 3587
rect 19432 3553 19466 3587
rect 10333 3485 10367 3519
rect 10793 3485 10827 3519
rect 11116 3485 11150 3519
rect 11299 3485 11333 3519
rect 11529 3485 11563 3519
rect 13048 3485 13082 3519
rect 13188 3485 13222 3519
rect 15577 3485 15611 3519
rect 17049 3485 17083 3519
rect 19165 3485 19199 3519
rect 5825 3417 5859 3451
rect 7573 3417 7607 3451
rect 9689 3417 9723 3451
rect 14565 3417 14599 3451
rect 9505 3349 9539 3383
rect 12633 3349 12667 3383
rect 18429 3349 18463 3383
rect 4445 3145 4479 3179
rect 8217 3145 8251 3179
rect 9689 3145 9723 3179
rect 15301 3145 15335 3179
rect 16957 3145 16991 3179
rect 20085 3145 20119 3179
rect 11713 3077 11747 3111
rect 18521 3077 18555 3111
rect 5089 3009 5123 3043
rect 11805 3009 11839 3043
rect 17417 3009 17451 3043
rect 17601 3009 17635 3043
rect 18705 3009 18739 3043
rect 4813 2941 4847 2975
rect 5273 2941 5307 2975
rect 5540 2941 5574 2975
rect 6837 2941 6871 2975
rect 8309 2941 8343 2975
rect 8576 2941 8610 2975
rect 10333 2941 10367 2975
rect 10600 2941 10634 2975
rect 12449 2941 12483 2975
rect 12716 2941 12750 2975
rect 13921 2941 13955 2975
rect 15485 2941 15519 2975
rect 18337 2941 18371 2975
rect 7104 2873 7138 2907
rect 14166 2873 14200 2907
rect 15730 2873 15764 2907
rect 17325 2873 17359 2907
rect 18972 2873 19006 2907
rect 4905 2805 4939 2839
rect 6653 2805 6687 2839
rect 13829 2805 13863 2839
rect 16865 2805 16899 2839
rect 6469 2601 6503 2635
rect 8309 2601 8343 2635
rect 8769 2601 8803 2635
rect 11621 2601 11655 2635
rect 12173 2601 12207 2635
rect 12633 2601 12667 2635
rect 13093 2601 13127 2635
rect 15301 2601 15335 2635
rect 17325 2601 17359 2635
rect 17417 2601 17451 2635
rect 19717 2601 19751 2635
rect 19809 2601 19843 2635
rect 20269 2601 20303 2635
rect 6377 2533 6411 2567
rect 10508 2533 10542 2567
rect 12081 2533 12115 2567
rect 13461 2533 13495 2567
rect 14188 2533 14222 2567
rect 16212 2533 16246 2567
rect 20177 2533 20211 2567
rect 6929 2465 6963 2499
rect 7196 2465 7230 2499
rect 10241 2465 10275 2499
rect 13001 2465 13035 2499
rect 13921 2465 13955 2499
rect 15945 2465 15979 2499
rect 17785 2465 17819 2499
rect 17877 2465 17911 2499
rect 18604 2465 18638 2499
rect 6653 2397 6687 2431
rect 8861 2397 8895 2431
rect 9045 2397 9079 2431
rect 12357 2397 12391 2431
rect 13277 2397 13311 2431
rect 18061 2397 18095 2431
rect 18337 2397 18371 2431
rect 20361 2397 20395 2431
rect 8401 2329 8435 2363
rect 5273 2261 5307 2295
rect 6009 2261 6043 2295
rect 11713 2261 11747 2295
<< metal1 >>
rect 9490 19660 9496 19712
rect 9548 19700 9554 19712
rect 15378 19700 15384 19712
rect 9548 19672 15384 19700
rect 9548 19660 9554 19672
rect 15378 19660 15384 19672
rect 15436 19660 15442 19712
rect 16022 19660 16028 19712
rect 16080 19700 16086 19712
rect 19702 19700 19708 19712
rect 16080 19672 19708 19700
rect 16080 19660 16086 19672
rect 19702 19660 19708 19672
rect 19760 19660 19766 19712
rect 1104 19610 20884 19632
rect 1104 19558 4280 19610
rect 4332 19558 4344 19610
rect 4396 19558 4408 19610
rect 4460 19558 4472 19610
rect 4524 19558 10878 19610
rect 10930 19558 10942 19610
rect 10994 19558 11006 19610
rect 11058 19558 11070 19610
rect 11122 19558 17475 19610
rect 17527 19558 17539 19610
rect 17591 19558 17603 19610
rect 17655 19558 17667 19610
rect 17719 19558 20884 19610
rect 1104 19536 20884 19558
rect 3896 19468 5028 19496
rect 2317 19363 2375 19369
rect 2317 19329 2329 19363
rect 2363 19360 2375 19363
rect 3145 19363 3203 19369
rect 3145 19360 3157 19363
rect 2363 19332 3157 19360
rect 2363 19329 2375 19332
rect 2317 19323 2375 19329
rect 3145 19329 3157 19332
rect 3191 19360 3203 19363
rect 3896 19360 3924 19468
rect 4890 19428 4896 19440
rect 3191 19332 3924 19360
rect 3988 19400 4896 19428
rect 3191 19329 3203 19332
rect 3145 19323 3203 19329
rect 1578 19252 1584 19304
rect 1636 19292 1642 19304
rect 2041 19295 2099 19301
rect 2041 19292 2053 19295
rect 1636 19264 2053 19292
rect 1636 19252 1642 19264
rect 2041 19261 2053 19264
rect 2087 19261 2099 19295
rect 2041 19255 2099 19261
rect 3329 19295 3387 19301
rect 3329 19261 3341 19295
rect 3375 19292 3387 19295
rect 3988 19292 4016 19400
rect 4890 19388 4896 19400
rect 4948 19388 4954 19440
rect 4709 19363 4767 19369
rect 4709 19329 4721 19363
rect 4755 19360 4767 19363
rect 5000 19360 5028 19468
rect 7466 19456 7472 19508
rect 7524 19496 7530 19508
rect 7653 19499 7711 19505
rect 7653 19496 7665 19499
rect 7524 19468 7665 19496
rect 7524 19456 7530 19468
rect 7653 19465 7665 19468
rect 7699 19465 7711 19499
rect 7653 19459 7711 19465
rect 9858 19456 9864 19508
rect 9916 19496 9922 19508
rect 12621 19499 12679 19505
rect 12621 19496 12633 19499
rect 9916 19468 12633 19496
rect 9916 19456 9922 19468
rect 12621 19465 12633 19468
rect 12667 19465 12679 19499
rect 12621 19459 12679 19465
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 15252 19468 18828 19496
rect 15252 19456 15258 19468
rect 14185 19431 14243 19437
rect 6656 19400 9536 19428
rect 5074 19360 5080 19372
rect 4755 19332 5080 19360
rect 4755 19329 4767 19332
rect 4709 19323 4767 19329
rect 5074 19320 5080 19332
rect 5132 19360 5138 19372
rect 5442 19360 5448 19372
rect 5132 19332 5448 19360
rect 5132 19320 5138 19332
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 6546 19360 6552 19372
rect 6380 19332 6552 19360
rect 3375 19264 4016 19292
rect 3375 19261 3387 19264
rect 3329 19255 3387 19261
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 6380 19301 6408 19332
rect 6546 19320 6552 19332
rect 6604 19320 6610 19372
rect 6656 19369 6684 19400
rect 9508 19372 9536 19400
rect 14185 19397 14197 19431
rect 14231 19397 14243 19431
rect 14185 19391 14243 19397
rect 6641 19363 6699 19369
rect 6641 19329 6653 19363
rect 6687 19329 6699 19363
rect 8202 19360 8208 19372
rect 8163 19332 8208 19360
rect 6641 19323 6699 19329
rect 8202 19320 8208 19332
rect 8260 19320 8266 19372
rect 9490 19360 9496 19372
rect 9451 19332 9496 19360
rect 9490 19320 9496 19332
rect 9548 19320 9554 19372
rect 10965 19363 11023 19369
rect 9600 19332 9904 19360
rect 6365 19295 6423 19301
rect 4212 19264 5764 19292
rect 4212 19252 4218 19264
rect 1486 19184 1492 19236
rect 1544 19224 1550 19236
rect 1544 19196 3556 19224
rect 1544 19184 1550 19196
rect 1670 19156 1676 19168
rect 1631 19128 1676 19156
rect 1670 19116 1676 19128
rect 1728 19116 1734 19168
rect 2130 19156 2136 19168
rect 2091 19128 2136 19156
rect 2130 19116 2136 19128
rect 2188 19116 2194 19168
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2590 19156 2596 19168
rect 2547 19128 2596 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 2866 19156 2872 19168
rect 2827 19128 2872 19156
rect 2866 19116 2872 19128
rect 2924 19116 2930 19168
rect 2961 19159 3019 19165
rect 2961 19125 2973 19159
rect 3007 19156 3019 19159
rect 3050 19156 3056 19168
rect 3007 19128 3056 19156
rect 3007 19125 3019 19128
rect 2961 19119 3019 19125
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3528 19165 3556 19196
rect 3602 19184 3608 19236
rect 3660 19224 3666 19236
rect 4525 19227 4583 19233
rect 4525 19224 4537 19227
rect 3660 19196 4537 19224
rect 3660 19184 3666 19196
rect 4525 19193 4537 19196
rect 4571 19193 4583 19227
rect 4525 19187 4583 19193
rect 4798 19184 4804 19236
rect 4856 19224 4862 19236
rect 5353 19227 5411 19233
rect 5353 19224 5365 19227
rect 4856 19196 5365 19224
rect 4856 19184 4862 19196
rect 5353 19193 5365 19196
rect 5399 19193 5411 19227
rect 5736 19224 5764 19264
rect 6365 19261 6377 19295
rect 6411 19261 6423 19295
rect 6365 19255 6423 19261
rect 6454 19252 6460 19304
rect 6512 19292 6518 19304
rect 6917 19295 6975 19301
rect 6917 19292 6929 19295
rect 6512 19264 6929 19292
rect 6512 19252 6518 19264
rect 6917 19261 6929 19264
rect 6963 19261 6975 19295
rect 6917 19255 6975 19261
rect 7285 19295 7343 19301
rect 7285 19261 7297 19295
rect 7331 19261 7343 19295
rect 7285 19255 7343 19261
rect 7300 19224 7328 19255
rect 7558 19252 7564 19304
rect 7616 19292 7622 19304
rect 8481 19295 8539 19301
rect 8481 19292 8493 19295
rect 7616 19264 8493 19292
rect 7616 19252 7622 19264
rect 8481 19261 8493 19264
rect 8527 19261 8539 19295
rect 8481 19255 8539 19261
rect 9217 19295 9275 19301
rect 9217 19261 9229 19295
rect 9263 19292 9275 19295
rect 9600 19292 9628 19332
rect 9263 19264 9628 19292
rect 9263 19261 9275 19264
rect 9217 19255 9275 19261
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 9775 19295 9833 19301
rect 9775 19292 9787 19295
rect 9732 19264 9787 19292
rect 9732 19252 9738 19264
rect 9775 19261 9787 19264
rect 9821 19261 9833 19295
rect 9876 19292 9904 19332
rect 10965 19329 10977 19363
rect 11011 19360 11023 19363
rect 11238 19360 11244 19372
rect 11011 19332 11244 19360
rect 11011 19329 11023 19332
rect 10965 19323 11023 19329
rect 11238 19320 11244 19332
rect 11296 19320 11302 19372
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19360 11851 19363
rect 12066 19360 12072 19372
rect 11839 19332 12072 19360
rect 11839 19329 11851 19332
rect 11793 19323 11851 19329
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 12250 19320 12256 19372
rect 12308 19360 12314 19372
rect 12308 19332 12848 19360
rect 12308 19320 12314 19332
rect 11974 19292 11980 19304
rect 9876 19264 11980 19292
rect 9775 19255 9833 19261
rect 11974 19252 11980 19264
rect 12032 19252 12038 19304
rect 12161 19295 12219 19301
rect 12161 19261 12173 19295
rect 12207 19292 12219 19295
rect 12434 19292 12440 19304
rect 12207 19264 12440 19292
rect 12207 19261 12219 19264
rect 12161 19255 12219 19261
rect 12434 19252 12440 19264
rect 12492 19252 12498 19304
rect 12710 19292 12716 19304
rect 12671 19264 12716 19292
rect 12710 19252 12716 19264
rect 12768 19252 12774 19304
rect 12820 19292 12848 19332
rect 14200 19304 14228 19391
rect 14829 19363 14887 19369
rect 14829 19329 14841 19363
rect 14875 19360 14887 19363
rect 14918 19360 14924 19372
rect 14875 19332 14924 19360
rect 14875 19329 14887 19332
rect 14829 19323 14887 19329
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 16942 19320 16948 19372
rect 17000 19360 17006 19372
rect 17678 19360 17684 19372
rect 17000 19332 17684 19360
rect 17000 19320 17006 19332
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 18800 19369 18828 19468
rect 18785 19363 18843 19369
rect 18785 19329 18797 19363
rect 18831 19329 18843 19363
rect 18966 19360 18972 19372
rect 18927 19332 18972 19360
rect 18785 19323 18843 19329
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 19702 19360 19708 19372
rect 19663 19332 19708 19360
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 12820 19264 13124 19292
rect 12986 19233 12992 19236
rect 12980 19224 12992 19233
rect 5736 19196 7236 19224
rect 7300 19196 12848 19224
rect 12947 19196 12992 19224
rect 5353 19187 5411 19193
rect 3513 19159 3571 19165
rect 3513 19125 3525 19159
rect 3559 19125 3571 19159
rect 4062 19156 4068 19168
rect 4023 19128 4068 19156
rect 3513 19119 3571 19125
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4433 19159 4491 19165
rect 4433 19156 4445 19159
rect 4212 19128 4445 19156
rect 4212 19116 4218 19128
rect 4433 19125 4445 19128
rect 4479 19125 4491 19159
rect 4433 19119 4491 19125
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 4893 19159 4951 19165
rect 4893 19156 4905 19159
rect 4764 19128 4905 19156
rect 4764 19116 4770 19128
rect 4893 19125 4905 19128
rect 4939 19125 4951 19159
rect 5258 19156 5264 19168
rect 5219 19128 5264 19156
rect 4893 19119 4951 19125
rect 5258 19116 5264 19128
rect 5316 19116 5322 19168
rect 5997 19159 6055 19165
rect 5997 19125 6009 19159
rect 6043 19156 6055 19159
rect 6270 19156 6276 19168
rect 6043 19128 6276 19156
rect 6043 19125 6055 19128
rect 5997 19119 6055 19125
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 6457 19159 6515 19165
rect 6457 19125 6469 19159
rect 6503 19156 6515 19159
rect 6822 19156 6828 19168
rect 6503 19128 6828 19156
rect 6503 19125 6515 19128
rect 6457 19119 6515 19125
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7098 19156 7104 19168
rect 7059 19128 7104 19156
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 7208 19156 7236 19196
rect 7469 19159 7527 19165
rect 7469 19156 7481 19159
rect 7208 19128 7481 19156
rect 7469 19125 7481 19128
rect 7515 19125 7527 19159
rect 8018 19156 8024 19168
rect 7979 19128 8024 19156
rect 7469 19119 7527 19125
rect 8018 19116 8024 19128
rect 8076 19116 8082 19168
rect 8110 19116 8116 19168
rect 8168 19156 8174 19168
rect 8168 19128 8213 19156
rect 8168 19116 8174 19128
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 8665 19159 8723 19165
rect 8665 19156 8677 19159
rect 8352 19128 8677 19156
rect 8352 19116 8358 19128
rect 8665 19125 8677 19128
rect 8711 19125 8723 19159
rect 8846 19156 8852 19168
rect 8807 19128 8852 19156
rect 8665 19119 8723 19125
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 9309 19159 9367 19165
rect 9309 19125 9321 19159
rect 9355 19156 9367 19159
rect 9858 19156 9864 19168
rect 9355 19128 9864 19156
rect 9355 19125 9367 19128
rect 9309 19119 9367 19125
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 9950 19116 9956 19168
rect 10008 19156 10014 19168
rect 10318 19156 10324 19168
rect 10008 19128 10053 19156
rect 10279 19128 10324 19156
rect 10008 19116 10014 19128
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 10502 19116 10508 19168
rect 10560 19156 10566 19168
rect 10689 19159 10747 19165
rect 10689 19156 10701 19159
rect 10560 19128 10701 19156
rect 10560 19116 10566 19128
rect 10689 19125 10701 19128
rect 10735 19125 10747 19159
rect 10689 19119 10747 19125
rect 10781 19159 10839 19165
rect 10781 19125 10793 19159
rect 10827 19156 10839 19159
rect 11054 19156 11060 19168
rect 10827 19128 11060 19156
rect 10827 19125 10839 19128
rect 10781 19119 10839 19125
rect 11054 19116 11060 19128
rect 11112 19116 11118 19168
rect 11146 19116 11152 19168
rect 11204 19156 11210 19168
rect 11514 19156 11520 19168
rect 11204 19128 11249 19156
rect 11475 19128 11520 19156
rect 11204 19116 11210 19128
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 11609 19159 11667 19165
rect 11609 19125 11621 19159
rect 11655 19156 11667 19159
rect 12250 19156 12256 19168
rect 11655 19128 12256 19156
rect 11655 19125 11667 19128
rect 11609 19119 11667 19125
rect 12250 19116 12256 19128
rect 12308 19116 12314 19168
rect 12345 19159 12403 19165
rect 12345 19125 12357 19159
rect 12391 19156 12403 19159
rect 12526 19156 12532 19168
rect 12391 19128 12532 19156
rect 12391 19125 12403 19128
rect 12345 19119 12403 19125
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 12618 19116 12624 19168
rect 12676 19156 12682 19168
rect 12820 19156 12848 19196
rect 12980 19187 12992 19196
rect 12986 19184 12992 19187
rect 13044 19184 13050 19236
rect 13096 19224 13124 19264
rect 14182 19252 14188 19304
rect 14240 19252 14246 19304
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15102 19292 15108 19304
rect 15059 19264 15108 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15562 19252 15568 19304
rect 15620 19292 15626 19304
rect 15664 19295 15722 19301
rect 15664 19292 15676 19295
rect 15620 19264 15676 19292
rect 15620 19252 15626 19264
rect 15664 19261 15676 19264
rect 15710 19261 15722 19295
rect 16206 19292 16212 19304
rect 15664 19255 15722 19261
rect 15764 19264 16212 19292
rect 15764 19224 15792 19264
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 16666 19252 16672 19304
rect 16724 19292 16730 19304
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 16724 19264 19625 19292
rect 16724 19252 16730 19264
rect 19613 19261 19625 19264
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 19981 19295 20039 19301
rect 19981 19261 19993 19295
rect 20027 19292 20039 19295
rect 20714 19292 20720 19304
rect 20027 19264 20720 19292
rect 20027 19261 20039 19264
rect 19981 19255 20039 19261
rect 20714 19252 20720 19264
rect 20772 19252 20778 19304
rect 13096 19196 15792 19224
rect 15838 19184 15844 19236
rect 15896 19233 15902 19236
rect 15896 19227 15960 19233
rect 15896 19193 15914 19227
rect 15948 19193 15960 19227
rect 16574 19224 16580 19236
rect 15896 19187 15960 19193
rect 16040 19196 16580 19224
rect 15896 19184 15902 19187
rect 13906 19156 13912 19168
rect 12676 19128 12721 19156
rect 12820 19128 13912 19156
rect 12676 19116 12682 19128
rect 13906 19116 13912 19128
rect 13964 19116 13970 19168
rect 13998 19116 14004 19168
rect 14056 19156 14062 19168
rect 14093 19159 14151 19165
rect 14093 19156 14105 19159
rect 14056 19128 14105 19156
rect 14056 19116 14062 19128
rect 14093 19125 14105 19128
rect 14139 19125 14151 19159
rect 14093 19119 14151 19125
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 14553 19159 14611 19165
rect 14553 19156 14565 19159
rect 14516 19128 14565 19156
rect 14516 19116 14522 19128
rect 14553 19125 14565 19128
rect 14599 19125 14611 19159
rect 14553 19119 14611 19125
rect 14642 19116 14648 19168
rect 14700 19156 14706 19168
rect 15197 19159 15255 19165
rect 14700 19128 14745 19156
rect 14700 19116 14706 19128
rect 15197 19125 15209 19159
rect 15243 19156 15255 19159
rect 16040 19156 16068 19196
rect 16574 19184 16580 19196
rect 16632 19184 16638 19236
rect 19521 19227 19579 19233
rect 19521 19224 19533 19227
rect 17144 19196 19533 19224
rect 15243 19128 16068 19156
rect 15243 19125 15255 19128
rect 15197 19119 15255 19125
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 17144 19165 17172 19196
rect 19521 19193 19533 19196
rect 19567 19193 19579 19227
rect 19521 19187 19579 19193
rect 17037 19159 17095 19165
rect 17037 19156 17049 19159
rect 16172 19128 17049 19156
rect 16172 19116 16178 19128
rect 17037 19125 17049 19128
rect 17083 19125 17095 19159
rect 17037 19119 17095 19125
rect 17129 19159 17187 19165
rect 17129 19125 17141 19159
rect 17175 19125 17187 19159
rect 17129 19119 17187 19125
rect 17310 19116 17316 19168
rect 17368 19156 17374 19168
rect 17497 19159 17555 19165
rect 17497 19156 17509 19159
rect 17368 19128 17509 19156
rect 17368 19116 17374 19128
rect 17497 19125 17509 19128
rect 17543 19125 17555 19159
rect 17497 19119 17555 19125
rect 17586 19116 17592 19168
rect 17644 19156 17650 19168
rect 17644 19128 17689 19156
rect 17644 19116 17650 19128
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 18325 19159 18383 19165
rect 18325 19156 18337 19159
rect 18104 19128 18337 19156
rect 18104 19116 18110 19128
rect 18325 19125 18337 19128
rect 18371 19125 18383 19159
rect 18690 19156 18696 19168
rect 18651 19128 18696 19156
rect 18325 19119 18383 19125
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 19150 19156 19156 19168
rect 19111 19128 19156 19156
rect 19150 19116 19156 19128
rect 19208 19116 19214 19168
rect 20165 19159 20223 19165
rect 20165 19125 20177 19159
rect 20211 19156 20223 19159
rect 20993 19159 21051 19165
rect 20993 19156 21005 19159
rect 20211 19128 21005 19156
rect 20211 19125 20223 19128
rect 20165 19119 20223 19125
rect 20993 19125 21005 19128
rect 21039 19125 21051 19159
rect 20993 19119 21051 19125
rect 1104 19066 20884 19088
rect 1104 19014 7579 19066
rect 7631 19014 7643 19066
rect 7695 19014 7707 19066
rect 7759 19014 7771 19066
rect 7823 19014 14176 19066
rect 14228 19014 14240 19066
rect 14292 19014 14304 19066
rect 14356 19014 14368 19066
rect 14420 19014 20884 19066
rect 1104 18992 20884 19014
rect 842 18912 848 18964
rect 900 18952 906 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 900 18924 1593 18952
rect 900 18912 906 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 1581 18915 1639 18921
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 3142 18952 3148 18964
rect 1728 18924 3148 18952
rect 1728 18912 1734 18924
rect 3142 18912 3148 18924
rect 3200 18912 3206 18964
rect 3513 18955 3571 18961
rect 3513 18921 3525 18955
rect 3559 18952 3571 18955
rect 3602 18952 3608 18964
rect 3559 18924 3608 18952
rect 3559 18921 3571 18924
rect 3513 18915 3571 18921
rect 3602 18912 3608 18924
rect 3660 18912 3666 18964
rect 3789 18955 3847 18961
rect 3789 18921 3801 18955
rect 3835 18952 3847 18955
rect 4614 18952 4620 18964
rect 3835 18924 4620 18952
rect 3835 18921 3847 18924
rect 3789 18915 3847 18921
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 4890 18912 4896 18964
rect 4948 18952 4954 18964
rect 7101 18955 7159 18961
rect 7101 18952 7113 18955
rect 4948 18924 7113 18952
rect 4948 18912 4954 18924
rect 7101 18921 7113 18924
rect 7147 18921 7159 18955
rect 7101 18915 7159 18921
rect 8018 18912 8024 18964
rect 8076 18952 8082 18964
rect 9122 18952 9128 18964
rect 8076 18924 9128 18952
rect 8076 18912 8082 18924
rect 9122 18912 9128 18924
rect 9180 18912 9186 18964
rect 9217 18955 9275 18961
rect 9217 18921 9229 18955
rect 9263 18952 9275 18955
rect 9677 18955 9735 18961
rect 9677 18952 9689 18955
rect 9263 18924 9689 18952
rect 9263 18921 9275 18924
rect 9217 18915 9275 18921
rect 9677 18921 9689 18924
rect 9723 18921 9735 18955
rect 9677 18915 9735 18921
rect 10318 18912 10324 18964
rect 10376 18912 10382 18964
rect 10505 18955 10563 18961
rect 10505 18921 10517 18955
rect 10551 18952 10563 18955
rect 10870 18952 10876 18964
rect 10551 18924 10876 18952
rect 10551 18921 10563 18924
rect 10505 18915 10563 18921
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 11606 18952 11612 18964
rect 11112 18924 11612 18952
rect 11112 18912 11118 18924
rect 11606 18912 11612 18924
rect 11664 18912 11670 18964
rect 12986 18912 12992 18964
rect 13044 18952 13050 18964
rect 13814 18952 13820 18964
rect 13044 18924 13820 18952
rect 13044 18912 13050 18924
rect 13814 18912 13820 18924
rect 13872 18952 13878 18964
rect 14001 18955 14059 18961
rect 14001 18952 14013 18955
rect 13872 18924 14013 18952
rect 13872 18912 13878 18924
rect 14001 18921 14013 18924
rect 14047 18921 14059 18955
rect 14001 18915 14059 18921
rect 14093 18955 14151 18961
rect 14093 18921 14105 18955
rect 14139 18952 14151 18955
rect 14642 18952 14648 18964
rect 14139 18924 14648 18952
rect 14139 18921 14151 18924
rect 14093 18915 14151 18921
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 15838 18912 15844 18964
rect 15896 18952 15902 18964
rect 15896 18924 16528 18952
rect 15896 18912 15902 18924
rect 10336 18884 10364 18912
rect 16500 18896 16528 18924
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 16942 18952 16948 18964
rect 16632 18924 16948 18952
rect 16632 18912 16638 18924
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 17126 18952 17132 18964
rect 17039 18924 17132 18952
rect 17126 18912 17132 18924
rect 17184 18952 17190 18964
rect 17586 18952 17592 18964
rect 17184 18924 17592 18952
rect 17184 18912 17190 18924
rect 17586 18912 17592 18924
rect 17644 18912 17650 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 17696 18924 19809 18952
rect 1412 18856 10364 18884
rect 10956 18887 11014 18893
rect 1412 18825 1440 18856
rect 10956 18853 10968 18887
rect 11002 18884 11014 18887
rect 11422 18884 11428 18896
rect 11002 18856 11428 18884
rect 11002 18853 11014 18856
rect 10956 18847 11014 18853
rect 11422 18844 11428 18856
rect 11480 18844 11486 18896
rect 11514 18844 11520 18896
rect 11572 18884 11578 18896
rect 14921 18887 14979 18893
rect 14921 18884 14933 18887
rect 11572 18856 12388 18884
rect 11572 18844 11578 18856
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18785 1455 18819
rect 1397 18779 1455 18785
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18785 1823 18819
rect 1765 18779 1823 18785
rect 2133 18819 2191 18825
rect 2133 18785 2145 18819
rect 2179 18816 2191 18819
rect 2222 18816 2228 18828
rect 2179 18788 2228 18816
rect 2179 18785 2191 18788
rect 2133 18779 2191 18785
rect 1780 18680 1808 18779
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 2406 18825 2412 18828
rect 2400 18816 2412 18825
rect 2367 18788 2412 18816
rect 2400 18779 2412 18788
rect 2406 18776 2412 18779
rect 2464 18776 2470 18828
rect 3602 18816 3608 18828
rect 3563 18788 3608 18816
rect 3602 18776 3608 18788
rect 3660 18776 3666 18828
rect 4329 18776 4335 18828
rect 4387 18816 4393 18828
rect 5804 18819 5862 18825
rect 5804 18816 5816 18819
rect 4387 18788 4432 18816
rect 5460 18788 5816 18816
rect 4387 18776 4393 18788
rect 4065 18751 4123 18757
rect 4065 18717 4077 18751
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 1780 18652 2176 18680
rect 290 18572 296 18624
rect 348 18612 354 18624
rect 1949 18615 2007 18621
rect 1949 18612 1961 18615
rect 348 18584 1961 18612
rect 348 18572 354 18584
rect 1949 18581 1961 18584
rect 1995 18581 2007 18615
rect 2148 18612 2176 18652
rect 3878 18612 3884 18624
rect 2148 18584 3884 18612
rect 1949 18575 2007 18581
rect 3878 18572 3884 18584
rect 3936 18572 3942 18624
rect 4080 18612 4108 18711
rect 5460 18689 5488 18788
rect 5804 18785 5816 18788
rect 5850 18816 5862 18819
rect 6270 18816 6276 18828
rect 5850 18788 6276 18816
rect 5850 18785 5862 18788
rect 5804 18779 5862 18785
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 7460 18819 7518 18825
rect 7460 18785 7472 18819
rect 7506 18816 7518 18819
rect 8018 18816 8024 18828
rect 7506 18788 8024 18816
rect 7506 18785 7518 18788
rect 7460 18779 7518 18785
rect 8018 18776 8024 18788
rect 8076 18776 8082 18828
rect 9125 18819 9183 18825
rect 9125 18785 9137 18819
rect 9171 18816 9183 18819
rect 9950 18816 9956 18828
rect 9171 18788 9956 18816
rect 9171 18785 9183 18788
rect 9125 18779 9183 18785
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18816 10103 18819
rect 10318 18816 10324 18828
rect 10091 18788 10324 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 10689 18819 10747 18825
rect 10689 18785 10701 18819
rect 10735 18816 10747 18819
rect 10778 18816 10784 18828
rect 10735 18788 10784 18816
rect 10735 18785 10747 18788
rect 10689 18779 10747 18785
rect 10778 18776 10784 18788
rect 10836 18776 10842 18828
rect 11330 18776 11336 18828
rect 11388 18816 11394 18828
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11388 18788 12173 18816
rect 11388 18776 11394 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12360 18816 12388 18856
rect 12452 18856 14933 18884
rect 12452 18816 12480 18856
rect 14921 18853 14933 18856
rect 14967 18853 14979 18887
rect 14921 18847 14979 18853
rect 16016 18887 16074 18893
rect 16016 18853 16028 18887
rect 16062 18884 16074 18887
rect 16114 18884 16120 18896
rect 16062 18856 16120 18884
rect 16062 18853 16074 18856
rect 16016 18847 16074 18853
rect 16114 18844 16120 18856
rect 16172 18844 16178 18896
rect 16482 18844 16488 18896
rect 16540 18884 16546 18896
rect 17696 18884 17724 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 20073 18955 20131 18961
rect 20073 18921 20085 18955
rect 20119 18952 20131 18955
rect 20990 18952 20996 18964
rect 20119 18924 20996 18952
rect 20119 18921 20131 18924
rect 20073 18915 20131 18921
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 16540 18856 17724 18884
rect 17957 18887 18015 18893
rect 16540 18844 16546 18856
rect 17957 18853 17969 18887
rect 18003 18884 18015 18887
rect 18003 18856 18644 18884
rect 18003 18853 18015 18856
rect 17957 18847 18015 18853
rect 12360 18788 12480 18816
rect 12161 18779 12219 18785
rect 12526 18776 12532 18828
rect 12584 18816 12590 18828
rect 12621 18819 12679 18825
rect 12621 18816 12633 18819
rect 12584 18788 12633 18816
rect 12584 18776 12590 18788
rect 12621 18785 12633 18788
rect 12667 18816 12679 18819
rect 12710 18816 12716 18828
rect 12667 18788 12716 18816
rect 12667 18785 12679 18788
rect 12621 18779 12679 18785
rect 12710 18776 12716 18788
rect 12768 18776 12774 18828
rect 12888 18819 12946 18825
rect 12888 18785 12900 18819
rect 12934 18816 12946 18819
rect 14274 18816 14280 18828
rect 12934 18788 14280 18816
rect 12934 18785 12946 18788
rect 12888 18779 12946 18785
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 14366 18776 14372 18828
rect 14424 18816 14430 18828
rect 14461 18819 14519 18825
rect 14461 18816 14473 18819
rect 14424 18788 14473 18816
rect 14424 18776 14430 18788
rect 14461 18785 14473 18788
rect 14507 18785 14519 18819
rect 14461 18779 14519 18785
rect 14734 18776 14740 18828
rect 14792 18816 14798 18828
rect 15289 18819 15347 18825
rect 15289 18816 15301 18819
rect 14792 18788 15301 18816
rect 14792 18776 14798 18788
rect 15289 18785 15301 18788
rect 15335 18785 15347 18819
rect 15473 18819 15531 18825
rect 15473 18816 15485 18819
rect 15289 18779 15347 18785
rect 15396 18788 15485 18816
rect 5537 18751 5595 18757
rect 5537 18717 5549 18751
rect 5583 18717 5595 18751
rect 5537 18711 5595 18717
rect 5445 18683 5503 18689
rect 5445 18649 5457 18683
rect 5491 18649 5503 18683
rect 5445 18643 5503 18649
rect 5258 18612 5264 18624
rect 4080 18584 5264 18612
rect 5258 18572 5264 18584
rect 5316 18612 5322 18624
rect 5552 18612 5580 18711
rect 7098 18708 7104 18760
rect 7156 18748 7162 18760
rect 7193 18751 7251 18757
rect 7193 18748 7205 18751
rect 7156 18720 7205 18748
rect 7156 18708 7162 18720
rect 7193 18717 7205 18720
rect 7239 18717 7251 18751
rect 9306 18748 9312 18760
rect 9267 18720 9312 18748
rect 7193 18711 7251 18717
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 10134 18748 10140 18760
rect 10095 18720 10140 18748
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10226 18708 10232 18760
rect 10284 18748 10290 18760
rect 10284 18720 10329 18748
rect 10284 18708 10290 18720
rect 13630 18708 13636 18760
rect 13688 18748 13694 18760
rect 14553 18751 14611 18757
rect 14553 18748 14565 18751
rect 13688 18720 14565 18748
rect 13688 18708 13694 18720
rect 14553 18717 14565 18720
rect 14599 18717 14611 18751
rect 14553 18711 14611 18717
rect 14645 18751 14703 18757
rect 14645 18717 14657 18751
rect 14691 18748 14703 18751
rect 14918 18748 14924 18760
rect 14691 18720 14924 18748
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 14918 18708 14924 18720
rect 14976 18708 14982 18760
rect 8757 18683 8815 18689
rect 8757 18680 8769 18683
rect 8128 18652 8769 18680
rect 5316 18584 5580 18612
rect 5316 18572 5322 18584
rect 6454 18572 6460 18624
rect 6512 18612 6518 18624
rect 6917 18615 6975 18621
rect 6917 18612 6929 18615
rect 6512 18584 6929 18612
rect 6512 18572 6518 18584
rect 6917 18581 6929 18584
rect 6963 18581 6975 18615
rect 6917 18575 6975 18581
rect 7101 18615 7159 18621
rect 7101 18581 7113 18615
rect 7147 18612 7159 18615
rect 8128 18612 8156 18652
rect 8757 18649 8769 18652
rect 8803 18680 8815 18683
rect 10410 18680 10416 18692
rect 8803 18652 10416 18680
rect 8803 18649 8815 18652
rect 8757 18643 8815 18649
rect 10410 18640 10416 18652
rect 10468 18640 10474 18692
rect 13814 18640 13820 18692
rect 13872 18680 13878 18692
rect 15396 18680 15424 18788
rect 15473 18785 15485 18788
rect 15519 18785 15531 18819
rect 16758 18816 16764 18828
rect 15473 18779 15531 18785
rect 15571 18788 16764 18816
rect 15571 18680 15599 18788
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 16942 18776 16948 18828
rect 17000 18816 17006 18828
rect 17221 18819 17279 18825
rect 17221 18816 17233 18819
rect 17000 18788 17233 18816
rect 17000 18776 17006 18788
rect 17221 18785 17233 18788
rect 17267 18785 17279 18819
rect 17221 18779 17279 18785
rect 17678 18776 17684 18828
rect 17736 18816 17742 18828
rect 18049 18819 18107 18825
rect 17736 18788 17816 18816
rect 17736 18776 17742 18788
rect 15654 18708 15660 18760
rect 15712 18748 15718 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 15712 18720 15761 18748
rect 15712 18708 15718 18720
rect 15749 18717 15761 18720
rect 15795 18717 15807 18751
rect 15749 18711 15807 18717
rect 16850 18708 16856 18760
rect 16908 18748 16914 18760
rect 17788 18748 17816 18788
rect 18049 18785 18061 18819
rect 18095 18816 18107 18819
rect 18322 18816 18328 18828
rect 18095 18788 18328 18816
rect 18095 18785 18107 18788
rect 18049 18779 18107 18785
rect 18322 18776 18328 18788
rect 18380 18776 18386 18828
rect 18616 18816 18644 18856
rect 18684 18819 18742 18825
rect 18684 18816 18696 18819
rect 18616 18788 18696 18816
rect 18684 18785 18696 18788
rect 18730 18816 18742 18819
rect 19426 18816 19432 18828
rect 18730 18788 19432 18816
rect 18730 18785 18742 18788
rect 18684 18779 18742 18785
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 19889 18819 19947 18825
rect 19889 18816 19901 18819
rect 19760 18788 19901 18816
rect 19760 18776 19766 18788
rect 19889 18785 19901 18788
rect 19935 18785 19947 18819
rect 19889 18779 19947 18785
rect 20257 18819 20315 18825
rect 20257 18785 20269 18819
rect 20303 18816 20315 18819
rect 20806 18816 20812 18828
rect 20303 18788 20812 18816
rect 20303 18785 20315 18788
rect 20257 18779 20315 18785
rect 20806 18776 20812 18788
rect 20864 18776 20870 18828
rect 18141 18751 18199 18757
rect 18141 18748 18153 18751
rect 16908 18720 17724 18748
rect 17788 18720 18153 18748
rect 16908 18708 16914 18720
rect 17589 18683 17647 18689
rect 17589 18680 17601 18683
rect 13872 18652 15424 18680
rect 15488 18652 15599 18680
rect 16684 18652 17601 18680
rect 13872 18640 13878 18652
rect 7147 18584 8156 18612
rect 7147 18581 7159 18584
rect 7101 18575 7159 18581
rect 8202 18572 8208 18624
rect 8260 18612 8266 18624
rect 8573 18615 8631 18621
rect 8573 18612 8585 18615
rect 8260 18584 8585 18612
rect 8260 18572 8266 18584
rect 8573 18581 8585 18584
rect 8619 18581 8631 18615
rect 8573 18575 8631 18581
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 10505 18615 10563 18621
rect 10505 18612 10517 18615
rect 9088 18584 10517 18612
rect 9088 18572 9094 18584
rect 10505 18581 10517 18584
rect 10551 18581 10563 18615
rect 12066 18612 12072 18624
rect 12027 18584 12072 18612
rect 10505 18575 10563 18581
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12158 18572 12164 18624
rect 12216 18612 12222 18624
rect 12345 18615 12403 18621
rect 12345 18612 12357 18615
rect 12216 18584 12357 18612
rect 12216 18572 12222 18584
rect 12345 18581 12357 18584
rect 12391 18581 12403 18615
rect 12345 18575 12403 18581
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 15488 18612 15516 18652
rect 15654 18612 15660 18624
rect 13320 18584 15516 18612
rect 15615 18584 15660 18612
rect 13320 18572 13326 18584
rect 15654 18572 15660 18584
rect 15712 18572 15718 18624
rect 15746 18572 15752 18624
rect 15804 18612 15810 18624
rect 16684 18612 16712 18652
rect 17589 18649 17601 18652
rect 17635 18649 17647 18683
rect 17696 18680 17724 18720
rect 18141 18717 18153 18720
rect 18187 18717 18199 18751
rect 18141 18711 18199 18717
rect 18230 18708 18236 18760
rect 18288 18748 18294 18760
rect 18417 18751 18475 18757
rect 18417 18748 18429 18751
rect 18288 18720 18429 18748
rect 18288 18708 18294 18720
rect 18417 18717 18429 18720
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 20441 18683 20499 18689
rect 17696 18652 18000 18680
rect 17589 18643 17647 18649
rect 15804 18584 16712 18612
rect 17405 18615 17463 18621
rect 15804 18572 15810 18584
rect 17405 18581 17417 18615
rect 17451 18612 17463 18615
rect 17862 18612 17868 18624
rect 17451 18584 17868 18612
rect 17451 18581 17463 18584
rect 17405 18575 17463 18581
rect 17862 18572 17868 18584
rect 17920 18572 17926 18624
rect 17972 18612 18000 18652
rect 20441 18649 20453 18683
rect 20487 18680 20499 18683
rect 21634 18680 21640 18692
rect 20487 18652 21640 18680
rect 20487 18649 20499 18652
rect 20441 18643 20499 18649
rect 21634 18640 21640 18652
rect 21692 18640 21698 18692
rect 19150 18612 19156 18624
rect 17972 18584 19156 18612
rect 19150 18572 19156 18584
rect 19208 18572 19214 18624
rect 1104 18522 20884 18544
rect 1104 18470 4280 18522
rect 4332 18470 4344 18522
rect 4396 18470 4408 18522
rect 4460 18470 4472 18522
rect 4524 18470 10878 18522
rect 10930 18470 10942 18522
rect 10994 18470 11006 18522
rect 11058 18470 11070 18522
rect 11122 18470 17475 18522
rect 17527 18470 17539 18522
rect 17591 18470 17603 18522
rect 17655 18470 17667 18522
rect 17719 18470 20884 18522
rect 1104 18448 20884 18470
rect 2406 18368 2412 18420
rect 2464 18408 2470 18420
rect 2777 18411 2835 18417
rect 2777 18408 2789 18411
rect 2464 18380 2789 18408
rect 2464 18368 2470 18380
rect 2777 18377 2789 18380
rect 2823 18377 2835 18411
rect 2777 18371 2835 18377
rect 3878 18368 3884 18420
rect 3936 18368 3942 18420
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 4341 18411 4399 18417
rect 4341 18408 4353 18411
rect 4212 18380 4353 18408
rect 4212 18368 4218 18380
rect 4341 18377 4353 18380
rect 4387 18377 4399 18411
rect 9030 18408 9036 18420
rect 4341 18371 4399 18377
rect 5276 18380 9036 18408
rect 3896 18340 3924 18368
rect 5276 18340 5304 18380
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 9217 18411 9275 18417
rect 9217 18377 9229 18411
rect 9263 18408 9275 18411
rect 10226 18408 10232 18420
rect 9263 18380 10232 18408
rect 9263 18377 9275 18380
rect 9217 18371 9275 18377
rect 3896 18312 5304 18340
rect 6641 18343 6699 18349
rect 6641 18309 6653 18343
rect 6687 18309 6699 18343
rect 6641 18303 6699 18309
rect 6825 18343 6883 18349
rect 6825 18309 6837 18343
rect 6871 18340 6883 18343
rect 7282 18340 7288 18352
rect 6871 18312 7288 18340
rect 6871 18309 6883 18312
rect 6825 18303 6883 18309
rect 5074 18272 5080 18284
rect 5035 18244 5080 18272
rect 5074 18232 5080 18244
rect 5132 18232 5138 18284
rect 5258 18272 5264 18284
rect 5219 18244 5264 18272
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 6362 18232 6368 18284
rect 6420 18272 6426 18284
rect 6656 18272 6684 18303
rect 7282 18300 7288 18312
rect 7340 18300 7346 18352
rect 6914 18272 6920 18284
rect 6420 18244 6592 18272
rect 6656 18244 6920 18272
rect 6420 18232 6426 18244
rect 1394 18204 1400 18216
rect 1307 18176 1400 18204
rect 1394 18164 1400 18176
rect 1452 18204 1458 18216
rect 2222 18204 2228 18216
rect 1452 18176 2228 18204
rect 1452 18164 1458 18176
rect 2222 18164 2228 18176
rect 2280 18204 2286 18216
rect 2961 18207 3019 18213
rect 2961 18204 2973 18207
rect 2280 18176 2973 18204
rect 2280 18164 2286 18176
rect 2961 18173 2973 18176
rect 3007 18173 3019 18207
rect 2961 18167 3019 18173
rect 3228 18207 3286 18213
rect 3228 18173 3240 18207
rect 3274 18204 3286 18207
rect 3510 18204 3516 18216
rect 3274 18176 3516 18204
rect 3274 18173 3286 18176
rect 3228 18167 3286 18173
rect 1664 18139 1722 18145
rect 1664 18105 1676 18139
rect 1710 18136 1722 18139
rect 2774 18136 2780 18148
rect 1710 18108 2780 18136
rect 1710 18105 1722 18108
rect 1664 18099 1722 18105
rect 2774 18096 2780 18108
rect 2832 18096 2838 18148
rect 2976 18136 3004 18167
rect 3510 18164 3516 18176
rect 3568 18164 3574 18216
rect 3602 18164 3608 18216
rect 3660 18204 3666 18216
rect 4893 18207 4951 18213
rect 4893 18204 4905 18207
rect 3660 18176 4905 18204
rect 3660 18164 3666 18176
rect 4893 18173 4905 18176
rect 4939 18173 4951 18207
rect 4893 18167 4951 18173
rect 5276 18136 5304 18232
rect 5528 18207 5586 18213
rect 5528 18173 5540 18207
rect 5574 18204 5586 18207
rect 6454 18204 6460 18216
rect 5574 18176 6460 18204
rect 5574 18173 5586 18176
rect 5528 18167 5586 18173
rect 6454 18164 6460 18176
rect 6512 18164 6518 18216
rect 6564 18204 6592 18244
rect 6914 18232 6920 18244
rect 6972 18272 6978 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 6972 18244 7389 18272
rect 6972 18232 6978 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 9324 18272 9352 18380
rect 10226 18368 10232 18380
rect 10284 18368 10290 18420
rect 11422 18368 11428 18420
rect 11480 18408 11486 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 11480 18380 12173 18408
rect 11480 18368 11486 18380
rect 12161 18377 12173 18380
rect 12207 18408 12219 18411
rect 12342 18408 12348 18420
rect 12207 18380 12348 18408
rect 12207 18377 12219 18380
rect 12161 18371 12219 18377
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 12452 18380 13400 18408
rect 9324 18244 9444 18272
rect 7377 18235 7435 18241
rect 7837 18207 7895 18213
rect 6564 18176 7788 18204
rect 2976 18108 5304 18136
rect 5718 18096 5724 18148
rect 5776 18136 5782 18148
rect 7285 18139 7343 18145
rect 7285 18136 7297 18139
rect 5776 18108 7297 18136
rect 5776 18096 5782 18108
rect 7285 18105 7297 18108
rect 7331 18105 7343 18139
rect 7285 18099 7343 18105
rect 4154 18028 4160 18080
rect 4212 18068 4218 18080
rect 4433 18071 4491 18077
rect 4433 18068 4445 18071
rect 4212 18040 4445 18068
rect 4212 18028 4218 18040
rect 4433 18037 4445 18040
rect 4479 18037 4491 18071
rect 4798 18068 4804 18080
rect 4759 18040 4804 18068
rect 4433 18031 4491 18037
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 4982 18028 4988 18080
rect 5040 18068 5046 18080
rect 7193 18071 7251 18077
rect 7193 18068 7205 18071
rect 5040 18040 7205 18068
rect 5040 18028 5046 18040
rect 7193 18037 7205 18040
rect 7239 18037 7251 18071
rect 7760 18068 7788 18176
rect 7837 18173 7849 18207
rect 7883 18204 7895 18207
rect 8478 18204 8484 18216
rect 7883 18176 8484 18204
rect 7883 18173 7895 18176
rect 7837 18167 7895 18173
rect 8478 18164 8484 18176
rect 8536 18204 8542 18216
rect 9030 18204 9036 18216
rect 8536 18176 9036 18204
rect 8536 18164 8542 18176
rect 9030 18164 9036 18176
rect 9088 18204 9094 18216
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 9088 18176 9321 18204
rect 9088 18164 9094 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9416 18204 9444 18244
rect 10410 18232 10416 18284
rect 10468 18272 10474 18284
rect 12452 18272 12480 18380
rect 13372 18340 13400 18380
rect 14274 18368 14280 18420
rect 14332 18408 14338 18420
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 14332 18380 14933 18408
rect 14332 18368 14338 18380
rect 14921 18377 14933 18380
rect 14967 18377 14979 18411
rect 19521 18411 19579 18417
rect 19521 18408 19533 18411
rect 14921 18371 14979 18377
rect 15580 18380 19533 18408
rect 15286 18340 15292 18352
rect 13372 18312 15292 18340
rect 15286 18300 15292 18312
rect 15344 18300 15350 18352
rect 14090 18272 14096 18284
rect 10468 18244 10916 18272
rect 10468 18232 10474 18244
rect 9565 18207 9623 18213
rect 9565 18204 9577 18207
rect 9416 18176 9577 18204
rect 9309 18167 9367 18173
rect 9565 18173 9577 18176
rect 9611 18173 9623 18207
rect 10778 18204 10784 18216
rect 10739 18176 10784 18204
rect 9565 18167 9623 18173
rect 10778 18164 10784 18176
rect 10836 18164 10842 18216
rect 10888 18204 10916 18244
rect 11808 18244 12480 18272
rect 13740 18244 14096 18272
rect 11808 18204 11836 18244
rect 10888 18176 11836 18204
rect 12437 18207 12495 18213
rect 12437 18173 12449 18207
rect 12483 18204 12495 18207
rect 12526 18204 12532 18216
rect 12483 18176 12532 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 12526 18164 12532 18176
rect 12584 18164 12590 18216
rect 12704 18207 12762 18213
rect 12704 18173 12716 18207
rect 12750 18204 12762 18207
rect 13740 18204 13768 18244
rect 14090 18232 14096 18244
rect 14148 18272 14154 18284
rect 15580 18281 15608 18380
rect 19521 18377 19533 18380
rect 19567 18377 19579 18411
rect 19521 18371 19579 18377
rect 15838 18300 15844 18352
rect 15896 18340 15902 18352
rect 17310 18340 17316 18352
rect 15896 18312 15976 18340
rect 17271 18312 17316 18340
rect 15896 18300 15902 18312
rect 15948 18281 15976 18312
rect 17310 18300 17316 18312
rect 17368 18300 17374 18352
rect 17770 18340 17776 18352
rect 17731 18312 17776 18340
rect 17770 18300 17776 18312
rect 17828 18300 17834 18352
rect 19426 18340 19432 18352
rect 19387 18312 19432 18340
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 20990 18340 20996 18352
rect 20951 18312 20996 18340
rect 20990 18300 20996 18312
rect 21048 18300 21054 18352
rect 14461 18275 14519 18281
rect 14461 18272 14473 18275
rect 14148 18244 14473 18272
rect 14148 18232 14154 18244
rect 14461 18241 14473 18244
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 15933 18275 15991 18281
rect 15703 18244 15884 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 12750 18176 13768 18204
rect 12750 18173 12762 18176
rect 12704 18167 12762 18173
rect 13998 18164 14004 18216
rect 14056 18204 14062 18216
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 14056 18176 14381 18204
rect 14056 18164 14062 18176
rect 14369 18173 14381 18176
rect 14415 18173 14427 18207
rect 14734 18204 14740 18216
rect 14695 18176 14740 18204
rect 14369 18167 14427 18173
rect 14734 18164 14740 18176
rect 14792 18204 14798 18216
rect 15194 18204 15200 18216
rect 14792 18176 15200 18204
rect 14792 18164 14798 18176
rect 15194 18164 15200 18176
rect 15252 18164 15258 18216
rect 15473 18207 15531 18213
rect 15473 18173 15485 18207
rect 15519 18204 15531 18207
rect 15746 18204 15752 18216
rect 15519 18176 15752 18204
rect 15519 18173 15531 18176
rect 15473 18167 15531 18173
rect 15746 18164 15752 18176
rect 15804 18164 15810 18216
rect 15856 18204 15884 18244
rect 15933 18241 15945 18275
rect 15979 18241 15991 18275
rect 20073 18275 20131 18281
rect 20073 18272 20085 18275
rect 15933 18235 15991 18241
rect 19076 18244 20085 18272
rect 16022 18204 16028 18216
rect 15856 18176 16028 18204
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 16200 18207 16258 18213
rect 16200 18173 16212 18207
rect 16246 18204 16258 18207
rect 17126 18204 17132 18216
rect 16246 18176 17132 18204
rect 16246 18173 16258 18176
rect 16200 18167 16258 18173
rect 17126 18164 17132 18176
rect 17184 18164 17190 18216
rect 17589 18207 17647 18213
rect 17589 18173 17601 18207
rect 17635 18204 17647 18207
rect 17862 18204 17868 18216
rect 17635 18176 17868 18204
rect 17635 18173 17647 18176
rect 17589 18167 17647 18173
rect 17862 18164 17868 18176
rect 17920 18164 17926 18216
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 18138 18204 18144 18216
rect 18095 18176 18144 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 8104 18139 8162 18145
rect 8104 18105 8116 18139
rect 8150 18136 8162 18139
rect 8202 18136 8208 18148
rect 8150 18108 8208 18136
rect 8150 18105 8162 18108
rect 8104 18099 8162 18105
rect 8202 18096 8208 18108
rect 8260 18096 8266 18148
rect 8846 18096 8852 18148
rect 8904 18136 8910 18148
rect 10870 18136 10876 18148
rect 8904 18108 10876 18136
rect 8904 18096 8910 18108
rect 10870 18096 10876 18108
rect 10928 18096 10934 18148
rect 11048 18139 11106 18145
rect 11048 18105 11060 18139
rect 11094 18136 11106 18139
rect 11238 18136 11244 18148
rect 11094 18108 11244 18136
rect 11094 18105 11106 18108
rect 11048 18099 11106 18105
rect 11238 18096 11244 18108
rect 11296 18096 11302 18148
rect 14274 18136 14280 18148
rect 14235 18108 14280 18136
rect 14274 18096 14280 18108
rect 14332 18096 14338 18148
rect 18322 18145 18328 18148
rect 18316 18136 18328 18145
rect 18283 18108 18328 18136
rect 18316 18099 18328 18108
rect 18322 18096 18328 18099
rect 18380 18096 18386 18148
rect 9214 18068 9220 18080
rect 7760 18040 9220 18068
rect 7193 18031 7251 18037
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 9306 18028 9312 18080
rect 9364 18068 9370 18080
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 9364 18040 10701 18068
rect 9364 18028 9370 18040
rect 10689 18037 10701 18040
rect 10735 18037 10747 18071
rect 10689 18031 10747 18037
rect 12894 18028 12900 18080
rect 12952 18068 12958 18080
rect 13538 18068 13544 18080
rect 12952 18040 13544 18068
rect 12952 18028 12958 18040
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 13814 18068 13820 18080
rect 13775 18040 13820 18068
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 15105 18071 15163 18077
rect 13964 18040 14009 18068
rect 13964 18028 13970 18040
rect 15105 18037 15117 18071
rect 15151 18068 15163 18071
rect 17218 18068 17224 18080
rect 15151 18040 17224 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 17218 18028 17224 18040
rect 17276 18028 17282 18080
rect 17678 18028 17684 18080
rect 17736 18068 17742 18080
rect 19076 18068 19104 18244
rect 20073 18241 20085 18244
rect 20119 18241 20131 18275
rect 20073 18235 20131 18241
rect 19242 18096 19248 18148
rect 19300 18136 19306 18148
rect 19981 18139 20039 18145
rect 19981 18136 19993 18139
rect 19300 18108 19993 18136
rect 19300 18096 19306 18108
rect 19981 18105 19993 18108
rect 20027 18105 20039 18139
rect 19981 18099 20039 18105
rect 17736 18040 19104 18068
rect 17736 18028 17742 18040
rect 19426 18028 19432 18080
rect 19484 18068 19490 18080
rect 19889 18071 19947 18077
rect 19889 18068 19901 18071
rect 19484 18040 19901 18068
rect 19484 18028 19490 18040
rect 19889 18037 19901 18040
rect 19935 18037 19947 18071
rect 19889 18031 19947 18037
rect 1104 17978 20884 18000
rect 1104 17926 7579 17978
rect 7631 17926 7643 17978
rect 7695 17926 7707 17978
rect 7759 17926 7771 17978
rect 7823 17926 14176 17978
rect 14228 17926 14240 17978
rect 14292 17926 14304 17978
rect 14356 17926 14368 17978
rect 14420 17926 20884 17978
rect 1104 17904 20884 17926
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 3513 17867 3571 17873
rect 2832 17836 2925 17864
rect 2832 17824 2838 17836
rect 3513 17833 3525 17867
rect 3559 17864 3571 17867
rect 4062 17864 4068 17876
rect 3559 17836 4068 17864
rect 3559 17833 3571 17836
rect 3513 17827 3571 17833
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 4890 17824 4896 17876
rect 4948 17864 4954 17876
rect 5721 17867 5779 17873
rect 5721 17864 5733 17867
rect 4948 17836 5733 17864
rect 4948 17824 4954 17836
rect 5721 17833 5733 17836
rect 5767 17833 5779 17867
rect 5721 17827 5779 17833
rect 6104 17836 9076 17864
rect 2792 17796 2820 17824
rect 3970 17796 3976 17808
rect 2792 17768 3976 17796
rect 3970 17756 3976 17768
rect 4028 17756 4034 17808
rect 4982 17796 4988 17808
rect 4080 17768 4988 17796
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 1670 17737 1676 17740
rect 1664 17728 1676 17737
rect 1631 17700 1676 17728
rect 1664 17691 1676 17700
rect 1670 17688 1676 17691
rect 1728 17688 1734 17740
rect 4080 17737 4108 17768
rect 4982 17756 4988 17768
rect 5040 17756 5046 17808
rect 6104 17805 6132 17836
rect 6089 17799 6147 17805
rect 6089 17765 6101 17799
rect 6135 17765 6147 17799
rect 6270 17796 6276 17808
rect 6231 17768 6276 17796
rect 6089 17759 6147 17765
rect 6270 17756 6276 17768
rect 6328 17756 6334 17808
rect 6457 17799 6515 17805
rect 6457 17765 6469 17799
rect 6503 17796 6515 17799
rect 6730 17796 6736 17808
rect 6503 17768 6736 17796
rect 6503 17765 6515 17768
rect 6457 17759 6515 17765
rect 6730 17756 6736 17768
rect 6788 17756 6794 17808
rect 6914 17805 6920 17808
rect 6908 17796 6920 17805
rect 6875 17768 6920 17796
rect 6908 17759 6920 17768
rect 6914 17756 6920 17759
rect 6972 17756 6978 17808
rect 7926 17756 7932 17808
rect 7984 17796 7990 17808
rect 9048 17796 9076 17836
rect 9122 17824 9128 17876
rect 9180 17864 9186 17876
rect 9309 17867 9367 17873
rect 9309 17864 9321 17867
rect 9180 17836 9321 17864
rect 9180 17824 9186 17836
rect 9309 17833 9321 17836
rect 9355 17833 9367 17867
rect 11238 17864 11244 17876
rect 11199 17836 11244 17864
rect 9309 17827 9367 17833
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 12805 17867 12863 17873
rect 12805 17864 12817 17867
rect 12492 17836 12817 17864
rect 12492 17824 12498 17836
rect 12805 17833 12817 17836
rect 12851 17833 12863 17867
rect 12805 17827 12863 17833
rect 13909 17867 13967 17873
rect 13909 17833 13921 17867
rect 13955 17864 13967 17867
rect 13998 17864 14004 17876
rect 13955 17836 14004 17864
rect 13955 17833 13967 17836
rect 13909 17827 13967 17833
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 15470 17864 15476 17876
rect 15120 17836 15476 17864
rect 9398 17796 9404 17808
rect 7984 17768 8984 17796
rect 9048 17768 9404 17796
rect 7984 17756 7990 17768
rect 3605 17731 3663 17737
rect 3605 17697 3617 17731
rect 3651 17728 3663 17731
rect 4065 17731 4123 17737
rect 3651 17700 4016 17728
rect 3651 17697 3663 17700
rect 3605 17691 3663 17697
rect 3789 17663 3847 17669
rect 3789 17629 3801 17663
rect 3835 17660 3847 17663
rect 3878 17660 3884 17672
rect 3835 17632 3884 17660
rect 3835 17629 3847 17632
rect 3789 17623 3847 17629
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 3988 17660 4016 17700
rect 4065 17697 4077 17731
rect 4111 17697 4123 17731
rect 4065 17691 4123 17697
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17728 4767 17731
rect 5629 17731 5687 17737
rect 4755 17700 4936 17728
rect 4755 17697 4767 17700
rect 4709 17691 4767 17697
rect 4614 17660 4620 17672
rect 3988 17632 4620 17660
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 4798 17660 4804 17672
rect 4759 17632 4804 17660
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 2406 17552 2412 17604
rect 2464 17592 2470 17604
rect 4908 17592 4936 17700
rect 5629 17697 5641 17731
rect 5675 17728 5687 17731
rect 5902 17728 5908 17740
rect 5675 17700 5908 17728
rect 5675 17697 5687 17700
rect 5629 17691 5687 17697
rect 4985 17663 5043 17669
rect 4985 17629 4997 17663
rect 5031 17660 5043 17663
rect 5534 17660 5540 17672
rect 5031 17632 5540 17660
rect 5031 17629 5043 17632
rect 4985 17623 5043 17629
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 5644 17592 5672 17691
rect 5902 17688 5908 17700
rect 5960 17688 5966 17740
rect 7282 17688 7288 17740
rect 7340 17728 7346 17740
rect 8481 17731 8539 17737
rect 8481 17728 8493 17731
rect 7340 17700 8493 17728
rect 7340 17688 7346 17700
rect 8481 17697 8493 17700
rect 8527 17697 8539 17731
rect 8481 17691 8539 17697
rect 8573 17731 8631 17737
rect 8573 17697 8585 17731
rect 8619 17728 8631 17731
rect 8846 17728 8852 17740
rect 8619 17700 8852 17728
rect 8619 17697 8631 17700
rect 8573 17691 8631 17697
rect 8846 17688 8852 17700
rect 8904 17688 8910 17740
rect 8956 17737 8984 17768
rect 9398 17756 9404 17768
rect 9456 17756 9462 17808
rect 10128 17799 10186 17805
rect 10128 17765 10140 17799
rect 10174 17796 10186 17799
rect 11330 17796 11336 17808
rect 10174 17768 11336 17796
rect 10174 17765 10186 17768
rect 10128 17759 10186 17765
rect 11330 17756 11336 17768
rect 11388 17756 11394 17808
rect 11600 17799 11658 17805
rect 11600 17765 11612 17799
rect 11646 17796 11658 17799
rect 12066 17796 12072 17808
rect 11646 17768 12072 17796
rect 11646 17765 11658 17768
rect 11600 17759 11658 17765
rect 12066 17756 12072 17768
rect 12124 17756 12130 17808
rect 12342 17756 12348 17808
rect 12400 17796 12406 17808
rect 12400 17768 13391 17796
rect 12400 17756 12406 17768
rect 8941 17731 8999 17737
rect 8941 17697 8953 17731
rect 8987 17697 8999 17731
rect 8941 17691 8999 17697
rect 9582 17688 9588 17740
rect 9640 17728 9646 17740
rect 13173 17731 13231 17737
rect 13173 17728 13185 17731
rect 9640 17700 13185 17728
rect 9640 17688 9646 17700
rect 13173 17697 13185 17700
rect 13219 17697 13231 17731
rect 13173 17691 13231 17697
rect 5810 17660 5816 17672
rect 5771 17632 5816 17660
rect 5810 17620 5816 17632
rect 5868 17620 5874 17672
rect 6638 17660 6644 17672
rect 6599 17632 6644 17660
rect 6638 17620 6644 17632
rect 6696 17620 6702 17672
rect 8665 17663 8723 17669
rect 8665 17660 8677 17663
rect 8036 17632 8677 17660
rect 8036 17604 8064 17632
rect 8665 17629 8677 17632
rect 8711 17629 8723 17663
rect 9674 17660 9680 17672
rect 8665 17623 8723 17629
rect 8864 17632 9680 17660
rect 8018 17592 8024 17604
rect 2464 17564 4936 17592
rect 5184 17564 5672 17592
rect 7979 17564 8024 17592
rect 2464 17552 2470 17564
rect 1578 17484 1584 17536
rect 1636 17524 1642 17536
rect 3145 17527 3203 17533
rect 3145 17524 3157 17527
rect 1636 17496 3157 17524
rect 1636 17484 1642 17496
rect 3145 17493 3157 17496
rect 3191 17493 3203 17527
rect 3145 17487 3203 17493
rect 4341 17527 4399 17533
rect 4341 17493 4353 17527
rect 4387 17524 4399 17527
rect 5184 17524 5212 17564
rect 8018 17552 8024 17564
rect 8076 17552 8082 17604
rect 8110 17552 8116 17604
rect 8168 17592 8174 17604
rect 8168 17564 8213 17592
rect 8168 17552 8174 17564
rect 4387 17496 5212 17524
rect 5261 17527 5319 17533
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 5261 17493 5273 17527
rect 5307 17524 5319 17527
rect 8864 17524 8892 17632
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 9861 17663 9919 17669
rect 9861 17629 9873 17663
rect 9907 17629 9919 17663
rect 9861 17623 9919 17629
rect 9030 17552 9036 17604
rect 9088 17592 9094 17604
rect 9876 17592 9904 17623
rect 11238 17620 11244 17672
rect 11296 17660 11302 17672
rect 11333 17663 11391 17669
rect 11333 17660 11345 17663
rect 11296 17632 11345 17660
rect 11296 17620 11302 17632
rect 11333 17629 11345 17632
rect 11379 17629 11391 17663
rect 11333 17623 11391 17629
rect 12986 17620 12992 17672
rect 13044 17660 13050 17672
rect 13363 17669 13391 17768
rect 14090 17756 14096 17808
rect 14148 17796 14154 17808
rect 14826 17796 14832 17808
rect 14148 17768 14832 17796
rect 14148 17756 14154 17768
rect 14826 17756 14832 17768
rect 14884 17756 14890 17808
rect 13725 17731 13783 17737
rect 13725 17697 13737 17731
rect 13771 17728 13783 17731
rect 14734 17728 14740 17740
rect 13771 17700 14504 17728
rect 14695 17700 14740 17728
rect 13771 17697 13783 17700
rect 13725 17691 13783 17697
rect 13265 17663 13323 17669
rect 13265 17660 13277 17663
rect 13044 17632 13277 17660
rect 13044 17620 13050 17632
rect 13265 17629 13277 17632
rect 13311 17629 13323 17663
rect 13265 17623 13323 17629
rect 13357 17663 13415 17669
rect 13357 17629 13369 17663
rect 13403 17629 13415 17663
rect 13357 17623 13415 17629
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13688 17632 14105 17660
rect 13688 17620 13694 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 12710 17592 12716 17604
rect 9088 17564 9904 17592
rect 12671 17564 12716 17592
rect 9088 17552 9094 17564
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 14476 17592 14504 17700
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 14829 17663 14887 17669
rect 14829 17660 14841 17663
rect 14608 17632 14841 17660
rect 14608 17620 14614 17632
rect 14829 17629 14841 17632
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17660 15071 17663
rect 15120 17660 15148 17836
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 15841 17867 15899 17873
rect 15841 17833 15853 17867
rect 15887 17864 15899 17867
rect 15930 17864 15936 17876
rect 15887 17836 15936 17864
rect 15887 17833 15899 17836
rect 15841 17827 15899 17833
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 16393 17867 16451 17873
rect 16393 17864 16405 17867
rect 16172 17836 16405 17864
rect 16172 17824 16178 17836
rect 16393 17833 16405 17836
rect 16439 17833 16451 17867
rect 16393 17827 16451 17833
rect 16482 17824 16488 17876
rect 16540 17864 16546 17876
rect 18046 17864 18052 17876
rect 16540 17836 16585 17864
rect 16684 17836 18052 17864
rect 16540 17824 16546 17836
rect 16684 17796 16712 17836
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 18322 17824 18328 17876
rect 18380 17864 18386 17876
rect 19337 17867 19395 17873
rect 19337 17864 19349 17867
rect 18380 17836 19349 17864
rect 18380 17824 18386 17836
rect 19337 17833 19349 17836
rect 19383 17833 19395 17867
rect 19337 17827 19395 17833
rect 15059 17632 15148 17660
rect 15212 17768 16712 17796
rect 17589 17799 17647 17805
rect 15059 17629 15071 17632
rect 15013 17623 15071 17629
rect 15212 17592 15240 17768
rect 17589 17765 17601 17799
rect 17635 17796 17647 17799
rect 17954 17796 17960 17808
rect 17635 17768 17960 17796
rect 17635 17765 17647 17768
rect 17589 17759 17647 17765
rect 17954 17756 17960 17768
rect 18012 17756 18018 17808
rect 18138 17756 18144 17808
rect 18196 17756 18202 17808
rect 19797 17799 19855 17805
rect 19797 17765 19809 17799
rect 19843 17796 19855 17799
rect 19886 17796 19892 17808
rect 19843 17768 19892 17796
rect 19843 17765 19855 17768
rect 19797 17759 19855 17765
rect 19886 17756 19892 17768
rect 19944 17756 19950 17808
rect 15289 17731 15347 17737
rect 15289 17697 15301 17731
rect 15335 17697 15347 17731
rect 15289 17691 15347 17697
rect 15657 17731 15715 17737
rect 15657 17697 15669 17731
rect 15703 17728 15715 17731
rect 16206 17728 16212 17740
rect 15703 17700 16212 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 15304 17660 15332 17691
rect 16206 17688 16212 17700
rect 16264 17688 16270 17740
rect 17497 17731 17555 17737
rect 17497 17697 17509 17731
rect 17543 17728 17555 17731
rect 17770 17728 17776 17740
rect 17543 17700 17776 17728
rect 17543 17697 17555 17700
rect 17497 17691 17555 17697
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 18156 17728 18184 17756
rect 17972 17700 18184 17728
rect 18224 17731 18282 17737
rect 15838 17660 15844 17672
rect 15304 17632 15844 17660
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16390 17660 16396 17672
rect 15948 17632 16396 17660
rect 14476 17564 15240 17592
rect 15473 17595 15531 17601
rect 15473 17561 15485 17595
rect 15519 17592 15531 17595
rect 15948 17592 15976 17632
rect 16390 17620 16396 17632
rect 16448 17620 16454 17672
rect 16574 17660 16580 17672
rect 16535 17632 16580 17660
rect 16574 17620 16580 17632
rect 16632 17660 16638 17672
rect 17678 17660 17684 17672
rect 16632 17632 17684 17660
rect 16632 17620 16638 17632
rect 17678 17620 17684 17632
rect 17736 17620 17742 17672
rect 17972 17669 18000 17700
rect 18224 17697 18236 17731
rect 18270 17728 18282 17731
rect 19426 17728 19432 17740
rect 18270 17700 19432 17728
rect 18270 17697 18282 17700
rect 18224 17691 18282 17697
rect 19426 17688 19432 17700
rect 19484 17688 19490 17740
rect 20254 17728 20260 17740
rect 20215 17700 20260 17728
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 17957 17663 18015 17669
rect 17957 17629 17969 17663
rect 18003 17629 18015 17663
rect 17957 17623 18015 17629
rect 19150 17620 19156 17672
rect 19208 17660 19214 17672
rect 19889 17663 19947 17669
rect 19889 17660 19901 17663
rect 19208 17632 19901 17660
rect 19208 17620 19214 17632
rect 19889 17629 19901 17632
rect 19935 17629 19947 17663
rect 20070 17660 20076 17672
rect 20031 17632 20076 17660
rect 19889 17623 19947 17629
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 15519 17564 15976 17592
rect 16025 17595 16083 17601
rect 15519 17561 15531 17564
rect 15473 17555 15531 17561
rect 16025 17561 16037 17595
rect 16071 17592 16083 17595
rect 16666 17592 16672 17604
rect 16071 17564 16672 17592
rect 16071 17561 16083 17564
rect 16025 17555 16083 17561
rect 16666 17552 16672 17564
rect 16724 17552 16730 17604
rect 19429 17595 19487 17601
rect 19429 17561 19441 17595
rect 19475 17592 19487 17595
rect 20990 17592 20996 17604
rect 19475 17564 20996 17592
rect 19475 17561 19487 17564
rect 19429 17555 19487 17561
rect 20990 17552 20996 17564
rect 21048 17552 21054 17604
rect 9122 17524 9128 17536
rect 5307 17496 8892 17524
rect 9083 17496 9128 17524
rect 5307 17493 5319 17496
rect 5261 17487 5319 17493
rect 9122 17484 9128 17496
rect 9180 17484 9186 17536
rect 14369 17527 14427 17533
rect 14369 17493 14381 17527
rect 14415 17524 14427 17527
rect 14826 17524 14832 17536
rect 14415 17496 14832 17524
rect 14415 17493 14427 17496
rect 14369 17487 14427 17493
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 17129 17527 17187 17533
rect 17129 17524 17141 17527
rect 16172 17496 17141 17524
rect 16172 17484 16178 17496
rect 17129 17493 17141 17496
rect 17175 17493 17187 17527
rect 17129 17487 17187 17493
rect 19150 17484 19156 17536
rect 19208 17524 19214 17536
rect 20441 17527 20499 17533
rect 20441 17524 20453 17527
rect 19208 17496 20453 17524
rect 19208 17484 19214 17496
rect 20441 17493 20453 17496
rect 20487 17493 20499 17527
rect 20441 17487 20499 17493
rect 1104 17434 20884 17456
rect 1104 17382 4280 17434
rect 4332 17382 4344 17434
rect 4396 17382 4408 17434
rect 4460 17382 4472 17434
rect 4524 17382 10878 17434
rect 10930 17382 10942 17434
rect 10994 17382 11006 17434
rect 11058 17382 11070 17434
rect 11122 17382 17475 17434
rect 17527 17382 17539 17434
rect 17591 17382 17603 17434
rect 17655 17382 17667 17434
rect 17719 17382 20884 17434
rect 1104 17360 20884 17382
rect 5718 17320 5724 17332
rect 5679 17292 5724 17320
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 5810 17280 5816 17332
rect 5868 17320 5874 17332
rect 8573 17323 8631 17329
rect 8573 17320 8585 17323
rect 5868 17292 8585 17320
rect 5868 17280 5874 17292
rect 8573 17289 8585 17292
rect 8619 17289 8631 17323
rect 8573 17283 8631 17289
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 11238 17320 11244 17332
rect 8720 17292 9812 17320
rect 8720 17280 8726 17292
rect 1581 17255 1639 17261
rect 1581 17221 1593 17255
rect 1627 17252 1639 17255
rect 1762 17252 1768 17264
rect 1627 17224 1768 17252
rect 1627 17221 1639 17224
rect 1581 17215 1639 17221
rect 1762 17212 1768 17224
rect 1820 17212 1826 17264
rect 3878 17184 3884 17196
rect 3839 17156 3884 17184
rect 3878 17144 3884 17156
rect 3936 17144 3942 17196
rect 4706 17184 4712 17196
rect 4619 17156 4712 17184
rect 4706 17144 4712 17156
rect 4764 17184 4770 17196
rect 4982 17184 4988 17196
rect 4764 17156 4988 17184
rect 4764 17144 4770 17156
rect 4982 17144 4988 17156
rect 5040 17184 5046 17196
rect 5350 17184 5356 17196
rect 5040 17156 5356 17184
rect 5040 17144 5046 17156
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17184 5503 17187
rect 5534 17184 5540 17196
rect 5491 17156 5540 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 5534 17144 5540 17156
rect 5592 17184 5598 17196
rect 5718 17184 5724 17196
rect 5592 17156 5724 17184
rect 5592 17144 5598 17156
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17184 6423 17187
rect 6454 17184 6460 17196
rect 6411 17156 6460 17184
rect 6411 17153 6423 17156
rect 6365 17147 6423 17153
rect 6454 17144 6460 17156
rect 6512 17144 6518 17196
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 6788 17156 7052 17184
rect 6788 17144 6794 17156
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 1397 17119 1455 17125
rect 1397 17116 1409 17119
rect 1360 17088 1409 17116
rect 1360 17076 1366 17088
rect 1397 17085 1409 17088
rect 1443 17085 1455 17119
rect 1397 17079 1455 17085
rect 1486 17076 1492 17128
rect 1544 17116 1550 17128
rect 1765 17119 1823 17125
rect 1765 17116 1777 17119
rect 1544 17088 1777 17116
rect 1544 17076 1550 17088
rect 1765 17085 1777 17088
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 3142 17076 3148 17128
rect 3200 17116 3206 17128
rect 3605 17119 3663 17125
rect 3605 17116 3617 17119
rect 3200 17088 3617 17116
rect 3200 17076 3206 17088
rect 3605 17085 3617 17088
rect 3651 17085 3663 17119
rect 3605 17079 3663 17085
rect 3697 17119 3755 17125
rect 3697 17085 3709 17119
rect 3743 17116 3755 17119
rect 4154 17116 4160 17128
rect 3743 17088 4160 17116
rect 3743 17085 3755 17088
rect 3697 17079 3755 17085
rect 4154 17076 4160 17088
rect 4212 17076 4218 17128
rect 4433 17119 4491 17125
rect 4433 17085 4445 17119
rect 4479 17116 4491 17119
rect 5074 17116 5080 17128
rect 4479 17088 5080 17116
rect 4479 17085 4491 17088
rect 4433 17079 4491 17085
rect 5074 17076 5080 17088
rect 5132 17076 5138 17128
rect 6638 17076 6644 17128
rect 6696 17116 6702 17128
rect 6914 17116 6920 17128
rect 6696 17088 6920 17116
rect 6696 17076 6702 17088
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 7024 17116 7052 17156
rect 7926 17144 7932 17196
rect 7984 17184 7990 17196
rect 7984 17156 8892 17184
rect 7984 17144 7990 17156
rect 8389 17119 8447 17125
rect 8389 17116 8401 17119
rect 7024 17088 8401 17116
rect 8389 17085 8401 17088
rect 8435 17085 8447 17119
rect 8389 17079 8447 17085
rect 8478 17076 8484 17128
rect 8536 17116 8542 17128
rect 8757 17119 8815 17125
rect 8757 17116 8769 17119
rect 8536 17088 8769 17116
rect 8536 17076 8542 17088
rect 8757 17085 8769 17088
rect 8803 17085 8815 17119
rect 8757 17079 8815 17085
rect 2032 17051 2090 17057
rect 2032 17017 2044 17051
rect 2078 17048 2090 17051
rect 2130 17048 2136 17060
rect 2078 17020 2136 17048
rect 2078 17017 2090 17020
rect 2032 17011 2090 17017
rect 2130 17008 2136 17020
rect 2188 17008 2194 17060
rect 2682 17008 2688 17060
rect 2740 17048 2746 17060
rect 3510 17048 3516 17060
rect 2740 17020 3516 17048
rect 2740 17008 2746 17020
rect 3510 17008 3516 17020
rect 3568 17008 3574 17060
rect 4338 17008 4344 17060
rect 4396 17048 4402 17060
rect 5261 17051 5319 17057
rect 5261 17048 5273 17051
rect 4396 17020 5273 17048
rect 4396 17008 4402 17020
rect 5261 17017 5273 17020
rect 5307 17017 5319 17051
rect 5261 17011 5319 17017
rect 7184 17051 7242 17057
rect 7184 17017 7196 17051
rect 7230 17048 7242 17051
rect 7466 17048 7472 17060
rect 7230 17020 7472 17048
rect 7230 17017 7242 17020
rect 7184 17011 7242 17017
rect 7466 17008 7472 17020
rect 7524 17048 7530 17060
rect 8864 17048 8892 17156
rect 9024 17119 9082 17125
rect 9024 17085 9036 17119
rect 9070 17116 9082 17119
rect 9306 17116 9312 17128
rect 9070 17088 9312 17116
rect 9070 17085 9082 17088
rect 9024 17079 9082 17085
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 9784 17116 9812 17292
rect 10888 17292 11244 17320
rect 10778 17212 10784 17264
rect 10836 17252 10842 17264
rect 10888 17252 10916 17292
rect 11238 17280 11244 17292
rect 11296 17320 11302 17332
rect 12526 17320 12532 17332
rect 11296 17292 12532 17320
rect 11296 17280 11302 17292
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 13262 17320 13268 17332
rect 13223 17292 13268 17320
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 17770 17320 17776 17332
rect 17731 17292 17776 17320
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 19426 17320 19432 17332
rect 17880 17292 19003 17320
rect 19387 17292 19432 17320
rect 10836 17224 10916 17252
rect 12544 17252 12572 17280
rect 12544 17224 14228 17252
rect 10836 17212 10842 17224
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10888 17193 10916 17224
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10008 17156 10609 17184
rect 10008 17144 10014 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17184 13139 17187
rect 13170 17184 13176 17196
rect 13127 17156 13176 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 13814 17184 13820 17196
rect 13775 17156 13820 17184
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 14200 17193 14228 17224
rect 15286 17212 15292 17264
rect 15344 17252 15350 17264
rect 15749 17255 15807 17261
rect 15749 17252 15761 17255
rect 15344 17224 15761 17252
rect 15344 17212 15350 17224
rect 15749 17221 15761 17224
rect 15795 17221 15807 17255
rect 17880 17252 17908 17292
rect 15749 17215 15807 17221
rect 15856 17224 17908 17252
rect 18975 17252 19003 17292
rect 19426 17280 19432 17292
rect 19484 17280 19490 17332
rect 19521 17323 19579 17329
rect 19521 17289 19533 17323
rect 19567 17320 19579 17323
rect 19794 17320 19800 17332
rect 19567 17292 19800 17320
rect 19567 17289 19579 17292
rect 19521 17283 19579 17289
rect 19794 17280 19800 17292
rect 19852 17280 19858 17332
rect 18975 17224 20116 17252
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 15194 17144 15200 17196
rect 15252 17184 15258 17196
rect 15856 17184 15884 17224
rect 16022 17184 16028 17196
rect 15252 17156 15884 17184
rect 15948 17156 16028 17184
rect 15252 17144 15258 17156
rect 10229 17119 10287 17125
rect 10229 17116 10241 17119
rect 9784 17088 10241 17116
rect 10229 17085 10241 17088
rect 10275 17085 10287 17119
rect 10229 17079 10287 17085
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17116 12863 17119
rect 13630 17116 13636 17128
rect 12851 17088 13492 17116
rect 13591 17088 13636 17116
rect 12851 17085 12863 17088
rect 12805 17079 12863 17085
rect 9858 17048 9864 17060
rect 7524 17020 8708 17048
rect 8864 17020 9864 17048
rect 7524 17008 7530 17020
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 3145 16983 3203 16989
rect 3145 16980 3157 16983
rect 1728 16952 3157 16980
rect 1728 16940 1734 16952
rect 3145 16949 3157 16952
rect 3191 16949 3203 16983
rect 3145 16943 3203 16949
rect 3234 16940 3240 16992
rect 3292 16980 3298 16992
rect 4062 16980 4068 16992
rect 3292 16952 3337 16980
rect 4023 16952 4068 16980
rect 3292 16940 3298 16952
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 4525 16983 4583 16989
rect 4525 16949 4537 16983
rect 4571 16980 4583 16983
rect 4614 16980 4620 16992
rect 4571 16952 4620 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 4614 16940 4620 16952
rect 4672 16940 4678 16992
rect 4893 16983 4951 16989
rect 4893 16949 4905 16983
rect 4939 16980 4951 16983
rect 4982 16980 4988 16992
rect 4939 16952 4988 16980
rect 4939 16949 4951 16952
rect 4893 16943 4951 16949
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 5353 16983 5411 16989
rect 5353 16949 5365 16983
rect 5399 16980 5411 16983
rect 5626 16980 5632 16992
rect 5399 16952 5632 16980
rect 5399 16949 5411 16952
rect 5353 16943 5411 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 6086 16980 6092 16992
rect 6047 16952 6092 16980
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 6181 16983 6239 16989
rect 6181 16949 6193 16983
rect 6227 16980 6239 16983
rect 7926 16980 7932 16992
rect 6227 16952 7932 16980
rect 6227 16949 6239 16952
rect 6181 16943 6239 16949
rect 7926 16940 7932 16952
rect 7984 16940 7990 16992
rect 8018 16940 8024 16992
rect 8076 16980 8082 16992
rect 8297 16983 8355 16989
rect 8297 16980 8309 16983
rect 8076 16952 8309 16980
rect 8076 16940 8082 16952
rect 8297 16949 8309 16952
rect 8343 16949 8355 16983
rect 8680 16980 8708 17020
rect 9858 17008 9864 17020
rect 9916 17008 9922 17060
rect 9950 17008 9956 17060
rect 10008 17048 10014 17060
rect 10594 17048 10600 17060
rect 10008 17020 10600 17048
rect 10008 17008 10014 17020
rect 10594 17008 10600 17020
rect 10652 17008 10658 17060
rect 11140 17051 11198 17057
rect 11140 17017 11152 17051
rect 11186 17048 11198 17051
rect 11422 17048 11428 17060
rect 11186 17020 11428 17048
rect 11186 17017 11198 17020
rect 11140 17011 11198 17017
rect 11422 17008 11428 17020
rect 11480 17008 11486 17060
rect 11514 17008 11520 17060
rect 11572 17048 11578 17060
rect 12986 17048 12992 17060
rect 11572 17020 12992 17048
rect 11572 17008 11578 17020
rect 12986 17008 12992 17020
rect 13044 17008 13050 17060
rect 13464 17048 13492 17088
rect 13630 17076 13636 17088
rect 13688 17076 13694 17128
rect 13725 17119 13783 17125
rect 13725 17085 13737 17119
rect 13771 17116 13783 17119
rect 13906 17116 13912 17128
rect 13771 17088 13912 17116
rect 13771 17085 13783 17088
rect 13725 17079 13783 17085
rect 13906 17076 13912 17088
rect 13964 17076 13970 17128
rect 15470 17076 15476 17128
rect 15528 17116 15534 17128
rect 15948 17116 15976 17156
rect 16022 17144 16028 17156
rect 16080 17184 16086 17196
rect 16301 17187 16359 17193
rect 16301 17184 16313 17187
rect 16080 17156 16313 17184
rect 16080 17144 16086 17156
rect 16301 17153 16313 17156
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 20088 17193 20116 17224
rect 17129 17187 17187 17193
rect 17129 17184 17141 17187
rect 16632 17156 17141 17184
rect 16632 17144 16638 17156
rect 17129 17153 17141 17156
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 16114 17116 16120 17128
rect 15528 17088 15976 17116
rect 16075 17088 16120 17116
rect 15528 17076 15534 17088
rect 16114 17076 16120 17088
rect 16172 17076 16178 17128
rect 16758 17076 16764 17128
rect 16816 17116 16822 17128
rect 17589 17119 17647 17125
rect 17589 17116 17601 17119
rect 16816 17088 17601 17116
rect 16816 17076 16822 17088
rect 17589 17085 17601 17088
rect 17635 17085 17647 17119
rect 17589 17079 17647 17085
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 18138 17116 18144 17128
rect 18095 17088 18144 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 18316 17119 18374 17125
rect 18316 17085 18328 17119
rect 18362 17116 18374 17119
rect 19242 17116 19248 17128
rect 18362 17088 19248 17116
rect 18362 17085 18374 17088
rect 18316 17079 18374 17085
rect 19242 17076 19248 17088
rect 19300 17076 19306 17128
rect 19518 17076 19524 17128
rect 19576 17116 19582 17128
rect 19889 17119 19947 17125
rect 19889 17116 19901 17119
rect 19576 17088 19901 17116
rect 19576 17076 19582 17088
rect 19889 17085 19901 17088
rect 19935 17085 19947 17119
rect 19889 17079 19947 17085
rect 14090 17048 14096 17060
rect 13464 17020 14096 17048
rect 14090 17008 14096 17020
rect 14148 17008 14154 17060
rect 14458 17057 14464 17060
rect 14452 17048 14464 17057
rect 14419 17020 14464 17048
rect 14452 17011 14464 17020
rect 14458 17008 14464 17011
rect 14516 17008 14522 17060
rect 19794 17008 19800 17060
rect 19852 17048 19858 17060
rect 19981 17051 20039 17057
rect 19981 17048 19993 17051
rect 19852 17020 19993 17048
rect 19852 17008 19858 17020
rect 19981 17017 19993 17020
rect 20027 17017 20039 17051
rect 19981 17011 20039 17017
rect 10137 16983 10195 16989
rect 10137 16980 10149 16983
rect 8680 16952 10149 16980
rect 8297 16943 8355 16949
rect 10137 16949 10149 16952
rect 10183 16949 10195 16983
rect 10137 16943 10195 16949
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10413 16983 10471 16989
rect 10413 16980 10425 16983
rect 10284 16952 10425 16980
rect 10284 16940 10290 16952
rect 10413 16949 10425 16952
rect 10459 16949 10471 16983
rect 10413 16943 10471 16949
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 11974 16980 11980 16992
rect 10744 16952 11980 16980
rect 10744 16940 10750 16952
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 12250 16980 12256 16992
rect 12211 16952 12256 16980
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 12342 16940 12348 16992
rect 12400 16980 12406 16992
rect 12437 16983 12495 16989
rect 12437 16980 12449 16983
rect 12400 16952 12449 16980
rect 12400 16940 12406 16952
rect 12437 16949 12449 16952
rect 12483 16949 12495 16983
rect 12437 16943 12495 16949
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 12952 16952 12997 16980
rect 12952 16940 12958 16952
rect 13998 16940 14004 16992
rect 14056 16980 14062 16992
rect 15470 16980 15476 16992
rect 14056 16952 15476 16980
rect 14056 16940 14062 16952
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 15565 16983 15623 16989
rect 15565 16949 15577 16983
rect 15611 16980 15623 16983
rect 15654 16980 15660 16992
rect 15611 16952 15660 16980
rect 15611 16949 15623 16952
rect 15565 16943 15623 16949
rect 15654 16940 15660 16952
rect 15712 16940 15718 16992
rect 16209 16983 16267 16989
rect 16209 16949 16221 16983
rect 16255 16980 16267 16983
rect 16577 16983 16635 16989
rect 16577 16980 16589 16983
rect 16255 16952 16589 16980
rect 16255 16949 16267 16952
rect 16209 16943 16267 16949
rect 16577 16949 16589 16952
rect 16623 16949 16635 16983
rect 16577 16943 16635 16949
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 16724 16952 16957 16980
rect 16724 16940 16730 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 16945 16943 17003 16949
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 17092 16952 17137 16980
rect 17092 16940 17098 16952
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 20070 16980 20076 16992
rect 17368 16952 20076 16980
rect 17368 16940 17374 16952
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 1104 16890 20884 16912
rect 1104 16838 7579 16890
rect 7631 16838 7643 16890
rect 7695 16838 7707 16890
rect 7759 16838 7771 16890
rect 7823 16838 14176 16890
rect 14228 16838 14240 16890
rect 14292 16838 14304 16890
rect 14356 16838 14368 16890
rect 14420 16838 20884 16890
rect 1104 16816 20884 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 2314 16776 2320 16788
rect 1627 16748 2320 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 2314 16736 2320 16748
rect 2372 16736 2378 16788
rect 3145 16779 3203 16785
rect 3145 16745 3157 16779
rect 3191 16745 3203 16779
rect 3145 16739 3203 16745
rect 3421 16779 3479 16785
rect 3421 16745 3433 16779
rect 3467 16776 3479 16779
rect 3510 16776 3516 16788
rect 3467 16748 3516 16776
rect 3467 16745 3479 16748
rect 3421 16739 3479 16745
rect 2038 16717 2044 16720
rect 2032 16708 2044 16717
rect 1999 16680 2044 16708
rect 2032 16671 2044 16680
rect 2038 16668 2044 16671
rect 2096 16668 2102 16720
rect 2130 16668 2136 16720
rect 2188 16668 2194 16720
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16609 1455 16643
rect 1397 16603 1455 16609
rect 1412 16572 1440 16603
rect 1486 16600 1492 16652
rect 1544 16640 1550 16652
rect 1765 16643 1823 16649
rect 1765 16640 1777 16643
rect 1544 16612 1777 16640
rect 1544 16600 1550 16612
rect 1765 16609 1777 16612
rect 1811 16640 1823 16643
rect 1854 16640 1860 16652
rect 1811 16612 1860 16640
rect 1811 16609 1823 16612
rect 1765 16603 1823 16609
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 2148 16640 2176 16668
rect 3160 16640 3188 16739
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 4338 16776 4344 16788
rect 4299 16748 4344 16776
rect 4338 16736 4344 16748
rect 4396 16736 4402 16788
rect 4525 16779 4583 16785
rect 4525 16745 4537 16779
rect 4571 16776 4583 16779
rect 5353 16779 5411 16785
rect 4571 16748 5304 16776
rect 4571 16745 4583 16748
rect 4525 16739 4583 16745
rect 3970 16708 3976 16720
rect 3252 16680 3976 16708
rect 3252 16649 3280 16680
rect 3970 16668 3976 16680
rect 4028 16668 4034 16720
rect 4890 16708 4896 16720
rect 4851 16680 4896 16708
rect 4890 16668 4896 16680
rect 4948 16668 4954 16720
rect 2148 16612 3188 16640
rect 3237 16643 3295 16649
rect 3237 16609 3249 16643
rect 3283 16609 3295 16643
rect 3237 16603 3295 16609
rect 3605 16643 3663 16649
rect 3605 16609 3617 16643
rect 3651 16640 3663 16643
rect 3694 16640 3700 16652
rect 3651 16612 3700 16640
rect 3651 16609 3663 16612
rect 3605 16603 3663 16609
rect 3694 16600 3700 16612
rect 3752 16600 3758 16652
rect 4154 16640 4160 16652
rect 4115 16612 4160 16640
rect 4154 16600 4160 16612
rect 4212 16600 4218 16652
rect 4985 16643 5043 16649
rect 4985 16640 4997 16643
rect 4632 16612 4997 16640
rect 1578 16572 1584 16584
rect 1412 16544 1584 16572
rect 1578 16532 1584 16544
rect 1636 16532 1642 16584
rect 3326 16464 3332 16516
rect 3384 16504 3390 16516
rect 3789 16507 3847 16513
rect 3789 16504 3801 16507
rect 3384 16476 3801 16504
rect 3384 16464 3390 16476
rect 3789 16473 3801 16476
rect 3835 16473 3847 16507
rect 4632 16504 4660 16612
rect 4985 16609 4997 16612
rect 5031 16609 5043 16643
rect 5276 16640 5304 16748
rect 5353 16745 5365 16779
rect 5399 16745 5411 16779
rect 5353 16739 5411 16745
rect 5368 16708 5396 16739
rect 5626 16736 5632 16788
rect 5684 16776 5690 16788
rect 6365 16779 6423 16785
rect 6365 16776 6377 16779
rect 5684 16748 6377 16776
rect 5684 16736 5690 16748
rect 6365 16745 6377 16748
rect 6411 16745 6423 16779
rect 6365 16739 6423 16745
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7098 16776 7104 16788
rect 6972 16748 7104 16776
rect 6972 16736 6978 16748
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 7282 16776 7288 16788
rect 7243 16748 7288 16776
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 8119 16779 8177 16785
rect 8119 16745 8131 16779
rect 8165 16776 8177 16779
rect 8386 16776 8392 16788
rect 8165 16748 8392 16776
rect 8165 16745 8177 16748
rect 8119 16739 8177 16745
rect 8386 16736 8392 16748
rect 8444 16776 8450 16788
rect 8662 16776 8668 16788
rect 8444 16748 8668 16776
rect 8444 16736 8450 16748
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 8846 16736 8852 16788
rect 8904 16776 8910 16788
rect 9493 16779 9551 16785
rect 9493 16776 9505 16779
rect 8904 16748 9505 16776
rect 8904 16736 8910 16748
rect 9493 16745 9505 16748
rect 9539 16745 9551 16779
rect 11606 16776 11612 16788
rect 9493 16739 9551 16745
rect 9600 16748 11100 16776
rect 11567 16748 11612 16776
rect 9600 16708 9628 16748
rect 5368 16680 6224 16708
rect 5721 16643 5779 16649
rect 5721 16640 5733 16643
rect 5276 16612 5733 16640
rect 4985 16603 5043 16609
rect 5721 16609 5733 16612
rect 5767 16609 5779 16643
rect 5721 16603 5779 16609
rect 5810 16600 5816 16652
rect 5868 16640 5874 16652
rect 6196 16649 6224 16680
rect 9508 16680 9628 16708
rect 11072 16708 11100 16748
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 11974 16776 11980 16788
rect 11935 16748 11980 16776
rect 11974 16736 11980 16748
rect 12032 16776 12038 16788
rect 12894 16776 12900 16788
rect 12032 16748 12900 16776
rect 12032 16736 12038 16748
rect 12894 16736 12900 16748
rect 12952 16736 12958 16788
rect 13538 16736 13544 16788
rect 13596 16776 13602 16788
rect 14001 16779 14059 16785
rect 13596 16748 13952 16776
rect 13596 16736 13602 16748
rect 11514 16708 11520 16720
rect 11072 16680 11520 16708
rect 6181 16643 6239 16649
rect 5868 16612 5913 16640
rect 5868 16600 5874 16612
rect 6181 16609 6193 16643
rect 6227 16609 6239 16643
rect 6181 16603 6239 16609
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 7098 16640 7104 16652
rect 6595 16612 7104 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 7098 16600 7104 16612
rect 7156 16600 7162 16652
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16640 7251 16643
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 7239 16612 8401 16640
rect 7239 16609 7251 16612
rect 7193 16603 7251 16609
rect 8389 16609 8401 16612
rect 8435 16640 8447 16643
rect 9508 16640 9536 16680
rect 11514 16668 11520 16680
rect 11572 16668 11578 16720
rect 12796 16711 12854 16717
rect 12796 16677 12808 16711
rect 12842 16708 12854 16711
rect 13814 16708 13820 16720
rect 12842 16680 13820 16708
rect 12842 16677 12854 16680
rect 12796 16671 12854 16677
rect 13814 16668 13820 16680
rect 13872 16668 13878 16720
rect 13924 16708 13952 16748
rect 14001 16745 14013 16779
rect 14047 16776 14059 16779
rect 14550 16776 14556 16788
rect 14047 16748 14556 16776
rect 14047 16745 14059 16748
rect 14001 16739 14059 16745
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 14734 16736 14740 16788
rect 14792 16776 14798 16788
rect 15289 16779 15347 16785
rect 15289 16776 15301 16779
rect 14792 16748 15301 16776
rect 14792 16736 14798 16748
rect 15289 16745 15301 16748
rect 15335 16745 15347 16779
rect 15289 16739 15347 16745
rect 15470 16736 15476 16788
rect 15528 16776 15534 16788
rect 17310 16776 17316 16788
rect 15528 16748 17316 16776
rect 15528 16736 15534 16748
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 17773 16779 17831 16785
rect 17773 16745 17785 16779
rect 17819 16776 17831 16779
rect 17954 16776 17960 16788
rect 17819 16748 17960 16776
rect 17819 16745 17831 16748
rect 17773 16739 17831 16745
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 19242 16776 19248 16788
rect 19203 16748 19248 16776
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 20346 16776 20352 16788
rect 20307 16748 20352 16776
rect 20346 16736 20352 16748
rect 20404 16736 20410 16788
rect 14369 16711 14427 16717
rect 13924 16680 14320 16708
rect 10413 16643 10471 16649
rect 8435 16612 9536 16640
rect 9600 16612 10180 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 9600 16584 9628 16612
rect 4706 16532 4712 16584
rect 4764 16572 4770 16584
rect 5077 16575 5135 16581
rect 5077 16572 5089 16575
rect 4764 16544 5089 16572
rect 4764 16532 4770 16544
rect 5077 16541 5089 16544
rect 5123 16541 5135 16575
rect 5994 16572 6000 16584
rect 5907 16544 6000 16572
rect 5077 16535 5135 16541
rect 5994 16532 6000 16544
rect 6052 16572 6058 16584
rect 7466 16572 7472 16584
rect 6052 16544 7328 16572
rect 7427 16544 7472 16572
rect 6052 16532 6058 16544
rect 7190 16504 7196 16516
rect 4632 16476 7196 16504
rect 3789 16467 3847 16473
rect 7190 16464 7196 16476
rect 7248 16464 7254 16516
rect 7300 16504 7328 16544
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 7653 16575 7711 16581
rect 7653 16541 7665 16575
rect 7699 16572 7711 16575
rect 8018 16572 8024 16584
rect 7699 16544 8024 16572
rect 7699 16541 7711 16544
rect 7653 16535 7711 16541
rect 8018 16532 8024 16544
rect 8076 16532 8082 16584
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 8168 16544 8213 16572
rect 8168 16532 8174 16544
rect 8294 16532 8300 16584
rect 8352 16572 8358 16584
rect 9582 16572 9588 16584
rect 8352 16544 9588 16572
rect 8352 16532 8358 16544
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 9677 16575 9735 16581
rect 9677 16541 9689 16575
rect 9723 16541 9735 16575
rect 9677 16535 9735 16541
rect 7300 16476 7420 16504
rect 2958 16396 2964 16448
rect 3016 16436 3022 16448
rect 6086 16436 6092 16448
rect 3016 16408 6092 16436
rect 3016 16396 3022 16408
rect 6086 16396 6092 16408
rect 6144 16396 6150 16448
rect 6825 16439 6883 16445
rect 6825 16405 6837 16439
rect 6871 16436 6883 16439
rect 7282 16436 7288 16448
rect 6871 16408 7288 16436
rect 6871 16405 6883 16408
rect 6825 16399 6883 16405
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 7392 16436 7420 16476
rect 9122 16436 9128 16448
rect 7392 16408 9128 16436
rect 9122 16396 9128 16408
rect 9180 16396 9186 16448
rect 9692 16436 9720 16535
rect 9858 16532 9864 16584
rect 9916 16572 9922 16584
rect 10152 16581 10180 16612
rect 10413 16609 10425 16643
rect 10459 16640 10471 16643
rect 12526 16640 12532 16652
rect 10459 16612 11560 16640
rect 12487 16612 12532 16640
rect 10459 16609 10471 16612
rect 10413 16603 10471 16609
rect 10000 16575 10058 16581
rect 10000 16572 10012 16575
rect 9916 16544 10012 16572
rect 9916 16532 9922 16544
rect 10000 16541 10012 16544
rect 10046 16541 10058 16575
rect 10000 16535 10058 16541
rect 10140 16575 10198 16581
rect 10140 16541 10152 16575
rect 10186 16541 10198 16575
rect 11532 16572 11560 16612
rect 12526 16600 12532 16612
rect 12584 16600 12590 16652
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 14292 16640 14320 16680
rect 14369 16677 14381 16711
rect 14415 16708 14427 16711
rect 14458 16708 14464 16720
rect 14415 16680 14464 16708
rect 14415 16677 14427 16680
rect 14369 16671 14427 16677
rect 14458 16668 14464 16680
rect 14516 16668 14522 16720
rect 16408 16680 17908 16708
rect 14826 16640 14832 16652
rect 12676 16612 13676 16640
rect 14292 16612 14596 16640
rect 14787 16612 14832 16640
rect 12676 16600 12682 16612
rect 12066 16572 12072 16584
rect 11532 16544 12072 16572
rect 10140 16535 10198 16541
rect 12066 16532 12072 16544
rect 12124 16532 12130 16584
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16541 12219 16575
rect 13648 16572 13676 16612
rect 13648 16544 13768 16572
rect 12161 16535 12219 16541
rect 11330 16464 11336 16516
rect 11388 16504 11394 16516
rect 12176 16504 12204 16535
rect 11388 16476 12204 16504
rect 11388 16464 11394 16476
rect 10318 16436 10324 16448
rect 9692 16408 10324 16436
rect 10318 16396 10324 16408
rect 10376 16396 10382 16448
rect 11514 16436 11520 16448
rect 11475 16408 11520 16436
rect 11514 16396 11520 16408
rect 11572 16396 11578 16448
rect 13740 16436 13768 16544
rect 13814 16532 13820 16584
rect 13872 16572 13878 16584
rect 14568 16581 14596 16612
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 15654 16640 15660 16652
rect 15615 16612 15660 16640
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 15804 16612 15849 16640
rect 15804 16600 15810 16612
rect 15930 16600 15936 16652
rect 15988 16640 15994 16652
rect 16408 16649 16436 16680
rect 16666 16649 16672 16652
rect 16393 16643 16451 16649
rect 16393 16640 16405 16643
rect 15988 16612 16405 16640
rect 15988 16600 15994 16612
rect 16393 16609 16405 16612
rect 16439 16609 16451 16643
rect 16660 16640 16672 16649
rect 16627 16612 16672 16640
rect 16393 16603 16451 16609
rect 16660 16603 16672 16612
rect 16666 16600 16672 16603
rect 16724 16600 16730 16652
rect 17880 16649 17908 16680
rect 18046 16668 18052 16720
rect 18104 16717 18110 16720
rect 18104 16711 18168 16717
rect 18104 16677 18122 16711
rect 18156 16677 18168 16711
rect 18104 16671 18168 16677
rect 18104 16668 18110 16671
rect 18230 16668 18236 16720
rect 18288 16668 18294 16720
rect 17865 16643 17923 16649
rect 17865 16609 17877 16643
rect 17911 16640 17923 16643
rect 18248 16640 18276 16668
rect 17911 16612 18276 16640
rect 17911 16609 17923 16612
rect 17865 16603 17923 16609
rect 19610 16600 19616 16652
rect 19668 16640 19674 16652
rect 19705 16643 19763 16649
rect 19705 16640 19717 16643
rect 19668 16612 19717 16640
rect 19668 16600 19674 16612
rect 19705 16609 19717 16612
rect 19751 16609 19763 16643
rect 19705 16603 19763 16609
rect 20165 16643 20223 16649
rect 20165 16609 20177 16643
rect 20211 16640 20223 16643
rect 20622 16640 20628 16652
rect 20211 16612 20628 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 14461 16575 14519 16581
rect 14461 16572 14473 16575
rect 13872 16544 14473 16572
rect 13872 16532 13878 16544
rect 14461 16541 14473 16544
rect 14507 16541 14519 16575
rect 14461 16535 14519 16541
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16572 14611 16575
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 14599 16544 15853 16572
rect 14599 16541 14611 16544
rect 14553 16535 14611 16541
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 13906 16504 13912 16516
rect 13819 16476 13912 16504
rect 13906 16464 13912 16476
rect 13964 16504 13970 16516
rect 14918 16504 14924 16516
rect 13964 16476 14924 16504
rect 13964 16464 13970 16476
rect 14918 16464 14924 16476
rect 14976 16464 14982 16516
rect 15013 16439 15071 16445
rect 15013 16436 15025 16439
rect 13740 16408 15025 16436
rect 15013 16405 15025 16408
rect 15059 16405 15071 16439
rect 15856 16436 15884 16535
rect 19426 16532 19432 16584
rect 19484 16572 19490 16584
rect 19797 16575 19855 16581
rect 19797 16572 19809 16575
rect 19484 16544 19809 16572
rect 19484 16532 19490 16544
rect 19797 16541 19809 16544
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16572 20039 16575
rect 20070 16572 20076 16584
rect 20027 16544 20076 16572
rect 20027 16541 20039 16544
rect 19981 16535 20039 16541
rect 20070 16532 20076 16544
rect 20128 16532 20134 16584
rect 18874 16464 18880 16516
rect 18932 16504 18938 16516
rect 19702 16504 19708 16516
rect 18932 16476 19708 16504
rect 18932 16464 18938 16476
rect 19702 16464 19708 16476
rect 19760 16464 19766 16516
rect 16574 16436 16580 16448
rect 15856 16408 16580 16436
rect 15013 16399 15071 16405
rect 16574 16396 16580 16408
rect 16632 16396 16638 16448
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 19392 16408 19437 16436
rect 19392 16396 19398 16408
rect 1104 16346 20884 16368
rect 1104 16294 4280 16346
rect 4332 16294 4344 16346
rect 4396 16294 4408 16346
rect 4460 16294 4472 16346
rect 4524 16294 10878 16346
rect 10930 16294 10942 16346
rect 10994 16294 11006 16346
rect 11058 16294 11070 16346
rect 11122 16294 17475 16346
rect 17527 16294 17539 16346
rect 17591 16294 17603 16346
rect 17655 16294 17667 16346
rect 17719 16294 20884 16346
rect 1104 16272 20884 16294
rect 3605 16235 3663 16241
rect 1504 16204 3556 16232
rect 1504 16037 1532 16204
rect 3237 16167 3295 16173
rect 3237 16133 3249 16167
rect 3283 16164 3295 16167
rect 3418 16164 3424 16176
rect 3283 16136 3424 16164
rect 3283 16133 3295 16136
rect 3237 16127 3295 16133
rect 3418 16124 3424 16136
rect 3476 16124 3482 16176
rect 3528 16164 3556 16204
rect 3605 16201 3617 16235
rect 3651 16232 3663 16235
rect 4154 16232 4160 16244
rect 3651 16204 4160 16232
rect 3651 16201 3663 16204
rect 3605 16195 3663 16201
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 4982 16232 4988 16244
rect 4816 16204 4988 16232
rect 4816 16164 4844 16204
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 5718 16192 5724 16244
rect 5776 16232 5782 16244
rect 6457 16235 6515 16241
rect 6457 16232 6469 16235
rect 5776 16204 6469 16232
rect 5776 16192 5782 16204
rect 6457 16201 6469 16204
rect 6503 16201 6515 16235
rect 6457 16195 6515 16201
rect 7285 16235 7343 16241
rect 7285 16201 7297 16235
rect 7331 16232 7343 16235
rect 7926 16232 7932 16244
rect 7331 16204 7932 16232
rect 7331 16201 7343 16204
rect 7285 16195 7343 16201
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 8754 16232 8760 16244
rect 8128 16204 8760 16232
rect 8128 16164 8156 16204
rect 8754 16192 8760 16204
rect 8812 16192 8818 16244
rect 9953 16235 10011 16241
rect 9953 16201 9965 16235
rect 9999 16232 10011 16235
rect 10134 16232 10140 16244
rect 9999 16204 10140 16232
rect 9999 16201 10011 16204
rect 9953 16195 10011 16201
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 12066 16192 12072 16244
rect 12124 16232 12130 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 12124 16204 12173 16232
rect 12124 16192 12130 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 13078 16232 13084 16244
rect 12161 16195 12219 16201
rect 12728 16204 13084 16232
rect 3528 16136 4844 16164
rect 6288 16136 8156 16164
rect 1854 16096 1860 16108
rect 1815 16068 1860 16096
rect 1854 16056 1860 16068
rect 1912 16056 1918 16108
rect 3602 16096 3608 16108
rect 3436 16068 3608 16096
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 15997 1547 16031
rect 1489 15991 1547 15997
rect 2124 16031 2182 16037
rect 2124 15997 2136 16031
rect 2170 16028 2182 16031
rect 3436 16028 3464 16068
rect 3602 16056 3608 16068
rect 3660 16056 3666 16108
rect 4062 16096 4068 16108
rect 4023 16068 4068 16096
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16065 4215 16099
rect 4157 16059 4215 16065
rect 2170 16000 3464 16028
rect 3513 16031 3571 16037
rect 2170 15997 2182 16000
rect 2124 15991 2182 15997
rect 3513 15997 3525 16031
rect 3559 16028 3571 16031
rect 3694 16028 3700 16040
rect 3559 16000 3700 16028
rect 3559 15997 3571 16000
rect 3513 15991 3571 15997
rect 3694 15988 3700 16000
rect 3752 15988 3758 16040
rect 3878 15988 3884 16040
rect 3936 16028 3942 16040
rect 4172 16028 4200 16059
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 4801 16099 4859 16105
rect 4801 16096 4813 16099
rect 4304 16068 4813 16096
rect 4304 16056 4310 16068
rect 4801 16065 4813 16068
rect 4847 16065 4859 16099
rect 4801 16059 4859 16065
rect 3936 16000 4200 16028
rect 3936 15988 3942 16000
rect 2590 15920 2596 15972
rect 2648 15960 2654 15972
rect 3973 15963 4031 15969
rect 3973 15960 3985 15963
rect 2648 15932 3985 15960
rect 2648 15920 2654 15932
rect 3973 15929 3985 15932
rect 4019 15929 4031 15963
rect 4172 15960 4200 16000
rect 4433 16031 4491 16037
rect 4433 15997 4445 16031
rect 4479 16028 4491 16031
rect 5534 16028 5540 16040
rect 4479 16000 5540 16028
rect 4479 15997 4491 16000
rect 4433 15991 4491 15997
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 6288 16037 6316 16136
rect 7282 16056 7288 16108
rect 7340 16096 7346 16108
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7340 16068 7757 16096
rect 7340 16056 7346 16068
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 8576 16099 8634 16105
rect 7892 16068 7937 16096
rect 7892 16056 7898 16068
rect 8576 16065 8588 16099
rect 8622 16065 8634 16099
rect 8846 16096 8852 16108
rect 8807 16068 8852 16096
rect 8576 16059 8634 16065
rect 6273 16031 6331 16037
rect 6273 15997 6285 16031
rect 6319 15997 6331 16031
rect 6273 15991 6331 15997
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 15997 6975 16031
rect 6917 15991 6975 15997
rect 5068 15963 5126 15969
rect 4172 15932 4844 15960
rect 3973 15923 4031 15929
rect 1673 15895 1731 15901
rect 1673 15861 1685 15895
rect 1719 15892 1731 15895
rect 2958 15892 2964 15904
rect 1719 15864 2964 15892
rect 1719 15861 1731 15864
rect 1673 15855 1731 15861
rect 2958 15852 2964 15864
rect 3016 15852 3022 15904
rect 3329 15895 3387 15901
rect 3329 15861 3341 15895
rect 3375 15892 3387 15895
rect 4062 15892 4068 15904
rect 3375 15864 4068 15892
rect 3375 15861 3387 15864
rect 3329 15855 3387 15861
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 4617 15895 4675 15901
rect 4617 15861 4629 15895
rect 4663 15892 4675 15895
rect 4706 15892 4712 15904
rect 4663 15864 4712 15892
rect 4663 15861 4675 15864
rect 4617 15855 4675 15861
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 4816 15892 4844 15932
rect 5068 15929 5080 15963
rect 5114 15960 5126 15963
rect 6822 15960 6828 15972
rect 5114 15932 6828 15960
rect 5114 15929 5126 15932
rect 5068 15923 5126 15929
rect 6822 15920 6828 15932
rect 6880 15920 6886 15972
rect 6932 15960 6960 15991
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 7653 16031 7711 16037
rect 7653 16028 7665 16031
rect 7156 16000 7665 16028
rect 7156 15988 7162 16000
rect 7653 15997 7665 16000
rect 7699 15997 7711 16031
rect 7653 15991 7711 15997
rect 8018 15988 8024 16040
rect 8076 16028 8082 16040
rect 8113 16031 8171 16037
rect 8113 16028 8125 16031
rect 8076 16000 8125 16028
rect 8076 15988 8082 16000
rect 8113 15997 8125 16000
rect 8159 15997 8171 16031
rect 8113 15991 8171 15997
rect 8386 15988 8392 16040
rect 8444 16037 8450 16040
rect 8444 16031 8494 16037
rect 8444 15997 8448 16031
rect 8482 15997 8494 16031
rect 8588 16028 8616 16059
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 10045 16099 10103 16105
rect 10045 16065 10057 16099
rect 10091 16096 10103 16099
rect 10502 16096 10508 16108
rect 10091 16068 10508 16096
rect 10091 16065 10103 16068
rect 10045 16059 10103 16065
rect 10502 16056 10508 16068
rect 10560 16056 10566 16108
rect 10778 16096 10784 16108
rect 10742 16068 10784 16096
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 11057 16099 11115 16105
rect 11057 16065 11069 16099
rect 11103 16096 11115 16099
rect 12618 16096 12624 16108
rect 11103 16068 12624 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 10226 16028 10232 16040
rect 8588 16000 10232 16028
rect 8444 15991 8494 15997
rect 8444 15988 8450 15991
rect 10226 15988 10232 16000
rect 10284 15988 10290 16040
rect 10318 15988 10324 16040
rect 10376 16028 10382 16040
rect 12437 16031 12495 16037
rect 10376 16000 10421 16028
rect 10376 15988 10382 16000
rect 12437 15997 12449 16031
rect 12483 16028 12495 16031
rect 12728 16028 12756 16204
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 13998 16192 14004 16244
rect 14056 16232 14062 16244
rect 14185 16235 14243 16241
rect 14185 16232 14197 16235
rect 14056 16204 14197 16232
rect 14056 16192 14062 16204
rect 14185 16201 14197 16204
rect 14231 16232 14243 16235
rect 14918 16232 14924 16244
rect 14231 16204 14924 16232
rect 14231 16201 14243 16204
rect 14185 16195 14243 16201
rect 14918 16192 14924 16204
rect 14976 16192 14982 16244
rect 15654 16192 15660 16244
rect 15712 16232 15718 16244
rect 15933 16235 15991 16241
rect 15933 16232 15945 16235
rect 15712 16204 15945 16232
rect 15712 16192 15718 16204
rect 15933 16201 15945 16204
rect 15979 16201 15991 16235
rect 15933 16195 15991 16201
rect 16666 16192 16672 16244
rect 16724 16232 16730 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 16724 16204 17417 16232
rect 16724 16192 16730 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 18046 16192 18052 16244
rect 18104 16232 18110 16244
rect 19429 16235 19487 16241
rect 19429 16232 19441 16235
rect 18104 16204 19441 16232
rect 18104 16192 18110 16204
rect 19429 16201 19441 16204
rect 19475 16201 19487 16235
rect 19429 16195 19487 16201
rect 17126 16124 17132 16176
rect 17184 16164 17190 16176
rect 17681 16167 17739 16173
rect 17681 16164 17693 16167
rect 17184 16136 17693 16164
rect 17184 16124 17190 16136
rect 17681 16133 17693 16136
rect 17727 16133 17739 16167
rect 17681 16127 17739 16133
rect 15930 16056 15936 16108
rect 15988 16096 15994 16108
rect 16025 16099 16083 16105
rect 16025 16096 16037 16099
rect 15988 16068 16037 16096
rect 15988 16056 15994 16068
rect 16025 16065 16037 16068
rect 16071 16065 16083 16099
rect 20070 16096 20076 16108
rect 20031 16068 20076 16096
rect 16025 16059 16083 16065
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 12483 16000 12756 16028
rect 12805 16031 12863 16037
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 12805 15997 12817 16031
rect 12851 15997 12863 16031
rect 12805 15991 12863 15997
rect 13072 16031 13130 16037
rect 13072 15997 13084 16031
rect 13118 16028 13130 16031
rect 13906 16028 13912 16040
rect 13118 16000 13912 16028
rect 13118 15997 13130 16000
rect 13072 15991 13130 15997
rect 7926 15960 7932 15972
rect 6932 15932 7932 15960
rect 7926 15920 7932 15932
rect 7984 15920 7990 15972
rect 12526 15920 12532 15972
rect 12584 15960 12590 15972
rect 12710 15960 12716 15972
rect 12584 15932 12716 15960
rect 12584 15920 12590 15932
rect 12710 15920 12716 15932
rect 12768 15960 12774 15972
rect 12820 15960 12848 15991
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 16028 14611 16031
rect 14820 16031 14878 16037
rect 14599 16000 14780 16028
rect 14599 15997 14611 16000
rect 14553 15991 14611 15997
rect 12986 15960 12992 15972
rect 12768 15932 12992 15960
rect 12768 15920 12774 15932
rect 12986 15920 12992 15932
rect 13044 15920 13050 15972
rect 14090 15920 14096 15972
rect 14148 15920 14154 15972
rect 14277 15963 14335 15969
rect 14277 15929 14289 15963
rect 14323 15960 14335 15963
rect 14642 15960 14648 15972
rect 14323 15932 14648 15960
rect 14323 15929 14335 15932
rect 14277 15923 14335 15929
rect 14642 15920 14648 15932
rect 14700 15920 14706 15972
rect 5994 15892 6000 15904
rect 4816 15864 6000 15892
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 6178 15892 6184 15904
rect 6139 15864 6184 15892
rect 6178 15852 6184 15864
rect 6236 15852 6242 15904
rect 7101 15895 7159 15901
rect 7101 15861 7113 15895
rect 7147 15892 7159 15895
rect 8386 15892 8392 15904
rect 7147 15864 8392 15892
rect 7147 15861 7159 15864
rect 7101 15855 7159 15861
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 8662 15852 8668 15904
rect 8720 15892 8726 15904
rect 9582 15892 9588 15904
rect 8720 15864 9588 15892
rect 8720 15852 8726 15864
rect 9582 15852 9588 15864
rect 9640 15892 9646 15904
rect 10787 15895 10845 15901
rect 10787 15892 10799 15895
rect 9640 15864 10799 15892
rect 9640 15852 9646 15864
rect 10787 15861 10799 15864
rect 10833 15861 10845 15895
rect 10787 15855 10845 15861
rect 12621 15895 12679 15901
rect 12621 15861 12633 15895
rect 12667 15892 12679 15895
rect 14108 15892 14136 15920
rect 12667 15864 14136 15892
rect 14752 15892 14780 16000
rect 14820 15997 14832 16031
rect 14866 16028 14878 16031
rect 15746 16028 15752 16040
rect 14866 16000 15752 16028
rect 14866 15997 14878 16000
rect 14820 15991 14878 15997
rect 15746 15988 15752 16000
rect 15804 15988 15810 16040
rect 16292 16031 16350 16037
rect 16292 15997 16304 16031
rect 16338 16028 16350 16031
rect 17034 16028 17040 16040
rect 16338 16000 17040 16028
rect 16338 15997 16350 16000
rect 16292 15991 16350 15997
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 17218 15988 17224 16040
rect 17276 16028 17282 16040
rect 17497 16031 17555 16037
rect 17497 16028 17509 16031
rect 17276 16000 17509 16028
rect 17276 15988 17282 16000
rect 17497 15997 17509 16000
rect 17543 15997 17555 16031
rect 17497 15991 17555 15997
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18138 16028 18144 16040
rect 18095 16000 18144 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18138 15988 18144 16000
rect 18196 15988 18202 16040
rect 18598 15988 18604 16040
rect 18656 16028 18662 16040
rect 20088 16028 20116 16056
rect 18656 16000 20116 16028
rect 18656 15988 18662 16000
rect 14918 15920 14924 15972
rect 14976 15960 14982 15972
rect 15562 15960 15568 15972
rect 14976 15932 15568 15960
rect 14976 15920 14982 15932
rect 15562 15920 15568 15932
rect 15620 15920 15626 15972
rect 17954 15920 17960 15972
rect 18012 15960 18018 15972
rect 18294 15963 18352 15969
rect 18294 15960 18306 15963
rect 18012 15932 18306 15960
rect 18012 15920 18018 15932
rect 18294 15929 18306 15932
rect 18340 15929 18352 15963
rect 18294 15923 18352 15929
rect 18690 15920 18696 15972
rect 18748 15960 18754 15972
rect 19889 15963 19947 15969
rect 18748 15932 19564 15960
rect 18748 15920 18754 15932
rect 15470 15892 15476 15904
rect 14752 15864 15476 15892
rect 12667 15861 12679 15864
rect 12621 15855 12679 15861
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 19536 15901 19564 15932
rect 19889 15929 19901 15963
rect 19935 15960 19947 15963
rect 20346 15960 20352 15972
rect 19935 15932 20352 15960
rect 19935 15929 19947 15932
rect 19889 15923 19947 15929
rect 20346 15920 20352 15932
rect 20404 15920 20410 15972
rect 19521 15895 19579 15901
rect 19521 15861 19533 15895
rect 19567 15861 19579 15895
rect 19521 15855 19579 15861
rect 19978 15852 19984 15904
rect 20036 15892 20042 15904
rect 20036 15864 20081 15892
rect 20036 15852 20042 15864
rect 1104 15802 20884 15824
rect 1104 15750 7579 15802
rect 7631 15750 7643 15802
rect 7695 15750 7707 15802
rect 7759 15750 7771 15802
rect 7823 15750 14176 15802
rect 14228 15750 14240 15802
rect 14292 15750 14304 15802
rect 14356 15750 14368 15802
rect 14420 15750 20884 15802
rect 1104 15728 20884 15750
rect 3421 15691 3479 15697
rect 3421 15657 3433 15691
rect 3467 15688 3479 15691
rect 4798 15688 4804 15700
rect 3467 15660 4804 15688
rect 3467 15657 3479 15660
rect 3421 15651 3479 15657
rect 4798 15648 4804 15660
rect 4856 15648 4862 15700
rect 6914 15688 6920 15700
rect 6748 15660 6920 15688
rect 2032 15623 2090 15629
rect 2032 15589 2044 15623
rect 2078 15620 2090 15623
rect 2866 15620 2872 15632
rect 2078 15592 2872 15620
rect 2078 15589 2090 15592
rect 2032 15583 2090 15589
rect 2866 15580 2872 15592
rect 2924 15580 2930 15632
rect 4332 15623 4390 15629
rect 4332 15589 4344 15623
rect 4378 15620 4390 15623
rect 4614 15620 4620 15632
rect 4378 15592 4620 15620
rect 4378 15589 4390 15592
rect 4332 15583 4390 15589
rect 4614 15580 4620 15592
rect 4672 15580 4678 15632
rect 5804 15623 5862 15629
rect 5804 15589 5816 15623
rect 5850 15620 5862 15623
rect 6178 15620 6184 15632
rect 5850 15592 6184 15620
rect 5850 15589 5862 15592
rect 5804 15583 5862 15589
rect 6178 15580 6184 15592
rect 6236 15580 6242 15632
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15552 1823 15555
rect 1854 15552 1860 15564
rect 1811 15524 1860 15552
rect 1811 15521 1823 15524
rect 1765 15515 1823 15521
rect 1854 15512 1860 15524
rect 1912 15552 1918 15564
rect 3234 15552 3240 15564
rect 1912 15524 3096 15552
rect 3195 15524 3240 15552
rect 1912 15512 1918 15524
rect 3068 15484 3096 15524
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 3605 15555 3663 15561
rect 3605 15521 3617 15555
rect 3651 15552 3663 15555
rect 5166 15552 5172 15564
rect 3651 15524 5172 15552
rect 3651 15521 3663 15524
rect 3605 15515 3663 15521
rect 5166 15512 5172 15524
rect 5224 15512 5230 15564
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15552 5595 15555
rect 6748 15552 6776 15660
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 8389 15691 8447 15697
rect 8389 15688 8401 15691
rect 7248 15660 8401 15688
rect 7248 15648 7254 15660
rect 8389 15657 8401 15660
rect 8435 15657 8447 15691
rect 8389 15651 8447 15657
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 10686 15688 10692 15700
rect 8527 15660 10692 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 11057 15691 11115 15697
rect 11057 15657 11069 15691
rect 11103 15688 11115 15691
rect 11330 15688 11336 15700
rect 11103 15660 11336 15688
rect 11103 15657 11115 15660
rect 11057 15651 11115 15657
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 12250 15688 12256 15700
rect 11440 15660 12256 15688
rect 11440 15632 11468 15660
rect 12250 15648 12256 15660
rect 12308 15648 12314 15700
rect 14369 15691 14427 15697
rect 14369 15657 14381 15691
rect 14415 15688 14427 15691
rect 14458 15688 14464 15700
rect 14415 15660 14464 15688
rect 14415 15657 14427 15660
rect 14369 15651 14427 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 14645 15691 14703 15697
rect 14645 15657 14657 15691
rect 14691 15688 14703 15691
rect 14734 15688 14740 15700
rect 14691 15660 14740 15688
rect 14691 15657 14703 15660
rect 14645 15651 14703 15657
rect 14734 15648 14740 15660
rect 14792 15648 14798 15700
rect 15470 15648 15476 15700
rect 15528 15688 15534 15700
rect 15930 15688 15936 15700
rect 15528 15660 15936 15688
rect 15528 15648 15534 15660
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 16853 15691 16911 15697
rect 16853 15657 16865 15691
rect 16899 15688 16911 15691
rect 17034 15688 17040 15700
rect 16899 15660 17040 15688
rect 16899 15657 16911 15660
rect 16853 15651 16911 15657
rect 17034 15648 17040 15660
rect 17092 15648 17098 15700
rect 18509 15691 18567 15697
rect 18509 15657 18521 15691
rect 18555 15688 18567 15691
rect 19426 15688 19432 15700
rect 18555 15660 19432 15688
rect 18555 15657 18567 15660
rect 18509 15651 18567 15657
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 19978 15688 19984 15700
rect 19939 15660 19984 15688
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 6822 15580 6828 15632
rect 6880 15620 6886 15632
rect 11422 15620 11428 15632
rect 6880 15592 11428 15620
rect 6880 15580 6886 15592
rect 11422 15580 11428 15592
rect 11480 15580 11486 15632
rect 12434 15620 12440 15632
rect 11532 15592 12440 15620
rect 5583 15524 6868 15552
rect 5583 15521 5595 15524
rect 5537 15515 5595 15521
rect 4062 15484 4068 15496
rect 3068 15456 4068 15484
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 6840 15484 6868 15524
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 7265 15555 7323 15561
rect 7265 15552 7277 15555
rect 6972 15524 7277 15552
rect 6972 15512 6978 15524
rect 7265 15521 7277 15524
rect 7311 15521 7323 15555
rect 7265 15515 7323 15521
rect 8849 15555 8907 15561
rect 8849 15521 8861 15555
rect 8895 15552 8907 15555
rect 9309 15555 9367 15561
rect 9309 15552 9321 15555
rect 8895 15524 9321 15552
rect 8895 15521 8907 15524
rect 8849 15515 8907 15521
rect 9309 15521 9321 15524
rect 9355 15521 9367 15555
rect 9766 15552 9772 15564
rect 9309 15515 9367 15521
rect 9600 15524 9772 15552
rect 7009 15487 7067 15493
rect 7009 15484 7021 15487
rect 6840 15456 7021 15484
rect 7009 15453 7021 15456
rect 7055 15453 7067 15487
rect 7009 15447 7067 15453
rect 3145 15419 3203 15425
rect 3145 15385 3157 15419
rect 3191 15416 3203 15419
rect 3602 15416 3608 15428
rect 3191 15388 3608 15416
rect 3191 15385 3203 15388
rect 3145 15379 3203 15385
rect 3602 15376 3608 15388
rect 3660 15376 3666 15428
rect 6822 15376 6828 15428
rect 6880 15416 6886 15428
rect 7024 15416 7052 15447
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8352 15456 8953 15484
rect 8352 15444 8358 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9600 15484 9628 15524
rect 9766 15512 9772 15524
rect 9824 15552 9830 15564
rect 9933 15555 9991 15561
rect 9933 15552 9945 15555
rect 9824 15524 9945 15552
rect 9824 15512 9830 15524
rect 9933 15521 9945 15524
rect 9979 15521 9991 15555
rect 9933 15515 9991 15521
rect 10226 15512 10232 15564
rect 10284 15552 10290 15564
rect 10410 15552 10416 15564
rect 10284 15524 10416 15552
rect 10284 15512 10290 15524
rect 10410 15512 10416 15524
rect 10468 15512 10474 15564
rect 11532 15561 11560 15592
rect 12434 15580 12440 15592
rect 12492 15580 12498 15632
rect 13722 15580 13728 15632
rect 13780 15620 13786 15632
rect 15010 15620 15016 15632
rect 13780 15592 15016 15620
rect 13780 15580 13786 15592
rect 15010 15580 15016 15592
rect 15068 15580 15074 15632
rect 15654 15580 15660 15632
rect 15712 15629 15718 15632
rect 15712 15623 15776 15629
rect 15712 15589 15730 15623
rect 15764 15589 15776 15623
rect 15948 15620 15976 15648
rect 15948 15592 17172 15620
rect 15712 15583 15776 15589
rect 15712 15580 15718 15583
rect 11790 15561 11796 15564
rect 11517 15555 11575 15561
rect 11517 15521 11529 15555
rect 11563 15521 11575 15555
rect 11784 15552 11796 15561
rect 11751 15524 11796 15552
rect 11517 15515 11575 15521
rect 11784 15515 11796 15524
rect 11790 15512 11796 15515
rect 11848 15512 11854 15564
rect 13256 15555 13314 15561
rect 13256 15552 13268 15555
rect 12912 15524 13268 15552
rect 9171 15456 9628 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 11238 15484 11244 15496
rect 9732 15456 9777 15484
rect 11199 15456 11244 15484
rect 9732 15444 9738 15456
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 12912 15425 12940 15524
rect 13256 15521 13268 15524
rect 13302 15552 13314 15555
rect 13814 15552 13820 15564
rect 13302 15524 13820 15552
rect 13302 15521 13314 15524
rect 13256 15515 13314 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 14461 15555 14519 15561
rect 14461 15521 14473 15555
rect 14507 15521 14519 15555
rect 14461 15515 14519 15521
rect 14829 15555 14887 15561
rect 14829 15521 14841 15555
rect 14875 15552 14887 15555
rect 15286 15552 15292 15564
rect 14875 15524 15292 15552
rect 14875 15521 14887 15524
rect 14829 15515 14887 15521
rect 12986 15444 12992 15496
rect 13044 15484 13050 15496
rect 14476 15484 14504 15515
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 16850 15552 16856 15564
rect 15396 15524 16856 15552
rect 15396 15484 15424 15524
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 17144 15561 17172 15592
rect 17310 15580 17316 15632
rect 17368 15629 17374 15632
rect 17368 15623 17432 15629
rect 17368 15589 17386 15623
rect 17420 15589 17432 15623
rect 17368 15583 17432 15589
rect 17368 15580 17374 15583
rect 17129 15555 17187 15561
rect 17129 15521 17141 15555
rect 17175 15521 17187 15555
rect 17129 15515 17187 15521
rect 18138 15512 18144 15564
rect 18196 15552 18202 15564
rect 18601 15555 18659 15561
rect 18601 15552 18613 15555
rect 18196 15524 18613 15552
rect 18196 15512 18202 15524
rect 18601 15521 18613 15524
rect 18647 15521 18659 15555
rect 18601 15515 18659 15521
rect 18868 15555 18926 15561
rect 18868 15521 18880 15555
rect 18914 15552 18926 15555
rect 19610 15552 19616 15564
rect 18914 15524 19616 15552
rect 18914 15521 18926 15524
rect 18868 15515 18926 15521
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 20070 15552 20076 15564
rect 20031 15524 20076 15552
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 13044 15456 13089 15484
rect 14476 15456 15424 15484
rect 13044 15444 13050 15456
rect 15470 15444 15476 15496
rect 15528 15484 15534 15496
rect 15528 15456 15573 15484
rect 15528 15444 15534 15456
rect 6880 15388 7052 15416
rect 6880 15376 6886 15388
rect 3786 15348 3792 15360
rect 3699 15320 3792 15348
rect 3786 15308 3792 15320
rect 3844 15348 3850 15360
rect 4798 15348 4804 15360
rect 3844 15320 4804 15348
rect 3844 15308 3850 15320
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 5074 15308 5080 15360
rect 5132 15348 5138 15360
rect 5445 15351 5503 15357
rect 5445 15348 5457 15351
rect 5132 15320 5457 15348
rect 5132 15308 5138 15320
rect 5445 15317 5457 15320
rect 5491 15317 5503 15351
rect 6914 15348 6920 15360
rect 6875 15320 6920 15348
rect 5445 15311 5503 15317
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 7024 15348 7052 15388
rect 12897 15419 12955 15425
rect 12897 15385 12909 15419
rect 12943 15385 12955 15419
rect 12897 15379 12955 15385
rect 7650 15348 7656 15360
rect 7024 15320 7656 15348
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 8018 15308 8024 15360
rect 8076 15348 8082 15360
rect 10318 15348 10324 15360
rect 8076 15320 10324 15348
rect 8076 15308 8082 15320
rect 10318 15308 10324 15320
rect 10376 15308 10382 15360
rect 12802 15308 12808 15360
rect 12860 15348 12866 15360
rect 15013 15351 15071 15357
rect 15013 15348 15025 15351
rect 12860 15320 15025 15348
rect 12860 15308 12866 15320
rect 15013 15317 15025 15320
rect 15059 15317 15071 15351
rect 15013 15311 15071 15317
rect 18874 15308 18880 15360
rect 18932 15348 18938 15360
rect 20257 15351 20315 15357
rect 20257 15348 20269 15351
rect 18932 15320 20269 15348
rect 18932 15308 18938 15320
rect 20257 15317 20269 15320
rect 20303 15317 20315 15351
rect 20257 15311 20315 15317
rect 1104 15258 20884 15280
rect 1104 15206 4280 15258
rect 4332 15206 4344 15258
rect 4396 15206 4408 15258
rect 4460 15206 4472 15258
rect 4524 15206 10878 15258
rect 10930 15206 10942 15258
rect 10994 15206 11006 15258
rect 11058 15206 11070 15258
rect 11122 15206 17475 15258
rect 17527 15206 17539 15258
rect 17591 15206 17603 15258
rect 17655 15206 17667 15258
rect 17719 15206 20884 15258
rect 1104 15184 20884 15206
rect 1854 15144 1860 15156
rect 1504 15116 1860 15144
rect 1394 14968 1400 15020
rect 1452 15008 1458 15020
rect 1504 15017 1532 15116
rect 1854 15104 1860 15116
rect 1912 15104 1918 15156
rect 2866 15144 2872 15156
rect 2827 15116 2872 15144
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 4062 15144 4068 15156
rect 3436 15116 4068 15144
rect 3436 15017 3464 15116
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 4212 15116 4384 15144
rect 4212 15104 4218 15116
rect 4356 15076 4384 15116
rect 4614 15104 4620 15156
rect 4672 15144 4678 15156
rect 4801 15147 4859 15153
rect 4801 15144 4813 15147
rect 4672 15116 4813 15144
rect 4672 15104 4678 15116
rect 4801 15113 4813 15116
rect 4847 15113 4859 15147
rect 4801 15107 4859 15113
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 5810 15144 5816 15156
rect 5767 15116 5816 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 5810 15104 5816 15116
rect 5868 15104 5874 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 5920 15116 8217 15144
rect 4890 15076 4896 15088
rect 4356 15048 4896 15076
rect 4890 15036 4896 15048
rect 4948 15076 4954 15088
rect 5920 15076 5948 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8205 15107 8263 15113
rect 9677 15147 9735 15153
rect 9677 15113 9689 15147
rect 9723 15144 9735 15147
rect 9766 15144 9772 15156
rect 9723 15116 9772 15144
rect 9723 15113 9735 15116
rect 9677 15107 9735 15113
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 9876 15116 11928 15144
rect 4948 15048 5948 15076
rect 6012 15048 6316 15076
rect 4948 15036 4954 15048
rect 1489 15011 1547 15017
rect 1489 15008 1501 15011
rect 1452 14980 1501 15008
rect 1452 14968 1458 14980
rect 1489 14977 1501 14980
rect 1535 14977 1547 15011
rect 1489 14971 1547 14977
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 5445 15011 5503 15017
rect 5445 14977 5457 15011
rect 5491 14977 5503 15011
rect 5445 14971 5503 14977
rect 1756 14943 1814 14949
rect 1756 14909 1768 14943
rect 1802 14940 1814 14943
rect 2958 14940 2964 14952
rect 1802 14912 2964 14940
rect 1802 14909 1814 14912
rect 1756 14903 1814 14909
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 3053 14943 3111 14949
rect 3053 14909 3065 14943
rect 3099 14940 3111 14943
rect 3326 14940 3332 14952
rect 3099 14912 3332 14940
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 3510 14900 3516 14952
rect 3568 14940 3574 14952
rect 5353 14943 5411 14949
rect 5353 14940 5365 14943
rect 3568 14912 5365 14940
rect 3568 14900 3574 14912
rect 5353 14909 5365 14912
rect 5399 14909 5411 14943
rect 5460 14940 5488 14971
rect 5534 14968 5540 15020
rect 5592 15008 5598 15020
rect 6012 15008 6040 15048
rect 6178 15008 6184 15020
rect 5592 14980 6040 15008
rect 6139 14980 6184 15008
rect 5592 14968 5598 14980
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 6288 15017 6316 15048
rect 9306 15036 9312 15088
rect 9364 15076 9370 15088
rect 9876 15076 9904 15116
rect 9364 15048 9904 15076
rect 9364 15036 9370 15048
rect 10778 15036 10784 15088
rect 10836 15076 10842 15088
rect 10873 15079 10931 15085
rect 10873 15076 10885 15079
rect 10836 15048 10885 15076
rect 10836 15036 10842 15048
rect 10873 15045 10885 15048
rect 10919 15045 10931 15079
rect 10873 15039 10931 15045
rect 6273 15011 6331 15017
rect 6273 14977 6285 15011
rect 6319 14977 6331 15011
rect 6273 14971 6331 14977
rect 6380 14980 6960 15008
rect 6380 14940 6408 14980
rect 6822 14940 6828 14952
rect 5460 14912 6408 14940
rect 6783 14912 6828 14940
rect 5353 14903 5411 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6932 14940 6960 14980
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 10413 15011 10471 15017
rect 9732 14980 10272 15008
rect 9732 14968 9738 14980
rect 7374 14940 7380 14952
rect 6932 14912 7380 14940
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 7650 14900 7656 14952
rect 7708 14940 7714 14952
rect 8202 14940 8208 14952
rect 7708 14912 8208 14940
rect 7708 14900 7714 14912
rect 8202 14900 8208 14912
rect 8260 14940 8266 14952
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 8260 14912 8309 14940
rect 8260 14900 8266 14912
rect 8297 14909 8309 14912
rect 8343 14940 8355 14943
rect 9692 14940 9720 14968
rect 10134 14940 10140 14952
rect 8343 14912 9720 14940
rect 10095 14912 10140 14940
rect 8343 14909 8355 14912
rect 8297 14903 8355 14909
rect 10134 14900 10140 14912
rect 10192 14900 10198 14952
rect 10244 14940 10272 14980
rect 10413 14977 10425 15011
rect 10459 15008 10471 15011
rect 10594 15008 10600 15020
rect 10459 14980 10600 15008
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 11422 15008 11428 15020
rect 11383 14980 11428 15008
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 11238 14940 11244 14952
rect 10244 14912 10916 14940
rect 11199 14912 11244 14940
rect 3688 14875 3746 14881
rect 3688 14841 3700 14875
rect 3734 14872 3746 14875
rect 4154 14872 4160 14884
rect 3734 14844 4160 14872
rect 3734 14841 3746 14844
rect 3688 14835 3746 14841
rect 4154 14832 4160 14844
rect 4212 14832 4218 14884
rect 5261 14875 5319 14881
rect 5261 14872 5273 14875
rect 4264 14844 5273 14872
rect 3237 14807 3295 14813
rect 3237 14773 3249 14807
rect 3283 14804 3295 14807
rect 4264 14804 4292 14844
rect 5261 14841 5273 14844
rect 5307 14841 5319 14875
rect 5261 14835 5319 14841
rect 6089 14875 6147 14881
rect 6089 14841 6101 14875
rect 6135 14872 6147 14875
rect 6914 14872 6920 14884
rect 6135 14844 6920 14872
rect 6135 14841 6147 14844
rect 6089 14835 6147 14841
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 7092 14875 7150 14881
rect 7092 14841 7104 14875
rect 7138 14872 7150 14875
rect 7190 14872 7196 14884
rect 7138 14844 7196 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 7190 14832 7196 14844
rect 7248 14832 7254 14884
rect 8564 14875 8622 14881
rect 8564 14841 8576 14875
rect 8610 14872 8622 14875
rect 8662 14872 8668 14884
rect 8610 14844 8668 14872
rect 8610 14841 8622 14844
rect 8564 14835 8622 14841
rect 8662 14832 8668 14844
rect 8720 14832 8726 14884
rect 9674 14832 9680 14884
rect 9732 14872 9738 14884
rect 10229 14875 10287 14881
rect 10229 14872 10241 14875
rect 9732 14844 10241 14872
rect 9732 14832 9738 14844
rect 10229 14841 10241 14844
rect 10275 14841 10287 14875
rect 10229 14835 10287 14841
rect 10888 14816 10916 14912
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 11900 14949 11928 15116
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12989 15147 13047 15153
rect 12492 15116 12537 15144
rect 12492 15104 12498 15116
rect 12989 15113 13001 15147
rect 13035 15144 13047 15147
rect 15197 15147 15255 15153
rect 13035 15116 15148 15144
rect 13035 15113 13047 15116
rect 12989 15107 13047 15113
rect 15120 15076 15148 15116
rect 15197 15113 15209 15147
rect 15243 15144 15255 15147
rect 15286 15144 15292 15156
rect 15243 15116 15292 15144
rect 15243 15113 15255 15116
rect 15197 15107 15255 15113
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 15381 15147 15439 15153
rect 15381 15113 15393 15147
rect 15427 15144 15439 15147
rect 16850 15144 16856 15156
rect 15427 15116 16856 15144
rect 15427 15113 15439 15116
rect 15381 15107 15439 15113
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 18138 15144 18144 15156
rect 17727 15116 18144 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 18138 15104 18144 15116
rect 18196 15104 18202 15156
rect 18156 15076 18184 15104
rect 15120 15048 16252 15076
rect 18156 15048 19196 15076
rect 12986 14968 12992 15020
rect 13044 15008 13050 15020
rect 13173 15011 13231 15017
rect 13173 15008 13185 15011
rect 13044 14980 13185 15008
rect 13044 14968 13050 14980
rect 13173 14977 13185 14980
rect 13219 14977 13231 15011
rect 14826 15008 14832 15020
rect 13173 14971 13231 14977
rect 14660 14980 14832 15008
rect 11885 14943 11943 14949
rect 11885 14909 11897 14943
rect 11931 14909 11943 14943
rect 11885 14903 11943 14909
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12618 14940 12624 14952
rect 12299 14912 12624 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 12805 14943 12863 14949
rect 12805 14909 12817 14943
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 13440 14943 13498 14949
rect 13440 14909 13452 14943
rect 13486 14940 13498 14943
rect 13998 14940 14004 14952
rect 13486 14912 14004 14940
rect 13486 14909 13498 14912
rect 13440 14903 13498 14909
rect 11333 14875 11391 14881
rect 11333 14841 11345 14875
rect 11379 14872 11391 14875
rect 12342 14872 12348 14884
rect 11379 14844 12348 14872
rect 11379 14841 11391 14844
rect 11333 14835 11391 14841
rect 12342 14832 12348 14844
rect 12400 14832 12406 14884
rect 12820 14872 12848 14903
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 14660 14949 14688 14980
rect 14826 14968 14832 14980
rect 14884 14968 14890 15020
rect 16022 15008 16028 15020
rect 15983 14980 16028 15008
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 16224 15008 16252 15048
rect 16224 14980 16344 15008
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14909 14703 14943
rect 15010 14940 15016 14952
rect 14971 14912 15016 14940
rect 14645 14903 14703 14909
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 16209 14943 16267 14949
rect 16209 14940 16221 14943
rect 15344 14912 16221 14940
rect 15344 14900 15350 14912
rect 16209 14909 16221 14912
rect 16255 14909 16267 14943
rect 16316 14940 16344 14980
rect 18414 14968 18420 15020
rect 18472 15008 18478 15020
rect 18969 15011 19027 15017
rect 18969 15008 18981 15011
rect 18472 14980 18981 15008
rect 18472 14968 18478 14980
rect 18969 14977 18981 14980
rect 19015 15008 19027 15011
rect 19058 15008 19064 15020
rect 19015 14980 19064 15008
rect 19015 14977 19027 14980
rect 18969 14971 19027 14977
rect 19058 14968 19064 14980
rect 19116 14968 19122 15020
rect 19168 15017 19196 15048
rect 19153 15011 19211 15017
rect 19153 14977 19165 15011
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 16316 14912 16896 14940
rect 16209 14903 16267 14909
rect 14918 14872 14924 14884
rect 12820 14844 14924 14872
rect 14918 14832 14924 14844
rect 14976 14832 14982 14884
rect 16482 14881 16488 14884
rect 15841 14875 15899 14881
rect 15841 14841 15853 14875
rect 15887 14872 15899 14875
rect 16476 14872 16488 14881
rect 15887 14844 16488 14872
rect 15887 14841 15899 14844
rect 15841 14835 15899 14841
rect 16476 14835 16488 14844
rect 16482 14832 16488 14835
rect 16540 14832 16546 14884
rect 16868 14872 16896 14912
rect 17034 14900 17040 14952
rect 17092 14940 17098 14952
rect 17865 14943 17923 14949
rect 17865 14940 17877 14943
rect 17092 14912 17877 14940
rect 17092 14900 17098 14912
rect 17865 14909 17877 14912
rect 17911 14909 17923 14943
rect 18690 14940 18696 14952
rect 18651 14912 18696 14940
rect 17865 14903 17923 14909
rect 18690 14900 18696 14912
rect 18748 14900 18754 14952
rect 19420 14943 19478 14949
rect 19420 14909 19432 14943
rect 19466 14940 19478 14943
rect 19978 14940 19984 14952
rect 19466 14912 19984 14940
rect 19466 14909 19478 14912
rect 19420 14903 19478 14909
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 18785 14875 18843 14881
rect 16868 14844 18460 14872
rect 3283 14776 4292 14804
rect 4893 14807 4951 14813
rect 3283 14773 3295 14776
rect 3237 14767 3295 14773
rect 4893 14773 4905 14807
rect 4939 14804 4951 14807
rect 7926 14804 7932 14816
rect 4939 14776 7932 14804
rect 4939 14773 4951 14776
rect 4893 14767 4951 14773
rect 7926 14764 7932 14776
rect 7984 14764 7990 14816
rect 9766 14764 9772 14816
rect 9824 14804 9830 14816
rect 9824 14776 9869 14804
rect 9824 14764 9830 14776
rect 10410 14764 10416 14816
rect 10468 14804 10474 14816
rect 10597 14807 10655 14813
rect 10597 14804 10609 14807
rect 10468 14776 10609 14804
rect 10468 14764 10474 14776
rect 10597 14773 10609 14776
rect 10643 14773 10655 14807
rect 10597 14767 10655 14773
rect 10870 14764 10876 14816
rect 10928 14804 10934 14816
rect 11701 14807 11759 14813
rect 11701 14804 11713 14807
rect 10928 14776 11713 14804
rect 10928 14764 10934 14776
rect 11701 14773 11713 14776
rect 11747 14773 11759 14807
rect 12066 14804 12072 14816
rect 11979 14776 12072 14804
rect 11701 14767 11759 14773
rect 12066 14764 12072 14776
rect 12124 14804 12130 14816
rect 13538 14804 13544 14816
rect 12124 14776 13544 14804
rect 12124 14764 12130 14776
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 14550 14804 14556 14816
rect 14511 14776 14556 14804
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 14826 14804 14832 14816
rect 14787 14776 14832 14804
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 15749 14807 15807 14813
rect 15749 14773 15761 14807
rect 15795 14804 15807 14807
rect 17310 14804 17316 14816
rect 15795 14776 17316 14804
rect 15795 14773 15807 14776
rect 15749 14767 15807 14773
rect 17310 14764 17316 14776
rect 17368 14804 17374 14816
rect 17589 14807 17647 14813
rect 17589 14804 17601 14807
rect 17368 14776 17601 14804
rect 17368 14764 17374 14776
rect 17589 14773 17601 14776
rect 17635 14773 17647 14807
rect 17589 14767 17647 14773
rect 17770 14764 17776 14816
rect 17828 14804 17834 14816
rect 18325 14807 18383 14813
rect 18325 14804 18337 14807
rect 17828 14776 18337 14804
rect 17828 14764 17834 14776
rect 18325 14773 18337 14776
rect 18371 14773 18383 14807
rect 18432 14804 18460 14844
rect 18785 14841 18797 14875
rect 18831 14872 18843 14875
rect 19334 14872 19340 14884
rect 18831 14844 19340 14872
rect 18831 14841 18843 14844
rect 18785 14835 18843 14841
rect 19334 14832 19340 14844
rect 19392 14832 19398 14884
rect 18966 14804 18972 14816
rect 18432 14776 18972 14804
rect 18325 14767 18383 14773
rect 18966 14764 18972 14776
rect 19024 14764 19030 14816
rect 20346 14764 20352 14816
rect 20404 14804 20410 14816
rect 20533 14807 20591 14813
rect 20533 14804 20545 14807
rect 20404 14776 20545 14804
rect 20404 14764 20410 14776
rect 20533 14773 20545 14776
rect 20579 14773 20591 14807
rect 20533 14767 20591 14773
rect 1104 14714 20884 14736
rect 1104 14662 7579 14714
rect 7631 14662 7643 14714
rect 7695 14662 7707 14714
rect 7759 14662 7771 14714
rect 7823 14662 14176 14714
rect 14228 14662 14240 14714
rect 14292 14662 14304 14714
rect 14356 14662 14368 14714
rect 14420 14662 20884 14714
rect 1104 14640 20884 14662
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14569 2835 14603
rect 2777 14563 2835 14569
rect 2869 14603 2927 14609
rect 2869 14569 2881 14603
rect 2915 14600 2927 14603
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 2915 14572 4445 14600
rect 2915 14569 2927 14572
rect 2869 14563 2927 14569
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 4433 14563 4491 14569
rect 4893 14603 4951 14609
rect 4893 14569 4905 14603
rect 4939 14569 4951 14603
rect 4893 14563 4951 14569
rect 7193 14603 7251 14609
rect 7193 14569 7205 14603
rect 7239 14569 7251 14603
rect 7193 14563 7251 14569
rect 9217 14603 9275 14609
rect 9217 14569 9229 14603
rect 9263 14600 9275 14603
rect 9766 14600 9772 14612
rect 9263 14572 9772 14600
rect 9263 14569 9275 14572
rect 9217 14563 9275 14569
rect 2792 14532 2820 14563
rect 3050 14532 3056 14544
rect 2792 14504 3056 14532
rect 3050 14492 3056 14504
rect 3108 14492 3114 14544
rect 3237 14535 3295 14541
rect 3237 14532 3249 14535
rect 3160 14504 3249 14532
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 1664 14467 1722 14473
rect 1664 14433 1676 14467
rect 1710 14464 1722 14467
rect 1710 14436 2728 14464
rect 1710 14433 1722 14436
rect 1664 14427 1722 14433
rect 2700 14396 2728 14436
rect 2700 14368 3004 14396
rect 2976 14328 3004 14368
rect 3050 14356 3056 14408
rect 3108 14396 3114 14408
rect 3160 14396 3188 14504
rect 3237 14501 3249 14504
rect 3283 14501 3295 14535
rect 3237 14495 3295 14501
rect 3326 14492 3332 14544
rect 3384 14532 3390 14544
rect 4908 14532 4936 14563
rect 3384 14504 4936 14532
rect 3384 14492 3390 14504
rect 4982 14492 4988 14544
rect 5040 14532 5046 14544
rect 5353 14535 5411 14541
rect 5353 14532 5365 14535
rect 5040 14504 5365 14532
rect 5040 14492 5046 14504
rect 5353 14501 5365 14504
rect 5399 14501 5411 14535
rect 6822 14532 6828 14544
rect 5353 14495 5411 14501
rect 5828 14504 6828 14532
rect 3786 14464 3792 14476
rect 3436 14436 3792 14464
rect 3326 14396 3332 14408
rect 3108 14368 3188 14396
rect 3287 14368 3332 14396
rect 3108 14356 3114 14368
rect 3326 14356 3332 14368
rect 3384 14356 3390 14408
rect 3436 14405 3464 14436
rect 3786 14424 3792 14436
rect 3844 14424 3850 14476
rect 3881 14467 3939 14473
rect 3881 14433 3893 14467
rect 3927 14464 3939 14467
rect 3970 14464 3976 14476
rect 3927 14436 3976 14464
rect 3927 14433 3939 14436
rect 3881 14427 3939 14433
rect 3970 14424 3976 14436
rect 4028 14424 4034 14476
rect 5074 14464 5080 14476
rect 4080 14436 5080 14464
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 4080 14396 4108 14436
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5258 14464 5264 14476
rect 5219 14436 5264 14464
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 5828 14473 5856 14504
rect 6822 14492 6828 14504
rect 6880 14532 6886 14544
rect 6880 14504 7052 14532
rect 6880 14492 6886 14504
rect 6086 14473 6092 14476
rect 5813 14467 5871 14473
rect 5368 14436 5580 14464
rect 3421 14359 3479 14365
rect 3534 14368 4108 14396
rect 3534 14328 3562 14368
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4525 14399 4583 14405
rect 4525 14396 4537 14399
rect 4212 14368 4537 14396
rect 4212 14356 4218 14368
rect 4525 14365 4537 14368
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 4672 14368 4717 14396
rect 4672 14356 4678 14368
rect 2976 14300 3562 14328
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 4065 14331 4123 14337
rect 4065 14328 4077 14331
rect 3660 14300 4077 14328
rect 3660 14288 3666 14300
rect 4065 14297 4077 14300
rect 4111 14297 4123 14331
rect 4632 14328 4660 14356
rect 5368 14328 5396 14436
rect 5552 14408 5580 14436
rect 5813 14433 5825 14467
rect 5859 14433 5871 14467
rect 5813 14427 5871 14433
rect 6080 14427 6092 14473
rect 6144 14464 6150 14476
rect 7024 14464 7052 14504
rect 7098 14492 7104 14544
rect 7156 14532 7162 14544
rect 7208 14532 7236 14563
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 11698 14560 11704 14612
rect 11756 14600 11762 14612
rect 12066 14600 12072 14612
rect 11756 14572 12072 14600
rect 11756 14560 11762 14572
rect 12066 14560 12072 14572
rect 12124 14560 12130 14612
rect 13173 14603 13231 14609
rect 13173 14569 13185 14603
rect 13219 14569 13231 14603
rect 13173 14563 13231 14569
rect 13265 14603 13323 14609
rect 13265 14569 13277 14603
rect 13311 14600 13323 14603
rect 19518 14600 19524 14612
rect 13311 14572 16712 14600
rect 13311 14569 13323 14572
rect 13265 14563 13323 14569
rect 10594 14541 10600 14544
rect 7530 14535 7588 14541
rect 7530 14532 7542 14535
rect 7156 14504 7542 14532
rect 7156 14492 7162 14504
rect 7530 14501 7542 14504
rect 7576 14501 7588 14535
rect 7530 14495 7588 14501
rect 9125 14535 9183 14541
rect 9125 14501 9137 14535
rect 9171 14532 9183 14535
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 9171 14504 10057 14532
rect 9171 14501 9183 14504
rect 9125 14495 9183 14501
rect 10045 14501 10057 14504
rect 10091 14501 10103 14535
rect 10045 14495 10103 14501
rect 10577 14535 10600 14541
rect 10577 14501 10589 14535
rect 10652 14532 10658 14544
rect 13188 14532 13216 14563
rect 16574 14532 16580 14544
rect 10652 14504 13216 14532
rect 15396 14504 16580 14532
rect 10577 14495 10600 14501
rect 10594 14492 10600 14495
rect 10652 14492 10658 14504
rect 7285 14467 7343 14473
rect 7285 14464 7297 14467
rect 6144 14436 6180 14464
rect 7024 14436 7297 14464
rect 6086 14424 6092 14427
rect 6144 14424 6150 14436
rect 7285 14433 7297 14436
rect 7331 14433 7343 14467
rect 7285 14427 7343 14433
rect 7834 14424 7840 14476
rect 7892 14464 7898 14476
rect 8294 14464 8300 14476
rect 7892 14436 8300 14464
rect 7892 14424 7898 14436
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8386 14424 8392 14476
rect 8444 14464 8450 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 8444 14436 9689 14464
rect 8444 14424 8450 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 10321 14467 10379 14473
rect 10321 14433 10333 14467
rect 10367 14464 10379 14467
rect 10870 14464 10876 14476
rect 10367 14436 10876 14464
rect 10367 14433 10379 14436
rect 10321 14427 10379 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 12066 14473 12072 14476
rect 11793 14467 11851 14473
rect 11793 14464 11805 14467
rect 11756 14436 11805 14464
rect 11756 14424 11762 14436
rect 11793 14433 11805 14436
rect 11839 14433 11851 14467
rect 11793 14427 11851 14433
rect 12060 14427 12072 14473
rect 12124 14464 12130 14476
rect 13808 14467 13866 14473
rect 12124 14436 12160 14464
rect 12066 14424 12072 14427
rect 12124 14424 12130 14436
rect 13808 14433 13820 14467
rect 13854 14464 13866 14467
rect 14550 14464 14556 14476
rect 13854 14436 14556 14464
rect 13854 14433 13866 14436
rect 13808 14427 13866 14433
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 15396 14473 15424 14504
rect 16574 14492 16580 14504
rect 16632 14492 16638 14544
rect 16684 14532 16712 14572
rect 17236 14572 19524 14600
rect 17236 14532 17264 14572
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 19610 14560 19616 14612
rect 19668 14600 19674 14612
rect 20073 14603 20131 14609
rect 20073 14600 20085 14603
rect 19668 14572 20085 14600
rect 19668 14560 19674 14572
rect 20073 14569 20085 14572
rect 20119 14569 20131 14603
rect 20073 14563 20131 14569
rect 18138 14532 18144 14544
rect 16684 14504 17264 14532
rect 17328 14504 18144 14532
rect 15381 14467 15439 14473
rect 15381 14433 15393 14467
rect 15427 14433 15439 14467
rect 15381 14427 15439 14433
rect 15562 14424 15568 14476
rect 15620 14464 15626 14476
rect 15749 14467 15807 14473
rect 15749 14464 15761 14467
rect 15620 14436 15761 14464
rect 15620 14424 15626 14436
rect 15749 14433 15761 14436
rect 15795 14433 15807 14467
rect 15749 14427 15807 14433
rect 16016 14467 16074 14473
rect 16016 14433 16028 14467
rect 16062 14464 16074 14467
rect 17221 14467 17279 14473
rect 16062 14436 17172 14464
rect 16062 14433 16074 14436
rect 16016 14427 16074 14433
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 9401 14399 9459 14405
rect 5592 14368 5685 14396
rect 5592 14356 5598 14368
rect 9401 14365 9413 14399
rect 9447 14365 9459 14399
rect 13538 14396 13544 14408
rect 13499 14368 13544 14396
rect 9401 14359 9459 14365
rect 9306 14328 9312 14340
rect 4632 14300 5396 14328
rect 8220 14300 9312 14328
rect 4065 14291 4123 14297
rect 3697 14263 3755 14269
rect 3697 14229 3709 14263
rect 3743 14260 3755 14263
rect 3786 14260 3792 14272
rect 3743 14232 3792 14260
rect 3743 14229 3755 14232
rect 3697 14223 3755 14229
rect 3786 14220 3792 14232
rect 3844 14260 3850 14272
rect 8220 14260 8248 14300
rect 9306 14288 9312 14300
rect 9364 14288 9370 14340
rect 9416 14328 9444 14359
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 9416 14300 10364 14328
rect 8662 14260 8668 14272
rect 3844 14232 8248 14260
rect 8623 14232 8668 14260
rect 3844 14220 3850 14232
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 8757 14263 8815 14269
rect 8757 14229 8769 14263
rect 8803 14260 8815 14263
rect 9214 14260 9220 14272
rect 8803 14232 9220 14260
rect 8803 14229 8815 14232
rect 8757 14223 8815 14229
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 9858 14260 9864 14272
rect 9819 14232 9864 14260
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 10336 14260 10364 14300
rect 14642 14288 14648 14340
rect 14700 14328 14706 14340
rect 14921 14331 14979 14337
rect 14921 14328 14933 14331
rect 14700 14300 14933 14328
rect 14700 14288 14706 14300
rect 14921 14297 14933 14300
rect 14967 14328 14979 14331
rect 15194 14328 15200 14340
rect 14967 14300 15200 14328
rect 14967 14297 14979 14300
rect 14921 14291 14979 14297
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 17144 14328 17172 14436
rect 17221 14433 17233 14467
rect 17267 14464 17279 14467
rect 17328 14464 17356 14504
rect 18138 14492 18144 14504
rect 18196 14532 18202 14544
rect 18960 14535 19018 14541
rect 18196 14504 18736 14532
rect 18196 14492 18202 14504
rect 17494 14473 17500 14476
rect 17267 14436 17356 14464
rect 17267 14433 17279 14436
rect 17221 14427 17279 14433
rect 17488 14427 17500 14473
rect 17552 14464 17558 14476
rect 18708 14473 18736 14504
rect 18960 14501 18972 14535
rect 19006 14532 19018 14535
rect 19426 14532 19432 14544
rect 19006 14504 19432 14532
rect 19006 14501 19018 14504
rect 18960 14495 19018 14501
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 20162 14532 20168 14544
rect 20123 14504 20168 14532
rect 20162 14492 20168 14504
rect 20220 14492 20226 14544
rect 18693 14467 18751 14473
rect 17552 14436 17588 14464
rect 17494 14424 17500 14427
rect 17552 14424 17558 14436
rect 18693 14433 18705 14467
rect 18739 14433 18751 14467
rect 18693 14427 18751 14433
rect 20349 14467 20407 14473
rect 20349 14433 20361 14467
rect 20395 14464 20407 14467
rect 20438 14464 20444 14476
rect 20395 14436 20444 14464
rect 20395 14433 20407 14436
rect 20349 14427 20407 14433
rect 20438 14424 20444 14436
rect 20496 14424 20502 14476
rect 17144 14300 17264 14328
rect 17236 14272 17264 14300
rect 11701 14263 11759 14269
rect 11701 14260 11713 14263
rect 10336 14232 11713 14260
rect 11701 14229 11713 14232
rect 11747 14260 11759 14263
rect 11790 14260 11796 14272
rect 11747 14232 11796 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 11790 14220 11796 14232
rect 11848 14220 11854 14272
rect 15565 14263 15623 14269
rect 15565 14229 15577 14263
rect 15611 14260 15623 14263
rect 16022 14260 16028 14272
rect 15611 14232 16028 14260
rect 15611 14229 15623 14232
rect 15565 14223 15623 14229
rect 16022 14220 16028 14232
rect 16080 14220 16086 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 17129 14263 17187 14269
rect 17129 14260 17141 14263
rect 16540 14232 17141 14260
rect 16540 14220 16546 14232
rect 17129 14229 17141 14232
rect 17175 14229 17187 14263
rect 17129 14223 17187 14229
rect 17218 14220 17224 14272
rect 17276 14260 17282 14272
rect 18601 14263 18659 14269
rect 18601 14260 18613 14263
rect 17276 14232 18613 14260
rect 17276 14220 17282 14232
rect 18601 14229 18613 14232
rect 18647 14229 18659 14263
rect 20530 14260 20536 14272
rect 20491 14232 20536 14260
rect 18601 14223 18659 14229
rect 20530 14220 20536 14232
rect 20588 14220 20594 14272
rect 1104 14170 20884 14192
rect 1104 14118 4280 14170
rect 4332 14118 4344 14170
rect 4396 14118 4408 14170
rect 4460 14118 4472 14170
rect 4524 14118 10878 14170
rect 10930 14118 10942 14170
rect 10994 14118 11006 14170
rect 11058 14118 11070 14170
rect 11122 14118 17475 14170
rect 17527 14118 17539 14170
rect 17591 14118 17603 14170
rect 17655 14118 17667 14170
rect 17719 14118 20884 14170
rect 1104 14096 20884 14118
rect 3050 14056 3056 14068
rect 3011 14028 3056 14056
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 3329 14059 3387 14065
rect 3329 14025 3341 14059
rect 3375 14056 3387 14059
rect 3510 14056 3516 14068
rect 3375 14028 3516 14056
rect 3375 14025 3387 14028
rect 3329 14019 3387 14025
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 4982 14056 4988 14068
rect 4943 14028 4988 14056
rect 4982 14016 4988 14028
rect 5040 14016 5046 14068
rect 5258 14016 5264 14068
rect 5316 14056 5322 14068
rect 5813 14059 5871 14065
rect 5813 14056 5825 14059
rect 5316 14028 5825 14056
rect 5316 14016 5322 14028
rect 5813 14025 5825 14028
rect 5859 14025 5871 14059
rect 5813 14019 5871 14025
rect 7469 14059 7527 14065
rect 7469 14025 7481 14059
rect 7515 14056 7527 14059
rect 7834 14056 7840 14068
rect 7515 14028 7840 14056
rect 7515 14025 7527 14028
rect 7469 14019 7527 14025
rect 7834 14016 7840 14028
rect 7892 14016 7898 14068
rect 9858 14056 9864 14068
rect 8036 14028 9864 14056
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 1673 13923 1731 13929
rect 1673 13920 1685 13923
rect 1452 13892 1685 13920
rect 1452 13880 1458 13892
rect 1673 13889 1685 13892
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 2958 13880 2964 13932
rect 3016 13920 3022 13932
rect 3513 13923 3571 13929
rect 3513 13920 3525 13923
rect 3016 13892 3525 13920
rect 3016 13880 3022 13892
rect 3513 13889 3525 13892
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 4982 13880 4988 13932
rect 5040 13920 5046 13932
rect 5537 13923 5595 13929
rect 5537 13920 5549 13923
rect 5040 13892 5549 13920
rect 5040 13880 5046 13892
rect 5537 13889 5549 13892
rect 5583 13920 5595 13923
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 5583 13892 6377 13920
rect 5583 13889 5595 13892
rect 5537 13883 5595 13889
rect 6365 13889 6377 13892
rect 6411 13889 6423 13923
rect 7006 13920 7012 13932
rect 6365 13883 6423 13889
rect 6932 13892 7012 13920
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13821 3203 13855
rect 3145 13815 3203 13821
rect 3780 13855 3838 13861
rect 3780 13821 3792 13855
rect 3826 13852 3838 13855
rect 4154 13852 4160 13864
rect 3826 13824 4160 13852
rect 3826 13821 3838 13824
rect 3780 13815 3838 13821
rect 1940 13787 1998 13793
rect 1940 13753 1952 13787
rect 1986 13753 1998 13787
rect 3160 13784 3188 13815
rect 4154 13812 4160 13824
rect 4212 13852 4218 13864
rect 5445 13855 5503 13861
rect 5445 13852 5457 13855
rect 4212 13824 5457 13852
rect 4212 13812 4218 13824
rect 5445 13821 5457 13824
rect 5491 13821 5503 13855
rect 5445 13815 5503 13821
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6932 13861 6960 13892
rect 7006 13880 7012 13892
rect 7064 13880 7070 13932
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13920 7987 13923
rect 8036 13920 8064 14028
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10597 14059 10655 14065
rect 10597 14025 10609 14059
rect 10643 14056 10655 14059
rect 11606 14056 11612 14068
rect 10643 14028 11612 14056
rect 10643 14025 10655 14028
rect 10597 14019 10655 14025
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 12618 14016 12624 14068
rect 12676 14056 12682 14068
rect 12805 14059 12863 14065
rect 12805 14056 12817 14059
rect 12676 14028 12817 14056
rect 12676 14016 12682 14028
rect 12805 14025 12817 14028
rect 12851 14025 12863 14059
rect 12805 14019 12863 14025
rect 13446 14016 13452 14068
rect 13504 14056 13510 14068
rect 13906 14056 13912 14068
rect 13504 14028 13912 14056
rect 13504 14016 13510 14028
rect 13906 14016 13912 14028
rect 13964 14016 13970 14068
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 15013 14059 15071 14065
rect 15013 14056 15025 14059
rect 14424 14028 15025 14056
rect 14424 14016 14430 14028
rect 15013 14025 15025 14028
rect 15059 14025 15071 14059
rect 15013 14019 15071 14025
rect 15289 14059 15347 14065
rect 15289 14025 15301 14059
rect 15335 14056 15347 14059
rect 15335 14028 18736 14056
rect 15335 14025 15347 14028
rect 15289 14019 15347 14025
rect 16853 13991 16911 13997
rect 16853 13957 16865 13991
rect 16899 13988 16911 13991
rect 16899 13960 17356 13988
rect 16899 13957 16911 13960
rect 16853 13951 16911 13957
rect 17328 13932 17356 13960
rect 7975 13892 8064 13920
rect 8113 13923 8171 13929
rect 7975 13889 7987 13892
rect 7929 13883 7987 13889
rect 8113 13889 8125 13923
rect 8159 13920 8171 13923
rect 8662 13920 8668 13932
rect 8159 13892 8668 13920
rect 8159 13889 8171 13892
rect 8113 13883 8171 13889
rect 8662 13880 8668 13892
rect 8720 13880 8726 13932
rect 9214 13880 9220 13932
rect 9272 13920 9278 13932
rect 9493 13923 9551 13929
rect 9272 13892 9317 13920
rect 9272 13880 9278 13892
rect 9493 13889 9505 13923
rect 9539 13920 9551 13923
rect 10134 13920 10140 13932
rect 9539 13892 10140 13920
rect 9539 13889 9551 13892
rect 9493 13883 9551 13889
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 13173 13923 13231 13929
rect 13173 13920 13185 13923
rect 12452 13892 13185 13920
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 6144 13824 6193 13852
rect 6144 13812 6150 13824
rect 6181 13821 6193 13824
rect 6227 13821 6239 13855
rect 6181 13815 6239 13821
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13821 6975 13855
rect 7098 13852 7104 13864
rect 7059 13824 7104 13852
rect 6917 13815 6975 13821
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 7285 13855 7343 13861
rect 7285 13821 7297 13855
rect 7331 13852 7343 13855
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 7331 13824 8309 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 8757 13855 8815 13861
rect 8757 13821 8769 13855
rect 8803 13852 8815 13855
rect 10318 13852 10324 13864
rect 8803 13824 10324 13852
rect 8803 13821 8815 13824
rect 8757 13815 8815 13821
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10686 13852 10692 13864
rect 10647 13824 10692 13852
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 10962 13861 10968 13864
rect 10956 13852 10968 13861
rect 10923 13824 10968 13852
rect 10956 13815 10968 13824
rect 10962 13812 10968 13815
rect 11020 13812 11026 13864
rect 12342 13812 12348 13864
rect 12400 13852 12406 13864
rect 12452 13852 12480 13892
rect 13173 13889 13185 13892
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 13679 13923 13737 13929
rect 13679 13889 13691 13923
rect 13725 13920 13737 13923
rect 14826 13920 14832 13932
rect 13725 13892 14832 13920
rect 13725 13889 13737 13892
rect 13679 13883 13737 13889
rect 14826 13880 14832 13892
rect 14884 13880 14890 13932
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 15473 13923 15531 13929
rect 15473 13920 15485 13923
rect 15344 13892 15485 13920
rect 15344 13880 15350 13892
rect 15473 13889 15485 13892
rect 15519 13889 15531 13923
rect 15473 13883 15531 13889
rect 16666 13880 16672 13932
rect 16724 13920 16730 13932
rect 17034 13920 17040 13932
rect 16724 13892 17040 13920
rect 16724 13880 16730 13892
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 17310 13880 17316 13932
rect 17368 13920 17374 13932
rect 17405 13923 17463 13929
rect 17405 13920 17417 13923
rect 17368 13892 17417 13920
rect 17368 13880 17374 13892
rect 17405 13889 17417 13892
rect 17451 13889 17463 13923
rect 17405 13883 17463 13889
rect 17494 13880 17500 13932
rect 17552 13920 17558 13932
rect 17589 13923 17647 13929
rect 17589 13920 17601 13923
rect 17552 13892 17601 13920
rect 17552 13880 17558 13892
rect 17589 13889 17601 13892
rect 17635 13920 17647 13923
rect 18598 13920 18604 13932
rect 17635 13892 18604 13920
rect 17635 13889 17647 13892
rect 17589 13883 17647 13889
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 18708 13929 18736 14028
rect 18693 13923 18751 13929
rect 18693 13889 18705 13923
rect 18739 13889 18751 13923
rect 18874 13920 18880 13932
rect 18835 13892 18880 13920
rect 18693 13883 18751 13889
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 12400 13824 12480 13852
rect 12989 13855 13047 13861
rect 12400 13812 12406 13824
rect 12989 13821 13001 13855
rect 13035 13852 13047 13855
rect 13814 13852 13820 13864
rect 13035 13824 13820 13852
rect 13035 13821 13047 13824
rect 12989 13815 13047 13821
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 13906 13812 13912 13864
rect 13964 13852 13970 13864
rect 15105 13855 15163 13861
rect 13964 13824 14009 13852
rect 13964 13812 13970 13824
rect 15105 13821 15117 13855
rect 15151 13852 15163 13855
rect 15740 13855 15798 13861
rect 15151 13824 15700 13852
rect 15151 13821 15163 13824
rect 15105 13815 15163 13821
rect 3602 13784 3608 13796
rect 3160 13756 3608 13784
rect 1940 13747 1998 13753
rect 1955 13716 1983 13747
rect 3602 13744 3608 13756
rect 3660 13744 3666 13796
rect 7837 13787 7895 13793
rect 7837 13753 7849 13787
rect 7883 13784 7895 13787
rect 8662 13784 8668 13796
rect 7883 13756 8668 13784
rect 7883 13753 7895 13756
rect 7837 13747 7895 13753
rect 8662 13744 8668 13756
rect 8720 13744 8726 13796
rect 15672 13784 15700 13824
rect 15740 13821 15752 13855
rect 15786 13852 15798 13855
rect 17126 13852 17132 13864
rect 15786 13824 17132 13852
rect 15786 13821 15798 13824
rect 15740 13815 15798 13821
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 19058 13852 19064 13864
rect 19019 13824 19064 13852
rect 19058 13812 19064 13824
rect 19116 13812 19122 13864
rect 19328 13855 19386 13861
rect 19328 13821 19340 13855
rect 19374 13852 19386 13855
rect 20346 13852 20352 13864
rect 19374 13824 20352 13852
rect 19374 13821 19386 13824
rect 19328 13815 19386 13821
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 16114 13784 16120 13796
rect 11440 13756 12664 13784
rect 15672 13756 16120 13784
rect 3326 13716 3332 13728
rect 1955 13688 3332 13716
rect 3326 13676 3332 13688
rect 3384 13676 3390 13728
rect 4706 13676 4712 13728
rect 4764 13716 4770 13728
rect 4893 13719 4951 13725
rect 4893 13716 4905 13719
rect 4764 13688 4905 13716
rect 4764 13676 4770 13688
rect 4893 13685 4905 13688
rect 4939 13716 4951 13719
rect 5353 13719 5411 13725
rect 5353 13716 5365 13719
rect 4939 13688 5365 13716
rect 4939 13685 4951 13688
rect 4893 13679 4951 13685
rect 5353 13685 5365 13688
rect 5399 13685 5411 13719
rect 6270 13716 6276 13728
rect 6231 13688 6276 13716
rect 5353 13679 5411 13685
rect 6270 13676 6276 13688
rect 6328 13676 6334 13728
rect 8481 13719 8539 13725
rect 8481 13685 8493 13719
rect 8527 13716 8539 13719
rect 8754 13716 8760 13728
rect 8527 13688 8760 13716
rect 8527 13685 8539 13688
rect 8481 13679 8539 13685
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 9223 13719 9281 13725
rect 9223 13685 9235 13719
rect 9269 13716 9281 13719
rect 9582 13716 9588 13728
rect 9269 13688 9588 13716
rect 9269 13685 9281 13688
rect 9223 13679 9281 13685
rect 9582 13676 9588 13688
rect 9640 13716 9646 13728
rect 11440 13716 11468 13756
rect 12636 13728 12664 13756
rect 16114 13744 16120 13756
rect 16172 13744 16178 13796
rect 16298 13744 16304 13796
rect 16356 13784 16362 13796
rect 16356 13756 17080 13784
rect 16356 13744 16362 13756
rect 9640 13688 11468 13716
rect 9640 13676 9646 13688
rect 11514 13676 11520 13728
rect 11572 13716 11578 13728
rect 12069 13719 12127 13725
rect 12069 13716 12081 13719
rect 11572 13688 12081 13716
rect 11572 13676 11578 13688
rect 12069 13685 12081 13688
rect 12115 13685 12127 13719
rect 12069 13679 12127 13685
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12492 13688 12537 13716
rect 12492 13676 12498 13688
rect 12618 13676 12624 13728
rect 12676 13716 12682 13728
rect 13639 13719 13697 13725
rect 13639 13716 13651 13719
rect 12676 13688 13651 13716
rect 12676 13676 12682 13688
rect 13639 13685 13651 13688
rect 13685 13685 13697 13719
rect 16942 13716 16948 13728
rect 16903 13688 16948 13716
rect 13639 13679 13697 13685
rect 16942 13676 16948 13688
rect 17000 13676 17006 13728
rect 17052 13716 17080 13756
rect 17218 13744 17224 13796
rect 17276 13784 17282 13796
rect 17313 13787 17371 13793
rect 17313 13784 17325 13787
rect 17276 13756 17325 13784
rect 17276 13744 17282 13756
rect 17313 13753 17325 13756
rect 17359 13753 17371 13787
rect 18414 13784 18420 13796
rect 17313 13747 17371 13753
rect 17420 13756 18420 13784
rect 17420 13716 17448 13756
rect 18414 13744 18420 13756
rect 18472 13744 18478 13796
rect 18230 13716 18236 13728
rect 17052 13688 17448 13716
rect 18191 13688 18236 13716
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 18506 13676 18512 13728
rect 18564 13716 18570 13728
rect 18601 13719 18659 13725
rect 18601 13716 18613 13719
rect 18564 13688 18613 13716
rect 18564 13676 18570 13688
rect 18601 13685 18613 13688
rect 18647 13685 18659 13719
rect 20438 13716 20444 13728
rect 20399 13688 20444 13716
rect 18601 13679 18659 13685
rect 20438 13676 20444 13688
rect 20496 13676 20502 13728
rect 1104 13626 20884 13648
rect 1104 13574 7579 13626
rect 7631 13574 7643 13626
rect 7695 13574 7707 13626
rect 7759 13574 7771 13626
rect 7823 13574 14176 13626
rect 14228 13574 14240 13626
rect 14292 13574 14304 13626
rect 14356 13574 14368 13626
rect 14420 13574 20884 13626
rect 1104 13552 20884 13574
rect 3142 13472 3148 13524
rect 3200 13512 3206 13524
rect 3694 13512 3700 13524
rect 3200 13484 3700 13512
rect 3200 13472 3206 13484
rect 3694 13472 3700 13484
rect 3752 13472 3758 13524
rect 4614 13512 4620 13524
rect 4612 13472 4620 13512
rect 4672 13472 4678 13524
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 6457 13515 6515 13521
rect 6457 13512 6469 13515
rect 6144 13484 6469 13512
rect 6144 13472 6150 13484
rect 6457 13481 6469 13484
rect 6503 13481 6515 13515
rect 6457 13475 6515 13481
rect 8205 13515 8263 13521
rect 8205 13481 8217 13515
rect 8251 13512 8263 13515
rect 8386 13512 8392 13524
rect 8251 13484 8392 13512
rect 8251 13481 8263 13484
rect 8205 13475 8263 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8662 13472 8668 13524
rect 8720 13512 8726 13524
rect 9217 13515 9275 13521
rect 9217 13512 9229 13515
rect 8720 13484 9229 13512
rect 8720 13472 8726 13484
rect 9217 13481 9229 13484
rect 9263 13481 9275 13515
rect 9217 13475 9275 13481
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 10100 13484 11827 13512
rect 10100 13472 10106 13484
rect 2498 13404 2504 13456
rect 2556 13444 2562 13456
rect 4612 13444 4640 13472
rect 2556 13416 4640 13444
rect 4709 13447 4767 13453
rect 2556 13404 2562 13416
rect 4709 13413 4721 13447
rect 4755 13444 4767 13447
rect 4798 13444 4804 13456
rect 4755 13416 4804 13444
rect 4755 13413 4767 13416
rect 4709 13407 4767 13413
rect 4798 13404 4804 13416
rect 4856 13404 4862 13456
rect 5344 13447 5402 13453
rect 5344 13413 5356 13447
rect 5390 13444 5402 13447
rect 5810 13444 5816 13456
rect 5390 13416 5816 13444
rect 5390 13413 5402 13416
rect 5344 13407 5402 13413
rect 5810 13404 5816 13416
rect 5868 13444 5874 13456
rect 6270 13444 6276 13456
rect 5868 13416 6276 13444
rect 5868 13404 5874 13416
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 7745 13447 7803 13453
rect 7745 13444 7757 13447
rect 7064 13416 7757 13444
rect 7064 13404 7070 13416
rect 7745 13413 7757 13416
rect 7791 13413 7803 13447
rect 7745 13407 7803 13413
rect 7926 13404 7932 13456
rect 7984 13444 7990 13456
rect 8573 13447 8631 13453
rect 8573 13444 8585 13447
rect 7984 13416 8585 13444
rect 7984 13404 7990 13416
rect 8573 13413 8585 13416
rect 8619 13413 8631 13447
rect 10226 13444 10232 13456
rect 8573 13407 8631 13413
rect 8680 13416 10232 13444
rect 1664 13379 1722 13385
rect 1664 13345 1676 13379
rect 1710 13376 1722 13379
rect 2866 13376 2872 13388
rect 1710 13348 2872 13376
rect 1710 13345 1722 13348
rect 1664 13339 1722 13345
rect 2866 13336 2872 13348
rect 2924 13376 2930 13388
rect 3237 13379 3295 13385
rect 3237 13376 3249 13379
rect 2924 13348 3249 13376
rect 2924 13336 2930 13348
rect 3237 13345 3249 13348
rect 3283 13345 3295 13379
rect 3237 13339 3295 13345
rect 3881 13379 3939 13385
rect 3881 13345 3893 13379
rect 3927 13376 3939 13379
rect 3970 13376 3976 13388
rect 3927 13348 3976 13376
rect 3927 13345 3939 13348
rect 3881 13339 3939 13345
rect 3970 13336 3976 13348
rect 4028 13336 4034 13388
rect 4614 13376 4620 13388
rect 4172 13348 4476 13376
rect 4575 13348 4620 13376
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 3326 13308 3332 13320
rect 3287 13280 3332 13308
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3510 13308 3516 13320
rect 3471 13280 3516 13308
rect 3510 13268 3516 13280
rect 3568 13308 3574 13320
rect 4172 13308 4200 13348
rect 3568 13280 4200 13308
rect 3568 13268 3574 13280
rect 4246 13268 4252 13320
rect 4304 13268 4310 13320
rect 4448 13308 4476 13348
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 4890 13336 4896 13388
rect 4948 13376 4954 13388
rect 6914 13376 6920 13388
rect 4948 13348 6132 13376
rect 6875 13348 6920 13376
rect 4948 13336 4954 13348
rect 4801 13311 4859 13317
rect 4801 13308 4813 13311
rect 4448 13280 4813 13308
rect 4801 13277 4813 13280
rect 4847 13308 4859 13311
rect 4982 13308 4988 13320
rect 4847 13280 4988 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 6104 13308 6132 13348
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 8680 13376 8708 13416
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 11514 13453 11520 13456
rect 11508 13444 11520 13453
rect 11475 13416 11520 13444
rect 11508 13407 11520 13416
rect 11514 13404 11520 13407
rect 11572 13404 11578 13456
rect 11698 13404 11704 13456
rect 11756 13404 11762 13456
rect 11799 13444 11827 13484
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 12621 13515 12679 13521
rect 12621 13512 12633 13515
rect 12124 13484 12633 13512
rect 12124 13472 12130 13484
rect 12621 13481 12633 13484
rect 12667 13481 12679 13515
rect 12621 13475 12679 13481
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14921 13515 14979 13521
rect 14921 13512 14933 13515
rect 13872 13484 14933 13512
rect 13872 13472 13878 13484
rect 14921 13481 14933 13484
rect 14967 13481 14979 13515
rect 14921 13475 14979 13481
rect 16025 13515 16083 13521
rect 16025 13481 16037 13515
rect 16071 13512 16083 13515
rect 16761 13515 16819 13521
rect 16761 13512 16773 13515
rect 16071 13484 16773 13512
rect 16071 13481 16083 13484
rect 16025 13475 16083 13481
rect 16761 13481 16773 13484
rect 16807 13481 16819 13515
rect 16761 13475 16819 13481
rect 14936 13444 14964 13475
rect 16942 13472 16948 13524
rect 17000 13512 17006 13524
rect 18049 13515 18107 13521
rect 18049 13512 18061 13515
rect 17000 13484 18061 13512
rect 17000 13472 17006 13484
rect 18049 13481 18061 13484
rect 18095 13481 18107 13515
rect 18049 13475 18107 13481
rect 17126 13444 17132 13456
rect 11799 13416 12756 13444
rect 8036 13348 8708 13376
rect 9033 13379 9091 13385
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 5132 13280 5177 13308
rect 6104 13280 7021 13308
rect 5132 13268 5138 13280
rect 7009 13277 7021 13280
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13308 7251 13311
rect 7282 13308 7288 13320
rect 7239 13280 7288 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 8036 13317 8064 13348
rect 9033 13345 9045 13379
rect 9079 13345 9091 13379
rect 9033 13339 9091 13345
rect 7837 13311 7895 13317
rect 7837 13308 7849 13311
rect 7432 13280 7849 13308
rect 7432 13268 7438 13280
rect 7837 13277 7849 13280
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13277 8723 13311
rect 8665 13271 8723 13277
rect 2869 13243 2927 13249
rect 2869 13209 2881 13243
rect 2915 13240 2927 13243
rect 4264 13240 4292 13268
rect 2915 13212 4292 13240
rect 6549 13243 6607 13249
rect 2915 13209 2927 13212
rect 2869 13203 2927 13209
rect 6549 13209 6561 13243
rect 6595 13240 6607 13243
rect 8680 13240 8708 13271
rect 8754 13268 8760 13320
rect 8812 13308 8818 13320
rect 8812 13280 8857 13308
rect 8812 13268 8818 13280
rect 9048 13240 9076 13339
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 9933 13379 9991 13385
rect 9933 13376 9945 13379
rect 9824 13348 9945 13376
rect 9824 13336 9830 13348
rect 9933 13345 9945 13348
rect 9979 13345 9991 13379
rect 9933 13339 9991 13345
rect 10686 13336 10692 13388
rect 10744 13376 10750 13388
rect 11241 13379 11299 13385
rect 11241 13376 11253 13379
rect 10744 13348 11253 13376
rect 10744 13336 10750 13348
rect 11241 13345 11253 13348
rect 11287 13376 11299 13379
rect 11716 13376 11744 13404
rect 12728 13385 12756 13416
rect 13096 13416 14872 13444
rect 14936 13416 16712 13444
rect 17087 13416 17132 13444
rect 13096 13385 13124 13416
rect 11287 13348 11744 13376
rect 12713 13379 12771 13385
rect 11287 13345 11299 13348
rect 11241 13339 11299 13345
rect 12713 13345 12725 13379
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 13081 13379 13139 13385
rect 13081 13345 13093 13379
rect 13127 13345 13139 13379
rect 13081 13339 13139 13345
rect 13449 13379 13507 13385
rect 13449 13345 13461 13379
rect 13495 13376 13507 13379
rect 13538 13376 13544 13388
rect 13495 13348 13544 13376
rect 13495 13345 13507 13348
rect 13449 13339 13507 13345
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 13716 13379 13774 13385
rect 13716 13345 13728 13379
rect 13762 13376 13774 13379
rect 14642 13376 14648 13388
rect 13762 13348 14648 13376
rect 13762 13345 13774 13348
rect 13716 13339 13774 13345
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9640 13280 9689 13308
rect 9640 13268 9646 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 14844 13308 14872 13416
rect 15010 13336 15016 13388
rect 15068 13376 15074 13388
rect 15105 13379 15163 13385
rect 15105 13376 15117 13379
rect 15068 13348 15117 13376
rect 15068 13336 15074 13348
rect 15105 13345 15117 13348
rect 15151 13345 15163 13379
rect 15105 13339 15163 13345
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 16574 13376 16580 13388
rect 15335 13348 16580 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 16574 13336 16580 13348
rect 16632 13336 16638 13388
rect 16684 13385 16712 13416
rect 17126 13404 17132 13416
rect 17184 13404 17190 13456
rect 19150 13404 19156 13456
rect 19208 13444 19214 13456
rect 19208 13416 19748 13444
rect 19208 13404 19214 13416
rect 16669 13379 16727 13385
rect 16669 13345 16681 13379
rect 16715 13345 16727 13379
rect 16669 13339 16727 13345
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 16908 13348 17969 13376
rect 16908 13336 16914 13348
rect 17957 13345 17969 13348
rect 18003 13345 18015 13379
rect 18414 13376 18420 13388
rect 17957 13339 18015 13345
rect 18248 13348 18420 13376
rect 15562 13308 15568 13320
rect 14844 13280 15568 13308
rect 9677 13271 9735 13277
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13277 16175 13311
rect 16298 13308 16304 13320
rect 16259 13280 16304 13308
rect 16117 13271 16175 13277
rect 6595 13212 9076 13240
rect 6595 13209 6607 13212
rect 6549 13203 6607 13209
rect 10962 13200 10968 13252
rect 11020 13200 11026 13252
rect 14734 13200 14740 13252
rect 14792 13240 14798 13252
rect 14829 13243 14887 13249
rect 14829 13240 14841 13243
rect 14792 13212 14841 13240
rect 14792 13200 14798 13212
rect 14829 13209 14841 13212
rect 14875 13209 14887 13243
rect 14829 13203 14887 13209
rect 15473 13243 15531 13249
rect 15473 13209 15485 13243
rect 15519 13240 15531 13243
rect 15930 13240 15936 13252
rect 15519 13212 15936 13240
rect 15519 13209 15531 13212
rect 15473 13203 15531 13209
rect 15930 13200 15936 13212
rect 15988 13200 15994 13252
rect 16132 13240 16160 13271
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 16482 13268 16488 13320
rect 16540 13308 16546 13320
rect 16540 13280 16896 13308
rect 16540 13268 16546 13280
rect 16758 13240 16764 13252
rect 16132 13212 16764 13240
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 16868 13240 16896 13280
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 17000 13280 17233 13308
rect 17000 13268 17006 13280
rect 17221 13277 17233 13280
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 17405 13311 17463 13317
rect 17405 13308 17417 13311
rect 17368 13280 17417 13308
rect 17368 13268 17374 13280
rect 17405 13277 17417 13280
rect 17451 13308 17463 13311
rect 17494 13308 17500 13320
rect 17451 13280 17500 13308
rect 17451 13277 17463 13280
rect 17405 13271 17463 13277
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 18248 13317 18276 13348
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 18598 13336 18604 13388
rect 18656 13376 18662 13388
rect 18785 13379 18843 13385
rect 18785 13376 18797 13379
rect 18656 13348 18797 13376
rect 18656 13336 18662 13348
rect 18785 13345 18797 13348
rect 18831 13345 18843 13379
rect 18785 13339 18843 13345
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 19613 13379 19671 13385
rect 19613 13376 19625 13379
rect 19392 13348 19625 13376
rect 19392 13336 19398 13348
rect 19613 13345 19625 13348
rect 19659 13345 19671 13379
rect 19720 13376 19748 13416
rect 20073 13379 20131 13385
rect 19720 13348 19840 13376
rect 19613 13339 19671 13345
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 18322 13268 18328 13320
rect 18380 13308 18386 13320
rect 18877 13311 18935 13317
rect 18877 13308 18889 13311
rect 18380 13280 18889 13308
rect 18380 13268 18386 13280
rect 18877 13277 18889 13280
rect 18923 13277 18935 13311
rect 18877 13271 18935 13277
rect 18966 13268 18972 13320
rect 19024 13308 19030 13320
rect 19702 13308 19708 13320
rect 19024 13280 19069 13308
rect 19663 13280 19708 13308
rect 19024 13268 19030 13280
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 19812 13317 19840 13348
rect 20073 13345 20085 13379
rect 20119 13376 20131 13379
rect 20530 13376 20536 13388
rect 20119 13348 20536 13376
rect 20119 13345 20131 13348
rect 20073 13339 20131 13345
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 17589 13243 17647 13249
rect 17589 13240 17601 13243
rect 16868 13212 17601 13240
rect 17589 13209 17601 13212
rect 17635 13209 17647 13243
rect 17589 13203 17647 13209
rect 18782 13200 18788 13252
rect 18840 13240 18846 13252
rect 20257 13243 20315 13249
rect 20257 13240 20269 13243
rect 18840 13212 20269 13240
rect 18840 13200 18846 13212
rect 20257 13209 20269 13212
rect 20303 13209 20315 13243
rect 20257 13203 20315 13209
rect 2777 13175 2835 13181
rect 2777 13141 2789 13175
rect 2823 13172 2835 13175
rect 3418 13172 3424 13184
rect 2823 13144 3424 13172
rect 2823 13141 2835 13144
rect 2777 13135 2835 13141
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 4249 13175 4307 13181
rect 4249 13141 4261 13175
rect 4295 13172 4307 13175
rect 6362 13172 6368 13184
rect 4295 13144 6368 13172
rect 4295 13141 4307 13144
rect 4249 13135 4307 13141
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 7377 13175 7435 13181
rect 7377 13141 7389 13175
rect 7423 13172 7435 13175
rect 9950 13172 9956 13184
rect 7423 13144 9956 13172
rect 7423 13141 7435 13144
rect 7377 13135 7435 13141
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10980 13172 11008 13200
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10100 13144 11069 13172
rect 10100 13132 10106 13144
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 12526 13132 12532 13184
rect 12584 13172 12590 13184
rect 12897 13175 12955 13181
rect 12897 13172 12909 13175
rect 12584 13144 12909 13172
rect 12584 13132 12590 13144
rect 12897 13141 12909 13144
rect 12943 13141 12955 13175
rect 12897 13135 12955 13141
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 13265 13175 13323 13181
rect 13265 13172 13277 13175
rect 13044 13144 13277 13172
rect 13044 13132 13050 13144
rect 13265 13141 13277 13144
rect 13311 13141 13323 13175
rect 15654 13172 15660 13184
rect 15615 13144 15660 13172
rect 13265 13135 13323 13141
rect 15654 13132 15660 13144
rect 15712 13132 15718 13184
rect 16482 13132 16488 13184
rect 16540 13172 16546 13184
rect 18414 13172 18420 13184
rect 16540 13144 16585 13172
rect 18375 13144 18420 13172
rect 16540 13132 16546 13144
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 19245 13175 19303 13181
rect 19245 13141 19257 13175
rect 19291 13172 19303 13175
rect 20070 13172 20076 13184
rect 19291 13144 20076 13172
rect 19291 13141 19303 13144
rect 19245 13135 19303 13141
rect 20070 13132 20076 13144
rect 20128 13132 20134 13184
rect 1104 13082 20884 13104
rect 1104 13030 4280 13082
rect 4332 13030 4344 13082
rect 4396 13030 4408 13082
rect 4460 13030 4472 13082
rect 4524 13030 10878 13082
rect 10930 13030 10942 13082
rect 10994 13030 11006 13082
rect 11058 13030 11070 13082
rect 11122 13030 17475 13082
rect 17527 13030 17539 13082
rect 17591 13030 17603 13082
rect 17655 13030 17667 13082
rect 17719 13030 20884 13082
rect 1104 13008 20884 13030
rect 2866 12968 2872 12980
rect 2827 12940 2872 12968
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 4341 12971 4399 12977
rect 4341 12968 4353 12971
rect 4212 12940 4353 12968
rect 4212 12928 4218 12940
rect 4341 12937 4353 12940
rect 4387 12937 4399 12971
rect 5074 12968 5080 12980
rect 4341 12931 4399 12937
rect 4448 12940 5080 12968
rect 4062 12860 4068 12912
rect 4120 12900 4126 12912
rect 4448 12900 4476 12940
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5810 12968 5816 12980
rect 5771 12940 5816 12968
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 5902 12928 5908 12980
rect 5960 12968 5966 12980
rect 5960 12940 6005 12968
rect 5960 12928 5966 12940
rect 6270 12928 6276 12980
rect 6328 12968 6334 12980
rect 6822 12968 6828 12980
rect 6328 12940 6828 12968
rect 6328 12928 6334 12940
rect 6822 12928 6828 12940
rect 6880 12968 6886 12980
rect 8110 12968 8116 12980
rect 6880 12940 8116 12968
rect 6880 12928 6886 12940
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 10318 12928 10324 12980
rect 10376 12968 10382 12980
rect 10594 12968 10600 12980
rect 10376 12940 10600 12968
rect 10376 12928 10382 12940
rect 10594 12928 10600 12940
rect 10652 12968 10658 12980
rect 10781 12971 10839 12977
rect 10781 12968 10793 12971
rect 10652 12940 10793 12968
rect 10652 12928 10658 12940
rect 10781 12937 10793 12940
rect 10827 12937 10839 12971
rect 10781 12931 10839 12937
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11882 12968 11888 12980
rect 11296 12940 11888 12968
rect 11296 12928 11302 12940
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 13538 12968 13544 12980
rect 12912 12940 13544 12968
rect 4120 12872 4476 12900
rect 4120 12860 4126 12872
rect 4448 12841 4476 12872
rect 5534 12860 5540 12912
rect 5592 12900 5598 12912
rect 9953 12903 10011 12909
rect 5592 12872 6500 12900
rect 5592 12860 5598 12872
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12801 4491 12835
rect 6362 12832 6368 12844
rect 4433 12795 4491 12801
rect 5460 12804 5948 12832
rect 6323 12804 6368 12832
rect 1394 12724 1400 12776
rect 1452 12764 1458 12776
rect 1489 12767 1547 12773
rect 1489 12764 1501 12767
rect 1452 12736 1501 12764
rect 1452 12724 1458 12736
rect 1489 12733 1501 12736
rect 1535 12764 1547 12767
rect 2958 12764 2964 12776
rect 1535 12736 2964 12764
rect 1535 12733 1547 12736
rect 1489 12727 1547 12733
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 3234 12773 3240 12776
rect 3228 12764 3240 12773
rect 3195 12736 3240 12764
rect 3228 12727 3240 12736
rect 3234 12724 3240 12727
rect 3292 12724 3298 12776
rect 4706 12773 4712 12776
rect 4700 12727 4712 12773
rect 4764 12764 4770 12776
rect 4764 12736 4800 12764
rect 4706 12724 4712 12727
rect 4764 12724 4770 12736
rect 1756 12699 1814 12705
rect 1756 12665 1768 12699
rect 1802 12696 1814 12699
rect 2774 12696 2780 12708
rect 1802 12668 2780 12696
rect 1802 12665 1814 12668
rect 1756 12659 1814 12665
rect 2774 12656 2780 12668
rect 2832 12696 2838 12708
rect 3326 12696 3332 12708
rect 2832 12668 3332 12696
rect 2832 12656 2838 12668
rect 3326 12656 3332 12668
rect 3384 12656 3390 12708
rect 4154 12656 4160 12708
rect 4212 12696 4218 12708
rect 5460 12696 5488 12804
rect 4212 12668 5488 12696
rect 5920 12696 5948 12804
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 6472 12841 6500 12872
rect 9953 12869 9965 12903
rect 9999 12900 10011 12903
rect 9999 12872 11744 12900
rect 9999 12869 10011 12872
rect 9953 12863 10011 12869
rect 6457 12835 6515 12841
rect 6457 12801 6469 12835
rect 6503 12801 6515 12835
rect 6822 12832 6828 12844
rect 6783 12804 6828 12832
rect 6457 12795 6515 12801
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 10502 12832 10508 12844
rect 8352 12804 8397 12832
rect 10463 12804 10508 12832
rect 8352 12792 8358 12804
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 10612 12804 11652 12832
rect 7092 12767 7150 12773
rect 7092 12733 7104 12767
rect 7138 12764 7150 12767
rect 7466 12764 7472 12776
rect 7138 12736 7472 12764
rect 7138 12733 7150 12736
rect 7092 12727 7150 12733
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 10612 12764 10640 12804
rect 10962 12764 10968 12776
rect 8303 12736 10640 12764
rect 10923 12736 10968 12764
rect 6273 12699 6331 12705
rect 6273 12696 6285 12699
rect 5920 12668 6285 12696
rect 4212 12656 4218 12668
rect 6273 12665 6285 12668
rect 6319 12665 6331 12699
rect 8303 12696 8331 12736
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 6273 12659 6331 12665
rect 7208 12668 8331 12696
rect 8564 12699 8622 12705
rect 1854 12588 1860 12640
rect 1912 12628 1918 12640
rect 7208 12628 7236 12668
rect 8564 12665 8576 12699
rect 8610 12696 8622 12699
rect 9030 12696 9036 12708
rect 8610 12668 9036 12696
rect 8610 12665 8622 12668
rect 8564 12659 8622 12665
rect 9030 12656 9036 12668
rect 9088 12656 9094 12708
rect 9950 12656 9956 12708
rect 10008 12696 10014 12708
rect 10413 12699 10471 12705
rect 10413 12696 10425 12699
rect 10008 12668 10425 12696
rect 10008 12656 10014 12668
rect 10413 12665 10425 12668
rect 10459 12696 10471 12699
rect 11054 12696 11060 12708
rect 10459 12668 10963 12696
rect 11015 12668 11060 12696
rect 10459 12665 10471 12668
rect 10413 12659 10471 12665
rect 1912 12600 7236 12628
rect 1912 12588 1918 12600
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 7340 12600 8217 12628
rect 7340 12588 7346 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8205 12591 8263 12597
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 9582 12628 9588 12640
rect 8352 12600 9588 12628
rect 8352 12588 8358 12600
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 9677 12631 9735 12637
rect 9677 12597 9689 12631
rect 9723 12628 9735 12631
rect 9766 12628 9772 12640
rect 9723 12600 9772 12628
rect 9723 12597 9735 12600
rect 9677 12591 9735 12597
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 10318 12628 10324 12640
rect 10279 12600 10324 12628
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 10935 12628 10963 12668
rect 11054 12656 11060 12668
rect 11112 12656 11118 12708
rect 11238 12696 11244 12708
rect 11199 12668 11244 12696
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 11330 12656 11336 12708
rect 11388 12696 11394 12708
rect 11388 12668 11560 12696
rect 11388 12656 11394 12668
rect 11146 12628 11152 12640
rect 10935 12600 11152 12628
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 11422 12628 11428 12640
rect 11383 12600 11428 12628
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 11532 12637 11560 12668
rect 11517 12631 11575 12637
rect 11517 12597 11529 12631
rect 11563 12597 11575 12631
rect 11624 12628 11652 12804
rect 11716 12696 11744 12872
rect 12066 12832 12072 12844
rect 12027 12804 12072 12832
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 12912 12841 12940 12940
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 14461 12971 14519 12977
rect 14461 12937 14473 12971
rect 14507 12968 14519 12971
rect 16758 12968 16764 12980
rect 14507 12940 16620 12968
rect 16719 12940 16764 12968
rect 14507 12937 14519 12940
rect 14461 12931 14519 12937
rect 14277 12903 14335 12909
rect 14277 12869 14289 12903
rect 14323 12900 14335 12903
rect 14918 12900 14924 12912
rect 14323 12872 14924 12900
rect 14323 12869 14335 12872
rect 14277 12863 14335 12869
rect 14918 12860 14924 12872
rect 14976 12860 14982 12912
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12832 15163 12835
rect 16592 12832 16620 12940
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17773 12971 17831 12977
rect 17092 12940 17540 12968
rect 17092 12928 17098 12940
rect 16669 12903 16727 12909
rect 16669 12869 16681 12903
rect 16715 12900 16727 12903
rect 17126 12900 17132 12912
rect 16715 12872 17132 12900
rect 16715 12869 16727 12872
rect 16669 12863 16727 12869
rect 17126 12860 17132 12872
rect 17184 12860 17190 12912
rect 17034 12832 17040 12844
rect 15151 12804 15424 12832
rect 16592 12804 17040 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 11885 12767 11943 12773
rect 11885 12733 11897 12767
rect 11931 12764 11943 12767
rect 12434 12764 12440 12776
rect 11931 12736 12440 12764
rect 11931 12733 11943 12736
rect 11885 12727 11943 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 13998 12764 14004 12776
rect 13096 12736 14004 12764
rect 13096 12696 13124 12736
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 15286 12764 15292 12776
rect 15247 12736 15292 12764
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 15396 12764 15424 12804
rect 17034 12792 17040 12804
rect 17092 12792 17098 12844
rect 17310 12832 17316 12844
rect 17271 12804 17316 12832
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 16298 12764 16304 12776
rect 15396 12736 16304 12764
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 16632 12736 17448 12764
rect 16632 12724 16638 12736
rect 11716 12668 13124 12696
rect 13164 12699 13222 12705
rect 13164 12665 13176 12699
rect 13210 12696 13222 12699
rect 14734 12696 14740 12708
rect 13210 12668 14740 12696
rect 13210 12665 13222 12668
rect 13164 12659 13222 12665
rect 14734 12656 14740 12668
rect 14792 12656 14798 12708
rect 14829 12699 14887 12705
rect 14829 12665 14841 12699
rect 14875 12696 14887 12699
rect 15194 12696 15200 12708
rect 14875 12668 15200 12696
rect 14875 12665 14887 12668
rect 14829 12659 14887 12665
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 15556 12699 15614 12705
rect 15556 12665 15568 12699
rect 15602 12696 15614 12699
rect 16942 12696 16948 12708
rect 15602 12668 16948 12696
rect 15602 12665 15614 12668
rect 15556 12659 15614 12665
rect 16942 12656 16948 12668
rect 17000 12656 17006 12708
rect 11977 12631 12035 12637
rect 11977 12628 11989 12631
rect 11624 12600 11989 12628
rect 11517 12591 11575 12597
rect 11977 12597 11989 12600
rect 12023 12597 12035 12631
rect 11977 12591 12035 12597
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12628 12495 12631
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12483 12600 12817 12628
rect 12483 12597 12495 12600
rect 12437 12591 12495 12597
rect 12805 12597 12817 12600
rect 12851 12628 12863 12631
rect 13078 12628 13084 12640
rect 12851 12600 13084 12628
rect 12851 12597 12863 12600
rect 12805 12591 12863 12597
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 14921 12631 14979 12637
rect 14921 12597 14933 12631
rect 14967 12628 14979 12631
rect 16298 12628 16304 12640
rect 14967 12600 16304 12628
rect 14967 12597 14979 12600
rect 14921 12591 14979 12597
rect 16298 12588 16304 12600
rect 16356 12588 16362 12640
rect 16758 12588 16764 12640
rect 16816 12628 16822 12640
rect 17129 12631 17187 12637
rect 17129 12628 17141 12631
rect 16816 12600 17141 12628
rect 16816 12588 16822 12600
rect 17129 12597 17141 12600
rect 17175 12597 17187 12631
rect 17129 12591 17187 12597
rect 17218 12588 17224 12640
rect 17276 12628 17282 12640
rect 17420 12628 17448 12736
rect 17512 12696 17540 12940
rect 17773 12937 17785 12971
rect 17819 12968 17831 12971
rect 18506 12968 18512 12980
rect 17819 12940 18512 12968
rect 17819 12937 17831 12940
rect 17773 12931 17831 12937
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 18782 12832 18788 12844
rect 18743 12804 18788 12832
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 19058 12832 19064 12844
rect 18932 12804 19064 12832
rect 18932 12792 18938 12804
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 17589 12767 17647 12773
rect 17589 12733 17601 12767
rect 17635 12764 17647 12767
rect 17770 12764 17776 12776
rect 17635 12736 17776 12764
rect 17635 12733 17647 12736
rect 17589 12727 17647 12733
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 18230 12724 18236 12776
rect 18288 12764 18294 12776
rect 18509 12767 18567 12773
rect 18509 12764 18521 12767
rect 18288 12736 18521 12764
rect 18288 12724 18294 12736
rect 18509 12733 18521 12736
rect 18555 12733 18567 12767
rect 18509 12727 18567 12733
rect 19328 12767 19386 12773
rect 19328 12733 19340 12767
rect 19374 12764 19386 12767
rect 20438 12764 20444 12776
rect 19374 12736 20444 12764
rect 19374 12733 19386 12736
rect 19328 12727 19386 12733
rect 20438 12724 20444 12736
rect 20496 12724 20502 12776
rect 19058 12696 19064 12708
rect 17512 12668 19064 12696
rect 19058 12656 19064 12668
rect 19116 12656 19122 12708
rect 17494 12628 17500 12640
rect 17276 12600 17321 12628
rect 17420 12600 17500 12628
rect 17276 12588 17282 12600
rect 17494 12588 17500 12600
rect 17552 12588 17558 12640
rect 18138 12628 18144 12640
rect 18099 12600 18144 12628
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 18506 12588 18512 12640
rect 18564 12628 18570 12640
rect 18601 12631 18659 12637
rect 18601 12628 18613 12631
rect 18564 12600 18613 12628
rect 18564 12588 18570 12600
rect 18601 12597 18613 12600
rect 18647 12597 18659 12631
rect 18601 12591 18659 12597
rect 19150 12588 19156 12640
rect 19208 12628 19214 12640
rect 20441 12631 20499 12637
rect 20441 12628 20453 12631
rect 19208 12600 20453 12628
rect 19208 12588 19214 12600
rect 20441 12597 20453 12600
rect 20487 12597 20499 12631
rect 20441 12591 20499 12597
rect 1104 12538 20884 12560
rect 1104 12486 7579 12538
rect 7631 12486 7643 12538
rect 7695 12486 7707 12538
rect 7759 12486 7771 12538
rect 7823 12486 14176 12538
rect 14228 12486 14240 12538
rect 14292 12486 14304 12538
rect 14356 12486 14368 12538
rect 14420 12486 20884 12538
rect 1104 12464 20884 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3145 12427 3203 12433
rect 2832 12396 2877 12424
rect 2832 12384 2838 12396
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 4154 12424 4160 12436
rect 3191 12396 4160 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 5537 12427 5595 12433
rect 5537 12393 5549 12427
rect 5583 12393 5595 12427
rect 5537 12387 5595 12393
rect 5813 12427 5871 12433
rect 5813 12393 5825 12427
rect 5859 12424 5871 12427
rect 6914 12424 6920 12436
rect 5859 12396 6920 12424
rect 5859 12393 5871 12396
rect 5813 12387 5871 12393
rect 1664 12359 1722 12365
rect 1664 12325 1676 12359
rect 1710 12356 1722 12359
rect 3513 12359 3571 12365
rect 3513 12356 3525 12359
rect 1710 12328 3525 12356
rect 1710 12325 1722 12328
rect 1664 12319 1722 12325
rect 3513 12325 3525 12328
rect 3559 12356 3571 12359
rect 5552 12356 5580 12387
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 7653 12427 7711 12433
rect 7653 12424 7665 12427
rect 7156 12396 7665 12424
rect 7156 12384 7162 12396
rect 7653 12393 7665 12396
rect 7699 12393 7711 12427
rect 8294 12424 8300 12436
rect 7653 12387 7711 12393
rect 8036 12396 8300 12424
rect 3559 12328 5580 12356
rect 6540 12359 6598 12365
rect 3559 12325 3571 12328
rect 3513 12319 3571 12325
rect 6540 12325 6552 12359
rect 6586 12356 6598 12359
rect 7282 12356 7288 12368
rect 6586 12328 7288 12356
rect 6586 12325 6598 12328
rect 6540 12319 6598 12325
rect 7282 12316 7288 12328
rect 7340 12316 7346 12368
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 3053 12291 3111 12297
rect 3053 12257 3065 12291
rect 3099 12288 3111 12291
rect 3142 12288 3148 12300
rect 3099 12260 3148 12288
rect 3099 12257 3111 12260
rect 3053 12251 3111 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 3605 12291 3663 12297
rect 3605 12257 3617 12291
rect 3651 12288 3663 12291
rect 4424 12291 4482 12297
rect 4424 12288 4436 12291
rect 3651 12260 4436 12288
rect 3651 12257 3663 12260
rect 3605 12251 3663 12257
rect 4424 12257 4436 12260
rect 4470 12288 4482 12291
rect 5350 12288 5356 12300
rect 4470 12260 5356 12288
rect 4470 12257 4482 12260
rect 4424 12251 4482 12257
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 5629 12291 5687 12297
rect 5629 12257 5641 12291
rect 5675 12288 5687 12291
rect 5902 12288 5908 12300
rect 5675 12260 5908 12288
rect 5675 12257 5687 12260
rect 5629 12251 5687 12257
rect 5902 12248 5908 12260
rect 5960 12248 5966 12300
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 6362 12288 6368 12300
rect 6227 12260 6368 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 6362 12248 6368 12260
rect 6420 12288 6426 12300
rect 8036 12297 8064 12396
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 9030 12384 9036 12436
rect 9088 12424 9094 12436
rect 9401 12427 9459 12433
rect 9401 12424 9413 12427
rect 9088 12396 9413 12424
rect 9088 12384 9094 12396
rect 9401 12393 9413 12396
rect 9447 12393 9459 12427
rect 9401 12387 9459 12393
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 10318 12424 10324 12436
rect 9723 12396 10324 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 10318 12384 10324 12396
rect 10376 12424 10382 12436
rect 13262 12424 13268 12436
rect 10376 12396 13268 12424
rect 10376 12384 10382 12396
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 13780 12396 14381 12424
rect 13780 12384 13786 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 15013 12427 15071 12433
rect 15013 12393 15025 12427
rect 15059 12424 15071 12427
rect 18598 12424 18604 12436
rect 15059 12396 17172 12424
rect 15059 12393 15071 12396
rect 15013 12387 15071 12393
rect 10134 12316 10140 12368
rect 10192 12356 10198 12368
rect 10192 12328 10732 12356
rect 10192 12316 10198 12328
rect 7929 12291 7987 12297
rect 6420 12260 7328 12288
rect 6420 12248 6426 12260
rect 3510 12180 3516 12232
rect 3568 12220 3574 12232
rect 3697 12223 3755 12229
rect 3697 12220 3709 12223
rect 3568 12192 3709 12220
rect 3568 12180 3574 12192
rect 3697 12189 3709 12192
rect 3743 12189 3755 12223
rect 3697 12183 3755 12189
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 4120 12192 4169 12220
rect 4120 12180 4126 12192
rect 4157 12189 4169 12192
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 6270 12220 6276 12232
rect 5592 12192 6276 12220
rect 5592 12180 5598 12192
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 2869 12155 2927 12161
rect 2869 12121 2881 12155
rect 2915 12152 2927 12155
rect 2958 12152 2964 12164
rect 2915 12124 2964 12152
rect 2915 12121 2927 12124
rect 2869 12115 2927 12121
rect 2958 12112 2964 12124
rect 3016 12152 3022 12164
rect 4080 12152 4108 12180
rect 3016 12124 4108 12152
rect 3016 12112 3022 12124
rect 3970 12044 3976 12096
rect 4028 12084 4034 12096
rect 5997 12087 6055 12093
rect 5997 12084 6009 12087
rect 4028 12056 6009 12084
rect 4028 12044 4034 12056
rect 5997 12053 6009 12056
rect 6043 12053 6055 12087
rect 6288 12084 6316 12180
rect 7300 12152 7328 12260
rect 7929 12257 7941 12291
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 8021 12291 8079 12297
rect 8021 12257 8033 12291
rect 8067 12257 8079 12291
rect 8021 12251 8079 12257
rect 7745 12155 7803 12161
rect 7745 12152 7757 12155
rect 7300 12124 7757 12152
rect 7745 12121 7757 12124
rect 7791 12121 7803 12155
rect 7745 12115 7803 12121
rect 6638 12084 6644 12096
rect 6288 12056 6644 12084
rect 5997 12047 6055 12053
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 7374 12084 7380 12096
rect 6972 12056 7380 12084
rect 6972 12044 6978 12056
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 7944 12084 7972 12251
rect 8110 12248 8116 12300
rect 8168 12288 8174 12300
rect 8277 12291 8335 12297
rect 8277 12288 8289 12291
rect 8168 12260 8289 12288
rect 8168 12248 8174 12260
rect 8277 12257 8289 12260
rect 8323 12257 8335 12291
rect 8277 12251 8335 12257
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 8628 12260 10057 12288
rect 8628 12248 8634 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10594 12288 10600 12300
rect 10555 12260 10600 12288
rect 10045 12251 10103 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9180 12192 10149 12220
rect 9180 12180 9186 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10704 12220 10732 12328
rect 14384 12328 14964 12356
rect 10962 12297 10968 12300
rect 10920 12291 10968 12297
rect 10920 12257 10932 12291
rect 10966 12257 10968 12291
rect 10920 12251 10968 12257
rect 10962 12248 10968 12251
rect 11020 12248 11026 12300
rect 12618 12248 12624 12300
rect 12676 12288 12682 12300
rect 12852 12291 12910 12297
rect 12852 12288 12864 12291
rect 12676 12260 12864 12288
rect 12676 12248 12682 12260
rect 12852 12257 12864 12260
rect 12898 12257 12910 12291
rect 12852 12251 12910 12257
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 13265 12291 13323 12297
rect 13265 12288 13277 12291
rect 13228 12260 13277 12288
rect 13228 12248 13234 12260
rect 13265 12257 13277 12260
rect 13311 12288 13323 12291
rect 14384 12288 14412 12328
rect 13311 12260 14412 12288
rect 14461 12291 14519 12297
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 14461 12257 14473 12291
rect 14507 12288 14519 12291
rect 14734 12288 14740 12300
rect 14507 12260 14740 12288
rect 14507 12257 14519 12260
rect 14461 12251 14519 12257
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 14829 12291 14887 12297
rect 14829 12257 14841 12291
rect 14875 12257 14887 12291
rect 14936 12288 14964 12328
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 17144 12356 17172 12396
rect 17687 12396 18092 12424
rect 18559 12396 18604 12424
rect 17687 12356 17715 12396
rect 15252 12328 16795 12356
rect 17144 12328 17715 12356
rect 15252 12316 15258 12328
rect 15378 12288 15384 12300
rect 14936 12260 15384 12288
rect 14829 12251 14887 12257
rect 11060 12223 11118 12229
rect 11060 12220 11072 12223
rect 10284 12192 10329 12220
rect 10704 12192 11072 12220
rect 10284 12180 10290 12192
rect 11060 12189 11072 12192
rect 11106 12189 11118 12223
rect 11060 12183 11118 12189
rect 11333 12223 11391 12229
rect 11333 12189 11345 12223
rect 11379 12220 11391 12223
rect 11698 12220 11704 12232
rect 11379 12192 11704 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 12492 12192 12541 12220
rect 12492 12180 12498 12192
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 12992 12223 13050 12229
rect 12992 12220 13004 12223
rect 12768 12192 13004 12220
rect 12768 12180 12774 12192
rect 12992 12189 13004 12192
rect 13038 12189 13050 12223
rect 12992 12183 13050 12189
rect 14642 12180 14648 12232
rect 14700 12220 14706 12232
rect 14844 12220 14872 12251
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 15556 12291 15614 12297
rect 15556 12257 15568 12291
rect 15602 12288 15614 12291
rect 16022 12288 16028 12300
rect 15602 12260 16028 12288
rect 15602 12257 15614 12260
rect 15556 12251 15614 12257
rect 16022 12248 16028 12260
rect 16080 12288 16086 12300
rect 16666 12288 16672 12300
rect 16080 12260 16672 12288
rect 16080 12248 16086 12260
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 16767 12288 16795 12328
rect 17770 12316 17776 12368
rect 17828 12356 17834 12368
rect 17957 12359 18015 12365
rect 17957 12356 17969 12359
rect 17828 12328 17969 12356
rect 17828 12316 17834 12328
rect 17957 12325 17969 12328
rect 18003 12325 18015 12359
rect 18064 12356 18092 12396
rect 18598 12384 18604 12396
rect 18656 12384 18662 12436
rect 19702 12424 19708 12436
rect 18699 12396 19708 12424
rect 18699 12356 18727 12396
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 19150 12365 19156 12368
rect 19144 12356 19156 12365
rect 18064 12328 18727 12356
rect 19111 12328 19156 12356
rect 17957 12319 18015 12325
rect 19144 12319 19156 12328
rect 19150 12316 19156 12319
rect 19208 12316 19214 12368
rect 19426 12316 19432 12368
rect 19484 12356 19490 12368
rect 20346 12356 20352 12368
rect 19484 12328 20352 12356
rect 19484 12316 19490 12328
rect 20346 12316 20352 12328
rect 20404 12316 20410 12368
rect 17126 12288 17132 12300
rect 16767 12260 16896 12288
rect 17087 12260 17132 12288
rect 15286 12220 15292 12232
rect 14700 12192 14872 12220
rect 15247 12192 15292 12220
rect 14700 12180 14706 12192
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 16298 12180 16304 12232
rect 16356 12220 16362 12232
rect 16356 12192 16804 12220
rect 16356 12180 16362 12192
rect 16776 12161 16804 12192
rect 16761 12155 16819 12161
rect 9324 12124 10640 12152
rect 9324 12084 9352 12124
rect 7944 12056 9352 12084
rect 10612 12084 10640 12124
rect 16761 12121 16773 12155
rect 16807 12121 16819 12155
rect 16761 12115 16819 12121
rect 11330 12084 11336 12096
rect 10612 12056 11336 12084
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 12437 12087 12495 12093
rect 12437 12053 12449 12087
rect 12483 12084 12495 12087
rect 12894 12084 12900 12096
rect 12483 12056 12900 12084
rect 12483 12053 12495 12056
rect 12437 12047 12495 12053
rect 12894 12044 12900 12056
rect 12952 12084 12958 12096
rect 13170 12084 13176 12096
rect 12952 12056 13176 12084
rect 12952 12044 12958 12056
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 14645 12087 14703 12093
rect 14645 12053 14657 12087
rect 14691 12084 14703 12087
rect 15194 12084 15200 12096
rect 14691 12056 15200 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 16666 12084 16672 12096
rect 16627 12056 16672 12084
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 16868 12084 16896 12260
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17310 12248 17316 12300
rect 17368 12288 17374 12300
rect 18417 12291 18475 12297
rect 18417 12288 18429 12291
rect 17368 12260 18429 12288
rect 17368 12248 17374 12260
rect 18417 12257 18429 12260
rect 18463 12257 18475 12291
rect 18417 12251 18475 12257
rect 17218 12220 17224 12232
rect 17179 12192 17224 12220
rect 17218 12180 17224 12192
rect 17276 12180 17282 12232
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12220 17463 12223
rect 17586 12220 17592 12232
rect 17451 12192 17592 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 17862 12180 17868 12232
rect 17920 12220 17926 12232
rect 18049 12223 18107 12229
rect 18049 12220 18061 12223
rect 17920 12192 18061 12220
rect 17920 12180 17926 12192
rect 18049 12189 18061 12192
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12189 18199 12223
rect 18874 12220 18880 12232
rect 18835 12192 18880 12220
rect 18141 12183 18199 12189
rect 17604 12152 17632 12180
rect 18156 12152 18184 12183
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 20162 12180 20168 12232
rect 20220 12220 20226 12232
rect 20349 12223 20407 12229
rect 20349 12220 20361 12223
rect 20220 12192 20361 12220
rect 20220 12180 20226 12192
rect 20349 12189 20361 12192
rect 20395 12189 20407 12223
rect 20349 12183 20407 12189
rect 17604 12124 18184 12152
rect 17589 12087 17647 12093
rect 17589 12084 17601 12087
rect 16868 12056 17601 12084
rect 17589 12053 17601 12056
rect 17635 12053 17647 12087
rect 17589 12047 17647 12053
rect 20257 12087 20315 12093
rect 20257 12053 20269 12087
rect 20303 12084 20315 12087
rect 20346 12084 20352 12096
rect 20303 12056 20352 12084
rect 20303 12053 20315 12056
rect 20257 12047 20315 12053
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 1104 11994 20884 12016
rect 1104 11942 4280 11994
rect 4332 11942 4344 11994
rect 4396 11942 4408 11994
rect 4460 11942 4472 11994
rect 4524 11942 10878 11994
rect 10930 11942 10942 11994
rect 10994 11942 11006 11994
rect 11058 11942 11070 11994
rect 11122 11942 17475 11994
rect 17527 11942 17539 11994
rect 17591 11942 17603 11994
rect 17655 11942 17667 11994
rect 17719 11942 20884 11994
rect 1104 11920 20884 11942
rect 3697 11883 3755 11889
rect 3697 11849 3709 11883
rect 3743 11880 3755 11883
rect 4890 11880 4896 11892
rect 3743 11852 4896 11880
rect 3743 11849 3755 11852
rect 3697 11843 3755 11849
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 5350 11880 5356 11892
rect 5311 11852 5356 11880
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 10502 11880 10508 11892
rect 5951 11852 8984 11880
rect 10463 11852 10508 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 1857 11815 1915 11821
rect 1857 11781 1869 11815
rect 1903 11812 1915 11815
rect 5721 11815 5779 11821
rect 1903 11784 3556 11812
rect 1903 11781 1915 11784
rect 1857 11775 1915 11781
rect 2498 11744 2504 11756
rect 2459 11716 2504 11744
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 3326 11744 3332 11756
rect 3287 11716 3332 11744
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 3528 11685 3556 11784
rect 5721 11781 5733 11815
rect 5767 11812 5779 11815
rect 6822 11812 6828 11824
rect 5767 11784 6828 11812
rect 5767 11781 5779 11784
rect 5721 11775 5779 11781
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 8297 11815 8355 11821
rect 8297 11812 8309 11815
rect 7852 11784 8309 11812
rect 6270 11704 6276 11756
rect 6328 11744 6334 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6328 11716 6561 11744
rect 6328 11704 6334 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 6656 11716 6960 11744
rect 3513 11679 3571 11685
rect 3513 11645 3525 11679
rect 3559 11645 3571 11679
rect 3970 11676 3976 11688
rect 3931 11648 3976 11676
rect 3513 11639 3571 11645
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11676 5595 11679
rect 6656 11676 6684 11716
rect 5583 11648 6684 11676
rect 5583 11645 5595 11648
rect 5537 11639 5595 11645
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 6832 11679 6890 11685
rect 6832 11676 6844 11679
rect 6788 11648 6844 11676
rect 6788 11636 6794 11648
rect 6832 11645 6844 11648
rect 6878 11645 6890 11679
rect 6932 11676 6960 11716
rect 7852 11676 7880 11784
rect 8297 11781 8309 11784
rect 8343 11781 8355 11815
rect 8297 11775 8355 11781
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8849 11747 8907 11753
rect 8849 11744 8861 11747
rect 8536 11716 8861 11744
rect 8536 11704 8542 11716
rect 8849 11713 8861 11716
rect 8895 11713 8907 11747
rect 8849 11707 8907 11713
rect 6932 11648 7880 11676
rect 6832 11639 6890 11645
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 7984 11648 8677 11676
rect 7984 11636 7990 11648
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 8956 11676 8984 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 14001 11883 14059 11889
rect 10744 11852 12296 11880
rect 10744 11840 10750 11852
rect 12268 11756 12296 11852
rect 14001 11849 14013 11883
rect 14047 11880 14059 11883
rect 14090 11880 14096 11892
rect 14047 11852 14096 11880
rect 14047 11849 14059 11852
rect 14001 11843 14059 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 16666 11840 16672 11892
rect 16724 11880 16730 11892
rect 17862 11880 17868 11892
rect 16724 11852 17448 11880
rect 17823 11852 17868 11880
rect 16724 11840 16730 11852
rect 16022 11772 16028 11824
rect 16080 11812 16086 11824
rect 16301 11815 16359 11821
rect 16301 11812 16313 11815
rect 16080 11784 16313 11812
rect 16080 11772 16086 11784
rect 16301 11781 16313 11784
rect 16347 11781 16359 11815
rect 17420 11812 17448 11852
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 19794 11880 19800 11892
rect 17972 11852 19800 11880
rect 17972 11812 18000 11852
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 17420 11784 18000 11812
rect 16301 11775 16359 11781
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 10686 11744 10692 11756
rect 9999 11716 10088 11744
rect 10647 11716 10692 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 8803 11648 8984 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 2225 11611 2283 11617
rect 2225 11577 2237 11611
rect 2271 11608 2283 11611
rect 3053 11611 3111 11617
rect 2271 11580 2728 11608
rect 2271 11577 2283 11580
rect 2225 11571 2283 11577
rect 2314 11540 2320 11552
rect 2275 11512 2320 11540
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 2700 11549 2728 11580
rect 3053 11577 3065 11611
rect 3099 11608 3111 11611
rect 4240 11611 4298 11617
rect 3099 11580 4200 11608
rect 3099 11577 3111 11580
rect 3053 11571 3111 11577
rect 4172 11552 4200 11580
rect 4240 11577 4252 11611
rect 4286 11608 4298 11611
rect 4614 11608 4620 11620
rect 4286 11580 4620 11608
rect 4286 11577 4298 11580
rect 4240 11571 4298 11577
rect 4614 11568 4620 11580
rect 4672 11608 4678 11620
rect 5442 11608 5448 11620
rect 4672 11580 5448 11608
rect 4672 11568 4678 11580
rect 5442 11568 5448 11580
rect 5500 11568 5506 11620
rect 7098 11617 7104 11620
rect 6273 11611 6331 11617
rect 6273 11577 6285 11611
rect 6319 11608 6331 11611
rect 7092 11608 7104 11617
rect 6319 11580 7104 11608
rect 6319 11577 6331 11580
rect 6273 11571 6331 11577
rect 7092 11571 7104 11580
rect 7098 11568 7104 11571
rect 7156 11568 7162 11620
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 9122 11608 9128 11620
rect 7248 11580 9128 11608
rect 7248 11568 7254 11580
rect 9122 11568 9128 11580
rect 9180 11568 9186 11620
rect 9398 11568 9404 11620
rect 9456 11608 9462 11620
rect 10060 11608 10088 11716
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 12250 11744 12256 11756
rect 12163 11716 12256 11744
rect 12250 11704 12256 11716
rect 12308 11744 12314 11756
rect 12529 11747 12587 11753
rect 12529 11744 12541 11747
rect 12308 11716 12541 11744
rect 12308 11704 12314 11716
rect 12529 11713 12541 11716
rect 12575 11713 12587 11747
rect 14550 11744 14556 11756
rect 14511 11716 14556 11744
rect 12529 11707 12587 11713
rect 14550 11704 14556 11716
rect 14608 11704 14614 11756
rect 16408 11716 16620 11744
rect 10321 11679 10379 11685
rect 10321 11645 10333 11679
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 10956 11679 11014 11685
rect 10956 11645 10968 11679
rect 11002 11676 11014 11679
rect 11238 11676 11244 11688
rect 11002 11648 11244 11676
rect 11002 11645 11014 11648
rect 10956 11639 11014 11645
rect 9456 11580 10088 11608
rect 10336 11608 10364 11639
rect 11238 11636 11244 11648
rect 11296 11636 11302 11688
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 14369 11679 14427 11685
rect 11388 11648 13952 11676
rect 11388 11636 11394 11648
rect 11422 11608 11428 11620
rect 10336 11580 11428 11608
rect 9456 11568 9462 11580
rect 2685 11543 2743 11549
rect 2685 11509 2697 11543
rect 2731 11509 2743 11543
rect 2685 11503 2743 11509
rect 3142 11500 3148 11552
rect 3200 11540 3206 11552
rect 3200 11512 3245 11540
rect 3200 11500 3206 11512
rect 4154 11500 4160 11552
rect 4212 11500 4218 11552
rect 6365 11543 6423 11549
rect 6365 11509 6377 11543
rect 6411 11540 6423 11543
rect 7282 11540 7288 11552
rect 6411 11512 7288 11540
rect 6411 11509 6423 11512
rect 6365 11503 6423 11509
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 8202 11540 8208 11552
rect 8163 11512 8208 11540
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 8352 11512 9321 11540
rect 8352 11500 8358 11512
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 9674 11540 9680 11552
rect 9635 11512 9680 11540
rect 9309 11503 9367 11509
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 10060 11540 10088 11580
rect 11422 11568 11428 11580
rect 11480 11568 11486 11620
rect 12526 11608 12532 11620
rect 11532 11580 12532 11608
rect 11532 11540 11560 11580
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 12796 11611 12854 11617
rect 12796 11577 12808 11611
rect 12842 11608 12854 11611
rect 13814 11608 13820 11620
rect 12842 11580 13820 11608
rect 12842 11577 12854 11580
rect 12796 11571 12854 11577
rect 13814 11568 13820 11580
rect 13872 11568 13878 11620
rect 13924 11608 13952 11648
rect 14369 11645 14381 11679
rect 14415 11676 14427 11679
rect 14826 11676 14832 11688
rect 14415 11648 14832 11676
rect 14415 11645 14427 11648
rect 14369 11639 14427 11645
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 15188 11679 15246 11685
rect 15188 11645 15200 11679
rect 15234 11676 15246 11679
rect 16408 11676 16436 11716
rect 15234 11648 16436 11676
rect 16485 11679 16543 11685
rect 15234 11645 15246 11648
rect 15188 11639 15246 11645
rect 16485 11645 16497 11679
rect 16531 11645 16543 11679
rect 16485 11639 16543 11645
rect 14642 11608 14648 11620
rect 13924 11580 14648 11608
rect 14642 11568 14648 11580
rect 14700 11568 14706 11620
rect 14936 11608 14964 11639
rect 15286 11608 15292 11620
rect 14936 11580 15292 11608
rect 15286 11568 15292 11580
rect 15344 11608 15350 11620
rect 16298 11608 16304 11620
rect 15344 11580 16304 11608
rect 15344 11568 15350 11580
rect 16298 11568 16304 11580
rect 16356 11608 16362 11620
rect 16500 11608 16528 11639
rect 16356 11580 16528 11608
rect 16356 11568 16362 11580
rect 9824 11512 9869 11540
rect 10060 11512 11560 11540
rect 9824 11500 9830 11512
rect 11974 11500 11980 11552
rect 12032 11540 12038 11552
rect 12069 11543 12127 11549
rect 12069 11540 12081 11543
rect 12032 11512 12081 11540
rect 12032 11500 12038 11512
rect 12069 11509 12081 11512
rect 12115 11509 12127 11543
rect 12069 11503 12127 11509
rect 12158 11500 12164 11552
rect 12216 11540 12222 11552
rect 13722 11540 13728 11552
rect 12216 11512 13728 11540
rect 12216 11500 12222 11512
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 13906 11540 13912 11552
rect 13867 11512 13912 11540
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 14458 11540 14464 11552
rect 14419 11512 14464 11540
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 16592 11540 16620 11716
rect 17770 11704 17776 11756
rect 17828 11744 17834 11756
rect 17828 11716 18184 11744
rect 17828 11704 17834 11716
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11645 18107 11679
rect 18156 11676 18184 11716
rect 20070 11704 20076 11756
rect 20128 11744 20134 11756
rect 20257 11747 20315 11753
rect 20257 11744 20269 11747
rect 20128 11716 20269 11744
rect 20128 11704 20134 11716
rect 20257 11713 20269 11716
rect 20303 11713 20315 11747
rect 20257 11707 20315 11713
rect 20346 11704 20352 11756
rect 20404 11744 20410 11756
rect 20404 11716 20449 11744
rect 20404 11704 20410 11716
rect 18305 11679 18363 11685
rect 18305 11676 18317 11679
rect 18156 11648 18317 11676
rect 18049 11639 18107 11645
rect 18305 11645 18317 11648
rect 18351 11645 18363 11679
rect 20162 11676 20168 11688
rect 20123 11648 20168 11676
rect 18305 11639 18363 11645
rect 16752 11611 16810 11617
rect 16752 11577 16764 11611
rect 16798 11608 16810 11611
rect 17126 11608 17132 11620
rect 16798 11580 17132 11608
rect 16798 11577 16810 11580
rect 16752 11571 16810 11577
rect 17126 11568 17132 11580
rect 17184 11568 17190 11620
rect 17402 11568 17408 11620
rect 17460 11608 17466 11620
rect 18064 11608 18092 11639
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 18874 11608 18880 11620
rect 17460 11580 18880 11608
rect 17460 11568 17466 11580
rect 18874 11568 18880 11580
rect 18932 11568 18938 11620
rect 16666 11540 16672 11552
rect 16592 11512 16672 11540
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 18414 11500 18420 11552
rect 18472 11540 18478 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 18472 11512 19441 11540
rect 18472 11500 18478 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19429 11503 19487 11509
rect 19797 11543 19855 11549
rect 19797 11509 19809 11543
rect 19843 11540 19855 11543
rect 19886 11540 19892 11552
rect 19843 11512 19892 11540
rect 19843 11509 19855 11512
rect 19797 11503 19855 11509
rect 19886 11500 19892 11512
rect 19944 11500 19950 11552
rect 1104 11450 20884 11472
rect 1104 11398 7579 11450
rect 7631 11398 7643 11450
rect 7695 11398 7707 11450
rect 7759 11398 7771 11450
rect 7823 11398 14176 11450
rect 14228 11398 14240 11450
rect 14292 11398 14304 11450
rect 14356 11398 14368 11450
rect 14420 11398 20884 11450
rect 1104 11376 20884 11398
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 2869 11339 2927 11345
rect 2869 11336 2881 11339
rect 2372 11308 2881 11336
rect 2372 11296 2378 11308
rect 2869 11305 2881 11308
rect 2915 11305 2927 11339
rect 2869 11299 2927 11305
rect 3697 11339 3755 11345
rect 3697 11305 3709 11339
rect 3743 11305 3755 11339
rect 5442 11336 5448 11348
rect 5403 11308 5448 11336
rect 3697 11299 3755 11305
rect 3326 11228 3332 11280
rect 3384 11228 3390 11280
rect 3712 11268 3740 11299
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 5905 11339 5963 11345
rect 5905 11305 5917 11339
rect 5951 11336 5963 11339
rect 7190 11336 7196 11348
rect 5951 11308 7196 11336
rect 5951 11305 5963 11308
rect 5905 11299 5963 11305
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 7929 11339 7987 11345
rect 7929 11305 7941 11339
rect 7975 11305 7987 11339
rect 8294 11336 8300 11348
rect 8255 11308 8300 11336
rect 7929 11299 7987 11305
rect 5534 11268 5540 11280
rect 3712 11240 5540 11268
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 7650 11268 7656 11280
rect 5736 11240 7656 11268
rect 1486 11160 1492 11212
rect 1544 11200 1550 11212
rect 1653 11203 1711 11209
rect 1653 11200 1665 11203
rect 1544 11172 1665 11200
rect 1544 11160 1550 11172
rect 1653 11169 1665 11172
rect 1699 11169 1711 11203
rect 3234 11200 3240 11212
rect 3195 11172 3240 11200
rect 1653 11163 1711 11169
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 3344 11200 3372 11228
rect 3344 11172 3464 11200
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 3436 11141 3464 11172
rect 3786 11160 3792 11212
rect 3844 11200 3850 11212
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3844 11172 3893 11200
rect 3844 11160 3850 11172
rect 3881 11169 3893 11172
rect 3927 11169 3939 11203
rect 3881 11163 3939 11169
rect 4332 11203 4390 11209
rect 4332 11169 4344 11203
rect 4378 11200 4390 11203
rect 4614 11200 4620 11212
rect 4378 11172 4620 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5736 11209 5764 11240
rect 7650 11228 7656 11240
rect 7708 11228 7714 11280
rect 5721 11203 5779 11209
rect 5721 11169 5733 11203
rect 5767 11169 5779 11203
rect 5721 11163 5779 11169
rect 6356 11203 6414 11209
rect 6356 11169 6368 11203
rect 6402 11200 6414 11203
rect 6638 11200 6644 11212
rect 6402 11172 6644 11200
rect 6402 11169 6414 11172
rect 6356 11163 6414 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 7944 11200 7972 11299
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8389 11339 8447 11345
rect 8389 11305 8401 11339
rect 8435 11336 8447 11339
rect 8757 11339 8815 11345
rect 8757 11336 8769 11339
rect 8435 11308 8769 11336
rect 8435 11305 8447 11308
rect 8389 11299 8447 11305
rect 8757 11305 8769 11308
rect 8803 11305 8815 11339
rect 8757 11299 8815 11305
rect 9600 11308 11192 11336
rect 8110 11228 8116 11280
rect 8168 11268 8174 11280
rect 9600 11268 9628 11308
rect 8168 11240 9628 11268
rect 8168 11228 8174 11240
rect 9674 11228 9680 11280
rect 9732 11268 9738 11280
rect 11164 11268 11192 11308
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 11333 11339 11391 11345
rect 11333 11336 11345 11339
rect 11296 11308 11345 11336
rect 11296 11296 11302 11308
rect 11333 11305 11345 11308
rect 11379 11305 11391 11339
rect 11333 11299 11391 11305
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 13630 11336 13636 11348
rect 12299 11308 13636 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 14458 11336 14464 11348
rect 13780 11308 14464 11336
rect 13780 11296 13786 11308
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 14737 11339 14795 11345
rect 14737 11305 14749 11339
rect 14783 11336 14795 11339
rect 14826 11336 14832 11348
rect 14783 11308 14832 11336
rect 14783 11305 14795 11308
rect 14737 11299 14795 11305
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 15194 11296 15200 11348
rect 15252 11336 15258 11348
rect 16669 11339 16727 11345
rect 15252 11308 16620 11336
rect 15252 11296 15258 11308
rect 11974 11268 11980 11280
rect 9732 11240 10088 11268
rect 11164 11240 11980 11268
rect 9732 11228 9738 11240
rect 7607 11172 7972 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 8846 11160 8852 11212
rect 8904 11200 8910 11212
rect 9125 11203 9183 11209
rect 9125 11200 9137 11203
rect 8904 11172 9137 11200
rect 8904 11160 8910 11172
rect 9125 11169 9137 11172
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 9953 11203 10011 11209
rect 9953 11200 9965 11203
rect 9640 11172 9965 11200
rect 9640 11160 9646 11172
rect 9953 11169 9965 11172
rect 9999 11169 10011 11203
rect 10060 11200 10088 11240
rect 11974 11228 11980 11240
rect 12032 11228 12038 11280
rect 12621 11271 12679 11277
rect 12621 11237 12633 11271
rect 12667 11268 12679 11271
rect 13348 11271 13406 11277
rect 13348 11268 13360 11271
rect 12667 11240 13360 11268
rect 12667 11237 12679 11240
rect 12621 11231 12679 11237
rect 13348 11237 13360 11240
rect 13394 11268 13406 11271
rect 13906 11268 13912 11280
rect 13394 11240 13912 11268
rect 13394 11237 13406 11240
rect 13348 11231 13406 11237
rect 13906 11228 13912 11240
rect 13964 11228 13970 11280
rect 16114 11268 16120 11280
rect 14568 11240 16120 11268
rect 10220 11203 10278 11209
rect 10220 11200 10232 11203
rect 10060 11172 10232 11200
rect 9953 11163 10011 11169
rect 10220 11169 10232 11172
rect 10266 11200 10278 11203
rect 11514 11200 11520 11212
rect 10266 11172 11520 11200
rect 10266 11169 10278 11172
rect 10220 11163 10278 11169
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11200 11851 11203
rect 12434 11200 12440 11212
rect 11839 11172 12440 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11200 12771 11203
rect 13814 11200 13820 11212
rect 12759 11172 13820 11200
rect 12759 11169 12771 11172
rect 12713 11163 12771 11169
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 14568 11209 14596 11240
rect 16114 11228 16120 11240
rect 16172 11228 16178 11280
rect 16592 11268 16620 11308
rect 16669 11305 16681 11339
rect 16715 11336 16727 11339
rect 16758 11336 16764 11348
rect 16715 11308 16764 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 16758 11296 16764 11308
rect 16816 11296 16822 11348
rect 17221 11339 17279 11345
rect 17221 11305 17233 11339
rect 17267 11336 17279 11339
rect 18322 11336 18328 11348
rect 17267 11308 18328 11336
rect 17267 11305 17279 11308
rect 17221 11299 17279 11305
rect 18322 11296 18328 11308
rect 18380 11296 18386 11348
rect 20070 11336 20076 11348
rect 19352 11308 20076 11336
rect 17672 11271 17730 11277
rect 16592 11240 17632 11268
rect 14553 11203 14611 11209
rect 14553 11169 14565 11203
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 15562 11209 15568 11212
rect 15105 11203 15163 11209
rect 15105 11200 15117 11203
rect 14700 11172 15117 11200
rect 14700 11160 14706 11172
rect 15105 11169 15117 11172
rect 15151 11169 15163 11203
rect 15105 11163 15163 11169
rect 15556 11163 15568 11209
rect 15620 11200 15626 11212
rect 15620 11172 15656 11200
rect 15562 11160 15568 11163
rect 15620 11160 15626 11172
rect 16574 11160 16580 11212
rect 16632 11200 16638 11212
rect 16945 11203 17003 11209
rect 16945 11200 16957 11203
rect 16632 11172 16957 11200
rect 16632 11160 16638 11172
rect 16945 11169 16957 11172
rect 16991 11169 17003 11203
rect 16945 11163 17003 11169
rect 17034 11160 17040 11212
rect 17092 11200 17098 11212
rect 17604 11200 17632 11240
rect 17672 11237 17684 11271
rect 17718 11268 17730 11271
rect 19352 11268 19380 11308
rect 20070 11296 20076 11308
rect 20128 11336 20134 11348
rect 20533 11339 20591 11345
rect 20533 11336 20545 11339
rect 20128 11308 20545 11336
rect 20128 11296 20134 11308
rect 20533 11305 20545 11308
rect 20579 11305 20591 11339
rect 20533 11299 20591 11305
rect 17718 11240 19380 11268
rect 19420 11271 19478 11277
rect 17718 11237 17730 11240
rect 17672 11231 17730 11237
rect 19420 11237 19432 11271
rect 19466 11268 19478 11271
rect 20346 11268 20352 11280
rect 19466 11240 20352 11268
rect 19466 11237 19478 11240
rect 19420 11231 19478 11237
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 19242 11200 19248 11212
rect 17092 11172 17137 11200
rect 17604 11172 19248 11200
rect 17092 11160 17098 11172
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 3329 11135 3387 11141
rect 3329 11132 3341 11135
rect 2792 11104 3341 11132
rect 2792 11076 2820 11104
rect 3329 11101 3341 11104
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11101 3479 11135
rect 3421 11095 3479 11101
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 2832 11036 2925 11064
rect 2832 11024 2838 11036
rect 4080 11008 4108 11095
rect 6104 11064 6132 11095
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 8110 11132 8116 11144
rect 7340 11104 8116 11132
rect 7340 11092 7346 11104
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8294 11092 8300 11144
rect 8352 11132 8358 11144
rect 8478 11132 8484 11144
rect 8352 11104 8484 11132
rect 8352 11092 8358 11104
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 9214 11132 9220 11144
rect 9175 11104 9220 11132
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 9398 11132 9404 11144
rect 9359 11104 9404 11132
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 9674 11132 9680 11144
rect 9635 11104 9680 11132
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 11882 11132 11888 11144
rect 11843 11104 11888 11132
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11132 12127 11135
rect 12802 11132 12808 11144
rect 12115 11104 12808 11132
rect 12115 11101 12127 11104
rect 12069 11095 12127 11101
rect 5000 11036 6132 11064
rect 4062 10996 4068 11008
rect 3975 10968 4068 10996
rect 4062 10956 4068 10968
rect 4120 10996 4126 11008
rect 5000 10996 5028 11036
rect 7098 11024 7104 11076
rect 7156 11064 7162 11076
rect 7745 11067 7803 11073
rect 7156 11036 7604 11064
rect 7156 11024 7162 11036
rect 4120 10968 5028 10996
rect 4120 10956 4126 10968
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 7469 10999 7527 11005
rect 7469 10996 7481 10999
rect 7248 10968 7481 10996
rect 7248 10956 7254 10968
rect 7469 10965 7481 10968
rect 7515 10965 7527 10999
rect 7576 10996 7604 11036
rect 7745 11033 7757 11067
rect 7791 11064 7803 11067
rect 8570 11064 8576 11076
rect 7791 11036 8576 11064
rect 7791 11033 7803 11036
rect 7745 11027 7803 11033
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 8662 11024 8668 11076
rect 8720 11064 8726 11076
rect 9416 11064 9444 11092
rect 12084 11064 12112 11095
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 13081 11135 13139 11141
rect 13081 11101 13093 11135
rect 13127 11101 13139 11135
rect 15286 11132 15292 11144
rect 15247 11104 15292 11132
rect 13081 11095 13139 11101
rect 8720 11036 9444 11064
rect 10888 11036 12112 11064
rect 8720 11024 8726 11036
rect 7926 10996 7932 11008
rect 7576 10968 7932 10996
rect 7469 10959 7527 10965
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 10888 10996 10916 11036
rect 12250 11024 12256 11076
rect 12308 11064 12314 11076
rect 13096 11064 13124 11095
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 17402 11132 17408 11144
rect 17315 11104 17408 11132
rect 17402 11092 17408 11104
rect 17460 11092 17466 11144
rect 18874 11132 18880 11144
rect 18835 11104 18880 11132
rect 18874 11092 18880 11104
rect 18932 11092 18938 11144
rect 18966 11092 18972 11144
rect 19024 11132 19030 11144
rect 19153 11135 19211 11141
rect 19153 11132 19165 11135
rect 19024 11104 19165 11132
rect 19024 11092 19030 11104
rect 19153 11101 19165 11104
rect 19199 11101 19211 11135
rect 19153 11095 19211 11101
rect 14458 11064 14464 11076
rect 12308 11036 13124 11064
rect 14371 11036 14464 11064
rect 12308 11024 12314 11036
rect 14458 11024 14464 11036
rect 14516 11064 14522 11076
rect 14516 11036 15332 11064
rect 14516 11024 14522 11036
rect 9364 10968 10916 10996
rect 9364 10956 9370 10968
rect 11422 10956 11428 11008
rect 11480 10996 11486 11008
rect 11480 10968 11525 10996
rect 11480 10956 11486 10968
rect 11606 10956 11612 11008
rect 11664 10996 11670 11008
rect 12342 10996 12348 11008
rect 11664 10968 12348 10996
rect 11664 10956 11670 10968
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 14918 10996 14924 11008
rect 14879 10968 14924 10996
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 15304 10996 15332 11036
rect 16298 11024 16304 11076
rect 16356 11064 16362 11076
rect 16761 11067 16819 11073
rect 16761 11064 16773 11067
rect 16356 11036 16773 11064
rect 16356 11024 16362 11036
rect 16761 11033 16773 11036
rect 16807 11064 16819 11067
rect 17420 11064 17448 11092
rect 16807 11036 17448 11064
rect 16807 11033 16819 11036
rect 16761 11027 16819 11033
rect 17310 10996 17316 11008
rect 15304 10968 17316 10996
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 18690 10956 18696 11008
rect 18748 10996 18754 11008
rect 18785 10999 18843 11005
rect 18785 10996 18797 10999
rect 18748 10968 18797 10996
rect 18748 10956 18754 10968
rect 18785 10965 18797 10968
rect 18831 10965 18843 10999
rect 18785 10959 18843 10965
rect 1104 10906 20884 10928
rect 1104 10854 4280 10906
rect 4332 10854 4344 10906
rect 4396 10854 4408 10906
rect 4460 10854 4472 10906
rect 4524 10854 10878 10906
rect 10930 10854 10942 10906
rect 10994 10854 11006 10906
rect 11058 10854 11070 10906
rect 11122 10854 17475 10906
rect 17527 10854 17539 10906
rect 17591 10854 17603 10906
rect 17655 10854 17667 10906
rect 17719 10854 20884 10906
rect 1104 10832 20884 10854
rect 2777 10795 2835 10801
rect 2777 10761 2789 10795
rect 2823 10792 2835 10795
rect 3234 10792 3240 10804
rect 2823 10764 3240 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 4249 10795 4307 10801
rect 4249 10792 4261 10795
rect 4212 10764 4261 10792
rect 4212 10752 4218 10764
rect 4249 10761 4261 10764
rect 4295 10761 4307 10795
rect 4249 10755 4307 10761
rect 4264 10656 4292 10755
rect 4614 10752 4620 10804
rect 4672 10792 4678 10804
rect 5721 10795 5779 10801
rect 5721 10792 5733 10795
rect 4672 10764 5733 10792
rect 4672 10752 4678 10764
rect 5721 10761 5733 10764
rect 5767 10761 5779 10795
rect 5721 10755 5779 10761
rect 6825 10795 6883 10801
rect 6825 10761 6837 10795
rect 6871 10792 6883 10795
rect 7098 10792 7104 10804
rect 6871 10764 7104 10792
rect 6871 10761 6883 10764
rect 6825 10755 6883 10761
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 7650 10792 7656 10804
rect 7611 10764 7656 10792
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 8018 10752 8024 10804
rect 8076 10792 8082 10804
rect 8076 10764 9720 10792
rect 8076 10752 8082 10764
rect 6546 10684 6552 10736
rect 6604 10724 6610 10736
rect 9692 10724 9720 10764
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 9824 10764 10057 10792
rect 9824 10752 9830 10764
rect 10045 10761 10057 10764
rect 10091 10792 10103 10795
rect 10318 10792 10324 10804
rect 10091 10764 10324 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11609 10795 11667 10801
rect 11609 10792 11621 10795
rect 11388 10764 11621 10792
rect 11388 10752 11394 10764
rect 11609 10761 11621 10764
rect 11655 10761 11667 10795
rect 11609 10755 11667 10761
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 13170 10792 13176 10804
rect 11848 10764 13176 10792
rect 11848 10752 11854 10764
rect 13170 10752 13176 10764
rect 13228 10752 13234 10804
rect 13814 10792 13820 10804
rect 13775 10764 13820 10792
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 15286 10792 15292 10804
rect 13924 10764 15292 10792
rect 12158 10724 12164 10736
rect 6604 10696 8524 10724
rect 9692 10696 12164 10724
rect 6604 10684 6610 10696
rect 4264 10628 4476 10656
rect 1394 10588 1400 10600
rect 1307 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 1664 10591 1722 10597
rect 1664 10557 1676 10591
rect 1710 10588 1722 10591
rect 2774 10588 2780 10600
rect 1710 10560 2780 10588
rect 1710 10557 1722 10560
rect 1664 10551 1722 10557
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 3142 10597 3148 10600
rect 2869 10591 2927 10597
rect 2869 10557 2881 10591
rect 2915 10557 2927 10591
rect 3136 10588 3148 10597
rect 3103 10560 3148 10588
rect 2869 10551 2927 10557
rect 3136 10551 3148 10560
rect 1412 10520 1440 10548
rect 2884 10520 2912 10551
rect 3142 10548 3148 10551
rect 3200 10548 3206 10600
rect 4062 10548 4068 10600
rect 4120 10588 4126 10600
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 4120 10560 4353 10588
rect 4120 10548 4126 10560
rect 4341 10557 4353 10560
rect 4387 10557 4399 10591
rect 4448 10588 4476 10628
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 5592 10628 6285 10656
rect 5592 10616 5598 10628
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 6454 10656 6460 10668
rect 6415 10628 6460 10656
rect 6273 10619 6331 10625
rect 6454 10616 6460 10628
rect 6512 10616 6518 10668
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 4597 10591 4655 10597
rect 4597 10588 4609 10591
rect 4448 10560 4609 10588
rect 4341 10551 4399 10557
rect 4597 10557 4609 10560
rect 4643 10557 4655 10591
rect 4597 10551 4655 10557
rect 5718 10548 5724 10600
rect 5776 10588 5782 10600
rect 7190 10588 7196 10600
rect 5776 10560 7196 10588
rect 5776 10548 5782 10560
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 4080 10520 4108 10548
rect 1412 10492 4108 10520
rect 4154 10480 4160 10532
rect 4212 10520 4218 10532
rect 7006 10520 7012 10532
rect 4212 10492 7012 10520
rect 4212 10480 4218 10492
rect 7006 10480 7012 10492
rect 7064 10480 7070 10532
rect 7374 10480 7380 10532
rect 7432 10520 7438 10532
rect 7484 10520 7512 10619
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 8352 10628 8397 10656
rect 8352 10616 8358 10628
rect 8202 10588 8208 10600
rect 7432 10492 7512 10520
rect 7668 10560 8208 10588
rect 7432 10480 7438 10492
rect 5810 10412 5816 10464
rect 5868 10452 5874 10464
rect 5868 10424 5913 10452
rect 5868 10412 5874 10424
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6181 10455 6239 10461
rect 6181 10452 6193 10455
rect 6052 10424 6193 10452
rect 6052 10412 6058 10424
rect 6181 10421 6193 10424
rect 6227 10421 6239 10455
rect 6181 10415 6239 10421
rect 6638 10412 6644 10464
rect 6696 10452 6702 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 6696 10424 7297 10452
rect 6696 10412 6702 10424
rect 7285 10421 7297 10424
rect 7331 10452 7343 10455
rect 7668 10452 7696 10560
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 7742 10480 7748 10532
rect 7800 10520 7806 10532
rect 8113 10523 8171 10529
rect 8113 10520 8125 10523
rect 7800 10492 8125 10520
rect 7800 10480 7806 10492
rect 8113 10489 8125 10492
rect 8159 10489 8171 10523
rect 8113 10483 8171 10489
rect 8018 10452 8024 10464
rect 7331 10424 7696 10452
rect 7979 10424 8024 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 8496 10452 8524 10696
rect 12158 10684 12164 10696
rect 12216 10684 12222 10736
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 13924 10665 13952 10764
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 16758 10792 16764 10804
rect 16080 10764 16620 10792
rect 16671 10764 16764 10792
rect 16080 10752 16086 10764
rect 16592 10724 16620 10764
rect 16758 10752 16764 10764
rect 16816 10792 16822 10804
rect 17218 10792 17224 10804
rect 16816 10764 17224 10792
rect 16816 10752 16822 10764
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 16592 10696 17448 10724
rect 12437 10659 12495 10665
rect 12437 10656 12449 10659
rect 12308 10628 12449 10656
rect 12308 10616 12314 10628
rect 12437 10625 12449 10628
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 13909 10659 13967 10665
rect 13909 10625 13921 10659
rect 13955 10625 13967 10659
rect 17310 10656 17316 10668
rect 17271 10628 17316 10656
rect 13909 10619 13967 10625
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 17420 10665 17448 10696
rect 17494 10684 17500 10736
rect 17552 10724 17558 10736
rect 17954 10724 17960 10736
rect 17552 10696 17960 10724
rect 17552 10684 17558 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 19334 10684 19340 10736
rect 19392 10724 19398 10736
rect 19429 10727 19487 10733
rect 19429 10724 19441 10727
rect 19392 10696 19441 10724
rect 19392 10684 19398 10696
rect 19429 10693 19441 10696
rect 19475 10693 19487 10727
rect 19429 10687 19487 10693
rect 17405 10659 17463 10665
rect 17405 10625 17417 10659
rect 17451 10625 17463 10659
rect 20070 10656 20076 10668
rect 20031 10628 20076 10656
rect 17405 10619 17463 10625
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 8665 10591 8723 10597
rect 8665 10588 8677 10591
rect 8628 10560 8677 10588
rect 8628 10548 8634 10560
rect 8665 10557 8677 10560
rect 8711 10557 8723 10591
rect 8665 10551 8723 10557
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 8812 10560 12480 10588
rect 8812 10548 8818 10560
rect 8846 10480 8852 10532
rect 8904 10529 8910 10532
rect 8904 10523 8968 10529
rect 8904 10489 8922 10523
rect 8956 10489 8968 10523
rect 8904 10483 8968 10489
rect 8904 10480 8910 10483
rect 10226 10480 10232 10532
rect 10284 10520 10290 10532
rect 10321 10523 10379 10529
rect 10321 10520 10333 10523
rect 10284 10492 10333 10520
rect 10284 10480 10290 10492
rect 10321 10489 10333 10492
rect 10367 10489 10379 10523
rect 10321 10483 10379 10489
rect 12250 10452 12256 10464
rect 8496 10424 12256 10452
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 12452 10452 12480 10560
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 12693 10591 12751 10597
rect 12693 10588 12705 10591
rect 12584 10560 12705 10588
rect 12584 10548 12590 10560
rect 12693 10557 12705 10560
rect 12739 10557 12751 10591
rect 12693 10551 12751 10557
rect 14176 10591 14234 10597
rect 14176 10557 14188 10591
rect 14222 10588 14234 10591
rect 15102 10588 15108 10600
rect 14222 10560 15108 10588
rect 14222 10557 14234 10560
rect 14176 10551 14234 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 15378 10588 15384 10600
rect 15339 10560 15384 10588
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 15488 10560 15783 10588
rect 15488 10520 15516 10560
rect 13731 10492 15516 10520
rect 15648 10523 15706 10529
rect 13731 10452 13759 10492
rect 15648 10489 15660 10523
rect 15694 10489 15706 10523
rect 15755 10520 15783 10560
rect 15930 10548 15936 10600
rect 15988 10588 15994 10600
rect 17221 10591 17279 10597
rect 17221 10588 17233 10591
rect 15988 10560 17233 10588
rect 15988 10548 15994 10560
rect 17221 10557 17233 10560
rect 17267 10557 17279 10591
rect 17221 10551 17279 10557
rect 17770 10548 17776 10600
rect 17828 10588 17834 10600
rect 17865 10591 17923 10597
rect 17865 10588 17877 10591
rect 17828 10560 17877 10588
rect 17828 10548 17834 10560
rect 17865 10557 17877 10560
rect 17911 10557 17923 10591
rect 18046 10588 18052 10600
rect 18007 10560 18052 10588
rect 17865 10551 17923 10557
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 20349 10591 20407 10597
rect 20349 10588 20361 10591
rect 18156 10560 20361 10588
rect 18156 10520 18184 10560
rect 20349 10557 20361 10560
rect 20395 10557 20407 10591
rect 20349 10551 20407 10557
rect 15755 10492 18184 10520
rect 18316 10523 18374 10529
rect 15648 10483 15706 10489
rect 18316 10489 18328 10523
rect 18362 10520 18374 10523
rect 18690 10520 18696 10532
rect 18362 10492 18696 10520
rect 18362 10489 18374 10492
rect 18316 10483 18374 10489
rect 15286 10452 15292 10464
rect 12452 10424 13759 10452
rect 15247 10424 15292 10452
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 15562 10412 15568 10464
rect 15620 10452 15626 10464
rect 15672 10452 15700 10483
rect 18690 10480 18696 10492
rect 18748 10480 18754 10532
rect 19702 10480 19708 10532
rect 19760 10520 19766 10532
rect 20806 10520 20812 10532
rect 19760 10492 20812 10520
rect 19760 10480 19766 10492
rect 20806 10480 20812 10492
rect 20864 10480 20870 10532
rect 15620 10424 15700 10452
rect 15620 10412 15626 10424
rect 15838 10412 15844 10464
rect 15896 10452 15902 10464
rect 16666 10452 16672 10464
rect 15896 10424 16672 10452
rect 15896 10412 15902 10424
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 16850 10452 16856 10464
rect 16811 10424 16856 10452
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 17681 10455 17739 10461
rect 17681 10452 17693 10455
rect 17276 10424 17693 10452
rect 17276 10412 17282 10424
rect 17681 10421 17693 10424
rect 17727 10452 17739 10455
rect 18046 10452 18052 10464
rect 17727 10424 18052 10452
rect 17727 10421 17739 10424
rect 17681 10415 17739 10421
rect 18046 10412 18052 10424
rect 18104 10452 18110 10464
rect 18506 10452 18512 10464
rect 18104 10424 18512 10452
rect 18104 10412 18110 10424
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 19518 10452 19524 10464
rect 19479 10424 19524 10452
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 19886 10452 19892 10464
rect 19847 10424 19892 10452
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 19978 10412 19984 10464
rect 20036 10452 20042 10464
rect 20036 10424 20081 10452
rect 20036 10412 20042 10424
rect 1104 10362 20884 10384
rect 1104 10310 7579 10362
rect 7631 10310 7643 10362
rect 7695 10310 7707 10362
rect 7759 10310 7771 10362
rect 7823 10310 14176 10362
rect 14228 10310 14240 10362
rect 14292 10310 14304 10362
rect 14356 10310 14368 10362
rect 14420 10310 20884 10362
rect 1104 10288 20884 10310
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 5534 10248 5540 10260
rect 5495 10220 5540 10248
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 6733 10251 6791 10257
rect 6733 10217 6745 10251
rect 6779 10248 6791 10251
rect 6914 10248 6920 10260
rect 6779 10220 6920 10248
rect 6779 10217 6791 10220
rect 6733 10211 6791 10217
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10248 7067 10251
rect 7466 10248 7472 10260
rect 7055 10220 7472 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 7837 10251 7895 10257
rect 7837 10217 7849 10251
rect 7883 10248 7895 10251
rect 8018 10248 8024 10260
rect 7883 10220 8024 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 8757 10251 8815 10257
rect 8352 10220 8423 10248
rect 8352 10208 8358 10220
rect 2032 10183 2090 10189
rect 2032 10149 2044 10183
rect 2078 10180 2090 10183
rect 3234 10180 3240 10192
rect 2078 10152 3240 10180
rect 2078 10149 2090 10152
rect 2032 10143 2090 10149
rect 3234 10140 3240 10152
rect 3292 10140 3298 10192
rect 4332 10183 4390 10189
rect 4332 10149 4344 10183
rect 4378 10180 4390 10183
rect 5718 10180 5724 10192
rect 4378 10152 5724 10180
rect 4378 10149 4390 10152
rect 4332 10143 4390 10149
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 8395 10180 8423 10220
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 8803 10220 10539 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 5868 10152 6592 10180
rect 8395 10152 9444 10180
rect 5868 10140 5874 10152
rect 1765 10115 1823 10121
rect 1765 10081 1777 10115
rect 1811 10112 1823 10115
rect 3881 10115 3939 10121
rect 1811 10084 3832 10112
rect 1811 10081 1823 10084
rect 1765 10075 1823 10081
rect 3804 10056 3832 10084
rect 3881 10081 3893 10115
rect 3927 10112 3939 10115
rect 4154 10112 4160 10124
rect 3927 10084 4160 10112
rect 3927 10081 3939 10084
rect 3881 10075 3939 10081
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 5902 10112 5908 10124
rect 5863 10084 5908 10112
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 6564 10121 6592 10152
rect 6549 10115 6607 10121
rect 6549 10081 6561 10115
rect 6595 10081 6607 10115
rect 7374 10112 7380 10124
rect 7335 10084 7380 10112
rect 6549 10075 6607 10081
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 8110 10072 8116 10124
rect 8168 10112 8174 10124
rect 8205 10115 8263 10121
rect 8205 10112 8217 10115
rect 8168 10084 8217 10112
rect 8168 10072 8174 10084
rect 8205 10081 8217 10084
rect 8251 10081 8263 10115
rect 8205 10075 8263 10081
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 9122 10112 9128 10124
rect 8352 10084 8397 10112
rect 9083 10084 9128 10112
rect 8352 10072 8358 10084
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10081 9275 10115
rect 9416 10112 9444 10152
rect 9582 10140 9588 10192
rect 9640 10180 9646 10192
rect 9640 10152 10272 10180
rect 9640 10140 9646 10152
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9416 10084 9689 10112
rect 9217 10075 9275 10081
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10112 9827 10115
rect 9950 10112 9956 10124
rect 9815 10084 9956 10112
rect 9815 10081 9827 10084
rect 9769 10075 9827 10081
rect 3786 10044 3792 10056
rect 3699 10016 3792 10044
rect 3786 10004 3792 10016
rect 3844 10044 3850 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 3844 10016 4077 10044
rect 3844 10004 3850 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5224 10016 6009 10044
rect 5224 10004 5230 10016
rect 5997 10013 6009 10016
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10044 6239 10047
rect 6270 10044 6276 10056
rect 6227 10016 6276 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 7466 10044 7472 10056
rect 7427 10016 7472 10044
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 7650 10004 7656 10056
rect 7708 10044 7714 10056
rect 8481 10047 8539 10053
rect 8481 10044 8493 10047
rect 7708 10016 8493 10044
rect 7708 10004 7714 10016
rect 8481 10013 8493 10016
rect 8527 10044 8539 10047
rect 8662 10044 8668 10056
rect 8527 10016 8668 10044
rect 8527 10013 8539 10016
rect 8481 10007 8539 10013
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 5092 9948 6776 9976
rect 3697 9911 3755 9917
rect 3697 9877 3709 9911
rect 3743 9908 3755 9911
rect 5092 9908 5120 9948
rect 3743 9880 5120 9908
rect 3743 9877 3755 9880
rect 3697 9871 3755 9877
rect 5166 9868 5172 9920
rect 5224 9908 5230 9920
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 5224 9880 5457 9908
rect 5224 9868 5230 9880
rect 5445 9877 5457 9880
rect 5491 9877 5503 9911
rect 6748 9908 6776 9948
rect 6822 9936 6828 9988
rect 6880 9976 6886 9988
rect 7926 9976 7932 9988
rect 6880 9948 7932 9976
rect 6880 9936 6886 9948
rect 7926 9936 7932 9948
rect 7984 9936 7990 9988
rect 7834 9908 7840 9920
rect 6748 9880 7840 9908
rect 5445 9871 5503 9877
rect 7834 9868 7840 9880
rect 7892 9908 7898 9920
rect 8386 9908 8392 9920
rect 7892 9880 8392 9908
rect 7892 9868 7898 9880
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 9238 9908 9266 10075
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 10244 10112 10272 10152
rect 10318 10140 10324 10192
rect 10376 10189 10382 10192
rect 10376 10183 10440 10189
rect 10376 10149 10394 10183
rect 10428 10149 10440 10183
rect 10511 10180 10539 10220
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11480 10220 11989 10248
rect 11480 10208 11486 10220
rect 11977 10217 11989 10220
rect 12023 10217 12035 10251
rect 11977 10211 12035 10217
rect 12158 10208 12164 10260
rect 12216 10248 12222 10260
rect 17034 10248 17040 10260
rect 12216 10220 17040 10248
rect 12216 10208 12222 10220
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 17126 10208 17132 10260
rect 17184 10248 17190 10260
rect 17405 10251 17463 10257
rect 17405 10248 17417 10251
rect 17184 10220 17417 10248
rect 17184 10208 17190 10220
rect 17405 10217 17417 10220
rect 17451 10217 17463 10251
rect 17405 10211 17463 10217
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 17552 10220 19288 10248
rect 17552 10208 17558 10220
rect 12069 10183 12127 10189
rect 12069 10180 12081 10183
rect 10511 10152 12081 10180
rect 10376 10143 10440 10149
rect 12069 10149 12081 10152
rect 12115 10149 12127 10183
rect 12986 10180 12992 10192
rect 12069 10143 12127 10149
rect 12176 10152 12992 10180
rect 10376 10140 10382 10143
rect 11790 10112 11796 10124
rect 10244 10084 11796 10112
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9306 9936 9312 9988
rect 9364 9976 9370 9988
rect 9416 9976 9444 10007
rect 9490 10004 9496 10056
rect 9548 10044 9554 10056
rect 12176 10053 12204 10152
rect 12986 10140 12992 10152
rect 13044 10180 13050 10192
rect 13354 10180 13360 10192
rect 13044 10152 13360 10180
rect 13044 10140 13050 10152
rect 13354 10140 13360 10152
rect 13412 10140 13418 10192
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 15654 10180 15660 10192
rect 15344 10152 15660 10180
rect 15344 10140 15350 10152
rect 15654 10140 15660 10152
rect 15712 10180 15718 10192
rect 15749 10183 15807 10189
rect 15749 10180 15761 10183
rect 15712 10152 15761 10180
rect 15712 10140 15718 10152
rect 15749 10149 15761 10152
rect 15795 10149 15807 10183
rect 15749 10143 15807 10149
rect 15933 10183 15991 10189
rect 15933 10149 15945 10183
rect 15979 10180 15991 10183
rect 15979 10152 17540 10180
rect 15979 10149 15991 10152
rect 15933 10143 15991 10149
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 12437 10115 12495 10121
rect 12437 10112 12449 10115
rect 12400 10084 12449 10112
rect 12400 10072 12406 10084
rect 12437 10081 12449 10084
rect 12483 10081 12495 10115
rect 12437 10075 12495 10081
rect 12710 10072 12716 10124
rect 12768 10112 12774 10124
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 12768 10084 12909 10112
rect 12768 10072 12774 10084
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 14056 10084 14749 10112
rect 14056 10072 14062 10084
rect 14737 10081 14749 10084
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 15470 10072 15476 10124
rect 15528 10112 15534 10124
rect 15565 10115 15623 10121
rect 15565 10112 15577 10115
rect 15528 10084 15577 10112
rect 15528 10072 15534 10084
rect 15565 10081 15577 10084
rect 15611 10081 15623 10115
rect 15565 10075 15623 10081
rect 16292 10115 16350 10121
rect 16292 10081 16304 10115
rect 16338 10112 16350 10115
rect 16758 10112 16764 10124
rect 16338 10084 16764 10112
rect 16338 10081 16350 10084
rect 16292 10075 16350 10081
rect 16758 10072 16764 10084
rect 16816 10072 16822 10124
rect 17512 10121 17540 10152
rect 17770 10140 17776 10192
rect 17828 10180 17834 10192
rect 19260 10180 19288 10220
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 20257 10251 20315 10257
rect 20257 10248 20269 10251
rect 19576 10220 20269 10248
rect 19576 10208 19582 10220
rect 20257 10217 20269 10220
rect 20303 10217 20315 10251
rect 20257 10211 20315 10217
rect 17828 10152 18000 10180
rect 19260 10152 20300 10180
rect 17828 10140 17834 10152
rect 17972 10124 18000 10152
rect 20272 10124 20300 10152
rect 17497 10115 17555 10121
rect 17497 10081 17509 10115
rect 17543 10081 17555 10115
rect 17865 10115 17923 10121
rect 17865 10112 17877 10115
rect 17497 10075 17555 10081
rect 17604 10084 17877 10112
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9548 10016 10149 10044
rect 9548 10004 9554 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 12802 10004 12808 10056
rect 12860 10044 12866 10056
rect 13630 10044 13636 10056
rect 12860 10016 13636 10044
rect 12860 10004 12866 10016
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 15286 10044 15292 10056
rect 15247 10016 15292 10044
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 16025 10047 16083 10053
rect 16025 10044 16037 10047
rect 15436 10016 16037 10044
rect 15436 10004 15442 10016
rect 16025 10013 16037 10016
rect 16071 10013 16083 10047
rect 16025 10007 16083 10013
rect 9364 9948 9444 9976
rect 9677 9979 9735 9985
rect 9364 9936 9370 9948
rect 9677 9945 9689 9979
rect 9723 9976 9735 9979
rect 9953 9979 10011 9985
rect 9953 9976 9965 9979
rect 9723 9948 9965 9976
rect 9723 9945 9735 9948
rect 9677 9939 9735 9945
rect 9953 9945 9965 9948
rect 9999 9945 10011 9979
rect 11514 9976 11520 9988
rect 11475 9948 11520 9976
rect 9953 9939 10011 9945
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 12526 9936 12532 9988
rect 12584 9976 12590 9988
rect 12621 9979 12679 9985
rect 12621 9976 12633 9979
rect 12584 9948 12633 9976
rect 12584 9936 12590 9948
rect 12621 9945 12633 9948
rect 12667 9945 12679 9979
rect 12621 9939 12679 9945
rect 13170 9936 13176 9988
rect 13228 9976 13234 9988
rect 14921 9979 14979 9985
rect 14921 9976 14933 9979
rect 13228 9948 14933 9976
rect 13228 9936 13234 9948
rect 14921 9945 14933 9948
rect 14967 9945 14979 9979
rect 14921 9939 14979 9945
rect 11422 9908 11428 9920
rect 9238 9880 11428 9908
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 11609 9911 11667 9917
rect 11609 9877 11621 9911
rect 11655 9908 11667 9911
rect 12986 9908 12992 9920
rect 11655 9880 12992 9908
rect 11655 9877 11667 9880
rect 11609 9871 11667 9877
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 13538 9868 13544 9920
rect 13596 9908 13602 9920
rect 14185 9911 14243 9917
rect 14185 9908 14197 9911
rect 13596 9880 14197 9908
rect 13596 9868 13602 9880
rect 14185 9877 14197 9880
rect 14231 9877 14243 9911
rect 14185 9871 14243 9877
rect 15102 9868 15108 9920
rect 15160 9908 15166 9920
rect 15930 9908 15936 9920
rect 15160 9880 15936 9908
rect 15160 9868 15166 9880
rect 15930 9868 15936 9880
rect 15988 9868 15994 9920
rect 16040 9908 16068 10007
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 17604 10044 17632 10084
rect 17865 10081 17877 10084
rect 17911 10081 17923 10115
rect 17865 10075 17923 10081
rect 17954 10072 17960 10124
rect 18012 10072 18018 10124
rect 18874 10072 18880 10124
rect 18932 10112 18938 10124
rect 20165 10115 20223 10121
rect 20165 10112 20177 10115
rect 18932 10084 20177 10112
rect 18932 10072 18938 10084
rect 20165 10081 20177 10084
rect 20211 10081 20223 10115
rect 20165 10075 20223 10081
rect 20254 10072 20260 10124
rect 20312 10072 20318 10124
rect 17092 10016 17632 10044
rect 17092 10004 17098 10016
rect 18046 10004 18052 10056
rect 18104 10044 18110 10056
rect 18414 10053 18420 10056
rect 18188 10047 18246 10053
rect 18188 10044 18200 10047
rect 18104 10016 18200 10044
rect 18104 10004 18110 10016
rect 18188 10013 18200 10016
rect 18234 10013 18246 10047
rect 18188 10007 18246 10013
rect 18371 10047 18420 10053
rect 18371 10013 18383 10047
rect 18417 10013 18420 10047
rect 18371 10007 18420 10013
rect 18414 10004 18420 10007
rect 18472 10004 18478 10056
rect 18598 10044 18604 10056
rect 18559 10016 18604 10044
rect 18598 10004 18604 10016
rect 18656 10004 18662 10056
rect 18690 10004 18696 10056
rect 18748 10044 18754 10056
rect 20349 10047 20407 10053
rect 20349 10044 20361 10047
rect 18748 10016 20361 10044
rect 18748 10004 18754 10016
rect 20349 10013 20361 10016
rect 20395 10013 20407 10047
rect 20349 10007 20407 10013
rect 19978 9976 19984 9988
rect 19260 9948 19984 9976
rect 17218 9908 17224 9920
rect 16040 9880 17224 9908
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 17681 9911 17739 9917
rect 17681 9877 17693 9911
rect 17727 9908 17739 9911
rect 17770 9908 17776 9920
rect 17727 9880 17776 9908
rect 17727 9877 17739 9880
rect 17681 9871 17739 9877
rect 17770 9868 17776 9880
rect 17828 9868 17834 9920
rect 18598 9868 18604 9920
rect 18656 9908 18662 9920
rect 19260 9908 19288 9948
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 19702 9908 19708 9920
rect 18656 9880 19288 9908
rect 19663 9880 19708 9908
rect 18656 9868 18662 9880
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 19797 9911 19855 9917
rect 19797 9877 19809 9911
rect 19843 9908 19855 9911
rect 20254 9908 20260 9920
rect 19843 9880 20260 9908
rect 19843 9877 19855 9880
rect 19797 9871 19855 9877
rect 20254 9868 20260 9880
rect 20312 9868 20318 9920
rect 1104 9818 20884 9840
rect 1104 9766 4280 9818
rect 4332 9766 4344 9818
rect 4396 9766 4408 9818
rect 4460 9766 4472 9818
rect 4524 9766 10878 9818
rect 10930 9766 10942 9818
rect 10994 9766 11006 9818
rect 11058 9766 11070 9818
rect 11122 9766 17475 9818
rect 17527 9766 17539 9818
rect 17591 9766 17603 9818
rect 17655 9766 17667 9818
rect 17719 9766 20884 9818
rect 1104 9744 20884 9766
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6052 9676 6837 9704
rect 6052 9664 6058 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 6825 9667 6883 9673
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 8754 9704 8760 9716
rect 7064 9676 8760 9704
rect 7064 9664 7070 9676
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 10689 9707 10747 9713
rect 10689 9704 10701 9707
rect 8904 9676 10701 9704
rect 8904 9664 8910 9676
rect 10689 9673 10701 9676
rect 10735 9673 10747 9707
rect 10689 9667 10747 9673
rect 11422 9664 11428 9716
rect 11480 9704 11486 9716
rect 12253 9707 12311 9713
rect 12253 9704 12265 9707
rect 11480 9676 12265 9704
rect 11480 9664 11486 9676
rect 12253 9673 12265 9676
rect 12299 9673 12311 9707
rect 12253 9667 12311 9673
rect 12342 9664 12348 9716
rect 12400 9704 12406 9716
rect 15102 9704 15108 9716
rect 12400 9676 14964 9704
rect 15063 9676 15108 9704
rect 12400 9664 12406 9676
rect 1765 9639 1823 9645
rect 1765 9605 1777 9639
rect 1811 9636 1823 9639
rect 1854 9636 1860 9648
rect 1811 9608 1860 9636
rect 1811 9605 1823 9608
rect 1765 9599 1823 9605
rect 1854 9596 1860 9608
rect 1912 9596 1918 9648
rect 2958 9636 2964 9648
rect 2919 9608 2964 9636
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 6641 9639 6699 9645
rect 6641 9605 6653 9639
rect 6687 9636 6699 9639
rect 6914 9636 6920 9648
rect 6687 9608 6920 9636
rect 6687 9605 6699 9608
rect 6641 9599 6699 9605
rect 6914 9596 6920 9608
rect 6972 9636 6978 9648
rect 7466 9636 7472 9648
rect 6972 9608 7472 9636
rect 6972 9596 6978 9608
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 9214 9636 9220 9648
rect 9175 9608 9220 9636
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 11882 9596 11888 9648
rect 11940 9596 11946 9648
rect 12158 9596 12164 9648
rect 12216 9636 12222 9648
rect 13449 9639 13507 9645
rect 13449 9636 13461 9639
rect 12216 9608 13461 9636
rect 12216 9596 12222 9608
rect 13449 9605 13461 9608
rect 13495 9605 13507 9639
rect 14936 9636 14964 9676
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 17862 9704 17868 9716
rect 15212 9676 17868 9704
rect 15212 9636 15240 9676
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 17678 9636 17684 9648
rect 14936 9608 15240 9636
rect 17236 9608 17684 9636
rect 13449 9599 13507 9605
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9537 2467 9571
rect 2409 9531 2467 9537
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 3651 9540 3924 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9500 2191 9503
rect 2424 9500 2452 9531
rect 3326 9500 3332 9512
rect 2179 9472 2360 9500
rect 2424 9472 3332 9500
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 2222 9432 2228 9444
rect 2183 9404 2228 9432
rect 2222 9392 2228 9404
rect 2280 9392 2286 9444
rect 2332 9432 2360 9472
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 3786 9500 3792 9512
rect 3747 9472 3792 9500
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 3896 9432 3924 9540
rect 4982 9528 4988 9580
rect 5040 9568 5046 9580
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 5040 9540 5273 9568
rect 5040 9528 5046 9540
rect 5261 9537 5273 9540
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 6328 9540 7389 9568
rect 6328 9528 6334 9540
rect 7377 9537 7389 9540
rect 7423 9568 7435 9571
rect 7650 9568 7656 9580
rect 7423 9540 7656 9568
rect 7423 9537 7435 9540
rect 7377 9531 7435 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7834 9568 7840 9580
rect 7795 9540 7840 9568
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 9232 9568 9260 9596
rect 9232 9540 9444 9568
rect 4056 9503 4114 9509
rect 4056 9469 4068 9503
rect 4102 9500 4114 9503
rect 5166 9500 5172 9512
rect 4102 9472 5172 9500
rect 4102 9469 4114 9472
rect 4056 9463 4114 9469
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 9309 9503 9367 9509
rect 5460 9472 7420 9500
rect 5460 9432 5488 9472
rect 2332 9404 3648 9432
rect 3896 9404 5488 9432
rect 5528 9435 5586 9441
rect 2869 9367 2927 9373
rect 2869 9333 2881 9367
rect 2915 9364 2927 9367
rect 3326 9364 3332 9376
rect 2915 9336 3332 9364
rect 2915 9333 2927 9336
rect 2869 9327 2927 9333
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3620 9364 3648 9404
rect 5528 9401 5540 9435
rect 5574 9432 5586 9435
rect 6270 9432 6276 9444
rect 5574 9404 6276 9432
rect 5574 9401 5586 9404
rect 5528 9395 5586 9401
rect 6270 9392 6276 9404
rect 6328 9432 6334 9444
rect 7193 9435 7251 9441
rect 7193 9432 7205 9435
rect 6328 9404 7205 9432
rect 6328 9392 6334 9404
rect 7193 9401 7205 9404
rect 7239 9401 7251 9435
rect 7193 9395 7251 9401
rect 5074 9364 5080 9376
rect 3476 9336 3521 9364
rect 3620 9336 5080 9364
rect 3476 9324 3482 9336
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5902 9364 5908 9376
rect 5215 9336 5908 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 6052 9336 7297 9364
rect 6052 9324 6058 9336
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7392 9364 7420 9472
rect 9309 9469 9321 9503
rect 9355 9469 9367 9503
rect 9416 9500 9444 9540
rect 9565 9503 9623 9509
rect 9565 9500 9577 9503
rect 9416 9472 9577 9500
rect 9309 9463 9367 9469
rect 9565 9469 9577 9472
rect 9611 9469 9623 9503
rect 9565 9463 9623 9469
rect 8110 9441 8116 9444
rect 8104 9432 8116 9441
rect 8071 9404 8116 9432
rect 8104 9395 8116 9404
rect 8110 9392 8116 9395
rect 8168 9392 8174 9444
rect 8478 9392 8484 9444
rect 8536 9432 8542 9444
rect 9324 9432 9352 9463
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 10781 9503 10839 9509
rect 10781 9500 10793 9503
rect 10744 9472 10793 9500
rect 10744 9460 10750 9472
rect 10781 9469 10793 9472
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 11330 9460 11336 9512
rect 11388 9500 11394 9512
rect 11900 9500 11928 9596
rect 17236 9580 17264 9608
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 18414 9636 18420 9648
rect 18375 9608 18420 9636
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 13081 9571 13139 9577
rect 12268 9540 12940 9568
rect 12158 9500 12164 9512
rect 11388 9472 12164 9500
rect 11388 9460 11394 9472
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 9398 9432 9404 9444
rect 8536 9404 9404 9432
rect 8536 9392 8542 9404
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 11048 9435 11106 9441
rect 11048 9432 11060 9435
rect 9732 9404 11060 9432
rect 9732 9392 9738 9404
rect 11048 9401 11060 9404
rect 11094 9432 11106 9435
rect 12268 9432 12296 9540
rect 12345 9503 12403 9509
rect 12345 9469 12357 9503
rect 12391 9500 12403 9503
rect 12618 9500 12624 9512
rect 12391 9472 12624 9500
rect 12391 9469 12403 9472
rect 12345 9463 12403 9469
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 12802 9460 12808 9512
rect 12860 9460 12866 9512
rect 12912 9500 12940 9540
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13354 9568 13360 9580
rect 13127 9540 13360 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 15102 9528 15108 9580
rect 15160 9568 15166 9580
rect 15378 9568 15384 9580
rect 15160 9540 15384 9568
rect 15160 9528 15166 9540
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 17218 9568 17224 9580
rect 16540 9540 17224 9568
rect 16540 9528 16546 9540
rect 17218 9528 17224 9540
rect 17276 9528 17282 9580
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9568 17555 9571
rect 17770 9568 17776 9580
rect 17543 9540 17776 9568
rect 17543 9537 17555 9540
rect 17497 9531 17555 9537
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 18506 9528 18512 9580
rect 18564 9568 18570 9580
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 18564 9540 18613 9568
rect 18564 9528 18570 9540
rect 18601 9537 18613 9540
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 13170 9500 13176 9512
rect 12912 9472 13176 9500
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 13262 9460 13268 9512
rect 13320 9500 13326 9512
rect 13320 9472 13365 9500
rect 13320 9460 13326 9472
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 13725 9503 13783 9509
rect 13725 9500 13737 9503
rect 13596 9472 13737 9500
rect 13596 9460 13602 9472
rect 13725 9469 13737 9472
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 13992 9503 14050 9509
rect 13992 9469 14004 9503
rect 14038 9500 14050 9503
rect 14458 9500 14464 9512
rect 14038 9472 14464 9500
rect 14038 9469 14050 9472
rect 13992 9463 14050 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 15654 9509 15660 9512
rect 15648 9500 15660 9509
rect 15615 9472 15660 9500
rect 15648 9463 15660 9472
rect 15654 9460 15660 9463
rect 15712 9460 15718 9512
rect 16850 9500 16856 9512
rect 15764 9472 16856 9500
rect 11094 9404 12296 9432
rect 12820 9432 12848 9460
rect 12897 9435 12955 9441
rect 12897 9432 12909 9435
rect 12820 9404 12909 9432
rect 11094 9401 11106 9404
rect 11048 9395 11106 9401
rect 12897 9401 12909 9404
rect 12943 9401 12955 9435
rect 12897 9395 12955 9401
rect 14550 9392 14556 9444
rect 14608 9432 14614 9444
rect 15764 9432 15792 9472
rect 16850 9460 16856 9472
rect 16908 9460 16914 9512
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 17865 9503 17923 9509
rect 17865 9500 17877 9503
rect 17000 9472 17877 9500
rect 17000 9460 17006 9472
rect 17865 9469 17877 9472
rect 17911 9469 17923 9503
rect 18230 9500 18236 9512
rect 18191 9472 18236 9500
rect 17865 9463 17923 9469
rect 18230 9460 18236 9472
rect 18288 9460 18294 9512
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 20073 9503 20131 9509
rect 20073 9500 20085 9503
rect 19300 9472 20085 9500
rect 19300 9460 19306 9472
rect 20073 9469 20085 9472
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 16666 9432 16672 9444
rect 14608 9404 15792 9432
rect 15856 9404 16672 9432
rect 14608 9392 14614 9404
rect 10778 9364 10784 9376
rect 7392 9336 10784 9364
rect 7285 9327 7343 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 11790 9364 11796 9376
rect 10928 9336 11796 9364
rect 10928 9324 10934 9336
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12158 9364 12164 9376
rect 12119 9336 12164 9364
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12250 9324 12256 9376
rect 12308 9364 12314 9376
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 12308 9336 12449 9364
rect 12308 9324 12314 9336
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12437 9327 12495 9333
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 12860 9336 12905 9364
rect 12860 9324 12866 9336
rect 15194 9324 15200 9376
rect 15252 9364 15258 9376
rect 15856 9364 15884 9404
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 18138 9432 18144 9444
rect 16776 9404 18144 9432
rect 16776 9376 16804 9404
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18598 9432 18604 9444
rect 18248 9404 18604 9432
rect 16758 9364 16764 9376
rect 15252 9336 15884 9364
rect 16671 9336 16764 9364
rect 15252 9324 15258 9336
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 17218 9364 17224 9376
rect 16908 9336 16953 9364
rect 17179 9336 17224 9364
rect 16908 9324 16914 9336
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 17313 9367 17371 9373
rect 17313 9333 17325 9367
rect 17359 9364 17371 9367
rect 17402 9364 17408 9376
rect 17359 9336 17408 9364
rect 17359 9333 17371 9336
rect 17313 9327 17371 9333
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 17681 9367 17739 9373
rect 17681 9333 17693 9367
rect 17727 9364 17739 9367
rect 18248 9364 18276 9404
rect 18598 9392 18604 9404
rect 18656 9392 18662 9444
rect 18782 9392 18788 9444
rect 18840 9441 18846 9444
rect 18840 9435 18904 9441
rect 18840 9401 18858 9435
rect 18892 9432 18904 9435
rect 19150 9432 19156 9444
rect 18892 9404 19156 9432
rect 18892 9401 18904 9404
rect 18840 9395 18904 9401
rect 18840 9392 18846 9395
rect 19150 9392 19156 9404
rect 19208 9392 19214 9444
rect 19260 9404 20300 9432
rect 17727 9336 18276 9364
rect 17727 9333 17739 9336
rect 17681 9327 17739 9333
rect 18690 9324 18696 9376
rect 18748 9364 18754 9376
rect 19260 9364 19288 9404
rect 18748 9336 19288 9364
rect 18748 9324 18754 9336
rect 19426 9324 19432 9376
rect 19484 9364 19490 9376
rect 20272 9373 20300 9404
rect 19981 9367 20039 9373
rect 19981 9364 19993 9367
rect 19484 9336 19993 9364
rect 19484 9324 19490 9336
rect 19981 9333 19993 9336
rect 20027 9333 20039 9367
rect 19981 9327 20039 9333
rect 20257 9367 20315 9373
rect 20257 9333 20269 9367
rect 20303 9333 20315 9367
rect 20257 9327 20315 9333
rect 1104 9274 20884 9296
rect 1104 9222 7579 9274
rect 7631 9222 7643 9274
rect 7695 9222 7707 9274
rect 7759 9222 7771 9274
rect 7823 9222 14176 9274
rect 14228 9222 14240 9274
rect 14292 9222 14304 9274
rect 14356 9222 14368 9274
rect 14420 9222 20884 9274
rect 1104 9200 20884 9222
rect 2682 9160 2688 9172
rect 2643 9132 2688 9160
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3844 9132 4077 9160
rect 3844 9120 3850 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 3605 9095 3663 9101
rect 3605 9061 3617 9095
rect 3651 9092 3663 9095
rect 3970 9092 3976 9104
rect 3651 9064 3976 9092
rect 3651 9061 3663 9064
rect 3605 9055 3663 9061
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 4080 9092 4108 9123
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 5350 9160 5356 9172
rect 4304 9132 5356 9160
rect 4304 9120 4310 9132
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 5721 9163 5779 9169
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 5994 9160 6000 9172
rect 5767 9132 6000 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9160 7251 9163
rect 7374 9160 7380 9172
rect 7239 9132 7380 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 8018 9160 8024 9172
rect 7484 9132 8024 9160
rect 4608 9095 4666 9101
rect 4080 9064 4384 9092
rect 2777 9027 2835 9033
rect 2777 8993 2789 9027
rect 2823 9024 2835 9027
rect 2958 9024 2964 9036
rect 2823 8996 2964 9024
rect 2823 8993 2835 8996
rect 2777 8987 2835 8993
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 3513 9027 3571 9033
rect 3513 8993 3525 9027
rect 3559 9024 3571 9027
rect 3559 8996 3740 9024
rect 3559 8993 3571 8996
rect 3513 8987 3571 8993
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 2682 8848 2688 8900
rect 2740 8888 2746 8900
rect 2884 8888 2912 8919
rect 2740 8860 2912 8888
rect 3712 8888 3740 8996
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4356 9033 4384 9064
rect 4608 9061 4620 9095
rect 4654 9092 4666 9095
rect 5902 9092 5908 9104
rect 4654 9064 5908 9092
rect 4654 9061 4666 9064
rect 4608 9055 4666 9061
rect 5902 9052 5908 9064
rect 5960 9052 5966 9104
rect 6080 9095 6138 9101
rect 6080 9061 6092 9095
rect 6126 9092 6138 9095
rect 6914 9092 6920 9104
rect 6126 9064 6920 9092
rect 6126 9061 6138 9064
rect 6080 9055 6138 9061
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 7006 9052 7012 9104
rect 7064 9092 7070 9104
rect 7484 9092 7512 9132
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8110 9120 8116 9172
rect 8168 9160 8174 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8168 9132 8677 9160
rect 8168 9120 8174 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 9858 9160 9864 9172
rect 8665 9123 8723 9129
rect 8772 9132 9864 9160
rect 7064 9064 7512 9092
rect 7552 9095 7610 9101
rect 7064 9052 7070 9064
rect 7552 9061 7564 9095
rect 7598 9092 7610 9095
rect 8202 9092 8208 9104
rect 7598 9064 8208 9092
rect 7598 9061 7610 9064
rect 7552 9055 7610 9061
rect 8202 9052 8208 9064
rect 8260 9052 8266 9104
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 4212 8996 4261 9024
rect 4212 8984 4218 8996
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 9024 4399 9027
rect 4982 9024 4988 9036
rect 4387 8996 4988 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 4982 8984 4988 8996
rect 5040 9024 5046 9036
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5040 8996 5825 9024
rect 5040 8984 5046 8996
rect 5813 8993 5825 8996
rect 5859 9024 5871 9027
rect 7285 9027 7343 9033
rect 7285 9024 7297 9027
rect 5859 8996 7297 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 6932 8968 6960 8996
rect 7285 8993 7297 8996
rect 7331 8993 7343 9027
rect 7285 8987 7343 8993
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 8772 9024 8800 9132
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 12434 9160 12440 9172
rect 10428 9132 11652 9160
rect 12395 9132 12440 9160
rect 10042 9092 10048 9104
rect 7892 8996 8800 9024
rect 8864 9064 10048 9092
rect 7892 8984 7898 8996
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8956 3847 8959
rect 3835 8928 4384 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 4246 8888 4252 8900
rect 3712 8860 4252 8888
rect 2740 8848 2746 8860
rect 4246 8848 4252 8860
rect 4304 8848 4310 8900
rect 2317 8823 2375 8829
rect 2317 8789 2329 8823
rect 2363 8820 2375 8823
rect 2866 8820 2872 8832
rect 2363 8792 2872 8820
rect 2363 8789 2375 8792
rect 2317 8783 2375 8789
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 3145 8823 3203 8829
rect 3145 8789 3157 8823
rect 3191 8820 3203 8823
rect 3970 8820 3976 8832
rect 3191 8792 3976 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 4356 8820 4384 8928
rect 6914 8916 6920 8968
rect 6972 8916 6978 8968
rect 8864 8888 8892 9064
rect 10042 9052 10048 9064
rect 10100 9052 10106 9104
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 9024 9183 9027
rect 9677 9027 9735 9033
rect 9171 8996 9628 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 8220 8860 8892 8888
rect 9232 8888 9260 8919
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 9600 8956 9628 8996
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 10428 9024 10456 9132
rect 10689 9095 10747 9101
rect 10689 9061 10701 9095
rect 10735 9092 10747 9095
rect 11624 9092 11652 9132
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 12544 9132 12940 9160
rect 12544 9092 12572 9132
rect 10735 9064 11560 9092
rect 11624 9064 12572 9092
rect 10735 9061 10747 9064
rect 10689 9055 10747 9061
rect 9723 8996 10456 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 11330 9033 11336 9036
rect 10597 9027 10655 9033
rect 10597 9024 10609 9027
rect 10560 8996 10609 9024
rect 10560 8984 10566 8996
rect 10597 8993 10609 8996
rect 10643 8993 10655 9027
rect 11057 9027 11115 9033
rect 11057 9024 11069 9027
rect 10597 8987 10655 8993
rect 10704 8996 11069 9024
rect 10704 8968 10732 8996
rect 11057 8993 11069 8996
rect 11103 8993 11115 9027
rect 11324 9024 11336 9033
rect 11291 8996 11336 9024
rect 11057 8987 11115 8993
rect 11324 8987 11336 8996
rect 11330 8984 11336 8987
rect 11388 8984 11394 9036
rect 11532 9024 11560 9064
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 12774 9095 12832 9101
rect 12774 9092 12786 9095
rect 12676 9064 12786 9092
rect 12676 9052 12682 9064
rect 12774 9061 12786 9064
rect 12820 9061 12832 9095
rect 12912 9092 12940 9132
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 13909 9163 13967 9169
rect 13909 9160 13921 9163
rect 13228 9132 13921 9160
rect 13228 9120 13234 9132
rect 13909 9129 13921 9132
rect 13955 9129 13967 9163
rect 13909 9123 13967 9129
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9160 14243 9163
rect 17957 9163 18015 9169
rect 17957 9160 17969 9163
rect 14231 9132 17969 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 17957 9129 17969 9132
rect 18003 9129 18015 9163
rect 17957 9123 18015 9129
rect 18049 9163 18107 9169
rect 18049 9129 18061 9163
rect 18095 9160 18107 9163
rect 18601 9163 18659 9169
rect 18601 9160 18613 9163
rect 18095 9132 18613 9160
rect 18095 9129 18107 9132
rect 18049 9123 18107 9129
rect 18601 9129 18613 9132
rect 18647 9129 18659 9163
rect 18601 9123 18659 9129
rect 15556 9095 15614 9101
rect 12912 9064 13952 9092
rect 12774 9055 12832 9061
rect 13078 9024 13084 9036
rect 11532 8996 13084 9024
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 10410 8956 10416 8968
rect 9364 8928 9409 8956
rect 9600 8928 10416 8956
rect 9364 8916 9370 8928
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10686 8916 10692 8968
rect 10744 8916 10750 8968
rect 10870 8956 10876 8968
rect 10831 8928 10876 8956
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 12250 8916 12256 8968
rect 12308 8956 12314 8968
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 12308 8928 12541 8956
rect 12308 8916 12314 8928
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 13924 8956 13952 9064
rect 14016 9064 15516 9092
rect 14016 9033 14044 9064
rect 14001 9027 14059 9033
rect 14001 8993 14013 9027
rect 14047 8993 14059 9027
rect 14734 9024 14740 9036
rect 14695 8996 14740 9024
rect 14001 8987 14059 8993
rect 14734 8984 14740 8996
rect 14792 8984 14798 9036
rect 14829 9027 14887 9033
rect 14829 8993 14841 9027
rect 14875 9024 14887 9027
rect 15378 9024 15384 9036
rect 14875 8996 15384 9024
rect 14875 8993 14887 8996
rect 14829 8987 14887 8993
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 15488 9024 15516 9064
rect 15556 9061 15568 9095
rect 15602 9092 15614 9095
rect 16758 9092 16764 9104
rect 15602 9064 16764 9092
rect 15602 9061 15614 9064
rect 15556 9055 15614 9061
rect 16758 9052 16764 9064
rect 16816 9052 16822 9104
rect 16850 9052 16856 9104
rect 16908 9092 16914 9104
rect 20530 9092 20536 9104
rect 16908 9064 18460 9092
rect 16908 9052 16914 9064
rect 17126 9024 17132 9036
rect 15488 8996 16344 9024
rect 17087 8996 17132 9024
rect 15010 8956 15016 8968
rect 13924 8928 14596 8956
rect 14971 8928 15016 8956
rect 12529 8919 12587 8925
rect 10042 8888 10048 8900
rect 9232 8860 10048 8888
rect 4614 8820 4620 8832
rect 4356 8792 4620 8820
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 8220 8820 8248 8860
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 14568 8888 14596 8928
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 15160 8928 15301 8956
rect 15160 8916 15166 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 15194 8888 15200 8900
rect 13464 8860 14504 8888
rect 14568 8860 15200 8888
rect 4764 8792 8248 8820
rect 8757 8823 8815 8829
rect 4764 8780 4770 8792
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 9766 8820 9772 8832
rect 8803 8792 9772 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 9861 8823 9919 8829
rect 9861 8789 9873 8823
rect 9907 8820 9919 8823
rect 9950 8820 9956 8832
rect 9907 8792 9956 8820
rect 9907 8789 9919 8792
rect 9861 8783 9919 8789
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 10229 8823 10287 8829
rect 10229 8789 10241 8823
rect 10275 8820 10287 8823
rect 12342 8820 12348 8832
rect 10275 8792 12348 8820
rect 10275 8789 10287 8792
rect 10229 8783 10287 8789
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 13464 8820 13492 8860
rect 14366 8820 14372 8832
rect 12584 8792 13492 8820
rect 14327 8792 14372 8820
rect 12584 8780 12590 8792
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 14476 8820 14504 8860
rect 15194 8848 15200 8860
rect 15252 8848 15258 8900
rect 16316 8888 16344 8996
rect 17126 8984 17132 8996
rect 17184 8984 17190 9036
rect 18432 9033 18460 9064
rect 18800 9064 20536 9092
rect 18800 9033 18828 9064
rect 20530 9052 20536 9064
rect 20588 9052 20594 9104
rect 19426 9033 19432 9036
rect 18417 9027 18475 9033
rect 18417 8993 18429 9027
rect 18463 8993 18475 9027
rect 18417 8987 18475 8993
rect 18785 9027 18843 9033
rect 18785 8993 18797 9027
rect 18831 8993 18843 9027
rect 19420 9024 19432 9033
rect 19387 8996 19432 9024
rect 18785 8987 18843 8993
rect 19420 8987 19432 8996
rect 19426 8984 19432 8987
rect 19484 8984 19490 9036
rect 16850 8916 16856 8968
rect 16908 8956 16914 8968
rect 17221 8959 17279 8965
rect 17221 8956 17233 8959
rect 16908 8928 17233 8956
rect 16908 8916 16914 8928
rect 17221 8925 17233 8928
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 18138 8956 18144 8968
rect 17368 8928 17413 8956
rect 18099 8928 18144 8956
rect 17368 8916 17374 8928
rect 18138 8916 18144 8928
rect 18196 8916 18202 8968
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 19153 8959 19211 8965
rect 19153 8956 19165 8959
rect 18564 8928 19165 8956
rect 18564 8916 18570 8928
rect 19153 8925 19165 8928
rect 19199 8925 19211 8959
rect 19153 8919 19211 8925
rect 16761 8891 16819 8897
rect 16761 8888 16773 8891
rect 16316 8860 16773 8888
rect 16761 8857 16773 8860
rect 16807 8888 16819 8891
rect 17402 8888 17408 8900
rect 16807 8860 17408 8888
rect 16807 8857 16819 8860
rect 16761 8851 16819 8857
rect 17402 8848 17408 8860
rect 17460 8848 17466 8900
rect 17494 8848 17500 8900
rect 17552 8888 17558 8900
rect 18414 8888 18420 8900
rect 17552 8860 18420 8888
rect 17552 8848 17558 8860
rect 18414 8848 18420 8860
rect 18472 8848 18478 8900
rect 15930 8820 15936 8832
rect 14476 8792 15936 8820
rect 15930 8780 15936 8792
rect 15988 8780 15994 8832
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 16080 8792 16681 8820
rect 16080 8780 16086 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16669 8783 16727 8789
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 17589 8823 17647 8829
rect 17589 8820 17601 8823
rect 17368 8792 17601 8820
rect 17368 8780 17374 8792
rect 17589 8789 17601 8792
rect 17635 8789 17647 8823
rect 17589 8783 17647 8789
rect 18138 8780 18144 8832
rect 18196 8820 18202 8832
rect 18969 8823 19027 8829
rect 18969 8820 18981 8823
rect 18196 8792 18981 8820
rect 18196 8780 18202 8792
rect 18969 8789 18981 8792
rect 19015 8789 19027 8823
rect 18969 8783 19027 8789
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 20533 8823 20591 8829
rect 20533 8820 20545 8823
rect 19576 8792 20545 8820
rect 19576 8780 19582 8792
rect 20533 8789 20545 8792
rect 20579 8789 20591 8823
rect 20533 8783 20591 8789
rect 1104 8730 20884 8752
rect 1104 8678 4280 8730
rect 4332 8678 4344 8730
rect 4396 8678 4408 8730
rect 4460 8678 4472 8730
rect 4524 8678 10878 8730
rect 10930 8678 10942 8730
rect 10994 8678 11006 8730
rect 11058 8678 11070 8730
rect 11122 8678 17475 8730
rect 17527 8678 17539 8730
rect 17591 8678 17603 8730
rect 17655 8678 17667 8730
rect 17719 8678 20884 8730
rect 1104 8656 20884 8678
rect 2406 8616 2412 8628
rect 2367 8588 2412 8616
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 3936 8588 4077 8616
rect 3936 8576 3942 8588
rect 4065 8585 4077 8588
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 4614 8576 4620 8628
rect 4672 8616 4678 8628
rect 6270 8616 6276 8628
rect 4672 8588 5856 8616
rect 6231 8588 6276 8616
rect 4672 8576 4678 8588
rect 3237 8551 3295 8557
rect 3237 8517 3249 8551
rect 3283 8548 3295 8551
rect 4890 8548 4896 8560
rect 3283 8520 4896 8548
rect 3283 8517 3295 8520
rect 3237 8511 3295 8517
rect 4890 8508 4896 8520
rect 4948 8508 4954 8560
rect 5828 8548 5856 8588
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 7834 8616 7840 8628
rect 6380 8588 7840 8616
rect 6380 8548 6408 8588
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8202 8576 8208 8628
rect 8260 8616 8266 8628
rect 8297 8619 8355 8625
rect 8297 8616 8309 8619
rect 8260 8588 8309 8616
rect 8260 8576 8266 8588
rect 8297 8585 8309 8588
rect 8343 8585 8355 8619
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 8297 8579 8355 8585
rect 8404 8588 10057 8616
rect 5828 8520 6408 8548
rect 6454 8508 6460 8560
rect 6512 8548 6518 8560
rect 6512 8520 6557 8548
rect 6512 8508 6518 8520
rect 2866 8480 2872 8492
rect 2827 8452 2872 8480
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3050 8480 3056 8492
rect 3011 8452 3056 8480
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 3878 8480 3884 8492
rect 3839 8452 3884 8480
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 3970 8440 3976 8492
rect 4028 8480 4034 8492
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 4028 8452 4537 8480
rect 4028 8440 4034 8452
rect 4525 8449 4537 8452
rect 4571 8449 4583 8483
rect 4706 8480 4712 8492
rect 4667 8452 4712 8480
rect 4525 8443 4583 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 3697 8415 3755 8421
rect 2832 8384 2877 8412
rect 2832 8372 2838 8384
rect 3697 8381 3709 8415
rect 3743 8412 3755 8415
rect 4062 8412 4068 8424
rect 3743 8384 4068 8412
rect 3743 8381 3755 8384
rect 3697 8375 3755 8381
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4798 8412 4804 8424
rect 4479 8384 4804 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8412 4951 8415
rect 4982 8412 4988 8424
rect 4939 8384 4988 8412
rect 4939 8381 4951 8384
rect 4893 8375 4951 8381
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 5160 8415 5218 8421
rect 5160 8381 5172 8415
rect 5206 8412 5218 8415
rect 5994 8412 6000 8424
rect 5206 8384 6000 8412
rect 5206 8381 5218 8384
rect 5160 8375 5218 8381
rect 5994 8372 6000 8384
rect 6052 8372 6058 8424
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 6420 8384 6653 8412
rect 6420 8372 6426 8384
rect 6641 8381 6653 8384
rect 6687 8381 6699 8415
rect 8404 8412 8432 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 12618 8616 12624 8628
rect 10560 8588 12624 8616
rect 10560 8576 10566 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12802 8576 12808 8628
rect 12860 8616 12866 8628
rect 13265 8619 13323 8625
rect 13265 8616 13277 8619
rect 12860 8588 13277 8616
rect 12860 8576 12866 8588
rect 13265 8585 13277 8588
rect 13311 8585 13323 8619
rect 13265 8579 13323 8585
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 14458 8616 14464 8628
rect 13872 8588 14464 8616
rect 13872 8576 13878 8588
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 15105 8619 15163 8625
rect 14792 8588 15056 8616
rect 14792 8576 14798 8588
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 11517 8551 11575 8557
rect 11517 8548 11529 8551
rect 11480 8520 11529 8548
rect 11480 8508 11486 8520
rect 11517 8517 11529 8520
rect 11563 8517 11575 8551
rect 11517 8511 11575 8517
rect 11974 8508 11980 8560
rect 12032 8508 12038 8560
rect 12161 8551 12219 8557
rect 12161 8517 12173 8551
rect 12207 8517 12219 8551
rect 12161 8511 12219 8517
rect 12437 8551 12495 8557
rect 12437 8517 12449 8551
rect 12483 8548 12495 8551
rect 12894 8548 12900 8560
rect 12483 8520 12900 8548
rect 12483 8517 12495 8520
rect 12437 8511 12495 8517
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 8536 8452 8581 8480
rect 8536 8440 8542 8452
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 9548 8452 10149 8480
rect 9548 8440 9554 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 11992 8480 12020 8508
rect 10137 8443 10195 8449
rect 11155 8452 12020 8480
rect 9950 8412 9956 8424
rect 6641 8375 6699 8381
rect 7116 8384 8432 8412
rect 8579 8384 9956 8412
rect 3605 8347 3663 8353
rect 3605 8313 3617 8347
rect 3651 8344 3663 8347
rect 7116 8344 7144 8384
rect 3651 8316 7144 8344
rect 7184 8347 7242 8353
rect 3651 8313 3663 8316
rect 3605 8307 3663 8313
rect 7184 8313 7196 8347
rect 7230 8344 7242 8347
rect 7374 8344 7380 8356
rect 7230 8316 7380 8344
rect 7230 8313 7242 8316
rect 7184 8307 7242 8313
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 7466 8304 7472 8356
rect 7524 8344 7530 8356
rect 8579 8344 8607 8384
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10045 8415 10103 8421
rect 10045 8381 10057 8415
rect 10091 8412 10103 8415
rect 11155 8412 11183 8452
rect 10091 8384 11183 8412
rect 11609 8415 11667 8421
rect 10091 8381 10103 8384
rect 10045 8375 10103 8381
rect 11609 8381 11621 8415
rect 11655 8381 11667 8415
rect 11974 8412 11980 8424
rect 11935 8384 11980 8412
rect 11609 8375 11667 8381
rect 7524 8316 8607 8344
rect 8748 8347 8806 8353
rect 7524 8304 7530 8316
rect 8748 8313 8760 8347
rect 8794 8344 8806 8347
rect 10134 8344 10140 8356
rect 8794 8316 10140 8344
rect 8794 8313 8806 8316
rect 8748 8307 8806 8313
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 10410 8353 10416 8356
rect 10404 8307 10416 8353
rect 10468 8344 10474 8356
rect 11624 8344 11652 8375
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12176 8412 12204 8511
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 13630 8548 13636 8560
rect 13096 8520 13636 8548
rect 13096 8489 13124 8520
rect 13630 8508 13636 8520
rect 13688 8548 13694 8560
rect 13688 8520 13860 8548
rect 13688 8508 13694 8520
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 13832 8489 13860 8520
rect 13906 8508 13912 8560
rect 13964 8548 13970 8560
rect 14093 8551 14151 8557
rect 14093 8548 14105 8551
rect 13964 8520 14105 8548
rect 13964 8508 13970 8520
rect 14093 8517 14105 8520
rect 14139 8517 14151 8551
rect 14093 8511 14151 8517
rect 14182 8508 14188 8560
rect 14240 8548 14246 8560
rect 15028 8548 15056 8588
rect 15105 8585 15117 8619
rect 15151 8616 15163 8619
rect 16850 8616 16856 8628
rect 15151 8588 16856 8616
rect 15151 8585 15163 8588
rect 15105 8579 15163 8585
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 16942 8576 16948 8628
rect 17000 8616 17006 8628
rect 19889 8619 19947 8625
rect 17000 8588 17045 8616
rect 17000 8576 17006 8588
rect 19889 8585 19901 8619
rect 19935 8616 19947 8619
rect 19978 8616 19984 8628
rect 19935 8588 19984 8616
rect 19935 8585 19947 8588
rect 19889 8579 19947 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 15381 8551 15439 8557
rect 15381 8548 15393 8551
rect 14240 8520 14964 8548
rect 15028 8520 15393 8548
rect 14240 8508 14246 8520
rect 13817 8483 13875 8489
rect 13412 8452 13768 8480
rect 13412 8440 13418 8452
rect 13740 8412 13768 8452
rect 13817 8449 13829 8483
rect 13863 8449 13875 8483
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 13817 8443 13875 8449
rect 13924 8452 14657 8480
rect 13924 8412 13952 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 12176 8384 13676 8412
rect 13740 8384 13952 8412
rect 14461 8415 14519 8421
rect 12434 8344 12440 8356
rect 10468 8316 10504 8344
rect 11624 8316 12440 8344
rect 10410 8304 10416 8307
rect 10468 8304 10474 8316
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 12802 8344 12808 8356
rect 12763 8316 12808 8344
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 13648 8344 13676 8384
rect 14461 8381 14473 8415
rect 14507 8412 14519 8415
rect 14550 8412 14556 8424
rect 14507 8384 14556 8412
rect 14507 8381 14519 8384
rect 14461 8375 14519 8381
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 14936 8421 14964 8520
rect 15381 8517 15393 8520
rect 15427 8517 15439 8551
rect 15381 8511 15439 8517
rect 16482 8508 16488 8560
rect 16540 8548 16546 8560
rect 17034 8548 17040 8560
rect 16540 8520 17040 8548
rect 16540 8508 16546 8520
rect 17034 8508 17040 8520
rect 17092 8548 17098 8560
rect 17092 8520 18092 8548
rect 17092 8508 17098 8520
rect 15194 8440 15200 8492
rect 15252 8480 15258 8492
rect 15470 8480 15476 8492
rect 15252 8452 15476 8480
rect 15252 8440 15258 8452
rect 15470 8440 15476 8452
rect 15528 8440 15534 8492
rect 18064 8489 18092 8520
rect 17497 8483 17555 8489
rect 17497 8480 17509 8483
rect 16500 8452 17509 8480
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 15740 8415 15798 8421
rect 15740 8381 15752 8415
rect 15786 8412 15798 8415
rect 16022 8412 16028 8424
rect 15786 8384 16028 8412
rect 15786 8381 15798 8384
rect 15740 8375 15798 8381
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 16206 8372 16212 8424
rect 16264 8412 16270 8424
rect 16500 8412 16528 8452
rect 17497 8449 17509 8452
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18512 8483 18570 8489
rect 18512 8480 18524 8483
rect 18288 8452 18524 8480
rect 18288 8440 18294 8452
rect 18512 8449 18524 8452
rect 18558 8449 18570 8483
rect 18512 8443 18570 8449
rect 16264 8384 16528 8412
rect 16264 8372 16270 8384
rect 16666 8372 16672 8424
rect 16724 8412 16730 8424
rect 17405 8415 17463 8421
rect 17405 8412 17417 8415
rect 16724 8384 17417 8412
rect 16724 8372 16730 8384
rect 17405 8381 17417 8384
rect 17451 8381 17463 8415
rect 18322 8412 18328 8424
rect 17405 8375 17463 8381
rect 18064 8384 18328 8412
rect 18064 8356 18092 8384
rect 18322 8372 18328 8384
rect 18380 8421 18386 8424
rect 18380 8415 18430 8421
rect 18380 8381 18384 8415
rect 18418 8381 18430 8415
rect 18782 8412 18788 8424
rect 18743 8384 18788 8412
rect 18380 8375 18430 8381
rect 18380 8372 18386 8375
rect 18782 8372 18788 8384
rect 18840 8372 18846 8424
rect 17126 8344 17132 8356
rect 13648 8316 17132 8344
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 18046 8304 18052 8356
rect 18104 8304 18110 8356
rect 20070 8304 20076 8356
rect 20128 8344 20134 8356
rect 20165 8347 20223 8353
rect 20165 8344 20177 8347
rect 20128 8316 20177 8344
rect 20128 8304 20134 8316
rect 20165 8313 20177 8316
rect 20211 8344 20223 8347
rect 20349 8347 20407 8353
rect 20349 8344 20361 8347
rect 20211 8316 20361 8344
rect 20211 8313 20223 8316
rect 20165 8307 20223 8313
rect 20349 8313 20361 8316
rect 20395 8313 20407 8347
rect 20349 8307 20407 8313
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 9674 8276 9680 8288
rect 5040 8248 9680 8276
rect 5040 8236 5046 8248
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 11793 8279 11851 8285
rect 11793 8245 11805 8279
rect 11839 8276 11851 8279
rect 12342 8276 12348 8288
rect 11839 8248 12348 8276
rect 11839 8245 11851 8248
rect 11793 8239 11851 8245
rect 12342 8236 12348 8248
rect 12400 8236 12406 8288
rect 12894 8276 12900 8288
rect 12855 8248 12900 8276
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 13630 8276 13636 8288
rect 13591 8248 13636 8276
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 13722 8236 13728 8288
rect 13780 8276 13786 8288
rect 13780 8248 13825 8276
rect 13780 8236 13786 8248
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 14553 8279 14611 8285
rect 14553 8276 14565 8279
rect 14516 8248 14565 8276
rect 14516 8236 14522 8248
rect 14553 8245 14565 8248
rect 14599 8245 14611 8279
rect 14553 8239 14611 8245
rect 15381 8279 15439 8285
rect 15381 8245 15393 8279
rect 15427 8276 15439 8279
rect 15838 8276 15844 8288
rect 15427 8248 15844 8276
rect 15427 8245 15439 8248
rect 15381 8239 15439 8245
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 16850 8276 16856 8288
rect 16811 8248 16856 8276
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 17218 8236 17224 8288
rect 17276 8276 17282 8288
rect 17313 8279 17371 8285
rect 17313 8276 17325 8279
rect 17276 8248 17325 8276
rect 17276 8236 17282 8248
rect 17313 8245 17325 8248
rect 17359 8245 17371 8279
rect 17313 8239 17371 8245
rect 1104 8186 20884 8208
rect 1104 8134 7579 8186
rect 7631 8134 7643 8186
rect 7695 8134 7707 8186
rect 7759 8134 7771 8186
rect 7823 8134 14176 8186
rect 14228 8134 14240 8186
rect 14292 8134 14304 8186
rect 14356 8134 14368 8186
rect 14420 8134 20884 8186
rect 1104 8112 20884 8134
rect 4890 8032 4896 8084
rect 4948 8072 4954 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4948 8044 5089 8072
rect 4948 8032 4954 8044
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5077 8035 5135 8041
rect 5445 8075 5503 8081
rect 5445 8041 5457 8075
rect 5491 8072 5503 8075
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 5491 8044 6745 8072
rect 5491 8041 5503 8044
rect 5445 8035 5503 8041
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 6733 8035 6791 8041
rect 7576 8044 9689 8072
rect 3513 8007 3571 8013
rect 3513 7973 3525 8007
rect 3559 8004 3571 8007
rect 5626 8004 5632 8016
rect 3559 7976 5632 8004
rect 3559 7973 3571 7976
rect 3513 7967 3571 7973
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 5813 8007 5871 8013
rect 5813 8004 5825 8007
rect 5736 7976 5825 8004
rect 5736 7948 5764 7976
rect 5813 7973 5825 7976
rect 5859 7973 5871 8007
rect 5813 7967 5871 7973
rect 5902 7964 5908 8016
rect 5960 8004 5966 8016
rect 7576 8004 7604 8044
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 9677 8035 9735 8041
rect 10410 8032 10416 8084
rect 10468 8072 10474 8084
rect 11149 8075 11207 8081
rect 11149 8072 11161 8075
rect 10468 8044 11161 8072
rect 10468 8032 10474 8044
rect 11149 8041 11161 8044
rect 11195 8041 11207 8075
rect 11149 8035 11207 8041
rect 11241 8075 11299 8081
rect 11241 8041 11253 8075
rect 11287 8072 11299 8075
rect 11974 8072 11980 8084
rect 11287 8044 11980 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 12069 8075 12127 8081
rect 12069 8041 12081 8075
rect 12115 8072 12127 8075
rect 13354 8072 13360 8084
rect 12115 8044 13360 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 13630 8072 13636 8084
rect 13591 8044 13636 8072
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 15105 8075 15163 8081
rect 15105 8041 15117 8075
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 5960 7976 7604 8004
rect 7653 8007 7711 8013
rect 5960 7964 5966 7976
rect 7653 7973 7665 8007
rect 7699 8004 7711 8007
rect 8846 8004 8852 8016
rect 7699 7976 8852 8004
rect 7699 7973 7711 7976
rect 7653 7967 7711 7973
rect 8846 7964 8852 7976
rect 8904 7964 8910 8016
rect 9766 7964 9772 8016
rect 9824 8004 9830 8016
rect 11609 8007 11667 8013
rect 11609 8004 11621 8007
rect 9824 7976 11621 8004
rect 9824 7964 9830 7976
rect 11609 7973 11621 7976
rect 11655 7973 11667 8007
rect 11609 7967 11667 7973
rect 12520 8007 12578 8013
rect 12520 7973 12532 8007
rect 12566 8004 12578 8007
rect 13722 8004 13728 8016
rect 12566 7976 13728 8004
rect 12566 7973 12578 7976
rect 12520 7967 12578 7973
rect 13722 7964 13728 7976
rect 13780 7964 13786 8016
rect 15120 8004 15148 8035
rect 15286 8032 15292 8084
rect 15344 8072 15350 8084
rect 15657 8075 15715 8081
rect 15657 8072 15669 8075
rect 15344 8044 15669 8072
rect 15344 8032 15350 8044
rect 15657 8041 15669 8044
rect 15703 8041 15715 8075
rect 15657 8035 15715 8041
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 16117 8075 16175 8081
rect 15804 8044 15849 8072
rect 15804 8032 15810 8044
rect 16117 8041 16129 8075
rect 16163 8072 16175 8075
rect 17034 8072 17040 8084
rect 16163 8044 17040 8072
rect 16163 8041 16175 8044
rect 16117 8035 16175 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 17126 8032 17132 8084
rect 17184 8072 17190 8084
rect 20533 8075 20591 8081
rect 20533 8072 20545 8075
rect 17184 8044 20545 8072
rect 17184 8032 17190 8044
rect 20533 8041 20545 8044
rect 20579 8072 20591 8075
rect 20993 8075 21051 8081
rect 20993 8072 21005 8075
rect 20579 8044 21005 8072
rect 20579 8041 20591 8044
rect 20533 8035 20591 8041
rect 20993 8041 21005 8044
rect 21039 8041 21051 8075
rect 20993 8035 21051 8041
rect 15562 8004 15568 8016
rect 15120 7976 15568 8004
rect 15562 7964 15568 7976
rect 15620 8004 15626 8016
rect 16206 8004 16212 8016
rect 15620 7976 16212 8004
rect 15620 7964 15626 7976
rect 16206 7964 16212 7976
rect 16264 7964 16270 8016
rect 18506 7964 18512 8016
rect 18564 8004 18570 8016
rect 18564 7976 19196 8004
rect 18564 7964 18570 7976
rect 3602 7896 3608 7948
rect 3660 7936 3666 7948
rect 4982 7936 4988 7948
rect 3660 7908 3705 7936
rect 4943 7908 4988 7936
rect 3660 7896 3666 7908
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 5718 7896 5724 7948
rect 5776 7896 5782 7948
rect 6638 7936 6644 7948
rect 5828 7908 6500 7936
rect 6599 7908 6644 7936
rect 3786 7868 3792 7880
rect 3747 7840 3792 7868
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5828 7868 5856 7908
rect 5307 7840 5856 7868
rect 5905 7871 5963 7877
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 5994 7868 6000 7880
rect 5951 7840 6000 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6135 7840 6408 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 5074 7760 5080 7812
rect 5132 7800 5138 7812
rect 6104 7800 6132 7831
rect 5132 7772 6132 7800
rect 5132 7760 5138 7772
rect 3145 7735 3203 7741
rect 3145 7701 3157 7735
rect 3191 7732 3203 7735
rect 4062 7732 4068 7744
rect 3191 7704 4068 7732
rect 3191 7701 3203 7704
rect 3145 7695 3203 7701
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 4617 7735 4675 7741
rect 4617 7701 4629 7735
rect 4663 7732 4675 7735
rect 5350 7732 5356 7744
rect 4663 7704 5356 7732
rect 4663 7701 4675 7704
rect 4617 7695 4675 7701
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 5994 7692 6000 7744
rect 6052 7732 6058 7744
rect 6273 7735 6331 7741
rect 6273 7732 6285 7735
rect 6052 7704 6285 7732
rect 6052 7692 6058 7704
rect 6273 7701 6285 7704
rect 6319 7701 6331 7735
rect 6380 7732 6408 7840
rect 6472 7800 6500 7908
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 7745 7939 7803 7945
rect 7745 7905 7757 7939
rect 7791 7936 7803 7939
rect 8018 7936 8024 7948
rect 7791 7908 8024 7936
rect 7791 7905 7803 7908
rect 7745 7899 7803 7905
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7936 8171 7939
rect 8202 7936 8208 7948
rect 8159 7908 8208 7936
rect 8159 7905 8171 7908
rect 8113 7899 8171 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8380 7939 8438 7945
rect 8380 7905 8392 7939
rect 8426 7936 8438 7939
rect 9858 7936 9864 7948
rect 8426 7908 9864 7936
rect 8426 7905 8438 7908
rect 8380 7899 8438 7905
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 10042 7945 10048 7948
rect 10036 7936 10048 7945
rect 10003 7908 10048 7936
rect 10036 7899 10048 7908
rect 10042 7896 10048 7899
rect 10100 7896 10106 7948
rect 13538 7936 13544 7948
rect 12268 7908 13544 7936
rect 12268 7880 12296 7908
rect 13538 7896 13544 7908
rect 13596 7936 13602 7948
rect 13992 7939 14050 7945
rect 13596 7908 13768 7936
rect 13596 7896 13602 7908
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7466 7868 7472 7880
rect 6871 7840 7472 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 7834 7800 7840 7812
rect 6472 7772 7840 7800
rect 7834 7760 7840 7772
rect 7892 7760 7898 7812
rect 6730 7732 6736 7744
rect 6380 7704 6736 7732
rect 6273 7695 6331 7701
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 7248 7704 7297 7732
rect 7248 7692 7254 7704
rect 7285 7701 7297 7704
rect 7331 7701 7343 7735
rect 7944 7732 7972 7831
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 9548 7840 9781 7868
rect 9548 7828 9554 7840
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 11296 7840 11713 7868
rect 11296 7828 11302 7840
rect 11701 7837 11713 7840
rect 11747 7837 11759 7871
rect 11701 7831 11759 7837
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7868 11943 7871
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11931 7840 12081 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12250 7868 12256 7880
rect 12211 7840 12256 7868
rect 12069 7831 12127 7837
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 13740 7877 13768 7908
rect 13992 7905 14004 7939
rect 14038 7936 14050 7939
rect 14458 7936 14464 7948
rect 14038 7908 14464 7936
rect 14038 7905 14050 7908
rect 13992 7899 14050 7905
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 16022 7936 16028 7948
rect 15948 7908 16028 7936
rect 15948 7877 15976 7908
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 16390 7936 16396 7948
rect 16351 7908 16396 7936
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 16716 7939 16774 7945
rect 16716 7905 16728 7939
rect 16762 7936 16774 7939
rect 17034 7936 17040 7948
rect 16762 7908 17040 7936
rect 16762 7905 16774 7908
rect 16716 7899 16774 7905
rect 17034 7896 17040 7908
rect 17092 7896 17098 7948
rect 17129 7939 17187 7945
rect 17129 7905 17141 7939
rect 17175 7936 17187 7939
rect 17218 7936 17224 7948
rect 17175 7908 17224 7936
rect 17175 7905 17187 7908
rect 17129 7899 17187 7905
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 17770 7896 17776 7948
rect 17828 7936 17834 7948
rect 19168 7945 19196 7976
rect 19426 7945 19432 7948
rect 18693 7939 18751 7945
rect 18693 7936 18705 7939
rect 17828 7908 18705 7936
rect 17828 7896 17834 7908
rect 18693 7905 18705 7908
rect 18739 7905 18751 7939
rect 18693 7899 18751 7905
rect 19153 7939 19211 7945
rect 19153 7905 19165 7939
rect 19199 7905 19211 7939
rect 19420 7936 19432 7945
rect 19387 7908 19432 7936
rect 19153 7899 19211 7905
rect 19420 7899 19432 7908
rect 19426 7896 19432 7899
rect 19484 7896 19490 7948
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 15933 7871 15991 7877
rect 15933 7837 15945 7871
rect 15979 7837 15991 7871
rect 15933 7831 15991 7837
rect 16899 7871 16957 7877
rect 16899 7837 16911 7871
rect 16945 7868 16957 7871
rect 17788 7868 17816 7896
rect 18782 7868 18788 7880
rect 16945 7840 17816 7868
rect 18248 7840 18788 7868
rect 16945 7837 16957 7840
rect 16899 7831 16957 7837
rect 8386 7732 8392 7744
rect 7944 7704 8392 7732
rect 7285 7695 7343 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 9490 7732 9496 7744
rect 9451 7704 9496 7732
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 9677 7735 9735 7741
rect 9677 7701 9689 7735
rect 9723 7732 9735 7735
rect 14918 7732 14924 7744
rect 9723 7704 14924 7732
rect 9723 7701 9735 7704
rect 9677 7695 9735 7701
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 15289 7735 15347 7741
rect 15289 7701 15301 7735
rect 15335 7732 15347 7735
rect 15746 7732 15752 7744
rect 15335 7704 15752 7732
rect 15335 7701 15347 7704
rect 15289 7695 15347 7701
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 18248 7741 18276 7840
rect 18782 7828 18788 7840
rect 18840 7828 18846 7880
rect 18874 7828 18880 7880
rect 18932 7868 18938 7880
rect 18932 7840 18977 7868
rect 18932 7828 18938 7840
rect 18233 7735 18291 7741
rect 18233 7732 18245 7735
rect 18104 7704 18245 7732
rect 18104 7692 18110 7704
rect 18233 7701 18245 7704
rect 18279 7701 18291 7735
rect 18233 7695 18291 7701
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 19886 7732 19892 7744
rect 18371 7704 19892 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 19886 7692 19892 7704
rect 19944 7692 19950 7744
rect 1104 7642 20884 7664
rect 1104 7590 4280 7642
rect 4332 7590 4344 7642
rect 4396 7590 4408 7642
rect 4460 7590 4472 7642
rect 4524 7590 10878 7642
rect 10930 7590 10942 7642
rect 10994 7590 11006 7642
rect 11058 7590 11070 7642
rect 11122 7590 17475 7642
rect 17527 7590 17539 7642
rect 17591 7590 17603 7642
rect 17655 7590 17667 7642
rect 17719 7590 20884 7642
rect 1104 7568 20884 7590
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 6638 7528 6644 7540
rect 4479 7500 6644 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 8294 7528 8300 7540
rect 6840 7500 8300 7528
rect 3602 7460 3608 7472
rect 3563 7432 3608 7460
rect 3602 7420 3608 7432
rect 3660 7420 3666 7472
rect 4062 7392 4068 7404
rect 4023 7364 4068 7392
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4246 7392 4252 7404
rect 4207 7364 4252 7392
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 5074 7392 5080 7404
rect 5035 7364 5080 7392
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 6840 7401 6868 7500
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 8573 7531 8631 7537
rect 8573 7497 8585 7531
rect 8619 7528 8631 7531
rect 11238 7528 11244 7540
rect 8619 7500 11244 7528
rect 8619 7497 8631 7500
rect 8573 7491 8631 7497
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12802 7528 12808 7540
rect 12299 7500 12808 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 13817 7531 13875 7537
rect 13817 7528 13829 7531
rect 13780 7500 13829 7528
rect 13780 7488 13786 7500
rect 13817 7497 13829 7500
rect 13863 7497 13875 7531
rect 13817 7491 13875 7497
rect 14918 7488 14924 7540
rect 14976 7528 14982 7540
rect 17770 7528 17776 7540
rect 14976 7500 17632 7528
rect 17731 7500 17776 7528
rect 14976 7488 14982 7500
rect 7834 7420 7840 7472
rect 7892 7460 7898 7472
rect 9030 7460 9036 7472
rect 7892 7432 9036 7460
rect 7892 7420 7898 7432
rect 9030 7420 9036 7432
rect 9088 7420 9094 7472
rect 15470 7420 15476 7472
rect 15528 7460 15534 7472
rect 17604 7460 17632 7500
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 18046 7460 18052 7472
rect 15528 7432 16160 7460
rect 17604 7432 18052 7460
rect 15528 7420 15534 7432
rect 16132 7404 16160 7432
rect 18046 7420 18052 7432
rect 18104 7420 18110 7472
rect 19058 7420 19064 7472
rect 19116 7460 19122 7472
rect 19521 7463 19579 7469
rect 19521 7460 19533 7463
rect 19116 7432 19533 7460
rect 19116 7420 19122 7432
rect 5261 7395 5319 7401
rect 5261 7392 5273 7395
rect 5224 7364 5273 7392
rect 5224 7352 5230 7364
rect 5261 7361 5273 7364
rect 5307 7361 5319 7395
rect 5261 7355 5319 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 9306 7392 9312 7404
rect 9263 7364 9312 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 9456 7364 9501 7392
rect 9456 7352 9462 7364
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 13998 7392 14004 7404
rect 13872 7364 14004 7392
rect 13872 7352 13878 7364
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 14507 7395 14565 7401
rect 14507 7361 14519 7395
rect 14553 7392 14565 7395
rect 16114 7392 16120 7404
rect 14553 7364 15792 7392
rect 16027 7364 16120 7392
rect 14553 7361 14565 7364
rect 14507 7355 14565 7361
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7324 4951 7327
rect 4939 7296 5571 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 3513 7259 3571 7265
rect 3513 7225 3525 7259
rect 3559 7256 3571 7259
rect 3970 7256 3976 7268
rect 3559 7228 3976 7256
rect 3559 7225 3571 7228
rect 3513 7219 3571 7225
rect 3970 7216 3976 7228
rect 4028 7216 4034 7268
rect 5543 7265 5571 7296
rect 6454 7284 6460 7336
rect 6512 7324 6518 7336
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 6512 7296 8493 7324
rect 6512 7284 6518 7296
rect 8481 7293 8493 7296
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9657 7327 9715 7333
rect 9657 7324 9669 7327
rect 9548 7296 9669 7324
rect 9548 7284 9554 7296
rect 9657 7293 9669 7296
rect 9703 7293 9715 7327
rect 9657 7287 9715 7293
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 10686 7324 10692 7336
rect 10468 7296 10692 7324
rect 10468 7284 10474 7296
rect 10686 7284 10692 7296
rect 10744 7324 10750 7336
rect 10873 7327 10931 7333
rect 10873 7324 10885 7327
rect 10744 7296 10885 7324
rect 10744 7284 10750 7296
rect 10873 7293 10885 7296
rect 10919 7324 10931 7327
rect 12250 7324 12256 7336
rect 10919 7296 12256 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 12250 7284 12256 7296
rect 12308 7324 12314 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12308 7296 12449 7324
rect 12308 7284 12314 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 14737 7327 14795 7333
rect 14737 7324 14749 7327
rect 12437 7287 12495 7293
rect 12535 7296 12940 7324
rect 5528 7259 5586 7265
rect 5528 7225 5540 7259
rect 5574 7256 5586 7259
rect 6270 7256 6276 7268
rect 5574 7228 6276 7256
rect 5574 7225 5586 7228
rect 5528 7219 5586 7225
rect 6270 7216 6276 7228
rect 6328 7216 6334 7268
rect 7070 7259 7128 7265
rect 7070 7256 7082 7259
rect 6656 7228 7082 7256
rect 4801 7191 4859 7197
rect 4801 7157 4813 7191
rect 4847 7188 4859 7191
rect 5166 7188 5172 7200
rect 4847 7160 5172 7188
rect 4847 7157 4859 7160
rect 4801 7151 4859 7157
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 6656 7197 6684 7228
rect 7070 7225 7082 7228
rect 7116 7225 7128 7259
rect 7070 7219 7128 7225
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7256 8999 7259
rect 9508 7256 9536 7284
rect 8987 7228 9536 7256
rect 11140 7259 11198 7265
rect 8987 7225 8999 7228
rect 8941 7219 8999 7225
rect 11140 7225 11152 7259
rect 11186 7256 11198 7259
rect 11422 7256 11428 7268
rect 11186 7228 11428 7256
rect 11186 7225 11198 7228
rect 11140 7219 11198 7225
rect 11422 7216 11428 7228
rect 11480 7256 11486 7268
rect 12535 7256 12563 7296
rect 12912 7268 12940 7296
rect 14108 7296 14749 7324
rect 11480 7228 12563 7256
rect 12704 7259 12762 7265
rect 11480 7216 11486 7228
rect 12704 7225 12716 7259
rect 12750 7256 12762 7259
rect 12802 7256 12808 7268
rect 12750 7228 12808 7256
rect 12750 7225 12762 7228
rect 12704 7219 12762 7225
rect 12802 7216 12808 7228
rect 12860 7216 12866 7268
rect 12894 7216 12900 7268
rect 12952 7216 12958 7268
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 14108 7256 14136 7296
rect 14737 7293 14749 7296
rect 14783 7324 14795 7327
rect 15654 7324 15660 7336
rect 14783 7296 15660 7324
rect 14783 7293 14795 7296
rect 14737 7287 14795 7293
rect 15654 7284 15660 7296
rect 15712 7284 15718 7336
rect 13872 7228 14136 7256
rect 15764 7256 15792 7364
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 17144 7364 18092 7392
rect 16384 7327 16442 7333
rect 16384 7293 16396 7327
rect 16430 7324 16442 7327
rect 16850 7324 16856 7336
rect 16430 7296 16856 7324
rect 16430 7293 16442 7296
rect 16384 7287 16442 7293
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 17144 7324 17172 7364
rect 17052 7296 17172 7324
rect 17589 7327 17647 7333
rect 17052 7268 17080 7296
rect 17589 7293 17601 7327
rect 17635 7324 17647 7327
rect 17862 7324 17868 7336
rect 17635 7296 17868 7324
rect 17635 7293 17647 7296
rect 17589 7287 17647 7293
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 18064 7333 18092 7364
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 18316 7327 18374 7333
rect 18316 7293 18328 7327
rect 18362 7324 18374 7327
rect 18874 7324 18880 7336
rect 18362 7296 18880 7324
rect 18362 7293 18374 7296
rect 18316 7287 18374 7293
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 16942 7256 16948 7268
rect 15764 7228 16948 7256
rect 13872 7216 13878 7228
rect 16942 7216 16948 7228
rect 17000 7216 17006 7268
rect 17034 7216 17040 7268
rect 17092 7216 17098 7268
rect 19352 7256 19380 7432
rect 19521 7429 19533 7432
rect 19567 7429 19579 7463
rect 19521 7423 19579 7429
rect 19886 7352 19892 7404
rect 19944 7392 19950 7404
rect 19981 7395 20039 7401
rect 19981 7392 19993 7395
rect 19944 7364 19993 7392
rect 19944 7352 19950 7364
rect 19981 7361 19993 7364
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 20073 7395 20131 7401
rect 20073 7361 20085 7395
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 20088 7324 20116 7355
rect 17880 7228 19380 7256
rect 19444 7296 20116 7324
rect 17880 7200 17908 7228
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 5408 7160 6653 7188
rect 5408 7148 5414 7160
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 8202 7188 8208 7200
rect 8163 7160 8208 7188
rect 6641 7151 6699 7157
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7188 8355 7191
rect 8754 7188 8760 7200
rect 8343 7160 8760 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 8754 7148 8760 7160
rect 8812 7148 8818 7200
rect 9033 7191 9091 7197
rect 9033 7157 9045 7191
rect 9079 7188 9091 7191
rect 9858 7188 9864 7200
rect 9079 7160 9864 7188
rect 9079 7157 9091 7160
rect 9033 7151 9091 7157
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10042 7148 10048 7200
rect 10100 7188 10106 7200
rect 10781 7191 10839 7197
rect 10781 7188 10793 7191
rect 10100 7160 10793 7188
rect 10100 7148 10106 7160
rect 10781 7157 10793 7160
rect 10827 7157 10839 7191
rect 10781 7151 10839 7157
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14467 7191 14525 7197
rect 14467 7188 14479 7191
rect 14056 7160 14479 7188
rect 14056 7148 14062 7160
rect 14467 7157 14479 7160
rect 14513 7157 14525 7191
rect 14467 7151 14525 7157
rect 15841 7191 15899 7197
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 17218 7188 17224 7200
rect 15887 7160 17224 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 17494 7188 17500 7200
rect 17455 7160 17500 7188
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 17862 7148 17868 7200
rect 17920 7148 17926 7200
rect 18598 7148 18604 7200
rect 18656 7188 18662 7200
rect 19444 7197 19472 7296
rect 19889 7259 19947 7265
rect 19889 7225 19901 7259
rect 19935 7256 19947 7259
rect 20349 7259 20407 7265
rect 20349 7256 20361 7259
rect 19935 7228 20361 7256
rect 19935 7225 19947 7228
rect 19889 7219 19947 7225
rect 20349 7225 20361 7228
rect 20395 7225 20407 7259
rect 20349 7219 20407 7225
rect 19429 7191 19487 7197
rect 19429 7188 19441 7191
rect 18656 7160 19441 7188
rect 18656 7148 18662 7160
rect 19429 7157 19441 7160
rect 19475 7157 19487 7191
rect 19429 7151 19487 7157
rect 1104 7098 20884 7120
rect 1104 7046 7579 7098
rect 7631 7046 7643 7098
rect 7695 7046 7707 7098
rect 7759 7046 7771 7098
rect 7823 7046 14176 7098
rect 14228 7046 14240 7098
rect 14292 7046 14304 7098
rect 14356 7046 14368 7098
rect 14420 7046 20884 7098
rect 1104 7024 20884 7046
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 6270 6984 6276 6996
rect 4304 6956 5948 6984
rect 6231 6956 6276 6984
rect 4304 6944 4310 6956
rect 5920 6916 5948 6956
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 8294 6984 8300 6996
rect 6380 6956 8300 6984
rect 6380 6916 6408 6956
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 8481 6987 8539 6993
rect 8481 6953 8493 6987
rect 8527 6953 8539 6987
rect 8481 6947 8539 6953
rect 9861 6987 9919 6993
rect 9861 6953 9873 6987
rect 9907 6984 9919 6987
rect 11422 6984 11428 6996
rect 9907 6956 9996 6984
rect 11383 6956 11428 6984
rect 9907 6953 9919 6956
rect 9861 6947 9919 6953
rect 7368 6919 7426 6925
rect 7368 6916 7380 6919
rect 5920 6888 6408 6916
rect 7300 6888 7380 6916
rect 5160 6851 5218 6857
rect 5160 6817 5172 6851
rect 5206 6848 5218 6851
rect 5718 6848 5724 6860
rect 5206 6820 5724 6848
rect 5206 6817 5218 6820
rect 5160 6811 5218 6817
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 6454 6808 6460 6860
rect 6512 6848 6518 6860
rect 6549 6851 6607 6857
rect 6549 6848 6561 6851
rect 6512 6820 6561 6848
rect 6512 6808 6518 6820
rect 6549 6817 6561 6820
rect 6595 6817 6607 6851
rect 6549 6811 6607 6817
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 6825 6851 6883 6857
rect 6696 6820 6741 6848
rect 6696 6808 6702 6820
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 7300 6848 7328 6888
rect 7368 6885 7380 6888
rect 7414 6916 7426 6919
rect 8202 6916 8208 6928
rect 7414 6888 8208 6916
rect 7414 6885 7426 6888
rect 7368 6879 7426 6885
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 8496 6916 8524 6947
rect 8570 6916 8576 6928
rect 8496 6888 8576 6916
rect 8570 6876 8576 6888
rect 8628 6876 8634 6928
rect 8754 6876 8760 6928
rect 8812 6916 8818 6928
rect 9030 6916 9036 6928
rect 8812 6888 9036 6916
rect 8812 6876 8818 6888
rect 9030 6876 9036 6888
rect 9088 6876 9094 6928
rect 9125 6919 9183 6925
rect 9125 6885 9137 6919
rect 9171 6916 9183 6919
rect 9968 6916 9996 6956
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 13357 6987 13415 6993
rect 13357 6984 13369 6987
rect 11532 6956 13369 6984
rect 10042 6916 10048 6928
rect 9171 6888 9904 6916
rect 9968 6888 10048 6916
rect 9171 6885 9183 6888
rect 9125 6879 9183 6885
rect 9876 6860 9904 6888
rect 10042 6876 10048 6888
rect 10100 6876 10106 6928
rect 11238 6876 11244 6928
rect 11296 6916 11302 6928
rect 11532 6916 11560 6956
rect 13357 6953 13369 6956
rect 13403 6984 13415 6987
rect 13722 6984 13728 6996
rect 13403 6956 13728 6984
rect 13403 6953 13415 6956
rect 13357 6947 13415 6953
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 15013 6987 15071 6993
rect 15013 6984 15025 6987
rect 14516 6956 15025 6984
rect 14516 6944 14522 6956
rect 15013 6953 15025 6956
rect 15059 6984 15071 6987
rect 15105 6987 15163 6993
rect 15105 6984 15117 6987
rect 15059 6956 15117 6984
rect 15059 6953 15071 6956
rect 15013 6947 15071 6953
rect 15105 6953 15117 6956
rect 15151 6953 15163 6987
rect 15746 6984 15752 6996
rect 15707 6956 15752 6984
rect 15105 6947 15163 6953
rect 15746 6944 15752 6956
rect 15804 6984 15810 6996
rect 16577 6987 16635 6993
rect 16577 6984 16589 6987
rect 15804 6956 16589 6984
rect 15804 6944 15810 6956
rect 16577 6953 16589 6956
rect 16623 6953 16635 6987
rect 16577 6947 16635 6953
rect 16669 6987 16727 6993
rect 16669 6953 16681 6987
rect 16715 6984 16727 6987
rect 17218 6984 17224 6996
rect 16715 6956 17224 6984
rect 16715 6953 16727 6956
rect 16669 6947 16727 6953
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 18417 6987 18475 6993
rect 18417 6953 18429 6987
rect 18463 6984 18475 6987
rect 18874 6984 18880 6996
rect 18463 6956 18880 6984
rect 18463 6953 18475 6956
rect 18417 6947 18475 6953
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 11296 6888 11560 6916
rect 15488 6888 15792 6916
rect 11296 6876 11302 6888
rect 6871 6820 7328 6848
rect 8665 6851 8723 6857
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 8665 6817 8677 6851
rect 8711 6848 8723 6851
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 8711 6820 9689 6848
rect 8711 6817 8723 6820
rect 8665 6811 8723 6817
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 9858 6808 9864 6860
rect 9916 6808 9922 6860
rect 10134 6848 10140 6860
rect 10060 6820 10140 6848
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4672 6752 4905 6780
rect 4672 6740 4678 6752
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 7098 6780 7104 6792
rect 7059 6752 7104 6780
rect 4893 6743 4951 6749
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 10060 6789 10088 6820
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10318 6857 10324 6860
rect 10312 6811 10324 6857
rect 10376 6848 10382 6860
rect 10376 6820 10412 6848
rect 10318 6808 10324 6811
rect 10376 6808 10382 6820
rect 10594 6808 10600 6860
rect 10652 6848 10658 6860
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 10652 6820 11529 6848
rect 10652 6808 10658 6820
rect 11517 6817 11529 6820
rect 11563 6817 11575 6851
rect 11773 6851 11831 6857
rect 11773 6848 11785 6851
rect 11517 6811 11575 6817
rect 11624 6820 11785 6848
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 8352 6752 9229 6780
rect 8352 6740 8358 6752
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 10045 6783 10103 6789
rect 9447 6752 9628 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 6365 6647 6423 6653
rect 6365 6644 6377 6647
rect 4212 6616 6377 6644
rect 4212 6604 4218 6616
rect 6365 6613 6377 6616
rect 6411 6613 6423 6647
rect 6365 6607 6423 6613
rect 7009 6647 7067 6653
rect 7009 6613 7021 6647
rect 7055 6644 7067 6647
rect 8665 6647 8723 6653
rect 8665 6644 8677 6647
rect 7055 6616 8677 6644
rect 7055 6613 7067 6616
rect 7009 6607 7067 6613
rect 8665 6613 8677 6616
rect 8711 6613 8723 6647
rect 8665 6607 8723 6613
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6644 8815 6647
rect 9490 6644 9496 6656
rect 8803 6616 9496 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 9600 6644 9628 6752
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 11624 6780 11652 6820
rect 11773 6817 11785 6820
rect 11819 6817 11831 6851
rect 11773 6811 11831 6817
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6848 13047 6851
rect 13035 6820 13492 6848
rect 13035 6817 13047 6820
rect 12989 6811 13047 6817
rect 10045 6743 10103 6749
rect 11532 6752 11652 6780
rect 11532 6644 11560 6752
rect 12897 6715 12955 6721
rect 12897 6681 12909 6715
rect 12943 6712 12955 6715
rect 13262 6712 13268 6724
rect 12943 6684 13268 6712
rect 12943 6681 12955 6684
rect 12897 6675 12955 6681
rect 13262 6672 13268 6684
rect 13320 6672 13326 6724
rect 11698 6644 11704 6656
rect 9600 6616 11704 6644
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 13173 6647 13231 6653
rect 13173 6644 13185 6647
rect 12676 6616 13185 6644
rect 12676 6604 12682 6616
rect 13173 6613 13185 6616
rect 13219 6613 13231 6647
rect 13464 6644 13492 6820
rect 13538 6808 13544 6860
rect 13596 6848 13602 6860
rect 13900 6851 13958 6857
rect 13596 6820 13641 6848
rect 13596 6808 13602 6820
rect 13900 6817 13912 6851
rect 13946 6848 13958 6851
rect 15488 6848 15516 6888
rect 15654 6848 15660 6860
rect 13946 6820 15516 6848
rect 15615 6820 15660 6848
rect 13946 6817 13958 6820
rect 13900 6811 13958 6817
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 15764 6848 15792 6888
rect 16114 6876 16120 6928
rect 16172 6916 16178 6928
rect 17034 6916 17040 6928
rect 16172 6888 17040 6916
rect 16172 6876 16178 6888
rect 17034 6876 17040 6888
rect 17092 6876 17098 6928
rect 17310 6925 17316 6928
rect 17304 6916 17316 6925
rect 17223 6888 17316 6916
rect 17304 6879 17316 6888
rect 17368 6916 17374 6928
rect 17494 6916 17500 6928
rect 17368 6888 17500 6916
rect 17310 6876 17316 6879
rect 17368 6876 17374 6888
rect 17494 6876 17500 6888
rect 17552 6876 17558 6928
rect 19521 6919 19579 6925
rect 19521 6885 19533 6919
rect 19567 6916 19579 6919
rect 19794 6916 19800 6928
rect 19567 6888 19800 6916
rect 19567 6885 19579 6888
rect 19521 6879 19579 6885
rect 19794 6876 19800 6888
rect 19852 6876 19858 6928
rect 20990 6916 20996 6928
rect 20951 6888 20996 6916
rect 20990 6876 20996 6888
rect 21048 6876 21054 6928
rect 18598 6848 18604 6860
rect 15764 6820 18604 6848
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 18693 6851 18751 6857
rect 18693 6817 18705 6851
rect 18739 6817 18751 6851
rect 18693 6811 18751 6817
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6749 13691 6783
rect 13633 6743 13691 6749
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6780 15163 6783
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15151 6752 15853 6780
rect 15151 6749 15163 6752
rect 15105 6743 15163 6749
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 16850 6780 16856 6792
rect 16811 6752 16856 6780
rect 15841 6743 15899 6749
rect 13538 6672 13544 6724
rect 13596 6712 13602 6724
rect 13648 6712 13676 6743
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 17034 6780 17040 6792
rect 16995 6752 17040 6780
rect 17034 6740 17040 6752
rect 17092 6740 17098 6792
rect 18506 6740 18512 6792
rect 18564 6780 18570 6792
rect 18708 6780 18736 6811
rect 18782 6808 18788 6860
rect 18840 6848 18846 6860
rect 19978 6848 19984 6860
rect 18840 6820 18885 6848
rect 19939 6820 19984 6848
rect 18840 6808 18846 6820
rect 19978 6808 19984 6820
rect 20036 6808 20042 6860
rect 19610 6780 19616 6792
rect 18564 6752 18736 6780
rect 19571 6752 19616 6780
rect 18564 6740 18570 6752
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 13596 6684 13676 6712
rect 15289 6715 15347 6721
rect 13596 6672 13602 6684
rect 15289 6681 15301 6715
rect 15335 6712 15347 6715
rect 16666 6712 16672 6724
rect 15335 6684 16672 6712
rect 15335 6681 15347 6684
rect 15289 6675 15347 6681
rect 16666 6672 16672 6684
rect 16724 6672 16730 6724
rect 18046 6672 18052 6724
rect 18104 6712 18110 6724
rect 19720 6712 19748 6743
rect 20165 6715 20223 6721
rect 20165 6712 20177 6715
rect 18104 6684 20177 6712
rect 18104 6672 18110 6684
rect 20165 6681 20177 6684
rect 20211 6712 20223 6715
rect 20993 6715 21051 6721
rect 20993 6712 21005 6715
rect 20211 6684 21005 6712
rect 20211 6681 20223 6684
rect 20165 6675 20223 6681
rect 20993 6681 21005 6684
rect 21039 6681 21051 6715
rect 20993 6675 21051 6681
rect 13906 6644 13912 6656
rect 13464 6616 13912 6644
rect 13173 6607 13231 6613
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 15654 6604 15660 6656
rect 15712 6644 15718 6656
rect 16114 6644 16120 6656
rect 15712 6616 16120 6644
rect 15712 6604 15718 6616
rect 16114 6604 16120 6616
rect 16172 6604 16178 6656
rect 16209 6647 16267 6653
rect 16209 6613 16221 6647
rect 16255 6644 16267 6647
rect 17034 6644 17040 6656
rect 16255 6616 17040 6644
rect 16255 6613 16267 6616
rect 16209 6607 16267 6613
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18509 6647 18567 6653
rect 18509 6644 18521 6647
rect 18012 6616 18521 6644
rect 18012 6604 18018 6616
rect 18509 6613 18521 6616
rect 18555 6644 18567 6647
rect 18598 6644 18604 6656
rect 18555 6616 18604 6644
rect 18555 6613 18567 6616
rect 18509 6607 18567 6613
rect 18598 6604 18604 6616
rect 18656 6604 18662 6656
rect 18966 6644 18972 6656
rect 18927 6616 18972 6644
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 19153 6647 19211 6653
rect 19153 6613 19165 6647
rect 19199 6644 19211 6647
rect 19426 6644 19432 6656
rect 19199 6616 19432 6644
rect 19199 6613 19211 6616
rect 19153 6607 19211 6613
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 1104 6554 20884 6576
rect 1104 6502 4280 6554
rect 4332 6502 4344 6554
rect 4396 6502 4408 6554
rect 4460 6502 4472 6554
rect 4524 6502 10878 6554
rect 10930 6502 10942 6554
rect 10994 6502 11006 6554
rect 11058 6502 11070 6554
rect 11122 6502 17475 6554
rect 17527 6502 17539 6554
rect 17591 6502 17603 6554
rect 17655 6502 17667 6554
rect 17719 6502 20884 6554
rect 1104 6480 20884 6502
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 5776 6412 5917 6440
rect 5776 6400 5782 6412
rect 5905 6409 5917 6412
rect 5951 6409 5963 6443
rect 5905 6403 5963 6409
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6440 6883 6443
rect 8294 6440 8300 6452
rect 6871 6412 8300 6440
rect 6871 6409 6883 6412
rect 6825 6403 6883 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 9490 6400 9496 6452
rect 9548 6440 9554 6452
rect 12526 6440 12532 6452
rect 9548 6412 12532 6440
rect 9548 6400 9554 6412
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 12621 6443 12679 6449
rect 12621 6409 12633 6443
rect 12667 6440 12679 6443
rect 13078 6440 13084 6452
rect 12667 6412 13084 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 18506 6440 18512 6452
rect 14700 6412 18512 6440
rect 14700 6400 14706 6412
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 20530 6440 20536 6452
rect 20491 6412 20536 6440
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 6549 6375 6607 6381
rect 6549 6341 6561 6375
rect 6595 6372 6607 6375
rect 6914 6372 6920 6384
rect 6595 6344 6920 6372
rect 6595 6341 6607 6344
rect 6549 6335 6607 6341
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 7650 6372 7656 6384
rect 7024 6344 7656 6372
rect 7024 6304 7052 6344
rect 7650 6332 7656 6344
rect 7708 6332 7714 6384
rect 11698 6332 11704 6384
rect 11756 6372 11762 6384
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 11756 6344 11989 6372
rect 11756 6332 11762 6344
rect 11977 6341 11989 6344
rect 12023 6341 12035 6375
rect 11977 6335 12035 6341
rect 12894 6332 12900 6384
rect 12952 6372 12958 6384
rect 13630 6372 13636 6384
rect 12952 6344 13636 6372
rect 12952 6332 12958 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 18417 6375 18475 6381
rect 18417 6341 18429 6375
rect 18463 6341 18475 6375
rect 18417 6335 18475 6341
rect 7466 6304 7472 6316
rect 5552 6276 7052 6304
rect 7427 6276 7472 6304
rect 4525 6239 4583 6245
rect 4525 6205 4537 6239
rect 4571 6236 4583 6239
rect 4614 6236 4620 6248
rect 4571 6208 4620 6236
rect 4571 6205 4583 6208
rect 4525 6199 4583 6205
rect 4614 6196 4620 6208
rect 4672 6196 4678 6248
rect 5074 6236 5080 6248
rect 4715 6208 5080 6236
rect 4246 6128 4252 6180
rect 4304 6168 4310 6180
rect 4715 6168 4743 6208
rect 5074 6196 5080 6208
rect 5132 6236 5138 6248
rect 5552 6236 5580 6276
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 13449 6307 13507 6313
rect 13449 6304 13461 6307
rect 11624 6276 13461 6304
rect 5994 6236 6000 6248
rect 5132 6208 5580 6236
rect 5955 6208 6000 6236
rect 5132 6196 5138 6208
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 6365 6239 6423 6245
rect 6365 6205 6377 6239
rect 6411 6236 6423 6239
rect 6822 6236 6828 6248
rect 6411 6208 6828 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 9122 6236 9128 6248
rect 7699 6208 9128 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 4304 6140 4743 6168
rect 4792 6171 4850 6177
rect 4304 6128 4310 6140
rect 4792 6137 4804 6171
rect 4838 6168 4850 6171
rect 5902 6168 5908 6180
rect 4838 6140 5908 6168
rect 4838 6137 4850 6140
rect 4792 6131 4850 6137
rect 5902 6128 5908 6140
rect 5960 6128 5966 6180
rect 7098 6128 7104 6180
rect 7156 6168 7162 6180
rect 7668 6168 7696 6199
rect 9122 6196 9128 6208
rect 9180 6236 9186 6248
rect 10134 6236 10140 6248
rect 9180 6208 10140 6236
rect 9180 6196 9186 6208
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 10594 6236 10600 6248
rect 10555 6208 10600 6236
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 11624 6236 11652 6276
rect 13449 6273 13461 6276
rect 13495 6304 13507 6307
rect 13538 6304 13544 6316
rect 13495 6276 13544 6304
rect 13495 6273 13507 6276
rect 13449 6267 13507 6273
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 15746 6304 15752 6316
rect 15707 6276 15752 6304
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 16482 6264 16488 6316
rect 16540 6304 16546 6316
rect 16577 6307 16635 6313
rect 16577 6304 16589 6307
rect 16540 6276 16589 6304
rect 16540 6264 16546 6276
rect 16577 6273 16589 6276
rect 16623 6273 16635 6307
rect 16577 6267 16635 6273
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 17405 6307 17463 6313
rect 17405 6304 17417 6307
rect 17368 6276 17417 6304
rect 17368 6264 17374 6276
rect 17405 6273 17417 6276
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17770 6264 17776 6316
rect 17828 6304 17834 6316
rect 18432 6304 18460 6335
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 17828 6276 18705 6304
rect 17828 6264 17834 6276
rect 18693 6273 18705 6276
rect 18739 6273 18751 6307
rect 18693 6267 18751 6273
rect 10796 6208 11652 6236
rect 7156 6140 7696 6168
rect 7156 6128 7162 6140
rect 6178 6100 6184 6112
rect 6139 6072 6184 6100
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 7190 6100 7196 6112
rect 7151 6072 7196 6100
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 7285 6103 7343 6109
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 7374 6100 7380 6112
rect 7331 6072 7380 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 7668 6100 7696 6140
rect 7920 6171 7978 6177
rect 7920 6137 7932 6171
rect 7966 6168 7978 6171
rect 8662 6168 8668 6180
rect 7966 6140 8668 6168
rect 7966 6137 7978 6140
rect 7920 6131 7978 6137
rect 8662 6128 8668 6140
rect 8720 6128 8726 6180
rect 9392 6171 9450 6177
rect 9392 6137 9404 6171
rect 9438 6168 9450 6171
rect 10796 6168 10824 6208
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 11848 6208 12081 6236
rect 11848 6196 11854 6208
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12986 6236 12992 6248
rect 12483 6208 12992 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13630 6236 13636 6248
rect 13412 6208 13636 6236
rect 13412 6196 13418 6208
rect 13630 6196 13636 6208
rect 13688 6196 13694 6248
rect 16393 6239 16451 6245
rect 16393 6236 16405 6239
rect 13731 6208 16405 6236
rect 10870 6177 10876 6180
rect 9438 6140 10824 6168
rect 9438 6137 9450 6140
rect 9392 6131 9450 6137
rect 10864 6131 10876 6177
rect 10928 6168 10934 6180
rect 10928 6140 10964 6168
rect 10870 6128 10876 6131
rect 10928 6128 10934 6140
rect 11606 6128 11612 6180
rect 11664 6168 11670 6180
rect 13731 6168 13759 6208
rect 16393 6205 16405 6208
rect 16439 6205 16451 6239
rect 16393 6199 16451 6205
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6205 18107 6239
rect 18598 6236 18604 6248
rect 18559 6208 18604 6236
rect 18049 6199 18107 6205
rect 11664 6140 13759 6168
rect 13900 6171 13958 6177
rect 11664 6128 11670 6140
rect 13900 6137 13912 6171
rect 13946 6168 13958 6171
rect 14550 6168 14556 6180
rect 13946 6140 14556 6168
rect 13946 6137 13958 6140
rect 13900 6131 13958 6137
rect 14550 6128 14556 6140
rect 14608 6128 14614 6180
rect 14660 6140 16068 6168
rect 8110 6100 8116 6112
rect 7668 6072 8116 6100
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 9033 6103 9091 6109
rect 9033 6100 9045 6103
rect 8444 6072 9045 6100
rect 8444 6060 8450 6072
rect 9033 6069 9045 6072
rect 9079 6069 9091 6103
rect 9033 6063 9091 6069
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 10134 6100 10140 6112
rect 9272 6072 10140 6100
rect 9272 6060 9278 6072
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10502 6100 10508 6112
rect 10463 6072 10508 6100
rect 10502 6060 10508 6072
rect 10560 6060 10566 6112
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 12986 6100 12992 6112
rect 12851 6072 12992 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 13170 6100 13176 6112
rect 13131 6072 13176 6100
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13265 6103 13323 6109
rect 13265 6069 13277 6103
rect 13311 6100 13323 6103
rect 14660 6100 14688 6140
rect 15010 6100 15016 6112
rect 13311 6072 14688 6100
rect 14971 6072 15016 6100
rect 13311 6069 13323 6072
rect 13265 6063 13323 6069
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 15194 6100 15200 6112
rect 15155 6072 15200 6100
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 15528 6072 15577 6100
rect 15528 6060 15534 6072
rect 15565 6069 15577 6072
rect 15611 6069 15623 6103
rect 15565 6063 15623 6069
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6100 15715 6103
rect 15930 6100 15936 6112
rect 15703 6072 15936 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16040 6109 16068 6140
rect 16114 6128 16120 6180
rect 16172 6168 16178 6180
rect 16485 6171 16543 6177
rect 16485 6168 16497 6171
rect 16172 6140 16497 6168
rect 16172 6128 16178 6140
rect 16485 6137 16497 6140
rect 16531 6137 16543 6171
rect 16485 6131 16543 6137
rect 17221 6171 17279 6177
rect 17221 6137 17233 6171
rect 17267 6168 17279 6171
rect 17681 6171 17739 6177
rect 17681 6168 17693 6171
rect 17267 6140 17693 6168
rect 17267 6137 17279 6140
rect 17221 6131 17279 6137
rect 17681 6137 17693 6140
rect 17727 6137 17739 6171
rect 18064 6168 18092 6199
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 19978 6236 19984 6248
rect 18892 6208 19984 6236
rect 18892 6168 18920 6208
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 20162 6236 20168 6248
rect 20123 6208 20168 6236
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 18064 6140 18920 6168
rect 18960 6171 19018 6177
rect 17681 6131 17739 6137
rect 18960 6137 18972 6171
rect 19006 6168 19018 6171
rect 19518 6168 19524 6180
rect 19006 6140 19524 6168
rect 19006 6137 19018 6140
rect 18960 6131 19018 6137
rect 19518 6128 19524 6140
rect 19576 6128 19582 6180
rect 20349 6171 20407 6177
rect 20349 6137 20361 6171
rect 20395 6137 20407 6171
rect 20349 6131 20407 6137
rect 16025 6103 16083 6109
rect 16025 6069 16037 6103
rect 16071 6069 16083 6103
rect 16025 6063 16083 6069
rect 16298 6060 16304 6112
rect 16356 6100 16362 6112
rect 16850 6100 16856 6112
rect 16356 6072 16856 6100
rect 16356 6060 16362 6072
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 17034 6060 17040 6112
rect 17092 6100 17098 6112
rect 17313 6103 17371 6109
rect 17313 6100 17325 6103
rect 17092 6072 17325 6100
rect 17092 6060 17098 6072
rect 17313 6069 17325 6072
rect 17359 6069 17371 6103
rect 18230 6100 18236 6112
rect 18191 6072 18236 6100
rect 17313 6063 17371 6069
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 19886 6060 19892 6112
rect 19944 6100 19950 6112
rect 20073 6103 20131 6109
rect 20073 6100 20085 6103
rect 19944 6072 20085 6100
rect 19944 6060 19950 6072
rect 20073 6069 20085 6072
rect 20119 6100 20131 6103
rect 20364 6100 20392 6131
rect 20119 6072 20392 6100
rect 20119 6069 20131 6072
rect 20073 6063 20131 6069
rect 1104 6010 20884 6032
rect 1104 5958 7579 6010
rect 7631 5958 7643 6010
rect 7695 5958 7707 6010
rect 7759 5958 7771 6010
rect 7823 5958 14176 6010
rect 14228 5958 14240 6010
rect 14292 5958 14304 6010
rect 14356 5958 14368 6010
rect 14420 5958 20884 6010
rect 1104 5936 20884 5958
rect 3602 5896 3608 5908
rect 3563 5868 3608 5896
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5896 4307 5899
rect 4614 5896 4620 5908
rect 4295 5868 4620 5896
rect 4295 5865 4307 5868
rect 4249 5859 4307 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5902 5896 5908 5908
rect 5863 5868 5908 5896
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 6178 5856 6184 5908
rect 6236 5896 6242 5908
rect 6733 5899 6791 5905
rect 6733 5896 6745 5899
rect 6236 5868 6745 5896
rect 6236 5856 6242 5868
rect 6733 5865 6745 5868
rect 6779 5865 6791 5899
rect 6733 5859 6791 5865
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 9493 5899 9551 5905
rect 9493 5896 9505 5899
rect 7524 5868 9505 5896
rect 7524 5856 7530 5868
rect 9493 5865 9505 5868
rect 9539 5896 9551 5899
rect 10870 5896 10876 5908
rect 9539 5868 10876 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 13078 5896 13084 5908
rect 11020 5868 13084 5896
rect 11020 5856 11026 5868
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 16482 5896 16488 5908
rect 13320 5868 16488 5896
rect 13320 5856 13326 5868
rect 16482 5856 16488 5868
rect 16540 5856 16546 5908
rect 16758 5856 16764 5908
rect 16816 5896 16822 5908
rect 17129 5899 17187 5905
rect 17129 5896 17141 5899
rect 16816 5868 17141 5896
rect 16816 5856 16822 5868
rect 17129 5865 17141 5868
rect 17175 5865 17187 5899
rect 19518 5896 19524 5908
rect 17129 5859 17187 5865
rect 17328 5868 19104 5896
rect 19479 5868 19524 5896
rect 3513 5831 3571 5837
rect 3513 5797 3525 5831
rect 3559 5828 3571 5831
rect 7282 5828 7288 5840
rect 3559 5800 5948 5828
rect 3559 5797 3571 5800
rect 3513 5791 3571 5797
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4212 5732 4445 5760
rect 4212 5720 4218 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 4525 5763 4583 5769
rect 4525 5729 4537 5763
rect 4571 5760 4583 5763
rect 4614 5760 4620 5772
rect 4571 5732 4620 5760
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 4792 5763 4850 5769
rect 4792 5729 4804 5763
rect 4838 5760 4850 5763
rect 5810 5760 5816 5772
rect 4838 5732 5816 5760
rect 4838 5729 4850 5732
rect 4792 5723 4850 5729
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 4246 5692 4252 5704
rect 3835 5664 4252 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 5920 5692 5948 5800
rect 6012 5800 7288 5828
rect 6012 5769 6040 5800
rect 7282 5788 7288 5800
rect 7340 5828 7346 5840
rect 7653 5831 7711 5837
rect 7653 5828 7665 5831
rect 7340 5800 7665 5828
rect 7340 5788 7346 5800
rect 7653 5797 7665 5800
rect 7699 5797 7711 5831
rect 10042 5828 10048 5840
rect 7653 5791 7711 5797
rect 7852 5800 10048 5828
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5729 6055 5763
rect 5997 5723 6055 5729
rect 6362 5720 6368 5772
rect 6420 5760 6426 5772
rect 7558 5760 7564 5772
rect 6420 5732 7564 5760
rect 6420 5720 6426 5732
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 6546 5692 6552 5704
rect 5920 5664 6552 5692
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 6822 5692 6828 5704
rect 6783 5664 6828 5692
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7852 5701 7880 5800
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 17221 5831 17279 5837
rect 17221 5828 17233 5831
rect 13188 5800 17233 5828
rect 8110 5760 8116 5772
rect 8071 5732 8116 5760
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 8386 5769 8392 5772
rect 8380 5760 8392 5769
rect 8347 5732 8392 5760
rect 8380 5723 8392 5732
rect 8386 5720 8392 5723
rect 8444 5720 8450 5772
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5760 10195 5763
rect 10778 5760 10784 5772
rect 10183 5732 10784 5760
rect 10183 5729 10195 5732
rect 10137 5723 10195 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 10962 5760 10968 5772
rect 10923 5732 10968 5760
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 12802 5720 12808 5772
rect 12860 5760 12866 5772
rect 13188 5760 13216 5800
rect 17221 5797 17233 5800
rect 17267 5797 17279 5831
rect 17221 5791 17279 5797
rect 13262 5769 13268 5772
rect 12860 5732 13216 5760
rect 12860 5720 12866 5732
rect 13256 5723 13268 5769
rect 13320 5760 13326 5772
rect 13320 5732 13356 5760
rect 13262 5720 13268 5723
rect 13320 5720 13326 5732
rect 13538 5720 13544 5772
rect 13596 5760 13602 5772
rect 14642 5760 14648 5772
rect 13596 5732 14412 5760
rect 14603 5732 14648 5760
rect 13596 5720 13602 5732
rect 7837 5695 7895 5701
rect 6972 5664 7017 5692
rect 6972 5652 6978 5664
rect 7837 5661 7849 5695
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 10229 5655 10287 5661
rect 3145 5627 3203 5633
rect 3145 5593 3157 5627
rect 3191 5624 3203 5627
rect 6181 5627 6239 5633
rect 3191 5596 4568 5624
rect 3191 5593 3203 5596
rect 3145 5587 3203 5593
rect 4540 5556 4568 5596
rect 6181 5593 6193 5627
rect 6227 5624 6239 5627
rect 8110 5624 8116 5636
rect 6227 5596 8116 5624
rect 6227 5593 6239 5596
rect 6181 5587 6239 5593
rect 8110 5584 8116 5596
rect 8168 5584 8174 5636
rect 10042 5624 10048 5636
rect 9692 5596 10048 5624
rect 6270 5556 6276 5568
rect 4540 5528 6276 5556
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 6362 5516 6368 5568
rect 6420 5556 6426 5568
rect 6420 5528 6465 5556
rect 6420 5516 6426 5528
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 7193 5559 7251 5565
rect 7193 5556 7205 5559
rect 6972 5528 7205 5556
rect 6972 5516 6978 5528
rect 7193 5525 7205 5528
rect 7239 5525 7251 5559
rect 7193 5519 7251 5525
rect 7374 5516 7380 5568
rect 7432 5556 7438 5568
rect 9692 5556 9720 5596
rect 10042 5584 10048 5596
rect 10100 5584 10106 5636
rect 10244 5624 10272 5655
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 11057 5695 11115 5701
rect 10376 5664 10421 5692
rect 10376 5652 10382 5664
rect 11057 5661 11069 5695
rect 11103 5692 11115 5695
rect 11238 5692 11244 5704
rect 11103 5664 11244 5692
rect 11103 5661 11115 5664
rect 11057 5655 11115 5661
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 11422 5701 11428 5704
rect 11380 5695 11428 5701
rect 11380 5661 11392 5695
rect 11426 5661 11428 5695
rect 11380 5655 11428 5661
rect 11422 5652 11428 5655
rect 11480 5652 11486 5704
rect 11606 5701 11612 5704
rect 11563 5695 11612 5701
rect 11563 5661 11575 5695
rect 11609 5661 11612 5695
rect 11563 5655 11612 5661
rect 11606 5652 11612 5655
rect 11664 5652 11670 5704
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12986 5692 12992 5704
rect 11848 5664 11893 5692
rect 12947 5664 12992 5692
rect 11848 5652 11854 5664
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 10244 5596 11100 5624
rect 7432 5528 9720 5556
rect 9769 5559 9827 5565
rect 7432 5516 7438 5528
rect 9769 5525 9781 5559
rect 9815 5556 9827 5559
rect 10134 5556 10140 5568
rect 9815 5528 10140 5556
rect 9815 5525 9827 5528
rect 9769 5519 9827 5525
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 10781 5559 10839 5565
rect 10781 5556 10793 5559
rect 10468 5528 10793 5556
rect 10468 5516 10474 5528
rect 10781 5525 10793 5528
rect 10827 5525 10839 5559
rect 11072 5556 11100 5596
rect 11330 5556 11336 5568
rect 11072 5528 11336 5556
rect 10781 5519 10839 5525
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 12894 5556 12900 5568
rect 12855 5528 12900 5556
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 14384 5565 14412 5732
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 14829 5763 14887 5769
rect 14829 5729 14841 5763
rect 14875 5760 14887 5763
rect 15194 5760 15200 5772
rect 14875 5732 15200 5760
rect 14875 5729 14887 5732
rect 14829 5723 14887 5729
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 15562 5769 15568 5772
rect 15556 5760 15568 5769
rect 15523 5732 15568 5760
rect 15556 5723 15568 5732
rect 15562 5720 15568 5723
rect 15620 5720 15626 5772
rect 15930 5720 15936 5772
rect 15988 5760 15994 5772
rect 17328 5760 17356 5868
rect 17954 5828 17960 5840
rect 15988 5732 17356 5760
rect 17512 5800 17960 5828
rect 15988 5720 15994 5732
rect 15286 5692 15292 5704
rect 15247 5664 15292 5692
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5692 17463 5695
rect 17512 5692 17540 5800
rect 17954 5788 17960 5800
rect 18012 5828 18018 5840
rect 18966 5828 18972 5840
rect 18012 5800 18972 5828
rect 18012 5788 18018 5800
rect 18966 5788 18972 5800
rect 19024 5788 19030 5840
rect 19076 5828 19104 5868
rect 19518 5856 19524 5868
rect 19576 5896 19582 5908
rect 19981 5899 20039 5905
rect 19981 5896 19993 5899
rect 19576 5868 19993 5896
rect 19576 5856 19582 5868
rect 19981 5865 19993 5868
rect 20027 5865 20039 5899
rect 19981 5859 20039 5865
rect 20714 5828 20720 5840
rect 19076 5800 20720 5828
rect 20714 5788 20720 5800
rect 20772 5788 20778 5840
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 18408 5763 18466 5769
rect 18408 5729 18420 5763
rect 18454 5760 18466 5763
rect 19334 5760 19340 5772
rect 18454 5732 19340 5760
rect 18454 5729 18466 5732
rect 18408 5723 18466 5729
rect 17451 5664 17540 5692
rect 17451 5661 17463 5664
rect 17405 5655 17463 5661
rect 16761 5627 16819 5633
rect 16761 5593 16773 5627
rect 16807 5624 16819 5627
rect 17604 5624 17632 5723
rect 19334 5720 19340 5732
rect 19392 5760 19398 5772
rect 20073 5763 20131 5769
rect 20073 5760 20085 5763
rect 19392 5732 20085 5760
rect 19392 5720 19398 5732
rect 20073 5729 20085 5732
rect 20119 5729 20131 5763
rect 20073 5723 20131 5729
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 18046 5692 18052 5704
rect 17828 5664 18052 5692
rect 17828 5652 17834 5664
rect 18046 5652 18052 5664
rect 18104 5692 18110 5704
rect 18141 5695 18199 5701
rect 18141 5692 18153 5695
rect 18104 5664 18153 5692
rect 18104 5652 18110 5664
rect 18141 5661 18153 5664
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 20257 5695 20315 5701
rect 20257 5661 20269 5695
rect 20303 5692 20315 5695
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 20303 5664 21005 5692
rect 20303 5661 20315 5664
rect 20257 5655 20315 5661
rect 20993 5661 21005 5664
rect 21039 5661 21051 5695
rect 20993 5655 21051 5661
rect 16807 5596 17632 5624
rect 16807 5593 16819 5596
rect 16761 5587 16819 5593
rect 14369 5559 14427 5565
rect 14369 5525 14381 5559
rect 14415 5525 14427 5559
rect 14369 5519 14427 5525
rect 14458 5516 14464 5568
rect 14516 5556 14522 5568
rect 15013 5559 15071 5565
rect 14516 5528 14561 5556
rect 14516 5516 14522 5528
rect 15013 5525 15025 5559
rect 15059 5556 15071 5559
rect 15562 5556 15568 5568
rect 15059 5528 15568 5556
rect 15059 5525 15071 5528
rect 15013 5519 15071 5525
rect 15562 5516 15568 5528
rect 15620 5516 15626 5568
rect 15930 5516 15936 5568
rect 15988 5556 15994 5568
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 15988 5528 16681 5556
rect 15988 5516 15994 5528
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 17770 5556 17776 5568
rect 17731 5528 17776 5556
rect 16669 5519 16727 5525
rect 17770 5516 17776 5528
rect 17828 5516 17834 5568
rect 19610 5516 19616 5568
rect 19668 5556 19674 5568
rect 19668 5528 19713 5556
rect 19668 5516 19674 5528
rect 1104 5466 20884 5488
rect 1104 5414 4280 5466
rect 4332 5414 4344 5466
rect 4396 5414 4408 5466
rect 4460 5414 4472 5466
rect 4524 5414 10878 5466
rect 10930 5414 10942 5466
rect 10994 5414 11006 5466
rect 11058 5414 11070 5466
rect 11122 5414 17475 5466
rect 17527 5414 17539 5466
rect 17591 5414 17603 5466
rect 17655 5414 17667 5466
rect 17719 5414 20884 5466
rect 1104 5392 20884 5414
rect 5810 5312 5816 5364
rect 5868 5352 5874 5364
rect 5997 5355 6055 5361
rect 5997 5352 6009 5355
rect 5868 5324 6009 5352
rect 5868 5312 5874 5324
rect 5997 5321 6009 5324
rect 6043 5352 6055 5355
rect 6270 5352 6276 5364
rect 6043 5324 6276 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 6822 5352 6828 5364
rect 6503 5324 6828 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7282 5352 7288 5364
rect 7243 5324 7288 5352
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 8076 5324 8125 5352
rect 8076 5312 8082 5324
rect 8113 5321 8125 5324
rect 8159 5321 8171 5355
rect 8113 5315 8171 5321
rect 8220 5324 10272 5352
rect 7190 5244 7196 5296
rect 7248 5284 7254 5296
rect 8220 5284 8248 5324
rect 7248 5256 8248 5284
rect 10244 5284 10272 5324
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 10689 5355 10747 5361
rect 10689 5352 10701 5355
rect 10376 5324 10701 5352
rect 10376 5312 10382 5324
rect 10689 5321 10701 5324
rect 10735 5321 10747 5355
rect 10689 5315 10747 5321
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 12437 5355 12495 5361
rect 12437 5352 12449 5355
rect 11388 5324 12449 5352
rect 11388 5312 11394 5324
rect 12437 5321 12449 5324
rect 12483 5321 12495 5355
rect 12437 5315 12495 5321
rect 13078 5312 13084 5364
rect 13136 5352 13142 5364
rect 14366 5352 14372 5364
rect 13136 5324 14372 5352
rect 13136 5312 13142 5324
rect 14366 5312 14372 5324
rect 14424 5352 14430 5364
rect 15102 5352 15108 5364
rect 14424 5324 15108 5352
rect 14424 5312 14430 5324
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 15672 5324 19288 5352
rect 10244 5256 10364 5284
rect 7248 5244 7254 5256
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7064 5188 7849 5216
rect 7064 5176 7070 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 8662 5216 8668 5228
rect 8623 5188 8668 5216
rect 7837 5179 7895 5185
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 9180 5188 9321 5216
rect 9180 5176 9186 5188
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 10336 5216 10364 5256
rect 11238 5244 11244 5296
rect 11296 5284 11302 5296
rect 12158 5284 12164 5296
rect 11296 5256 12164 5284
rect 11296 5244 11302 5256
rect 12158 5244 12164 5256
rect 12216 5244 12222 5296
rect 15672 5284 15700 5324
rect 15028 5256 15700 5284
rect 19260 5284 19288 5324
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 19392 5324 19441 5352
rect 19392 5312 19398 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 19429 5315 19487 5321
rect 19521 5355 19579 5361
rect 19521 5321 19533 5355
rect 19567 5352 19579 5355
rect 19978 5352 19984 5364
rect 19567 5324 19984 5352
rect 19567 5321 19579 5324
rect 19521 5315 19579 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 19886 5284 19892 5296
rect 19260 5256 19892 5284
rect 10778 5216 10784 5228
rect 10336 5188 10640 5216
rect 10739 5188 10784 5216
rect 9309 5179 9367 5185
rect 4614 5148 4620 5160
rect 4575 5120 4620 5148
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6273 5151 6331 5157
rect 6273 5148 6285 5151
rect 6052 5120 6285 5148
rect 6052 5108 6058 5120
rect 6273 5117 6285 5120
rect 6319 5117 6331 5151
rect 6914 5148 6920 5160
rect 6875 5120 6920 5148
rect 6273 5111 6331 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7558 5108 7564 5160
rect 7616 5148 7622 5160
rect 8941 5151 8999 5157
rect 8941 5148 8953 5151
rect 7616 5120 8953 5148
rect 7616 5108 7622 5120
rect 8941 5117 8953 5120
rect 8987 5117 8999 5151
rect 8941 5111 8999 5117
rect 9576 5151 9634 5157
rect 9576 5117 9588 5151
rect 9622 5148 9634 5151
rect 10502 5148 10508 5160
rect 9622 5120 10508 5148
rect 9622 5117 9634 5120
rect 9576 5111 9634 5117
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 10612 5148 10640 5188
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 11698 5176 11704 5228
rect 11756 5216 11762 5228
rect 11977 5219 12035 5225
rect 11977 5216 11989 5219
rect 11756 5188 11989 5216
rect 11756 5176 11762 5188
rect 11977 5185 11989 5188
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 12308 5188 13001 5216
rect 12308 5176 12314 5188
rect 12989 5185 13001 5188
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 13170 5176 13176 5228
rect 13228 5216 13234 5228
rect 13265 5219 13323 5225
rect 13265 5216 13277 5219
rect 13228 5188 13277 5216
rect 13228 5176 13234 5188
rect 13265 5185 13277 5188
rect 13311 5185 13323 5219
rect 13265 5179 13323 5185
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 10612 5120 12909 5148
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 13538 5108 13544 5160
rect 13596 5148 13602 5160
rect 13633 5151 13691 5157
rect 13633 5148 13645 5151
rect 13596 5120 13645 5148
rect 13596 5108 13602 5120
rect 13633 5117 13645 5120
rect 13679 5117 13691 5151
rect 13633 5111 13691 5117
rect 13900 5151 13958 5157
rect 13900 5117 13912 5151
rect 13946 5148 13958 5151
rect 15028 5148 15056 5256
rect 19886 5244 19892 5256
rect 19944 5244 19950 5296
rect 17681 5219 17739 5225
rect 17681 5185 17693 5219
rect 17727 5216 17739 5219
rect 17727 5188 18184 5216
rect 17727 5185 17739 5188
rect 17681 5179 17739 5185
rect 13946 5120 15056 5148
rect 15105 5151 15163 5157
rect 13946 5117 13958 5120
rect 13900 5111 13958 5117
rect 15105 5117 15117 5151
rect 15151 5117 15163 5151
rect 15105 5111 15163 5117
rect 4884 5083 4942 5089
rect 4884 5049 4896 5083
rect 4930 5080 4942 5083
rect 5810 5080 5816 5092
rect 4930 5052 5816 5080
rect 4930 5049 4942 5052
rect 4884 5043 4942 5049
rect 5810 5040 5816 5052
rect 5868 5040 5874 5092
rect 8573 5083 8631 5089
rect 8573 5080 8585 5083
rect 7116 5052 8585 5080
rect 7116 5021 7144 5052
rect 8573 5049 8585 5052
rect 8619 5049 8631 5083
rect 11514 5080 11520 5092
rect 8573 5043 8631 5049
rect 9140 5052 11520 5080
rect 7101 5015 7159 5021
rect 7101 4981 7113 5015
rect 7147 4981 7159 5015
rect 7101 4975 7159 4981
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 7653 5015 7711 5021
rect 7653 5012 7665 5015
rect 7524 4984 7665 5012
rect 7524 4972 7530 4984
rect 7653 4981 7665 4984
rect 7699 4981 7711 5015
rect 7653 4975 7711 4981
rect 7745 5015 7803 5021
rect 7745 4981 7757 5015
rect 7791 5012 7803 5015
rect 7926 5012 7932 5024
rect 7791 4984 7932 5012
rect 7791 4981 7803 4984
rect 7745 4975 7803 4981
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 8110 4972 8116 5024
rect 8168 5012 8174 5024
rect 9140 5021 9168 5052
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 11885 5083 11943 5089
rect 11885 5049 11897 5083
rect 11931 5080 11943 5083
rect 12526 5080 12532 5092
rect 11931 5052 12532 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 15120 5080 15148 5111
rect 15286 5108 15292 5160
rect 15344 5148 15350 5160
rect 15657 5151 15715 5157
rect 15657 5148 15669 5151
rect 15344 5120 15669 5148
rect 15344 5108 15350 5120
rect 15657 5117 15669 5120
rect 15703 5148 15715 5151
rect 15746 5148 15752 5160
rect 15703 5120 15752 5148
rect 15703 5117 15715 5120
rect 15657 5111 15715 5117
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 15930 5157 15936 5160
rect 15924 5148 15936 5157
rect 15891 5120 15936 5148
rect 15924 5111 15936 5120
rect 15930 5108 15936 5111
rect 15988 5108 15994 5160
rect 17589 5151 17647 5157
rect 17589 5117 17601 5151
rect 17635 5148 17647 5151
rect 17770 5148 17776 5160
rect 17635 5120 17776 5148
rect 17635 5117 17647 5120
rect 17589 5111 17647 5117
rect 17770 5108 17776 5120
rect 17828 5108 17834 5160
rect 18046 5148 18052 5160
rect 17959 5120 18052 5148
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 18156 5148 18184 5188
rect 19426 5176 19432 5228
rect 19484 5216 19490 5228
rect 19981 5219 20039 5225
rect 19981 5216 19993 5219
rect 19484 5188 19993 5216
rect 19484 5176 19490 5188
rect 19981 5185 19993 5188
rect 20027 5185 20039 5219
rect 19981 5179 20039 5185
rect 20073 5219 20131 5225
rect 20073 5185 20085 5219
rect 20119 5185 20131 5219
rect 20073 5179 20131 5185
rect 18690 5148 18696 5160
rect 18156 5120 18696 5148
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 19610 5108 19616 5160
rect 19668 5148 19674 5160
rect 19889 5151 19947 5157
rect 19889 5148 19901 5151
rect 19668 5120 19901 5148
rect 19668 5108 19674 5120
rect 19889 5117 19901 5120
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 16022 5080 16028 5092
rect 15120 5052 16028 5080
rect 16022 5040 16028 5052
rect 16080 5080 16086 5092
rect 18064 5080 18092 5108
rect 16080 5052 17172 5080
rect 16080 5040 16086 5052
rect 8481 5015 8539 5021
rect 8481 5012 8493 5015
rect 8168 4984 8493 5012
rect 8168 4972 8174 4984
rect 8481 4981 8493 4984
rect 8527 4981 8539 5015
rect 8481 4975 8539 4981
rect 9125 5015 9183 5021
rect 9125 4981 9137 5015
rect 9171 4981 9183 5015
rect 11422 5012 11428 5024
rect 11383 4984 11428 5012
rect 9125 4975 9183 4981
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 11606 4972 11612 5024
rect 11664 5012 11670 5024
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 11664 4984 11805 5012
rect 11664 4972 11670 4984
rect 11793 4981 11805 4984
rect 11839 5012 11851 5015
rect 12066 5012 12072 5024
rect 11839 4984 12072 5012
rect 11839 4981 11851 4984
rect 11793 4975 11851 4981
rect 12066 4972 12072 4984
rect 12124 4972 12130 5024
rect 12802 5012 12808 5024
rect 12715 4984 12808 5012
rect 12802 4972 12808 4984
rect 12860 5012 12866 5024
rect 14642 5012 14648 5024
rect 12860 4984 14648 5012
rect 12860 4972 12866 4984
rect 14642 4972 14648 4984
rect 14700 4972 14706 5024
rect 15013 5015 15071 5021
rect 15013 4981 15025 5015
rect 15059 5012 15071 5015
rect 15194 5012 15200 5024
rect 15059 4984 15200 5012
rect 15059 4981 15071 4984
rect 15013 4975 15071 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15289 5015 15347 5021
rect 15289 4981 15301 5015
rect 15335 5012 15347 5015
rect 15654 5012 15660 5024
rect 15335 4984 15660 5012
rect 15335 4981 15347 4984
rect 15289 4975 15347 4981
rect 15654 4972 15660 4984
rect 15712 4972 15718 5024
rect 16390 4972 16396 5024
rect 16448 5012 16454 5024
rect 17144 5021 17172 5052
rect 17604 5052 18092 5080
rect 18316 5083 18374 5089
rect 17604 5024 17632 5052
rect 18316 5049 18328 5083
rect 18362 5080 18374 5083
rect 19334 5080 19340 5092
rect 18362 5052 19340 5080
rect 18362 5049 18374 5052
rect 18316 5043 18374 5049
rect 19334 5040 19340 5052
rect 19392 5040 19398 5092
rect 17037 5015 17095 5021
rect 17037 5012 17049 5015
rect 16448 4984 17049 5012
rect 16448 4972 16454 4984
rect 17037 4981 17049 4984
rect 17083 4981 17095 5015
rect 17037 4975 17095 4981
rect 17129 5015 17187 5021
rect 17129 4981 17141 5015
rect 17175 4981 17187 5015
rect 17129 4975 17187 4981
rect 17218 4972 17224 5024
rect 17276 5012 17282 5024
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 17276 4984 17509 5012
rect 17276 4972 17282 4984
rect 17497 4981 17509 4984
rect 17543 4981 17555 5015
rect 17497 4975 17555 4981
rect 17586 4972 17592 5024
rect 17644 4972 17650 5024
rect 18966 4972 18972 5024
rect 19024 5012 19030 5024
rect 20088 5012 20116 5179
rect 19024 4984 20116 5012
rect 19024 4972 19030 4984
rect 1104 4922 20884 4944
rect 1104 4870 7579 4922
rect 7631 4870 7643 4922
rect 7695 4870 7707 4922
rect 7759 4870 7771 4922
rect 7823 4870 14176 4922
rect 14228 4870 14240 4922
rect 14292 4870 14304 4922
rect 14356 4870 14368 4922
rect 14420 4870 20884 4922
rect 1104 4848 20884 4870
rect 5994 4808 6000 4820
rect 5955 4780 6000 4808
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6457 4811 6515 4817
rect 6457 4777 6469 4811
rect 6503 4808 6515 4811
rect 6825 4811 6883 4817
rect 6825 4808 6837 4811
rect 6503 4780 6837 4808
rect 6503 4777 6515 4780
rect 6457 4771 6515 4777
rect 6825 4777 6837 4780
rect 6871 4777 6883 4811
rect 7190 4808 7196 4820
rect 7151 4780 7196 4808
rect 6825 4771 6883 4777
rect 7190 4768 7196 4780
rect 7248 4768 7254 4820
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7524 4780 7849 4808
rect 7524 4768 7530 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 8389 4811 8447 4817
rect 8389 4777 8401 4811
rect 8435 4808 8447 4811
rect 9766 4808 9772 4820
rect 8435 4780 9772 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 11330 4808 11336 4820
rect 10100 4780 11336 4808
rect 10100 4768 10106 4780
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 12069 4811 12127 4817
rect 12069 4808 12081 4811
rect 11480 4780 12081 4808
rect 11480 4768 11486 4780
rect 12069 4777 12081 4780
rect 12115 4777 12127 4811
rect 12618 4808 12624 4820
rect 12579 4780 12624 4808
rect 12069 4771 12127 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 12989 4811 13047 4817
rect 12989 4777 13001 4811
rect 13035 4808 13047 4811
rect 15010 4808 15016 4820
rect 13035 4780 15016 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 15010 4768 15016 4780
rect 15068 4768 15074 4820
rect 15654 4808 15660 4820
rect 15615 4780 15660 4808
rect 15654 4768 15660 4780
rect 15712 4768 15718 4820
rect 15838 4768 15844 4820
rect 15896 4808 15902 4820
rect 17497 4811 17555 4817
rect 17497 4808 17509 4811
rect 15896 4780 17509 4808
rect 15896 4768 15902 4780
rect 17497 4777 17509 4780
rect 17543 4777 17555 4811
rect 17497 4771 17555 4777
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19794 4808 19800 4820
rect 19392 4780 19800 4808
rect 19392 4768 19398 4780
rect 19794 4768 19800 4780
rect 19852 4808 19858 4820
rect 20533 4811 20591 4817
rect 20533 4808 20545 4811
rect 19852 4780 20545 4808
rect 19852 4768 19858 4780
rect 20533 4777 20545 4780
rect 20579 4777 20591 4811
rect 20533 4771 20591 4777
rect 4792 4743 4850 4749
rect 4792 4709 4804 4743
rect 4838 4740 4850 4743
rect 6086 4740 6092 4752
rect 4838 4712 6092 4740
rect 4838 4709 4850 4712
rect 4792 4703 4850 4709
rect 6086 4700 6092 4712
rect 6144 4740 6150 4752
rect 7285 4743 7343 4749
rect 7285 4740 7297 4743
rect 6144 4712 7297 4740
rect 6144 4700 6150 4712
rect 7285 4709 7297 4712
rect 7331 4709 7343 4743
rect 7285 4703 7343 4709
rect 8481 4743 8539 4749
rect 8481 4709 8493 4743
rect 8527 4740 8539 4743
rect 9674 4740 9680 4752
rect 8527 4712 9680 4740
rect 8527 4709 8539 4712
rect 8481 4703 8539 4709
rect 9674 4700 9680 4712
rect 9732 4700 9738 4752
rect 12802 4740 12808 4752
rect 11440 4712 12808 4740
rect 4525 4675 4583 4681
rect 4525 4641 4537 4675
rect 4571 4672 4583 4675
rect 4614 4672 4620 4684
rect 4571 4644 4620 4672
rect 4571 4641 4583 4644
rect 4525 4635 4583 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 7650 4672 7656 4684
rect 6656 4644 7512 4672
rect 7611 4644 7656 4672
rect 6656 4613 6684 4644
rect 7484 4616 7512 4644
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 8846 4672 8852 4684
rect 8807 4644 8852 4672
rect 8846 4632 8852 4644
rect 8904 4632 8910 4684
rect 9030 4632 9036 4684
rect 9088 4672 9094 4684
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 9088 4644 9321 4672
rect 9088 4632 9094 4644
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 10000 4675 10058 4681
rect 10000 4672 10012 4675
rect 9548 4644 10012 4672
rect 9548 4632 9554 4644
rect 10000 4641 10012 4644
rect 10046 4641 10058 4675
rect 10000 4635 10058 4641
rect 10413 4675 10471 4681
rect 10413 4641 10425 4675
rect 10459 4672 10471 4675
rect 11440 4672 11468 4712
rect 12802 4700 12808 4712
rect 12860 4700 12866 4752
rect 13081 4743 13139 4749
rect 13081 4709 13093 4743
rect 13127 4740 13139 4743
rect 14182 4740 14188 4752
rect 13127 4712 14188 4740
rect 13127 4709 13139 4712
rect 13081 4703 13139 4709
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 15562 4700 15568 4752
rect 15620 4740 15626 4752
rect 15749 4743 15807 4749
rect 15749 4740 15761 4743
rect 15620 4712 15761 4740
rect 15620 4700 15626 4712
rect 15749 4709 15761 4712
rect 15795 4709 15807 4743
rect 15749 4703 15807 4709
rect 19420 4743 19478 4749
rect 19420 4709 19432 4743
rect 19466 4740 19478 4743
rect 19702 4740 19708 4752
rect 19466 4712 19708 4740
rect 19466 4709 19478 4712
rect 19420 4703 19478 4709
rect 19702 4700 19708 4712
rect 19760 4700 19766 4752
rect 11974 4672 11980 4684
rect 10459 4644 11468 4672
rect 11935 4644 11980 4672
rect 10459 4641 10471 4644
rect 10413 4635 10471 4641
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 12066 4632 12072 4684
rect 12124 4672 12130 4684
rect 12986 4672 12992 4684
rect 12124 4644 12992 4672
rect 12124 4632 12130 4644
rect 12986 4632 12992 4644
rect 13044 4672 13050 4684
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 13044 4644 13461 4672
rect 13044 4632 13050 4644
rect 13449 4641 13461 4644
rect 13495 4672 13507 4675
rect 13538 4672 13544 4684
rect 13495 4644 13544 4672
rect 13495 4641 13507 4644
rect 13449 4635 13507 4641
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 6822 4564 6828 4616
rect 6880 4604 6886 4616
rect 7377 4607 7435 4613
rect 7377 4604 7389 4607
rect 6880 4576 7389 4604
rect 6880 4564 6886 4576
rect 7377 4573 7389 4576
rect 7423 4573 7435 4607
rect 7377 4567 7435 4573
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 8665 4607 8723 4613
rect 8665 4604 8677 4607
rect 7524 4576 8677 4604
rect 7524 4564 7530 4576
rect 8665 4573 8677 4576
rect 8711 4604 8723 4607
rect 9582 4604 9588 4616
rect 8711 4576 9588 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4604 9735 4607
rect 9723 4573 9745 4604
rect 9677 4567 9745 4573
rect 5902 4536 5908 4548
rect 5815 4508 5908 4536
rect 5902 4496 5908 4508
rect 5960 4536 5966 4548
rect 7190 4536 7196 4548
rect 5960 4508 7196 4536
rect 5960 4496 5966 4508
rect 7190 4496 7196 4508
rect 7248 4496 7254 4548
rect 9122 4536 9128 4548
rect 9083 4508 9128 4536
rect 9122 4496 9128 4508
rect 9180 4496 9186 4548
rect 8018 4468 8024 4480
rect 7979 4440 8024 4468
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 9717 4468 9745 4567
rect 10134 4564 10140 4616
rect 10192 4604 10198 4616
rect 10192 4576 10237 4604
rect 10192 4564 10198 4576
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 11940 4576 12173 4604
rect 11940 4564 11946 4576
rect 12161 4573 12173 4576
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 13173 4607 13231 4613
rect 13173 4604 13185 4607
rect 12492 4576 13185 4604
rect 12492 4564 12498 4576
rect 13173 4573 13185 4576
rect 13219 4604 13231 4607
rect 13354 4604 13360 4616
rect 13219 4576 13360 4604
rect 13219 4573 13231 4576
rect 13173 4567 13231 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 11609 4539 11667 4545
rect 11609 4536 11621 4539
rect 11388 4508 11621 4536
rect 11388 4496 11394 4508
rect 11609 4505 11621 4508
rect 11655 4505 11667 4539
rect 11609 4499 11667 4505
rect 11238 4468 11244 4480
rect 9717 4440 11244 4468
rect 11238 4428 11244 4440
rect 11296 4428 11302 4480
rect 11422 4428 11428 4480
rect 11480 4468 11486 4480
rect 11517 4471 11575 4477
rect 11517 4468 11529 4471
rect 11480 4440 11529 4468
rect 11480 4428 11486 4440
rect 11517 4437 11529 4440
rect 11563 4468 11575 4471
rect 11790 4468 11796 4480
rect 11563 4440 11796 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 11790 4428 11796 4440
rect 11848 4428 11854 4480
rect 13464 4468 13492 4635
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 13716 4675 13774 4681
rect 13716 4641 13728 4675
rect 13762 4672 13774 4675
rect 15102 4672 15108 4684
rect 13762 4644 14872 4672
rect 15063 4644 15108 4672
rect 13762 4641 13774 4644
rect 13716 4635 13774 4641
rect 14844 4604 14872 4644
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 16390 4681 16396 4684
rect 16373 4675 16396 4681
rect 16373 4672 16385 4675
rect 16040 4644 16385 4672
rect 15194 4604 15200 4616
rect 14844 4576 15200 4604
rect 15194 4564 15200 4576
rect 15252 4604 15258 4616
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15252 4576 15853 4604
rect 15252 4564 15258 4576
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 14921 4539 14979 4545
rect 14921 4536 14933 4539
rect 14384 4508 14933 4536
rect 14384 4468 14412 4508
rect 14921 4505 14933 4508
rect 14967 4505 14979 4539
rect 14921 4499 14979 4505
rect 15378 4496 15384 4548
rect 15436 4536 15442 4548
rect 16040 4536 16068 4644
rect 16373 4641 16385 4644
rect 16448 4672 16454 4684
rect 16448 4644 16521 4672
rect 16373 4635 16396 4641
rect 16390 4632 16396 4635
rect 16448 4632 16454 4644
rect 17310 4632 17316 4684
rect 17368 4672 17374 4684
rect 17845 4675 17903 4681
rect 17845 4672 17857 4675
rect 17368 4644 17857 4672
rect 17368 4632 17374 4644
rect 17845 4641 17857 4644
rect 17891 4641 17903 4675
rect 17845 4635 17903 4641
rect 18138 4632 18144 4684
rect 18196 4672 18202 4684
rect 20530 4672 20536 4684
rect 18196 4644 20536 4672
rect 18196 4632 18202 4644
rect 20530 4632 20536 4644
rect 20588 4632 20594 4684
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4573 16175 4607
rect 17586 4604 17592 4616
rect 17499 4576 17592 4604
rect 16117 4567 16175 4573
rect 15436 4508 16068 4536
rect 15436 4496 15442 4508
rect 14826 4468 14832 4480
rect 13464 4440 14412 4468
rect 14787 4440 14832 4468
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 15286 4468 15292 4480
rect 15247 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 15746 4428 15752 4480
rect 15804 4468 15810 4480
rect 16132 4468 16160 4567
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 19150 4604 19156 4616
rect 19111 4576 19156 4604
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 17604 4536 17632 4564
rect 17052 4508 17632 4536
rect 17052 4480 17080 4508
rect 17034 4468 17040 4480
rect 15804 4440 17040 4468
rect 15804 4428 15810 4440
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 18598 4428 18604 4480
rect 18656 4468 18662 4480
rect 18969 4471 19027 4477
rect 18969 4468 18981 4471
rect 18656 4440 18981 4468
rect 18656 4428 18662 4440
rect 18969 4437 18981 4440
rect 19015 4437 19027 4471
rect 18969 4431 19027 4437
rect 1104 4378 20884 4400
rect 1104 4326 4280 4378
rect 4332 4326 4344 4378
rect 4396 4326 4408 4378
rect 4460 4326 4472 4378
rect 4524 4326 10878 4378
rect 10930 4326 10942 4378
rect 10994 4326 11006 4378
rect 11058 4326 11070 4378
rect 11122 4326 17475 4378
rect 17527 4326 17539 4378
rect 17591 4326 17603 4378
rect 17655 4326 17667 4378
rect 17719 4326 20884 4378
rect 1104 4304 20884 4326
rect 5810 4264 5816 4276
rect 5771 4236 5816 4264
rect 5810 4224 5816 4236
rect 5868 4224 5874 4276
rect 5905 4267 5963 4273
rect 5905 4233 5917 4267
rect 5951 4264 5963 4267
rect 6362 4264 6368 4276
rect 5951 4236 6368 4264
rect 5951 4233 5963 4236
rect 5905 4227 5963 4233
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 6825 4267 6883 4273
rect 6825 4233 6837 4267
rect 6871 4264 6883 4267
rect 7650 4264 7656 4276
rect 6871 4236 7656 4264
rect 6871 4233 6883 4236
rect 6825 4227 6883 4233
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 7837 4267 7895 4273
rect 7837 4233 7849 4267
rect 7883 4264 7895 4267
rect 7926 4264 7932 4276
rect 7883 4236 7932 4264
rect 7883 4233 7895 4236
rect 7837 4227 7895 4233
rect 7926 4224 7932 4236
rect 7984 4224 7990 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 11333 4267 11391 4273
rect 11333 4264 11345 4267
rect 9732 4236 11345 4264
rect 9732 4224 9738 4236
rect 11333 4233 11345 4236
rect 11379 4233 11391 4267
rect 11333 4227 11391 4233
rect 12618 4224 12624 4276
rect 12676 4264 12682 4276
rect 14182 4264 14188 4276
rect 12676 4236 13400 4264
rect 14143 4236 14188 4264
rect 12676 4224 12682 4236
rect 5828 4128 5856 4224
rect 6730 4196 6736 4208
rect 6564 4168 6736 4196
rect 6564 4137 6592 4168
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 7466 4196 7472 4208
rect 7392 4168 7472 4196
rect 7392 4137 7420 4168
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 9769 4199 9827 4205
rect 9769 4165 9781 4199
rect 9815 4165 9827 4199
rect 9769 4159 9827 4165
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5828 4100 6377 4128
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9784 4128 9812 4159
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 13372 4196 13400 4236
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 15013 4267 15071 4273
rect 15013 4264 15025 4267
rect 14292 4236 15025 4264
rect 14292 4196 14320 4236
rect 15013 4233 15025 4236
rect 15059 4233 15071 4267
rect 15013 4227 15071 4233
rect 16117 4267 16175 4273
rect 16117 4233 16129 4267
rect 16163 4264 16175 4267
rect 17218 4264 17224 4276
rect 16163 4236 17224 4264
rect 16163 4233 16175 4236
rect 16117 4227 16175 4233
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 19794 4224 19800 4276
rect 19852 4264 19858 4276
rect 20533 4267 20591 4273
rect 20533 4264 20545 4267
rect 19852 4236 20545 4264
rect 19852 4224 19858 4236
rect 20533 4233 20545 4236
rect 20579 4233 20591 4267
rect 20533 4227 20591 4233
rect 10928 4168 12020 4196
rect 13372 4168 14320 4196
rect 10928 4156 10934 4168
rect 9456 4100 9996 4128
rect 9456 4088 9462 4100
rect 4430 4060 4436 4072
rect 4391 4032 4436 4060
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 4700 4063 4758 4069
rect 4700 4029 4712 4063
rect 4746 4060 4758 4063
rect 5902 4060 5908 4072
rect 4746 4032 5908 4060
rect 4746 4029 4758 4032
rect 4700 4023 4758 4029
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 6270 4060 6276 4072
rect 6231 4032 6276 4060
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4060 7711 4063
rect 8018 4060 8024 4072
rect 7699 4032 8024 4060
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 8018 4020 8024 4032
rect 8076 4020 8082 4072
rect 8110 4020 8116 4072
rect 8168 4060 8174 4072
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 8168 4032 8401 4060
rect 8168 4020 8174 4032
rect 8389 4029 8401 4032
rect 8435 4060 8447 4063
rect 9122 4060 9128 4072
rect 8435 4032 9128 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 9122 4020 9128 4032
rect 9180 4060 9186 4072
rect 9858 4060 9864 4072
rect 9180 4032 9864 4060
rect 9180 4020 9186 4032
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 9968 4060 9996 4100
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 11790 4128 11796 4140
rect 11112 4100 11796 4128
rect 11112 4088 11118 4100
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 11992 4137 12020 4168
rect 14826 4156 14832 4208
rect 14884 4196 14890 4208
rect 17954 4196 17960 4208
rect 14884 4168 15608 4196
rect 14884 4156 14890 4168
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4128 12035 4131
rect 12342 4128 12348 4140
rect 12023 4100 12348 4128
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4128 14795 4131
rect 15102 4128 15108 4140
rect 14783 4100 15108 4128
rect 14783 4097 14795 4100
rect 14737 4091 14795 4097
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 15286 4088 15292 4140
rect 15344 4128 15350 4140
rect 15580 4137 15608 4168
rect 16960 4168 17960 4196
rect 16960 4137 16988 4168
rect 17788 4137 17816 4168
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 18049 4199 18107 4205
rect 18049 4165 18061 4199
rect 18095 4165 18107 4199
rect 18690 4196 18696 4208
rect 18049 4159 18107 4165
rect 18616 4168 18696 4196
rect 15473 4131 15531 4137
rect 15473 4128 15485 4131
rect 15344 4100 15485 4128
rect 15344 4088 15350 4100
rect 15473 4097 15485 4100
rect 15519 4097 15531 4131
rect 15473 4091 15531 4097
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4097 15623 4131
rect 16945 4131 17003 4137
rect 15565 4091 15623 4097
rect 15672 4100 16436 4128
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 9968 4032 11713 4060
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 12066 4020 12072 4072
rect 12124 4060 12130 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12124 4032 12449 4060
rect 12124 4020 12130 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 12704 4063 12762 4069
rect 12704 4029 12716 4063
rect 12750 4060 12762 4063
rect 14826 4060 14832 4072
rect 12750 4032 14832 4060
rect 12750 4029 12762 4032
rect 12704 4023 12762 4029
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 14918 4020 14924 4072
rect 14976 4060 14982 4072
rect 15672 4060 15700 4100
rect 14976 4032 15700 4060
rect 15933 4063 15991 4069
rect 14976 4020 14982 4032
rect 15488 4004 15516 4032
rect 15933 4029 15945 4063
rect 15979 4060 15991 4063
rect 16408 4060 16436 4100
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 17773 4131 17831 4137
rect 17773 4097 17785 4131
rect 17819 4097 17831 4131
rect 17773 4091 17831 4097
rect 18064 4060 18092 4159
rect 18616 4137 18644 4168
rect 18690 4156 18696 4168
rect 18748 4156 18754 4208
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 18601 4091 18659 4097
rect 15979 4032 16344 4060
rect 16408 4032 18092 4060
rect 15979 4029 15991 4032
rect 15933 4023 15991 4029
rect 8656 3995 8714 4001
rect 8656 3961 8668 3995
rect 8702 3992 8714 3995
rect 10128 3995 10186 4001
rect 8702 3964 10088 3992
rect 8702 3961 8714 3964
rect 8656 3955 8714 3961
rect 7190 3924 7196 3936
rect 7151 3896 7196 3924
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 7285 3927 7343 3933
rect 7285 3893 7297 3927
rect 7331 3924 7343 3927
rect 8386 3924 8392 3936
rect 7331 3896 8392 3924
rect 7331 3893 7343 3896
rect 7285 3887 7343 3893
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 10060 3924 10088 3964
rect 10128 3961 10140 3995
rect 10174 3992 10186 3995
rect 11054 3992 11060 4004
rect 10174 3964 11060 3992
rect 10174 3961 10186 3964
rect 10128 3955 10186 3961
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 11793 3995 11851 4001
rect 11793 3992 11805 3995
rect 11256 3964 11805 3992
rect 11256 3933 11284 3964
rect 11793 3961 11805 3964
rect 11839 3961 11851 3995
rect 11793 3955 11851 3961
rect 13909 3995 13967 4001
rect 13909 3961 13921 3995
rect 13955 3992 13967 3995
rect 15381 3995 15439 4001
rect 15381 3992 15393 3995
rect 13955 3964 15393 3992
rect 13955 3961 13967 3964
rect 13909 3955 13967 3961
rect 15381 3961 15393 3964
rect 15427 3961 15439 3995
rect 15381 3955 15439 3961
rect 15470 3952 15476 4004
rect 15528 3952 15534 4004
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 10060 3896 11253 3924
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 11241 3887 11299 3893
rect 13262 3884 13268 3936
rect 13320 3924 13326 3936
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 13320 3896 13829 3924
rect 13320 3884 13326 3896
rect 13817 3893 13829 3896
rect 13863 3893 13875 3927
rect 14550 3924 14556 3936
rect 14511 3896 14556 3924
rect 13817 3887 13875 3893
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 16316 3933 16344 4032
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 18288 4032 18429 4060
rect 18288 4020 18294 4032
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 19150 4060 19156 4072
rect 19111 4032 19156 4060
rect 18417 4023 18475 4029
rect 19150 4020 19156 4032
rect 19208 4020 19214 4072
rect 17497 3995 17555 4001
rect 17497 3961 17509 3995
rect 17543 3992 17555 3995
rect 19420 3995 19478 4001
rect 17543 3964 19380 3992
rect 17543 3961 17555 3964
rect 17497 3955 17555 3961
rect 16301 3927 16359 3933
rect 14700 3896 14745 3924
rect 14700 3884 14706 3896
rect 16301 3893 16313 3927
rect 16347 3893 16359 3927
rect 16666 3924 16672 3936
rect 16627 3896 16672 3924
rect 16301 3887 16359 3893
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 17126 3924 17132 3936
rect 16816 3896 16861 3924
rect 17087 3896 17132 3924
rect 16816 3884 16822 3896
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17589 3927 17647 3933
rect 17589 3893 17601 3927
rect 17635 3924 17647 3927
rect 17770 3924 17776 3936
rect 17635 3896 17776 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18509 3927 18567 3933
rect 18509 3893 18521 3927
rect 18555 3924 18567 3927
rect 18690 3924 18696 3936
rect 18555 3896 18696 3924
rect 18555 3893 18567 3896
rect 18509 3887 18567 3893
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 19352 3924 19380 3964
rect 19420 3961 19432 3995
rect 19466 3992 19478 3995
rect 20438 3992 20444 4004
rect 19466 3964 20444 3992
rect 19466 3961 19478 3964
rect 19420 3955 19478 3961
rect 20438 3952 20444 3964
rect 20496 3952 20502 4004
rect 19794 3924 19800 3936
rect 19352 3896 19800 3924
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 1104 3834 20884 3856
rect 1104 3782 7579 3834
rect 7631 3782 7643 3834
rect 7695 3782 7707 3834
rect 7759 3782 7771 3834
rect 7823 3782 14176 3834
rect 14228 3782 14240 3834
rect 14292 3782 14304 3834
rect 14356 3782 14368 3834
rect 14420 3782 20884 3834
rect 1104 3760 20884 3782
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 4856 3692 12204 3720
rect 4856 3680 4862 3692
rect 4700 3655 4758 3661
rect 4700 3621 4712 3655
rect 4746 3652 4758 3655
rect 6362 3652 6368 3664
rect 4746 3624 6368 3652
rect 4746 3621 4758 3624
rect 4700 3615 4758 3621
rect 6362 3612 6368 3624
rect 6420 3652 6426 3664
rect 8380 3655 8438 3661
rect 6420 3624 6592 3652
rect 6420 3612 6426 3624
rect 4430 3584 4436 3596
rect 4343 3556 4436 3584
rect 4430 3544 4436 3556
rect 4488 3584 4494 3596
rect 6181 3587 6239 3593
rect 6181 3584 6193 3587
rect 4488 3556 6193 3584
rect 4488 3544 4494 3556
rect 6181 3553 6193 3556
rect 6227 3584 6239 3587
rect 6270 3584 6276 3596
rect 6227 3556 6276 3584
rect 6227 3553 6239 3556
rect 6181 3547 6239 3553
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 6454 3593 6460 3596
rect 6448 3584 6460 3593
rect 6415 3556 6460 3584
rect 6448 3547 6460 3556
rect 6454 3544 6460 3547
rect 6512 3544 6518 3596
rect 6564 3584 6592 3624
rect 8380 3621 8392 3655
rect 8426 3652 8438 3655
rect 9674 3652 9680 3664
rect 8426 3624 9680 3652
rect 8426 3621 8438 3624
rect 8380 3615 8438 3621
rect 9674 3612 9680 3624
rect 9732 3652 9738 3664
rect 10137 3655 10195 3661
rect 10137 3652 10149 3655
rect 9732 3624 10149 3652
rect 9732 3612 9738 3624
rect 10137 3621 10149 3624
rect 10183 3621 10195 3655
rect 12176 3652 12204 3692
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 12308 3692 14504 3720
rect 12308 3680 12314 3692
rect 12342 3652 12348 3664
rect 12176 3624 12348 3652
rect 10137 3615 10195 3621
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 14476 3652 14504 3692
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14608 3692 15025 3720
rect 14608 3680 14614 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15013 3683 15071 3689
rect 15654 3680 15660 3732
rect 15712 3720 15718 3732
rect 16945 3723 17003 3729
rect 16945 3720 16957 3723
rect 15712 3692 16957 3720
rect 15712 3680 15718 3692
rect 16945 3689 16957 3692
rect 16991 3689 17003 3723
rect 18690 3720 18696 3732
rect 18651 3692 18696 3720
rect 16945 3683 17003 3689
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 20438 3680 20444 3732
rect 20496 3720 20502 3732
rect 20533 3723 20591 3729
rect 20533 3720 20545 3723
rect 20496 3692 20545 3720
rect 20496 3680 20502 3692
rect 20533 3689 20545 3692
rect 20579 3689 20591 3723
rect 20533 3683 20591 3689
rect 16758 3652 16764 3664
rect 14476 3624 16764 3652
rect 16758 3612 16764 3624
rect 16816 3612 16822 3664
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 17184 3624 18552 3652
rect 17184 3612 17190 3624
rect 8110 3584 8116 3596
rect 6564 3556 7227 3584
rect 8071 3556 8116 3584
rect 5813 3451 5871 3457
rect 5813 3417 5825 3451
rect 5859 3448 5871 3451
rect 6086 3448 6092 3460
rect 5859 3420 6092 3448
rect 5859 3417 5871 3420
rect 5813 3411 5871 3417
rect 6086 3408 6092 3420
rect 6144 3408 6150 3460
rect 7199 3448 7227 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 9306 3544 9312 3596
rect 9364 3584 9370 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9364 3556 10057 3584
rect 9364 3544 9370 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10152 3556 11652 3584
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 10152 3516 10180 3556
rect 10318 3516 10324 3528
rect 9640 3488 10180 3516
rect 10231 3488 10324 3516
rect 9640 3476 9646 3488
rect 10318 3476 10324 3488
rect 10376 3516 10382 3528
rect 10686 3516 10692 3528
rect 10376 3488 10692 3516
rect 10376 3476 10382 3488
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 10778 3476 10784 3528
rect 10836 3516 10842 3528
rect 11146 3525 11152 3528
rect 11104 3519 11152 3525
rect 10836 3488 10881 3516
rect 10836 3476 10842 3488
rect 11104 3485 11116 3519
rect 11150 3485 11152 3519
rect 11104 3479 11152 3485
rect 11146 3476 11152 3479
rect 11204 3476 11210 3528
rect 11330 3525 11336 3528
rect 11287 3519 11336 3525
rect 11287 3485 11299 3519
rect 11333 3485 11336 3519
rect 11287 3479 11336 3485
rect 11330 3476 11336 3479
rect 11388 3476 11394 3528
rect 11514 3516 11520 3528
rect 11475 3488 11520 3516
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 11624 3516 11652 3556
rect 12158 3544 12164 3596
rect 12216 3584 12222 3596
rect 12713 3587 12771 3593
rect 12713 3584 12725 3587
rect 12216 3556 12725 3584
rect 12216 3544 12222 3556
rect 12713 3553 12725 3556
rect 12759 3553 12771 3587
rect 13403 3587 13461 3593
rect 12713 3547 12771 3553
rect 12820 3556 13308 3584
rect 12820 3516 12848 3556
rect 11624 3488 12848 3516
rect 12986 3476 12992 3528
rect 13044 3525 13050 3528
rect 13044 3519 13094 3525
rect 13044 3485 13048 3519
rect 13082 3485 13094 3519
rect 13170 3516 13176 3528
rect 13134 3488 13176 3516
rect 13044 3479 13094 3485
rect 13044 3476 13050 3479
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 13280 3516 13308 3556
rect 13403 3553 13415 3587
rect 13449 3584 13461 3587
rect 13538 3584 13544 3596
rect 13449 3556 13544 3584
rect 13449 3553 13461 3556
rect 13403 3547 13461 3553
rect 13538 3544 13544 3556
rect 13596 3544 13602 3596
rect 14829 3587 14887 3593
rect 14829 3553 14841 3587
rect 14875 3584 14887 3587
rect 14918 3584 14924 3596
rect 14875 3556 14924 3584
rect 14875 3553 14887 3556
rect 14829 3547 14887 3553
rect 14918 3544 14924 3556
rect 14976 3544 14982 3596
rect 15010 3544 15016 3596
rect 15068 3584 15074 3596
rect 15838 3593 15844 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 15068 3556 15301 3584
rect 15068 3544 15074 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15832 3584 15844 3593
rect 15799 3556 15844 3584
rect 15289 3547 15347 3553
rect 15832 3547 15844 3556
rect 15838 3544 15844 3547
rect 15896 3544 15902 3596
rect 17310 3593 17316 3596
rect 17304 3547 17316 3593
rect 17368 3584 17374 3596
rect 18524 3593 18552 3624
rect 18509 3587 18567 3593
rect 17368 3556 17404 3584
rect 17310 3544 17316 3547
rect 17368 3544 17374 3556
rect 18509 3553 18521 3587
rect 18555 3553 18567 3587
rect 18509 3547 18567 3553
rect 19420 3587 19478 3593
rect 19420 3553 19432 3587
rect 19466 3584 19478 3587
rect 19978 3584 19984 3596
rect 19466 3556 19984 3584
rect 19466 3553 19478 3556
rect 19420 3547 19478 3553
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 15470 3516 15476 3528
rect 13280 3488 15476 3516
rect 15470 3476 15476 3488
rect 15528 3476 15534 3528
rect 15562 3476 15568 3528
rect 15620 3516 15626 3528
rect 17034 3516 17040 3528
rect 15620 3488 15665 3516
rect 16776 3488 17040 3516
rect 15620 3476 15626 3488
rect 7561 3451 7619 3457
rect 7561 3448 7573 3451
rect 7199 3420 7573 3448
rect 7561 3417 7573 3420
rect 7607 3417 7619 3451
rect 7561 3411 7619 3417
rect 9122 3408 9128 3460
rect 9180 3448 9186 3460
rect 9677 3451 9735 3457
rect 9180 3420 9608 3448
rect 9180 3408 9186 3420
rect 6546 3340 6552 3392
rect 6604 3380 6610 3392
rect 9306 3380 9312 3392
rect 6604 3352 9312 3380
rect 6604 3340 6610 3352
rect 9306 3340 9312 3352
rect 9364 3380 9370 3392
rect 9493 3383 9551 3389
rect 9493 3380 9505 3383
rect 9364 3352 9505 3380
rect 9364 3340 9370 3352
rect 9493 3349 9505 3352
rect 9539 3349 9551 3383
rect 9580 3380 9608 3420
rect 9677 3417 9689 3451
rect 9723 3448 9735 3451
rect 9766 3448 9772 3460
rect 9723 3420 9772 3448
rect 9723 3417 9735 3420
rect 9677 3411 9735 3417
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 14553 3451 14611 3457
rect 14553 3417 14565 3451
rect 14599 3448 14611 3451
rect 14642 3448 14648 3460
rect 14599 3420 14648 3448
rect 14599 3417 14611 3420
rect 14553 3411 14611 3417
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 12250 3380 12256 3392
rect 9580 3352 12256 3380
rect 9493 3343 9551 3349
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 12621 3383 12679 3389
rect 12621 3349 12633 3383
rect 12667 3380 12679 3383
rect 12894 3380 12900 3392
rect 12667 3352 12900 3380
rect 12667 3349 12679 3352
rect 12621 3343 12679 3349
rect 12894 3340 12900 3352
rect 12952 3380 12958 3392
rect 13538 3380 13544 3392
rect 12952 3352 13544 3380
rect 12952 3340 12958 3352
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 15562 3340 15568 3392
rect 15620 3380 15626 3392
rect 16776 3380 16804 3488
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 18690 3476 18696 3528
rect 18748 3516 18754 3528
rect 19150 3516 19156 3528
rect 18748 3488 19156 3516
rect 18748 3476 18754 3488
rect 19150 3476 19156 3488
rect 19208 3476 19214 3528
rect 15620 3352 16804 3380
rect 15620 3340 15626 3352
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 18417 3383 18475 3389
rect 18417 3380 18429 3383
rect 17276 3352 18429 3380
rect 17276 3340 17282 3352
rect 18417 3349 18429 3352
rect 18463 3349 18475 3383
rect 18417 3343 18475 3349
rect 1104 3290 20884 3312
rect 1104 3238 4280 3290
rect 4332 3238 4344 3290
rect 4396 3238 4408 3290
rect 4460 3238 4472 3290
rect 4524 3238 10878 3290
rect 10930 3238 10942 3290
rect 10994 3238 11006 3290
rect 11058 3238 11070 3290
rect 11122 3238 17475 3290
rect 17527 3238 17539 3290
rect 17591 3238 17603 3290
rect 17655 3238 17667 3290
rect 17719 3238 20884 3290
rect 1104 3216 20884 3238
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 4706 3176 4712 3188
rect 4479 3148 4712 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 6512 3148 8217 3176
rect 6512 3136 6518 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 9490 3176 9496 3188
rect 9088 3148 9496 3176
rect 9088 3136 9094 3148
rect 9490 3136 9496 3148
rect 9548 3136 9554 3188
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 11238 3176 11244 3188
rect 10336 3148 11244 3176
rect 9508 3108 9536 3136
rect 10336 3108 10364 3148
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 12434 3176 12440 3188
rect 11532 3148 12440 3176
rect 9508 3080 10364 3108
rect 5074 3040 5080 3052
rect 5035 3012 5080 3040
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 6328 3012 6776 3040
rect 6328 3000 6334 3012
rect 6748 2984 6776 3012
rect 8128 3012 8432 3040
rect 4798 2972 4804 2984
rect 4759 2944 4804 2972
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 5261 2975 5319 2981
rect 5261 2941 5273 2975
rect 5307 2941 5319 2975
rect 5261 2935 5319 2941
rect 5528 2975 5586 2981
rect 5528 2941 5540 2975
rect 5574 2972 5586 2975
rect 6546 2972 6552 2984
rect 5574 2944 6552 2972
rect 5574 2941 5586 2944
rect 5528 2935 5586 2941
rect 5276 2904 5304 2935
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 6730 2932 6736 2984
rect 6788 2932 6794 2984
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2972 6883 2975
rect 6914 2972 6920 2984
rect 6871 2944 6920 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 8128 2972 8156 3012
rect 7024 2944 8156 2972
rect 6270 2904 6276 2916
rect 5276 2876 6276 2904
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 7024 2904 7052 2944
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 8260 2944 8309 2972
rect 8260 2932 8266 2944
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 6564 2876 7052 2904
rect 7092 2907 7150 2913
rect 4893 2839 4951 2845
rect 4893 2805 4905 2839
rect 4939 2836 4951 2839
rect 6564 2836 6592 2876
rect 7092 2873 7104 2907
rect 7138 2904 7150 2907
rect 7138 2876 8340 2904
rect 7138 2873 7150 2876
rect 7092 2867 7150 2873
rect 8312 2848 8340 2876
rect 4939 2808 6592 2836
rect 6641 2839 6699 2845
rect 4939 2805 4951 2808
rect 4893 2799 4951 2805
rect 6641 2805 6653 2839
rect 6687 2836 6699 2839
rect 7006 2836 7012 2848
rect 6687 2808 7012 2836
rect 6687 2805 6699 2808
rect 6641 2799 6699 2805
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 8294 2796 8300 2848
rect 8352 2796 8358 2848
rect 8404 2836 8432 3012
rect 8564 2975 8622 2981
rect 8564 2941 8576 2975
rect 8610 2972 8622 2975
rect 9398 2972 9404 2984
rect 8610 2944 9404 2972
rect 8610 2941 8622 2944
rect 8564 2935 8622 2941
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2941 10379 2975
rect 10321 2935 10379 2941
rect 10588 2975 10646 2981
rect 10588 2941 10600 2975
rect 10634 2972 10646 2975
rect 11532 2972 11560 3148
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 12676 3148 15056 3176
rect 12676 3136 12682 3148
rect 11698 3108 11704 3120
rect 11659 3080 11704 3108
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3040 11851 3043
rect 11974 3040 11980 3052
rect 11839 3012 11980 3040
rect 11839 3009 11851 3012
rect 11793 3003 11851 3009
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 15028 3040 15056 3148
rect 15102 3136 15108 3188
rect 15160 3176 15166 3188
rect 15289 3179 15347 3185
rect 15289 3176 15301 3179
rect 15160 3148 15301 3176
rect 15160 3136 15166 3148
rect 15289 3145 15301 3148
rect 15335 3145 15347 3179
rect 15289 3139 15347 3145
rect 15470 3136 15476 3188
rect 15528 3176 15534 3188
rect 15528 3148 16436 3176
rect 15528 3136 15534 3148
rect 16408 3108 16436 3148
rect 16666 3136 16672 3188
rect 16724 3176 16730 3188
rect 16945 3179 17003 3185
rect 16945 3176 16957 3179
rect 16724 3148 16957 3176
rect 16724 3136 16730 3148
rect 16945 3145 16957 3148
rect 16991 3145 17003 3179
rect 16945 3139 17003 3145
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20073 3179 20131 3185
rect 20073 3176 20085 3179
rect 20036 3148 20085 3176
rect 20036 3136 20042 3148
rect 20073 3145 20085 3148
rect 20119 3145 20131 3179
rect 20073 3139 20131 3145
rect 18509 3111 18567 3117
rect 18509 3108 18521 3111
rect 16408 3080 18521 3108
rect 18509 3077 18521 3080
rect 18555 3077 18567 3111
rect 18509 3071 18567 3077
rect 15028 3012 15608 3040
rect 12066 2972 12072 2984
rect 10634 2944 11560 2972
rect 11624 2944 12072 2972
rect 10634 2941 10646 2944
rect 10588 2935 10646 2941
rect 10336 2904 10364 2935
rect 10686 2904 10692 2916
rect 10336 2876 10692 2904
rect 10686 2864 10692 2876
rect 10744 2904 10750 2916
rect 11624 2904 11652 2944
rect 12066 2932 12072 2944
rect 12124 2972 12130 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12124 2944 12449 2972
rect 12124 2932 12130 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12704 2975 12762 2981
rect 12704 2941 12716 2975
rect 12750 2972 12762 2975
rect 13262 2972 13268 2984
rect 12750 2944 13268 2972
rect 12750 2941 12762 2944
rect 12704 2935 12762 2941
rect 10744 2876 11652 2904
rect 12452 2904 12480 2935
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13906 2972 13912 2984
rect 13372 2944 13912 2972
rect 13372 2904 13400 2944
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 15470 2972 15476 2984
rect 15431 2944 15476 2972
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 15580 2972 15608 3012
rect 17310 3000 17316 3052
rect 17368 3040 17374 3052
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 17368 3012 17417 3040
rect 17368 3000 17374 3012
rect 17405 3009 17417 3012
rect 17451 3009 17463 3043
rect 17586 3040 17592 3052
rect 17547 3012 17592 3040
rect 17405 3003 17463 3009
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 18690 3040 18696 3052
rect 17696 3012 18696 3040
rect 17696 2984 17724 3012
rect 18690 3000 18696 3012
rect 18748 3000 18754 3052
rect 16206 2972 16212 2984
rect 15580 2944 16212 2972
rect 16206 2932 16212 2944
rect 16264 2932 16270 2984
rect 17034 2932 17040 2984
rect 17092 2972 17098 2984
rect 17678 2972 17684 2984
rect 17092 2944 17684 2972
rect 17092 2932 17098 2944
rect 17678 2932 17684 2944
rect 17736 2932 17742 2984
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 19242 2972 19248 2984
rect 18371 2944 19248 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 19242 2932 19248 2944
rect 19300 2972 19306 2984
rect 20070 2972 20076 2984
rect 19300 2944 20076 2972
rect 19300 2932 19306 2944
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 14154 2907 14212 2913
rect 14154 2904 14166 2907
rect 12452 2876 13400 2904
rect 13832 2876 14166 2904
rect 10744 2864 10750 2876
rect 11514 2836 11520 2848
rect 8404 2808 11520 2836
rect 11514 2796 11520 2808
rect 11572 2796 11578 2848
rect 13078 2796 13084 2848
rect 13136 2836 13142 2848
rect 13832 2845 13860 2876
rect 14154 2873 14166 2876
rect 14200 2873 14212 2907
rect 14154 2867 14212 2873
rect 15654 2864 15660 2916
rect 15712 2913 15718 2916
rect 15712 2907 15776 2913
rect 15712 2873 15730 2907
rect 15764 2873 15776 2907
rect 15712 2867 15776 2873
rect 15712 2864 15718 2867
rect 17218 2864 17224 2916
rect 17276 2904 17282 2916
rect 17313 2907 17371 2913
rect 17313 2904 17325 2907
rect 17276 2876 17325 2904
rect 17276 2864 17282 2876
rect 17313 2873 17325 2876
rect 17359 2873 17371 2907
rect 17313 2867 17371 2873
rect 17586 2864 17592 2916
rect 17644 2904 17650 2916
rect 18046 2904 18052 2916
rect 17644 2876 18052 2904
rect 17644 2864 17650 2876
rect 18046 2864 18052 2876
rect 18104 2864 18110 2916
rect 18966 2913 18972 2916
rect 18960 2867 18972 2913
rect 19024 2904 19030 2916
rect 19024 2876 19060 2904
rect 18966 2864 18972 2867
rect 19024 2864 19030 2876
rect 13817 2839 13875 2845
rect 13817 2836 13829 2839
rect 13136 2808 13829 2836
rect 13136 2796 13142 2808
rect 13817 2805 13829 2808
rect 13863 2805 13875 2839
rect 13817 2799 13875 2805
rect 16206 2796 16212 2848
rect 16264 2836 16270 2848
rect 16853 2839 16911 2845
rect 16853 2836 16865 2839
rect 16264 2808 16865 2836
rect 16264 2796 16270 2808
rect 16853 2805 16865 2808
rect 16899 2805 16911 2839
rect 16853 2799 16911 2805
rect 1104 2746 20884 2768
rect 1104 2694 7579 2746
rect 7631 2694 7643 2746
rect 7695 2694 7707 2746
rect 7759 2694 7771 2746
rect 7823 2694 14176 2746
rect 14228 2694 14240 2746
rect 14292 2694 14304 2746
rect 14356 2694 14368 2746
rect 14420 2694 20884 2746
rect 1104 2672 20884 2694
rect 6454 2632 6460 2644
rect 6415 2604 6460 2632
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 6822 2592 6828 2644
rect 6880 2632 6886 2644
rect 8294 2632 8300 2644
rect 6880 2604 8156 2632
rect 8255 2604 8300 2632
rect 6880 2592 6886 2604
rect 6362 2564 6368 2576
rect 6323 2536 6368 2564
rect 6362 2524 6368 2536
rect 6420 2524 6426 2576
rect 6840 2564 6868 2592
rect 6656 2536 6868 2564
rect 6656 2437 6684 2536
rect 7006 2524 7012 2576
rect 7064 2564 7070 2576
rect 7064 2536 7144 2564
rect 7064 2524 7070 2536
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 6914 2496 6920 2508
rect 6788 2468 6920 2496
rect 6788 2456 6794 2468
rect 6914 2456 6920 2468
rect 6972 2496 6978 2508
rect 7116 2496 7144 2536
rect 7184 2499 7242 2505
rect 7184 2496 7196 2499
rect 6972 2468 7065 2496
rect 7116 2468 7196 2496
rect 6972 2456 6978 2468
rect 7184 2465 7196 2468
rect 7230 2496 7242 2499
rect 8128 2496 8156 2604
rect 8294 2592 8300 2604
rect 8352 2632 8358 2644
rect 8757 2635 8815 2641
rect 8757 2632 8769 2635
rect 8352 2604 8769 2632
rect 8352 2592 8358 2604
rect 8757 2601 8769 2604
rect 8803 2601 8815 2635
rect 8757 2595 8815 2601
rect 11609 2635 11667 2641
rect 11609 2601 11621 2635
rect 11655 2632 11667 2635
rect 11882 2632 11888 2644
rect 11655 2604 11888 2632
rect 11655 2601 11667 2604
rect 11609 2595 11667 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12161 2635 12219 2641
rect 12161 2601 12173 2635
rect 12207 2632 12219 2635
rect 12621 2635 12679 2641
rect 12621 2632 12633 2635
rect 12207 2604 12633 2632
rect 12207 2601 12219 2604
rect 12161 2595 12219 2601
rect 12621 2601 12633 2604
rect 12667 2601 12679 2635
rect 12621 2595 12679 2601
rect 12894 2592 12900 2644
rect 12952 2632 12958 2644
rect 13081 2635 13139 2641
rect 13081 2632 13093 2635
rect 12952 2604 13093 2632
rect 12952 2592 12958 2604
rect 13081 2601 13093 2604
rect 13127 2601 13139 2635
rect 13081 2595 13139 2601
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 15289 2635 15347 2641
rect 15289 2632 15301 2635
rect 13412 2604 15301 2632
rect 13412 2592 13418 2604
rect 15289 2601 15301 2604
rect 15335 2601 15347 2635
rect 17310 2632 17316 2644
rect 17271 2604 17316 2632
rect 15289 2595 15347 2601
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17405 2635 17463 2641
rect 17405 2601 17417 2635
rect 17451 2632 17463 2635
rect 17770 2632 17776 2644
rect 17451 2604 17776 2632
rect 17451 2601 17463 2604
rect 17405 2595 17463 2601
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 18966 2592 18972 2644
rect 19024 2632 19030 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 19024 2604 19717 2632
rect 19024 2592 19030 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 19705 2595 19763 2601
rect 19794 2592 19800 2644
rect 19852 2632 19858 2644
rect 19852 2604 19897 2632
rect 19852 2592 19858 2604
rect 19978 2592 19984 2644
rect 20036 2632 20042 2644
rect 20257 2635 20315 2641
rect 20257 2632 20269 2635
rect 20036 2604 20269 2632
rect 20036 2592 20042 2604
rect 20257 2601 20269 2604
rect 20303 2601 20315 2635
rect 20257 2595 20315 2601
rect 10496 2567 10554 2573
rect 10496 2533 10508 2567
rect 10542 2564 10554 2567
rect 11698 2564 11704 2576
rect 10542 2536 11704 2564
rect 10542 2533 10554 2536
rect 10496 2527 10554 2533
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 12069 2567 12127 2573
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 13449 2567 13507 2573
rect 13449 2564 13461 2567
rect 12115 2536 13461 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 13449 2533 13461 2536
rect 13495 2533 13507 2567
rect 13449 2527 13507 2533
rect 14176 2567 14234 2573
rect 14176 2533 14188 2567
rect 14222 2564 14234 2567
rect 15102 2564 15108 2576
rect 14222 2536 15108 2564
rect 14222 2533 14234 2536
rect 14176 2527 14234 2533
rect 15102 2524 15108 2536
rect 15160 2524 15166 2576
rect 16206 2573 16212 2576
rect 16200 2564 16212 2573
rect 16167 2536 16212 2564
rect 16200 2527 16212 2536
rect 16206 2524 16212 2527
rect 16264 2524 16270 2576
rect 18984 2564 19012 2592
rect 17788 2536 19012 2564
rect 20165 2567 20223 2573
rect 7230 2468 7972 2496
rect 8128 2468 9076 2496
rect 7230 2465 7242 2468
rect 7184 2459 7242 2465
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2397 6699 2431
rect 7944 2428 7972 2468
rect 9048 2437 9076 2468
rect 9858 2456 9864 2508
rect 9916 2496 9922 2508
rect 10229 2499 10287 2505
rect 10229 2496 10241 2499
rect 9916 2468 10241 2496
rect 9916 2456 9922 2468
rect 10229 2465 10241 2468
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 10318 2456 10324 2508
rect 10376 2456 10382 2508
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12989 2499 13047 2505
rect 12989 2496 13001 2499
rect 12584 2468 13001 2496
rect 12584 2456 12590 2468
rect 12989 2465 13001 2468
rect 13035 2465 13047 2499
rect 13906 2496 13912 2508
rect 13867 2468 13912 2496
rect 12989 2459 13047 2465
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 15470 2456 15476 2508
rect 15528 2496 15534 2508
rect 17788 2505 17816 2536
rect 20165 2533 20177 2567
rect 20211 2564 20223 2567
rect 20438 2564 20444 2576
rect 20211 2536 20444 2564
rect 20211 2533 20223 2536
rect 20165 2527 20223 2533
rect 20438 2524 20444 2536
rect 20496 2524 20502 2576
rect 18598 2505 18604 2508
rect 15933 2499 15991 2505
rect 15933 2496 15945 2499
rect 15528 2468 15945 2496
rect 15528 2456 15534 2468
rect 15933 2465 15945 2468
rect 15979 2465 15991 2499
rect 15933 2459 15991 2465
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2465 17831 2499
rect 17773 2459 17831 2465
rect 17865 2499 17923 2505
rect 17865 2465 17877 2499
rect 17911 2496 17923 2499
rect 18592 2496 18604 2505
rect 17911 2468 18604 2496
rect 17911 2465 17923 2468
rect 17865 2459 17923 2465
rect 18592 2459 18604 2468
rect 18598 2456 18604 2459
rect 18656 2456 18662 2508
rect 8849 2431 8907 2437
rect 8849 2428 8861 2431
rect 7944 2400 8861 2428
rect 6641 2391 6699 2397
rect 8849 2397 8861 2400
rect 8895 2397 8907 2431
rect 8849 2391 8907 2397
rect 9033 2431 9091 2437
rect 9033 2397 9045 2431
rect 9079 2428 9091 2431
rect 10336 2428 10364 2456
rect 9079 2400 10364 2428
rect 12345 2431 12403 2437
rect 9079 2397 9091 2400
rect 9033 2391 9091 2397
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 13078 2428 13084 2440
rect 12391 2400 13084 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 13262 2428 13268 2440
rect 13223 2400 13268 2428
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 18046 2428 18052 2440
rect 18007 2400 18052 2428
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 18325 2431 18383 2437
rect 18325 2397 18337 2431
rect 18371 2397 18383 2431
rect 20349 2431 20407 2437
rect 20349 2428 20361 2431
rect 18325 2391 18383 2397
rect 19352 2400 20361 2428
rect 8386 2360 8392 2372
rect 8347 2332 8392 2360
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 17678 2320 17684 2372
rect 17736 2360 17742 2372
rect 18340 2360 18368 2391
rect 17736 2332 18368 2360
rect 17736 2320 17742 2332
rect 5261 2295 5319 2301
rect 5261 2261 5273 2295
rect 5307 2292 5319 2295
rect 5350 2292 5356 2304
rect 5307 2264 5356 2292
rect 5307 2261 5319 2264
rect 5261 2255 5319 2261
rect 5350 2252 5356 2264
rect 5408 2252 5414 2304
rect 5997 2295 6055 2301
rect 5997 2261 6009 2295
rect 6043 2292 6055 2295
rect 7190 2292 7196 2304
rect 6043 2264 7196 2292
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 11698 2292 11704 2304
rect 11659 2264 11704 2292
rect 11698 2252 11704 2264
rect 11756 2252 11762 2304
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 19352 2292 19380 2400
rect 20349 2397 20361 2400
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 18104 2264 19380 2292
rect 18104 2252 18110 2264
rect 1104 2202 20884 2224
rect 1104 2150 4280 2202
rect 4332 2150 4344 2202
rect 4396 2150 4408 2202
rect 4460 2150 4472 2202
rect 4524 2150 10878 2202
rect 10930 2150 10942 2202
rect 10994 2150 11006 2202
rect 11058 2150 11070 2202
rect 11122 2150 17475 2202
rect 17527 2150 17539 2202
rect 17591 2150 17603 2202
rect 17655 2150 17667 2202
rect 17719 2150 20884 2202
rect 1104 2128 20884 2150
rect 1762 1232 1768 1284
rect 1820 1272 1826 1284
rect 9582 1272 9588 1284
rect 1820 1244 9588 1272
rect 1820 1232 1826 1244
rect 9582 1232 9588 1244
rect 9640 1232 9646 1284
<< via1 >>
rect 9496 19660 9548 19712
rect 15384 19660 15436 19712
rect 16028 19660 16080 19712
rect 19708 19660 19760 19712
rect 4280 19558 4332 19610
rect 4344 19558 4396 19610
rect 4408 19558 4460 19610
rect 4472 19558 4524 19610
rect 10878 19558 10930 19610
rect 10942 19558 10994 19610
rect 11006 19558 11058 19610
rect 11070 19558 11122 19610
rect 17475 19558 17527 19610
rect 17539 19558 17591 19610
rect 17603 19558 17655 19610
rect 17667 19558 17719 19610
rect 1584 19252 1636 19304
rect 4896 19388 4948 19440
rect 7472 19456 7524 19508
rect 9864 19456 9916 19508
rect 15200 19456 15252 19508
rect 5080 19320 5132 19372
rect 5448 19363 5500 19372
rect 5448 19329 5457 19363
rect 5457 19329 5491 19363
rect 5491 19329 5500 19363
rect 5448 19320 5500 19329
rect 4160 19252 4212 19304
rect 6552 19320 6604 19372
rect 8208 19363 8260 19372
rect 8208 19329 8217 19363
rect 8217 19329 8251 19363
rect 8251 19329 8260 19363
rect 8208 19320 8260 19329
rect 9496 19363 9548 19372
rect 9496 19329 9505 19363
rect 9505 19329 9539 19363
rect 9539 19329 9548 19363
rect 9496 19320 9548 19329
rect 1492 19184 1544 19236
rect 1676 19159 1728 19168
rect 1676 19125 1685 19159
rect 1685 19125 1719 19159
rect 1719 19125 1728 19159
rect 1676 19116 1728 19125
rect 2136 19159 2188 19168
rect 2136 19125 2145 19159
rect 2145 19125 2179 19159
rect 2179 19125 2188 19159
rect 2136 19116 2188 19125
rect 2596 19116 2648 19168
rect 2872 19159 2924 19168
rect 2872 19125 2881 19159
rect 2881 19125 2915 19159
rect 2915 19125 2924 19159
rect 2872 19116 2924 19125
rect 3056 19116 3108 19168
rect 3608 19184 3660 19236
rect 4804 19184 4856 19236
rect 6460 19252 6512 19304
rect 7564 19252 7616 19304
rect 9680 19252 9732 19304
rect 11244 19320 11296 19372
rect 12072 19320 12124 19372
rect 12256 19320 12308 19372
rect 11980 19252 12032 19304
rect 12440 19252 12492 19304
rect 12716 19295 12768 19304
rect 12716 19261 12725 19295
rect 12725 19261 12759 19295
rect 12759 19261 12768 19295
rect 12716 19252 12768 19261
rect 14924 19320 14976 19372
rect 16948 19320 17000 19372
rect 17684 19363 17736 19372
rect 17684 19329 17693 19363
rect 17693 19329 17727 19363
rect 17727 19329 17736 19363
rect 17684 19320 17736 19329
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 19708 19363 19760 19372
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 12992 19227 13044 19236
rect 4068 19159 4120 19168
rect 4068 19125 4077 19159
rect 4077 19125 4111 19159
rect 4111 19125 4120 19159
rect 4068 19116 4120 19125
rect 4160 19116 4212 19168
rect 4712 19116 4764 19168
rect 5264 19159 5316 19168
rect 5264 19125 5273 19159
rect 5273 19125 5307 19159
rect 5307 19125 5316 19159
rect 5264 19116 5316 19125
rect 6276 19116 6328 19168
rect 6828 19116 6880 19168
rect 7104 19159 7156 19168
rect 7104 19125 7113 19159
rect 7113 19125 7147 19159
rect 7147 19125 7156 19159
rect 7104 19116 7156 19125
rect 8024 19159 8076 19168
rect 8024 19125 8033 19159
rect 8033 19125 8067 19159
rect 8067 19125 8076 19159
rect 8024 19116 8076 19125
rect 8116 19159 8168 19168
rect 8116 19125 8125 19159
rect 8125 19125 8159 19159
rect 8159 19125 8168 19159
rect 8116 19116 8168 19125
rect 8300 19116 8352 19168
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 9864 19116 9916 19168
rect 9956 19159 10008 19168
rect 9956 19125 9965 19159
rect 9965 19125 9999 19159
rect 9999 19125 10008 19159
rect 10324 19159 10376 19168
rect 9956 19116 10008 19125
rect 10324 19125 10333 19159
rect 10333 19125 10367 19159
rect 10367 19125 10376 19159
rect 10324 19116 10376 19125
rect 10508 19116 10560 19168
rect 11060 19116 11112 19168
rect 11152 19159 11204 19168
rect 11152 19125 11161 19159
rect 11161 19125 11195 19159
rect 11195 19125 11204 19159
rect 11520 19159 11572 19168
rect 11152 19116 11204 19125
rect 11520 19125 11529 19159
rect 11529 19125 11563 19159
rect 11563 19125 11572 19159
rect 11520 19116 11572 19125
rect 12256 19116 12308 19168
rect 12532 19116 12584 19168
rect 12624 19159 12676 19168
rect 12624 19125 12633 19159
rect 12633 19125 12667 19159
rect 12667 19125 12676 19159
rect 12992 19193 13026 19227
rect 13026 19193 13044 19227
rect 12992 19184 13044 19193
rect 14188 19252 14240 19304
rect 15108 19252 15160 19304
rect 15568 19252 15620 19304
rect 16212 19252 16264 19304
rect 16672 19252 16724 19304
rect 20720 19252 20772 19304
rect 15844 19184 15896 19236
rect 12624 19116 12676 19125
rect 13912 19116 13964 19168
rect 14004 19116 14056 19168
rect 14464 19116 14516 19168
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 16580 19184 16632 19236
rect 16120 19116 16172 19168
rect 17316 19116 17368 19168
rect 17592 19159 17644 19168
rect 17592 19125 17601 19159
rect 17601 19125 17635 19159
rect 17635 19125 17644 19159
rect 17592 19116 17644 19125
rect 18052 19116 18104 19168
rect 18696 19159 18748 19168
rect 18696 19125 18705 19159
rect 18705 19125 18739 19159
rect 18739 19125 18748 19159
rect 18696 19116 18748 19125
rect 19156 19159 19208 19168
rect 19156 19125 19165 19159
rect 19165 19125 19199 19159
rect 19199 19125 19208 19159
rect 19156 19116 19208 19125
rect 7579 19014 7631 19066
rect 7643 19014 7695 19066
rect 7707 19014 7759 19066
rect 7771 19014 7823 19066
rect 14176 19014 14228 19066
rect 14240 19014 14292 19066
rect 14304 19014 14356 19066
rect 14368 19014 14420 19066
rect 848 18912 900 18964
rect 1676 18912 1728 18964
rect 3148 18912 3200 18964
rect 3608 18912 3660 18964
rect 4620 18912 4672 18964
rect 4896 18912 4948 18964
rect 8024 18912 8076 18964
rect 9128 18912 9180 18964
rect 10324 18912 10376 18964
rect 10876 18912 10928 18964
rect 11060 18912 11112 18964
rect 11612 18912 11664 18964
rect 12992 18912 13044 18964
rect 13820 18912 13872 18964
rect 14648 18912 14700 18964
rect 15844 18912 15896 18964
rect 16580 18912 16632 18964
rect 16948 18912 17000 18964
rect 17132 18955 17184 18964
rect 17132 18921 17141 18955
rect 17141 18921 17175 18955
rect 17175 18921 17184 18955
rect 17132 18912 17184 18921
rect 17592 18912 17644 18964
rect 11428 18844 11480 18896
rect 11520 18844 11572 18896
rect 2228 18776 2280 18828
rect 2412 18819 2464 18828
rect 2412 18785 2446 18819
rect 2446 18785 2464 18819
rect 2412 18776 2464 18785
rect 3608 18819 3660 18828
rect 3608 18785 3617 18819
rect 3617 18785 3651 18819
rect 3651 18785 3660 18819
rect 3608 18776 3660 18785
rect 4335 18819 4387 18828
rect 4335 18785 4344 18819
rect 4344 18785 4378 18819
rect 4378 18785 4387 18819
rect 4335 18776 4387 18785
rect 296 18572 348 18624
rect 3884 18572 3936 18624
rect 6276 18776 6328 18828
rect 8024 18776 8076 18828
rect 9956 18776 10008 18828
rect 10324 18776 10376 18828
rect 10784 18776 10836 18828
rect 11336 18776 11388 18828
rect 16120 18844 16172 18896
rect 16488 18844 16540 18896
rect 20996 18912 21048 18964
rect 12532 18776 12584 18828
rect 12716 18776 12768 18828
rect 14280 18776 14332 18828
rect 14372 18776 14424 18828
rect 14740 18776 14792 18828
rect 5264 18572 5316 18624
rect 7104 18708 7156 18760
rect 9312 18751 9364 18760
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 10140 18751 10192 18760
rect 10140 18717 10149 18751
rect 10149 18717 10183 18751
rect 10183 18717 10192 18751
rect 10140 18708 10192 18717
rect 10232 18751 10284 18760
rect 10232 18717 10241 18751
rect 10241 18717 10275 18751
rect 10275 18717 10284 18751
rect 10232 18708 10284 18717
rect 13636 18708 13688 18760
rect 14924 18708 14976 18760
rect 6460 18572 6512 18624
rect 10416 18640 10468 18692
rect 13820 18640 13872 18692
rect 16764 18776 16816 18828
rect 16948 18776 17000 18828
rect 17684 18776 17736 18828
rect 15660 18708 15712 18760
rect 16856 18708 16908 18760
rect 18328 18776 18380 18828
rect 19432 18776 19484 18828
rect 19708 18776 19760 18828
rect 20812 18776 20864 18828
rect 8208 18572 8260 18624
rect 9036 18572 9088 18624
rect 12072 18615 12124 18624
rect 12072 18581 12081 18615
rect 12081 18581 12115 18615
rect 12115 18581 12124 18615
rect 12072 18572 12124 18581
rect 12164 18572 12216 18624
rect 13268 18572 13320 18624
rect 15660 18615 15712 18624
rect 15660 18581 15669 18615
rect 15669 18581 15703 18615
rect 15703 18581 15712 18615
rect 15660 18572 15712 18581
rect 15752 18572 15804 18624
rect 18236 18708 18288 18760
rect 17868 18572 17920 18624
rect 21640 18640 21692 18692
rect 19156 18572 19208 18624
rect 4280 18470 4332 18522
rect 4344 18470 4396 18522
rect 4408 18470 4460 18522
rect 4472 18470 4524 18522
rect 10878 18470 10930 18522
rect 10942 18470 10994 18522
rect 11006 18470 11058 18522
rect 11070 18470 11122 18522
rect 17475 18470 17527 18522
rect 17539 18470 17591 18522
rect 17603 18470 17655 18522
rect 17667 18470 17719 18522
rect 2412 18368 2464 18420
rect 3884 18368 3936 18420
rect 4160 18368 4212 18420
rect 9036 18368 9088 18420
rect 5080 18275 5132 18284
rect 5080 18241 5089 18275
rect 5089 18241 5123 18275
rect 5123 18241 5132 18275
rect 5080 18232 5132 18241
rect 5264 18275 5316 18284
rect 5264 18241 5273 18275
rect 5273 18241 5307 18275
rect 5307 18241 5316 18275
rect 5264 18232 5316 18241
rect 6368 18232 6420 18284
rect 7288 18300 7340 18352
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 2228 18164 2280 18216
rect 2780 18096 2832 18148
rect 3516 18164 3568 18216
rect 3608 18164 3660 18216
rect 6460 18164 6512 18216
rect 6920 18232 6972 18284
rect 10232 18368 10284 18420
rect 11428 18368 11480 18420
rect 12348 18368 12400 18420
rect 5724 18096 5776 18148
rect 4160 18028 4212 18080
rect 4804 18071 4856 18080
rect 4804 18037 4813 18071
rect 4813 18037 4847 18071
rect 4847 18037 4856 18071
rect 4804 18028 4856 18037
rect 4988 18028 5040 18080
rect 8484 18164 8536 18216
rect 9036 18164 9088 18216
rect 10416 18232 10468 18284
rect 14280 18368 14332 18420
rect 15292 18300 15344 18352
rect 10784 18207 10836 18216
rect 10784 18173 10793 18207
rect 10793 18173 10827 18207
rect 10827 18173 10836 18207
rect 10784 18164 10836 18173
rect 12532 18164 12584 18216
rect 14096 18232 14148 18284
rect 15844 18300 15896 18352
rect 17316 18343 17368 18352
rect 17316 18309 17325 18343
rect 17325 18309 17359 18343
rect 17359 18309 17368 18343
rect 17316 18300 17368 18309
rect 17776 18343 17828 18352
rect 17776 18309 17785 18343
rect 17785 18309 17819 18343
rect 17819 18309 17828 18343
rect 17776 18300 17828 18309
rect 19432 18343 19484 18352
rect 19432 18309 19441 18343
rect 19441 18309 19475 18343
rect 19475 18309 19484 18343
rect 19432 18300 19484 18309
rect 20996 18343 21048 18352
rect 20996 18309 21005 18343
rect 21005 18309 21039 18343
rect 21039 18309 21048 18343
rect 20996 18300 21048 18309
rect 14004 18164 14056 18216
rect 14740 18207 14792 18216
rect 14740 18173 14749 18207
rect 14749 18173 14783 18207
rect 14783 18173 14792 18207
rect 14740 18164 14792 18173
rect 15200 18164 15252 18216
rect 15752 18164 15804 18216
rect 16028 18164 16080 18216
rect 17132 18164 17184 18216
rect 17868 18164 17920 18216
rect 18144 18164 18196 18216
rect 8208 18096 8260 18148
rect 8852 18096 8904 18148
rect 10876 18096 10928 18148
rect 11244 18096 11296 18148
rect 14280 18139 14332 18148
rect 14280 18105 14289 18139
rect 14289 18105 14323 18139
rect 14323 18105 14332 18139
rect 14280 18096 14332 18105
rect 18328 18139 18380 18148
rect 18328 18105 18362 18139
rect 18362 18105 18380 18139
rect 18328 18096 18380 18105
rect 9220 18028 9272 18080
rect 9312 18028 9364 18080
rect 12900 18028 12952 18080
rect 13544 18028 13596 18080
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 13912 18071 13964 18080
rect 13912 18037 13921 18071
rect 13921 18037 13955 18071
rect 13955 18037 13964 18071
rect 13912 18028 13964 18037
rect 17224 18028 17276 18080
rect 17684 18028 17736 18080
rect 19248 18096 19300 18148
rect 19432 18028 19484 18080
rect 7579 17926 7631 17978
rect 7643 17926 7695 17978
rect 7707 17926 7759 17978
rect 7771 17926 7823 17978
rect 14176 17926 14228 17978
rect 14240 17926 14292 17978
rect 14304 17926 14356 17978
rect 14368 17926 14420 17978
rect 2780 17867 2832 17876
rect 2780 17833 2789 17867
rect 2789 17833 2823 17867
rect 2823 17833 2832 17867
rect 2780 17824 2832 17833
rect 4068 17824 4120 17876
rect 4896 17824 4948 17876
rect 3976 17756 4028 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 1676 17731 1728 17740
rect 1676 17697 1710 17731
rect 1710 17697 1728 17731
rect 1676 17688 1728 17697
rect 4988 17756 5040 17808
rect 6276 17799 6328 17808
rect 6276 17765 6285 17799
rect 6285 17765 6319 17799
rect 6319 17765 6328 17799
rect 6276 17756 6328 17765
rect 6736 17756 6788 17808
rect 6920 17799 6972 17808
rect 6920 17765 6954 17799
rect 6954 17765 6972 17799
rect 6920 17756 6972 17765
rect 7932 17756 7984 17808
rect 9128 17824 9180 17876
rect 11244 17867 11296 17876
rect 11244 17833 11253 17867
rect 11253 17833 11287 17867
rect 11287 17833 11296 17867
rect 11244 17824 11296 17833
rect 12440 17824 12492 17876
rect 14004 17824 14056 17876
rect 3884 17620 3936 17672
rect 4620 17620 4672 17672
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 2412 17552 2464 17604
rect 5540 17620 5592 17672
rect 5908 17688 5960 17740
rect 7288 17688 7340 17740
rect 8852 17688 8904 17740
rect 9404 17756 9456 17808
rect 11336 17756 11388 17808
rect 12072 17756 12124 17808
rect 12348 17756 12400 17808
rect 9588 17688 9640 17740
rect 5816 17663 5868 17672
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 6644 17663 6696 17672
rect 6644 17629 6653 17663
rect 6653 17629 6687 17663
rect 6687 17629 6696 17663
rect 6644 17620 6696 17629
rect 8024 17595 8076 17604
rect 1584 17484 1636 17536
rect 8024 17561 8033 17595
rect 8033 17561 8067 17595
rect 8067 17561 8076 17595
rect 8024 17552 8076 17561
rect 8116 17595 8168 17604
rect 8116 17561 8125 17595
rect 8125 17561 8159 17595
rect 8159 17561 8168 17595
rect 8116 17552 8168 17561
rect 9680 17620 9732 17672
rect 9036 17552 9088 17604
rect 11244 17620 11296 17672
rect 12992 17620 13044 17672
rect 14096 17756 14148 17808
rect 14832 17756 14884 17808
rect 14740 17731 14792 17740
rect 13636 17620 13688 17672
rect 12716 17595 12768 17604
rect 12716 17561 12725 17595
rect 12725 17561 12759 17595
rect 12759 17561 12768 17595
rect 12716 17552 12768 17561
rect 14740 17697 14749 17731
rect 14749 17697 14783 17731
rect 14783 17697 14792 17731
rect 14740 17688 14792 17697
rect 14556 17620 14608 17672
rect 15476 17824 15528 17876
rect 15936 17824 15988 17876
rect 16120 17824 16172 17876
rect 16488 17867 16540 17876
rect 16488 17833 16497 17867
rect 16497 17833 16531 17867
rect 16531 17833 16540 17867
rect 16488 17824 16540 17833
rect 18052 17824 18104 17876
rect 18328 17824 18380 17876
rect 17960 17756 18012 17808
rect 18144 17756 18196 17808
rect 19892 17756 19944 17808
rect 16212 17688 16264 17740
rect 17776 17688 17828 17740
rect 15844 17620 15896 17672
rect 16396 17620 16448 17672
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 17684 17663 17736 17672
rect 16580 17620 16632 17629
rect 17684 17629 17693 17663
rect 17693 17629 17727 17663
rect 17727 17629 17736 17663
rect 17684 17620 17736 17629
rect 19432 17688 19484 17740
rect 20260 17731 20312 17740
rect 20260 17697 20269 17731
rect 20269 17697 20303 17731
rect 20303 17697 20312 17731
rect 20260 17688 20312 17697
rect 19156 17620 19208 17672
rect 20076 17663 20128 17672
rect 20076 17629 20085 17663
rect 20085 17629 20119 17663
rect 20119 17629 20128 17663
rect 20076 17620 20128 17629
rect 16672 17552 16724 17604
rect 20996 17552 21048 17604
rect 9128 17527 9180 17536
rect 9128 17493 9137 17527
rect 9137 17493 9171 17527
rect 9171 17493 9180 17527
rect 9128 17484 9180 17493
rect 14832 17484 14884 17536
rect 16120 17484 16172 17536
rect 19156 17484 19208 17536
rect 4280 17382 4332 17434
rect 4344 17382 4396 17434
rect 4408 17382 4460 17434
rect 4472 17382 4524 17434
rect 10878 17382 10930 17434
rect 10942 17382 10994 17434
rect 11006 17382 11058 17434
rect 11070 17382 11122 17434
rect 17475 17382 17527 17434
rect 17539 17382 17591 17434
rect 17603 17382 17655 17434
rect 17667 17382 17719 17434
rect 5724 17323 5776 17332
rect 5724 17289 5733 17323
rect 5733 17289 5767 17323
rect 5767 17289 5776 17323
rect 5724 17280 5776 17289
rect 5816 17280 5868 17332
rect 8668 17280 8720 17332
rect 1768 17212 1820 17264
rect 3884 17187 3936 17196
rect 3884 17153 3893 17187
rect 3893 17153 3927 17187
rect 3927 17153 3936 17187
rect 3884 17144 3936 17153
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 4988 17144 5040 17196
rect 5356 17144 5408 17196
rect 5540 17144 5592 17196
rect 5724 17144 5776 17196
rect 6460 17144 6512 17196
rect 6736 17144 6788 17196
rect 1308 17076 1360 17128
rect 1492 17076 1544 17128
rect 3148 17076 3200 17128
rect 4160 17076 4212 17128
rect 5080 17076 5132 17128
rect 6644 17076 6696 17128
rect 6920 17119 6972 17128
rect 6920 17085 6929 17119
rect 6929 17085 6963 17119
rect 6963 17085 6972 17119
rect 6920 17076 6972 17085
rect 7932 17144 7984 17196
rect 8484 17076 8536 17128
rect 2136 17008 2188 17060
rect 2688 17008 2740 17060
rect 3516 17008 3568 17060
rect 4344 17008 4396 17060
rect 7472 17008 7524 17060
rect 9312 17076 9364 17128
rect 10784 17212 10836 17264
rect 11244 17280 11296 17332
rect 12532 17280 12584 17332
rect 13268 17323 13320 17332
rect 13268 17289 13277 17323
rect 13277 17289 13311 17323
rect 13311 17289 13320 17323
rect 13268 17280 13320 17289
rect 17776 17323 17828 17332
rect 17776 17289 17785 17323
rect 17785 17289 17819 17323
rect 17819 17289 17828 17323
rect 17776 17280 17828 17289
rect 19432 17323 19484 17332
rect 9956 17144 10008 17196
rect 13176 17144 13228 17196
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 15292 17212 15344 17264
rect 19432 17289 19441 17323
rect 19441 17289 19475 17323
rect 19475 17289 19484 17323
rect 19432 17280 19484 17289
rect 19800 17280 19852 17332
rect 15200 17144 15252 17196
rect 13636 17119 13688 17128
rect 1676 16940 1728 16992
rect 3240 16983 3292 16992
rect 3240 16949 3249 16983
rect 3249 16949 3283 16983
rect 3283 16949 3292 16983
rect 4068 16983 4120 16992
rect 3240 16940 3292 16949
rect 4068 16949 4077 16983
rect 4077 16949 4111 16983
rect 4111 16949 4120 16983
rect 4068 16940 4120 16949
rect 4620 16940 4672 16992
rect 4988 16940 5040 16992
rect 5632 16940 5684 16992
rect 6092 16983 6144 16992
rect 6092 16949 6101 16983
rect 6101 16949 6135 16983
rect 6135 16949 6144 16983
rect 6092 16940 6144 16949
rect 7932 16940 7984 16992
rect 8024 16940 8076 16992
rect 9864 17008 9916 17060
rect 9956 17008 10008 17060
rect 10600 17008 10652 17060
rect 11428 17008 11480 17060
rect 11520 17008 11572 17060
rect 12992 17008 13044 17060
rect 13636 17085 13645 17119
rect 13645 17085 13679 17119
rect 13679 17085 13688 17119
rect 13636 17076 13688 17085
rect 13912 17076 13964 17128
rect 15476 17076 15528 17128
rect 16028 17144 16080 17196
rect 16580 17144 16632 17196
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 16764 17076 16816 17128
rect 18144 17076 18196 17128
rect 19248 17076 19300 17128
rect 19524 17076 19576 17128
rect 14096 17008 14148 17060
rect 14464 17051 14516 17060
rect 14464 17017 14498 17051
rect 14498 17017 14516 17051
rect 14464 17008 14516 17017
rect 19800 17008 19852 17060
rect 10232 16940 10284 16992
rect 10692 16940 10744 16992
rect 11980 16940 12032 16992
rect 12256 16983 12308 16992
rect 12256 16949 12265 16983
rect 12265 16949 12299 16983
rect 12299 16949 12308 16983
rect 12256 16940 12308 16949
rect 12348 16940 12400 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 14004 16940 14056 16992
rect 15476 16940 15528 16992
rect 15660 16940 15712 16992
rect 16672 16940 16724 16992
rect 17040 16983 17092 16992
rect 17040 16949 17049 16983
rect 17049 16949 17083 16983
rect 17083 16949 17092 16983
rect 17040 16940 17092 16949
rect 17316 16940 17368 16992
rect 20076 16940 20128 16992
rect 7579 16838 7631 16890
rect 7643 16838 7695 16890
rect 7707 16838 7759 16890
rect 7771 16838 7823 16890
rect 14176 16838 14228 16890
rect 14240 16838 14292 16890
rect 14304 16838 14356 16890
rect 14368 16838 14420 16890
rect 2320 16736 2372 16788
rect 2044 16711 2096 16720
rect 2044 16677 2078 16711
rect 2078 16677 2096 16711
rect 2044 16668 2096 16677
rect 2136 16668 2188 16720
rect 1492 16600 1544 16652
rect 1860 16600 1912 16652
rect 3516 16736 3568 16788
rect 4344 16779 4396 16788
rect 4344 16745 4353 16779
rect 4353 16745 4387 16779
rect 4387 16745 4396 16779
rect 4344 16736 4396 16745
rect 3976 16668 4028 16720
rect 4896 16711 4948 16720
rect 4896 16677 4905 16711
rect 4905 16677 4939 16711
rect 4939 16677 4948 16711
rect 4896 16668 4948 16677
rect 3700 16600 3752 16652
rect 4160 16643 4212 16652
rect 4160 16609 4169 16643
rect 4169 16609 4203 16643
rect 4203 16609 4212 16643
rect 4160 16600 4212 16609
rect 1584 16532 1636 16584
rect 3332 16464 3384 16516
rect 5632 16736 5684 16788
rect 6920 16736 6972 16788
rect 7104 16736 7156 16788
rect 7288 16779 7340 16788
rect 7288 16745 7297 16779
rect 7297 16745 7331 16779
rect 7331 16745 7340 16779
rect 7288 16736 7340 16745
rect 8392 16736 8444 16788
rect 8668 16736 8720 16788
rect 8852 16736 8904 16788
rect 11612 16779 11664 16788
rect 5816 16643 5868 16652
rect 5816 16609 5825 16643
rect 5825 16609 5859 16643
rect 5859 16609 5868 16643
rect 11612 16745 11621 16779
rect 11621 16745 11655 16779
rect 11655 16745 11664 16779
rect 11612 16736 11664 16745
rect 11980 16779 12032 16788
rect 11980 16745 11989 16779
rect 11989 16745 12023 16779
rect 12023 16745 12032 16779
rect 11980 16736 12032 16745
rect 12900 16736 12952 16788
rect 13544 16736 13596 16788
rect 5816 16600 5868 16609
rect 7104 16600 7156 16652
rect 11520 16668 11572 16720
rect 13820 16668 13872 16720
rect 14556 16736 14608 16788
rect 14740 16736 14792 16788
rect 15476 16736 15528 16788
rect 17316 16736 17368 16788
rect 17960 16736 18012 16788
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 4712 16532 4764 16584
rect 6000 16575 6052 16584
rect 6000 16541 6009 16575
rect 6009 16541 6043 16575
rect 6043 16541 6052 16575
rect 7472 16575 7524 16584
rect 6000 16532 6052 16541
rect 7196 16464 7248 16516
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 8024 16532 8076 16584
rect 8116 16575 8168 16584
rect 8116 16541 8128 16575
rect 8128 16541 8162 16575
rect 8162 16541 8168 16575
rect 8116 16532 8168 16541
rect 8300 16532 8352 16584
rect 9588 16532 9640 16584
rect 2964 16396 3016 16448
rect 6092 16396 6144 16448
rect 7288 16396 7340 16448
rect 9128 16396 9180 16448
rect 9864 16532 9916 16584
rect 12532 16643 12584 16652
rect 12532 16609 12541 16643
rect 12541 16609 12575 16643
rect 12575 16609 12584 16643
rect 12532 16600 12584 16609
rect 12624 16600 12676 16652
rect 14464 16668 14516 16720
rect 14832 16643 14884 16652
rect 12072 16575 12124 16584
rect 12072 16541 12081 16575
rect 12081 16541 12115 16575
rect 12115 16541 12124 16575
rect 12072 16532 12124 16541
rect 11336 16464 11388 16516
rect 10324 16396 10376 16448
rect 11520 16439 11572 16448
rect 11520 16405 11529 16439
rect 11529 16405 11563 16439
rect 11563 16405 11572 16439
rect 11520 16396 11572 16405
rect 13820 16532 13872 16584
rect 14832 16609 14841 16643
rect 14841 16609 14875 16643
rect 14875 16609 14884 16643
rect 14832 16600 14884 16609
rect 15660 16643 15712 16652
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 15936 16600 15988 16652
rect 16672 16643 16724 16652
rect 16672 16609 16706 16643
rect 16706 16609 16724 16643
rect 16672 16600 16724 16609
rect 18052 16668 18104 16720
rect 18236 16668 18288 16720
rect 19616 16600 19668 16652
rect 20628 16600 20680 16652
rect 13912 16507 13964 16516
rect 13912 16473 13921 16507
rect 13921 16473 13955 16507
rect 13955 16473 13964 16507
rect 13912 16464 13964 16473
rect 14924 16464 14976 16516
rect 19432 16532 19484 16584
rect 20076 16532 20128 16584
rect 18880 16464 18932 16516
rect 19708 16464 19760 16516
rect 16580 16396 16632 16448
rect 19340 16439 19392 16448
rect 19340 16405 19349 16439
rect 19349 16405 19383 16439
rect 19383 16405 19392 16439
rect 19340 16396 19392 16405
rect 4280 16294 4332 16346
rect 4344 16294 4396 16346
rect 4408 16294 4460 16346
rect 4472 16294 4524 16346
rect 10878 16294 10930 16346
rect 10942 16294 10994 16346
rect 11006 16294 11058 16346
rect 11070 16294 11122 16346
rect 17475 16294 17527 16346
rect 17539 16294 17591 16346
rect 17603 16294 17655 16346
rect 17667 16294 17719 16346
rect 3424 16124 3476 16176
rect 4160 16192 4212 16244
rect 4988 16192 5040 16244
rect 5724 16192 5776 16244
rect 7932 16192 7984 16244
rect 8760 16192 8812 16244
rect 10140 16192 10192 16244
rect 12072 16192 12124 16244
rect 1860 16099 1912 16108
rect 1860 16065 1869 16099
rect 1869 16065 1903 16099
rect 1903 16065 1912 16099
rect 1860 16056 1912 16065
rect 3608 16056 3660 16108
rect 4068 16099 4120 16108
rect 4068 16065 4077 16099
rect 4077 16065 4111 16099
rect 4111 16065 4120 16099
rect 4068 16056 4120 16065
rect 3700 15988 3752 16040
rect 3884 15988 3936 16040
rect 4252 16056 4304 16108
rect 2596 15920 2648 15972
rect 5540 15988 5592 16040
rect 7288 16056 7340 16108
rect 7840 16099 7892 16108
rect 7840 16065 7849 16099
rect 7849 16065 7883 16099
rect 7883 16065 7892 16099
rect 7840 16056 7892 16065
rect 8852 16099 8904 16108
rect 2964 15852 3016 15904
rect 4068 15852 4120 15904
rect 4712 15852 4764 15904
rect 6828 15920 6880 15972
rect 7104 15988 7156 16040
rect 8024 15988 8076 16040
rect 8392 15988 8444 16040
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 10508 16056 10560 16108
rect 10784 16099 10836 16108
rect 10784 16065 10796 16099
rect 10796 16065 10830 16099
rect 10830 16065 10836 16099
rect 10784 16056 10836 16065
rect 12624 16056 12676 16108
rect 10232 15988 10284 16040
rect 10324 16031 10376 16040
rect 10324 15997 10333 16031
rect 10333 15997 10367 16031
rect 10367 15997 10376 16031
rect 10324 15988 10376 15997
rect 13084 16192 13136 16244
rect 14004 16192 14056 16244
rect 14924 16192 14976 16244
rect 15660 16192 15712 16244
rect 16672 16192 16724 16244
rect 18052 16192 18104 16244
rect 17132 16124 17184 16176
rect 15936 16056 15988 16108
rect 20076 16099 20128 16108
rect 20076 16065 20085 16099
rect 20085 16065 20119 16099
rect 20119 16065 20128 16099
rect 20076 16056 20128 16065
rect 7932 15920 7984 15972
rect 12532 15920 12584 15972
rect 12716 15920 12768 15972
rect 13912 15988 13964 16040
rect 12992 15920 13044 15972
rect 14096 15920 14148 15972
rect 14648 15920 14700 15972
rect 6000 15852 6052 15904
rect 6184 15895 6236 15904
rect 6184 15861 6193 15895
rect 6193 15861 6227 15895
rect 6227 15861 6236 15895
rect 6184 15852 6236 15861
rect 8392 15852 8444 15904
rect 8668 15852 8720 15904
rect 9588 15852 9640 15904
rect 15752 15988 15804 16040
rect 17040 15988 17092 16040
rect 17224 15988 17276 16040
rect 18144 15988 18196 16040
rect 18604 15988 18656 16040
rect 14924 15920 14976 15972
rect 15568 15920 15620 15972
rect 17960 15920 18012 15972
rect 18696 15920 18748 15972
rect 15476 15852 15528 15904
rect 20352 15920 20404 15972
rect 19984 15895 20036 15904
rect 19984 15861 19993 15895
rect 19993 15861 20027 15895
rect 20027 15861 20036 15895
rect 19984 15852 20036 15861
rect 7579 15750 7631 15802
rect 7643 15750 7695 15802
rect 7707 15750 7759 15802
rect 7771 15750 7823 15802
rect 14176 15750 14228 15802
rect 14240 15750 14292 15802
rect 14304 15750 14356 15802
rect 14368 15750 14420 15802
rect 4804 15648 4856 15700
rect 2872 15580 2924 15632
rect 4620 15580 4672 15632
rect 6184 15580 6236 15632
rect 1860 15512 1912 15564
rect 3240 15555 3292 15564
rect 3240 15521 3249 15555
rect 3249 15521 3283 15555
rect 3283 15521 3292 15555
rect 3240 15512 3292 15521
rect 5172 15512 5224 15564
rect 6920 15648 6972 15700
rect 7196 15648 7248 15700
rect 10692 15648 10744 15700
rect 11336 15648 11388 15700
rect 12256 15648 12308 15700
rect 14464 15648 14516 15700
rect 14740 15648 14792 15700
rect 15476 15648 15528 15700
rect 15936 15648 15988 15700
rect 17040 15648 17092 15700
rect 19432 15648 19484 15700
rect 19984 15691 20036 15700
rect 19984 15657 19993 15691
rect 19993 15657 20027 15691
rect 20027 15657 20036 15691
rect 19984 15648 20036 15657
rect 6828 15580 6880 15632
rect 11428 15580 11480 15632
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 6920 15512 6972 15564
rect 3608 15376 3660 15428
rect 6828 15376 6880 15428
rect 8300 15444 8352 15496
rect 9772 15512 9824 15564
rect 10232 15512 10284 15564
rect 10416 15512 10468 15564
rect 12440 15580 12492 15632
rect 13728 15580 13780 15632
rect 15016 15580 15068 15632
rect 15660 15580 15712 15632
rect 11796 15555 11848 15564
rect 11796 15521 11830 15555
rect 11830 15521 11848 15555
rect 11796 15512 11848 15521
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 11244 15487 11296 15496
rect 9680 15444 9732 15453
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 11244 15444 11296 15453
rect 13820 15512 13872 15564
rect 12992 15487 13044 15496
rect 12992 15453 13001 15487
rect 13001 15453 13035 15487
rect 13035 15453 13044 15487
rect 15292 15512 15344 15564
rect 16856 15512 16908 15564
rect 17316 15580 17368 15632
rect 18144 15512 18196 15564
rect 19616 15512 19668 15564
rect 20076 15555 20128 15564
rect 20076 15521 20085 15555
rect 20085 15521 20119 15555
rect 20119 15521 20128 15555
rect 20076 15512 20128 15521
rect 12992 15444 13044 15453
rect 15476 15487 15528 15496
rect 15476 15453 15485 15487
rect 15485 15453 15519 15487
rect 15519 15453 15528 15487
rect 15476 15444 15528 15453
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 4804 15308 4856 15360
rect 5080 15308 5132 15360
rect 6920 15351 6972 15360
rect 6920 15317 6929 15351
rect 6929 15317 6963 15351
rect 6963 15317 6972 15351
rect 6920 15308 6972 15317
rect 7656 15308 7708 15360
rect 8024 15308 8076 15360
rect 10324 15308 10376 15360
rect 12808 15308 12860 15360
rect 18880 15308 18932 15360
rect 4280 15206 4332 15258
rect 4344 15206 4396 15258
rect 4408 15206 4460 15258
rect 4472 15206 4524 15258
rect 10878 15206 10930 15258
rect 10942 15206 10994 15258
rect 11006 15206 11058 15258
rect 11070 15206 11122 15258
rect 17475 15206 17527 15258
rect 17539 15206 17591 15258
rect 17603 15206 17655 15258
rect 17667 15206 17719 15258
rect 1400 14968 1452 15020
rect 1860 15104 1912 15156
rect 2872 15147 2924 15156
rect 2872 15113 2881 15147
rect 2881 15113 2915 15147
rect 2915 15113 2924 15147
rect 2872 15104 2924 15113
rect 4068 15104 4120 15156
rect 4160 15104 4212 15156
rect 4620 15104 4672 15156
rect 5816 15104 5868 15156
rect 4896 15036 4948 15088
rect 9772 15104 9824 15156
rect 2964 14900 3016 14952
rect 3332 14900 3384 14952
rect 3516 14900 3568 14952
rect 5540 14968 5592 15020
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 9312 15036 9364 15088
rect 10784 15036 10836 15088
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 9680 14968 9732 15020
rect 7380 14900 7432 14952
rect 7656 14900 7708 14952
rect 8208 14900 8260 14952
rect 10140 14943 10192 14952
rect 10140 14909 10149 14943
rect 10149 14909 10183 14943
rect 10183 14909 10192 14943
rect 10140 14900 10192 14909
rect 10600 14968 10652 15020
rect 11428 15011 11480 15020
rect 11428 14977 11437 15011
rect 11437 14977 11471 15011
rect 11471 14977 11480 15011
rect 11428 14968 11480 14977
rect 11244 14943 11296 14952
rect 4160 14832 4212 14884
rect 6920 14832 6972 14884
rect 7196 14832 7248 14884
rect 8668 14832 8720 14884
rect 9680 14832 9732 14884
rect 11244 14909 11253 14943
rect 11253 14909 11287 14943
rect 11287 14909 11296 14943
rect 11244 14900 11296 14909
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 12440 15104 12492 15113
rect 15292 15104 15344 15156
rect 16856 15104 16908 15156
rect 18144 15104 18196 15156
rect 12992 14968 13044 15020
rect 12624 14943 12676 14952
rect 12624 14909 12633 14943
rect 12633 14909 12667 14943
rect 12667 14909 12676 14943
rect 12624 14900 12676 14909
rect 12348 14832 12400 14884
rect 14004 14900 14056 14952
rect 14832 14968 14884 15020
rect 16028 15011 16080 15020
rect 16028 14977 16037 15011
rect 16037 14977 16071 15011
rect 16071 14977 16080 15011
rect 16028 14968 16080 14977
rect 15016 14943 15068 14952
rect 15016 14909 15025 14943
rect 15025 14909 15059 14943
rect 15059 14909 15068 14943
rect 15016 14900 15068 14909
rect 15292 14900 15344 14952
rect 18420 14968 18472 15020
rect 19064 14968 19116 15020
rect 14924 14832 14976 14884
rect 16488 14875 16540 14884
rect 16488 14841 16522 14875
rect 16522 14841 16540 14875
rect 16488 14832 16540 14841
rect 17040 14900 17092 14952
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 19984 14900 20036 14952
rect 7932 14764 7984 14816
rect 9772 14807 9824 14816
rect 9772 14773 9781 14807
rect 9781 14773 9815 14807
rect 9815 14773 9824 14807
rect 9772 14764 9824 14773
rect 10416 14764 10468 14816
rect 10876 14764 10928 14816
rect 12072 14807 12124 14816
rect 12072 14773 12081 14807
rect 12081 14773 12115 14807
rect 12115 14773 12124 14807
rect 12072 14764 12124 14773
rect 13544 14764 13596 14816
rect 14556 14807 14608 14816
rect 14556 14773 14565 14807
rect 14565 14773 14599 14807
rect 14599 14773 14608 14807
rect 14556 14764 14608 14773
rect 14832 14807 14884 14816
rect 14832 14773 14841 14807
rect 14841 14773 14875 14807
rect 14875 14773 14884 14807
rect 14832 14764 14884 14773
rect 17316 14764 17368 14816
rect 17776 14764 17828 14816
rect 19340 14832 19392 14884
rect 18972 14764 19024 14816
rect 20352 14764 20404 14816
rect 7579 14662 7631 14714
rect 7643 14662 7695 14714
rect 7707 14662 7759 14714
rect 7771 14662 7823 14714
rect 14176 14662 14228 14714
rect 14240 14662 14292 14714
rect 14304 14662 14356 14714
rect 14368 14662 14420 14714
rect 3056 14492 3108 14544
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 3056 14356 3108 14408
rect 3332 14492 3384 14544
rect 4988 14492 5040 14544
rect 3332 14399 3384 14408
rect 3332 14365 3341 14399
rect 3341 14365 3375 14399
rect 3375 14365 3384 14399
rect 3332 14356 3384 14365
rect 3792 14424 3844 14476
rect 3976 14424 4028 14476
rect 5080 14424 5132 14476
rect 5264 14467 5316 14476
rect 5264 14433 5273 14467
rect 5273 14433 5307 14467
rect 5307 14433 5316 14467
rect 5264 14424 5316 14433
rect 6828 14492 6880 14544
rect 4160 14356 4212 14408
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 3608 14288 3660 14340
rect 6092 14467 6144 14476
rect 6092 14433 6126 14467
rect 6126 14433 6144 14467
rect 7104 14492 7156 14544
rect 9772 14560 9824 14612
rect 11704 14560 11756 14612
rect 12072 14560 12124 14612
rect 10600 14535 10652 14544
rect 10600 14501 10623 14535
rect 10623 14501 10652 14535
rect 10600 14492 10652 14501
rect 6092 14424 6144 14433
rect 7840 14424 7892 14476
rect 8300 14424 8352 14476
rect 8392 14424 8444 14476
rect 10876 14424 10928 14476
rect 11704 14424 11756 14476
rect 12072 14467 12124 14476
rect 12072 14433 12106 14467
rect 12106 14433 12124 14467
rect 12072 14424 12124 14433
rect 14556 14424 14608 14476
rect 16580 14492 16632 14544
rect 19524 14560 19576 14612
rect 19616 14560 19668 14612
rect 15568 14424 15620 14476
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 13544 14399 13596 14408
rect 3792 14220 3844 14272
rect 9312 14288 9364 14340
rect 13544 14365 13553 14399
rect 13553 14365 13587 14399
rect 13587 14365 13596 14399
rect 13544 14356 13596 14365
rect 8668 14263 8720 14272
rect 8668 14229 8677 14263
rect 8677 14229 8711 14263
rect 8711 14229 8720 14263
rect 8668 14220 8720 14229
rect 9220 14220 9272 14272
rect 9864 14263 9916 14272
rect 9864 14229 9873 14263
rect 9873 14229 9907 14263
rect 9907 14229 9916 14263
rect 9864 14220 9916 14229
rect 14648 14288 14700 14340
rect 15200 14288 15252 14340
rect 18144 14492 18196 14544
rect 17500 14467 17552 14476
rect 17500 14433 17534 14467
rect 17534 14433 17552 14467
rect 19432 14492 19484 14544
rect 20168 14535 20220 14544
rect 20168 14501 20177 14535
rect 20177 14501 20211 14535
rect 20211 14501 20220 14535
rect 20168 14492 20220 14501
rect 17500 14424 17552 14433
rect 20444 14424 20496 14476
rect 11796 14220 11848 14272
rect 16028 14220 16080 14272
rect 16488 14220 16540 14272
rect 17224 14220 17276 14272
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 4280 14118 4332 14170
rect 4344 14118 4396 14170
rect 4408 14118 4460 14170
rect 4472 14118 4524 14170
rect 10878 14118 10930 14170
rect 10942 14118 10994 14170
rect 11006 14118 11058 14170
rect 11070 14118 11122 14170
rect 17475 14118 17527 14170
rect 17539 14118 17591 14170
rect 17603 14118 17655 14170
rect 17667 14118 17719 14170
rect 3056 14059 3108 14068
rect 3056 14025 3065 14059
rect 3065 14025 3099 14059
rect 3099 14025 3108 14059
rect 3056 14016 3108 14025
rect 3516 14016 3568 14068
rect 4988 14059 5040 14068
rect 4988 14025 4997 14059
rect 4997 14025 5031 14059
rect 5031 14025 5040 14059
rect 4988 14016 5040 14025
rect 5264 14016 5316 14068
rect 7840 14016 7892 14068
rect 1400 13880 1452 13932
rect 2964 13880 3016 13932
rect 4988 13880 5040 13932
rect 4160 13812 4212 13864
rect 6092 13812 6144 13864
rect 7012 13880 7064 13932
rect 9864 14016 9916 14068
rect 11612 14016 11664 14068
rect 12624 14016 12676 14068
rect 13452 14016 13504 14068
rect 13912 14016 13964 14068
rect 14372 14016 14424 14068
rect 8668 13880 8720 13932
rect 9220 13923 9272 13932
rect 9220 13889 9232 13923
rect 9232 13889 9266 13923
rect 9266 13889 9272 13923
rect 9220 13880 9272 13889
rect 10140 13880 10192 13932
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 10324 13812 10376 13864
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 10968 13855 11020 13864
rect 10968 13821 11002 13855
rect 11002 13821 11020 13855
rect 10968 13812 11020 13821
rect 12348 13812 12400 13864
rect 14832 13880 14884 13932
rect 15292 13880 15344 13932
rect 16672 13880 16724 13932
rect 17040 13880 17092 13932
rect 17316 13880 17368 13932
rect 17500 13880 17552 13932
rect 18604 13880 18656 13932
rect 18880 13923 18932 13932
rect 18880 13889 18889 13923
rect 18889 13889 18923 13923
rect 18923 13889 18932 13923
rect 18880 13880 18932 13889
rect 13820 13812 13872 13864
rect 13912 13855 13964 13864
rect 13912 13821 13921 13855
rect 13921 13821 13955 13855
rect 13955 13821 13964 13855
rect 13912 13812 13964 13821
rect 3608 13744 3660 13796
rect 8668 13744 8720 13796
rect 17132 13812 17184 13864
rect 19064 13855 19116 13864
rect 19064 13821 19073 13855
rect 19073 13821 19107 13855
rect 19107 13821 19116 13855
rect 19064 13812 19116 13821
rect 20352 13812 20404 13864
rect 3332 13676 3384 13728
rect 4712 13676 4764 13728
rect 6276 13719 6328 13728
rect 6276 13685 6285 13719
rect 6285 13685 6319 13719
rect 6319 13685 6328 13719
rect 6276 13676 6328 13685
rect 8760 13676 8812 13728
rect 9588 13676 9640 13728
rect 16120 13744 16172 13796
rect 16304 13744 16356 13796
rect 11520 13676 11572 13728
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 12624 13676 12676 13728
rect 16948 13719 17000 13728
rect 16948 13685 16957 13719
rect 16957 13685 16991 13719
rect 16991 13685 17000 13719
rect 16948 13676 17000 13685
rect 17224 13744 17276 13796
rect 18420 13744 18472 13796
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 18512 13676 18564 13728
rect 20444 13719 20496 13728
rect 20444 13685 20453 13719
rect 20453 13685 20487 13719
rect 20487 13685 20496 13719
rect 20444 13676 20496 13685
rect 7579 13574 7631 13626
rect 7643 13574 7695 13626
rect 7707 13574 7759 13626
rect 7771 13574 7823 13626
rect 14176 13574 14228 13626
rect 14240 13574 14292 13626
rect 14304 13574 14356 13626
rect 14368 13574 14420 13626
rect 3148 13472 3200 13524
rect 3700 13515 3752 13524
rect 3700 13481 3709 13515
rect 3709 13481 3743 13515
rect 3743 13481 3752 13515
rect 3700 13472 3752 13481
rect 4620 13472 4672 13524
rect 6092 13472 6144 13524
rect 8392 13472 8444 13524
rect 8668 13472 8720 13524
rect 10048 13472 10100 13524
rect 2504 13404 2556 13456
rect 4804 13404 4856 13456
rect 5816 13404 5868 13456
rect 6276 13404 6328 13456
rect 7012 13404 7064 13456
rect 7932 13404 7984 13456
rect 2872 13336 2924 13388
rect 3976 13336 4028 13388
rect 4620 13379 4672 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 3332 13311 3384 13320
rect 3332 13277 3341 13311
rect 3341 13277 3375 13311
rect 3375 13277 3384 13311
rect 3332 13268 3384 13277
rect 3516 13311 3568 13320
rect 3516 13277 3525 13311
rect 3525 13277 3559 13311
rect 3559 13277 3568 13311
rect 3516 13268 3568 13277
rect 4252 13268 4304 13320
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 4896 13336 4948 13388
rect 6920 13379 6972 13388
rect 4988 13268 5040 13320
rect 5080 13311 5132 13320
rect 5080 13277 5089 13311
rect 5089 13277 5123 13311
rect 5123 13277 5132 13311
rect 6920 13345 6929 13379
rect 6929 13345 6963 13379
rect 6963 13345 6972 13379
rect 6920 13336 6972 13345
rect 10232 13404 10284 13456
rect 11520 13447 11572 13456
rect 11520 13413 11554 13447
rect 11554 13413 11572 13447
rect 11520 13404 11572 13413
rect 11704 13404 11756 13456
rect 12072 13472 12124 13524
rect 13820 13472 13872 13524
rect 16948 13472 17000 13524
rect 17132 13447 17184 13456
rect 5080 13268 5132 13277
rect 7288 13268 7340 13320
rect 7380 13268 7432 13320
rect 8760 13311 8812 13320
rect 8760 13277 8769 13311
rect 8769 13277 8803 13311
rect 8803 13277 8812 13311
rect 8760 13268 8812 13277
rect 9772 13336 9824 13388
rect 10692 13336 10744 13388
rect 13544 13336 13596 13388
rect 14648 13336 14700 13388
rect 9588 13268 9640 13320
rect 15016 13336 15068 13388
rect 16580 13336 16632 13388
rect 17132 13413 17141 13447
rect 17141 13413 17175 13447
rect 17175 13413 17184 13447
rect 17132 13404 17184 13413
rect 19156 13404 19208 13456
rect 16856 13336 16908 13388
rect 15568 13268 15620 13320
rect 16304 13311 16356 13320
rect 10968 13200 11020 13252
rect 14740 13200 14792 13252
rect 15936 13200 15988 13252
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 16488 13268 16540 13320
rect 16764 13200 16816 13252
rect 16948 13268 17000 13320
rect 17316 13268 17368 13320
rect 17500 13268 17552 13320
rect 18420 13336 18472 13388
rect 18604 13336 18656 13388
rect 19340 13336 19392 13388
rect 18328 13268 18380 13320
rect 18972 13311 19024 13320
rect 18972 13277 18981 13311
rect 18981 13277 19015 13311
rect 19015 13277 19024 13311
rect 19708 13311 19760 13320
rect 18972 13268 19024 13277
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 20536 13336 20588 13388
rect 18788 13200 18840 13252
rect 3424 13132 3476 13184
rect 6368 13132 6420 13184
rect 9956 13132 10008 13184
rect 10048 13132 10100 13184
rect 12532 13132 12584 13184
rect 12992 13132 13044 13184
rect 15660 13175 15712 13184
rect 15660 13141 15669 13175
rect 15669 13141 15703 13175
rect 15703 13141 15712 13175
rect 15660 13132 15712 13141
rect 16488 13175 16540 13184
rect 16488 13141 16497 13175
rect 16497 13141 16531 13175
rect 16531 13141 16540 13175
rect 18420 13175 18472 13184
rect 16488 13132 16540 13141
rect 18420 13141 18429 13175
rect 18429 13141 18463 13175
rect 18463 13141 18472 13175
rect 18420 13132 18472 13141
rect 20076 13132 20128 13184
rect 4280 13030 4332 13082
rect 4344 13030 4396 13082
rect 4408 13030 4460 13082
rect 4472 13030 4524 13082
rect 10878 13030 10930 13082
rect 10942 13030 10994 13082
rect 11006 13030 11058 13082
rect 11070 13030 11122 13082
rect 17475 13030 17527 13082
rect 17539 13030 17591 13082
rect 17603 13030 17655 13082
rect 17667 13030 17719 13082
rect 2872 12971 2924 12980
rect 2872 12937 2881 12971
rect 2881 12937 2915 12971
rect 2915 12937 2924 12971
rect 2872 12928 2924 12937
rect 4160 12928 4212 12980
rect 4068 12860 4120 12912
rect 5080 12928 5132 12980
rect 5816 12971 5868 12980
rect 5816 12937 5825 12971
rect 5825 12937 5859 12971
rect 5859 12937 5868 12971
rect 5816 12928 5868 12937
rect 5908 12971 5960 12980
rect 5908 12937 5917 12971
rect 5917 12937 5951 12971
rect 5951 12937 5960 12971
rect 5908 12928 5960 12937
rect 6276 12928 6328 12980
rect 6828 12928 6880 12980
rect 8116 12928 8168 12980
rect 10324 12928 10376 12980
rect 10600 12928 10652 12980
rect 11244 12928 11296 12980
rect 11888 12928 11940 12980
rect 5540 12860 5592 12912
rect 6368 12835 6420 12844
rect 1400 12724 1452 12776
rect 2964 12767 3016 12776
rect 2964 12733 2973 12767
rect 2973 12733 3007 12767
rect 3007 12733 3016 12767
rect 2964 12724 3016 12733
rect 3240 12767 3292 12776
rect 3240 12733 3274 12767
rect 3274 12733 3292 12767
rect 3240 12724 3292 12733
rect 4712 12767 4764 12776
rect 4712 12733 4746 12767
rect 4746 12733 4764 12767
rect 4712 12724 4764 12733
rect 2780 12656 2832 12708
rect 3332 12656 3384 12708
rect 4160 12656 4212 12708
rect 6368 12801 6377 12835
rect 6377 12801 6411 12835
rect 6411 12801 6420 12835
rect 6368 12792 6420 12801
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 8300 12835 8352 12844
rect 8300 12801 8309 12835
rect 8309 12801 8343 12835
rect 8343 12801 8352 12835
rect 10508 12835 10560 12844
rect 8300 12792 8352 12801
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 7472 12724 7524 12776
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 1860 12588 1912 12640
rect 9036 12656 9088 12708
rect 9956 12656 10008 12708
rect 11060 12699 11112 12708
rect 7288 12588 7340 12640
rect 8300 12588 8352 12640
rect 9588 12588 9640 12640
rect 9772 12588 9824 12640
rect 10324 12631 10376 12640
rect 10324 12597 10333 12631
rect 10333 12597 10367 12631
rect 10367 12597 10376 12631
rect 10324 12588 10376 12597
rect 11060 12665 11069 12699
rect 11069 12665 11103 12699
rect 11103 12665 11112 12699
rect 11060 12656 11112 12665
rect 11244 12699 11296 12708
rect 11244 12665 11253 12699
rect 11253 12665 11287 12699
rect 11287 12665 11296 12699
rect 11244 12656 11296 12665
rect 11336 12656 11388 12708
rect 11152 12588 11204 12640
rect 11428 12631 11480 12640
rect 11428 12597 11437 12631
rect 11437 12597 11471 12631
rect 11471 12597 11480 12631
rect 11428 12588 11480 12597
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 13544 12928 13596 12980
rect 16764 12971 16816 12980
rect 14924 12860 14976 12912
rect 16764 12937 16773 12971
rect 16773 12937 16807 12971
rect 16807 12937 16816 12971
rect 16764 12928 16816 12937
rect 17040 12928 17092 12980
rect 17132 12860 17184 12912
rect 12440 12724 12492 12776
rect 14004 12724 14056 12776
rect 15292 12767 15344 12776
rect 15292 12733 15301 12767
rect 15301 12733 15335 12767
rect 15335 12733 15344 12767
rect 15292 12724 15344 12733
rect 17040 12792 17092 12844
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 16304 12724 16356 12776
rect 16580 12724 16632 12776
rect 14740 12656 14792 12708
rect 15200 12656 15252 12708
rect 16948 12656 17000 12708
rect 13084 12588 13136 12640
rect 16304 12588 16356 12640
rect 16764 12588 16816 12640
rect 17224 12631 17276 12640
rect 17224 12597 17233 12631
rect 17233 12597 17267 12631
rect 17267 12597 17276 12631
rect 18512 12928 18564 12980
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 18880 12792 18932 12844
rect 19064 12835 19116 12844
rect 19064 12801 19073 12835
rect 19073 12801 19107 12835
rect 19107 12801 19116 12835
rect 19064 12792 19116 12801
rect 17776 12724 17828 12776
rect 18236 12724 18288 12776
rect 20444 12724 20496 12776
rect 19064 12656 19116 12708
rect 17224 12588 17276 12597
rect 17500 12588 17552 12640
rect 18144 12631 18196 12640
rect 18144 12597 18153 12631
rect 18153 12597 18187 12631
rect 18187 12597 18196 12631
rect 18144 12588 18196 12597
rect 18512 12588 18564 12640
rect 19156 12588 19208 12640
rect 7579 12486 7631 12538
rect 7643 12486 7695 12538
rect 7707 12486 7759 12538
rect 7771 12486 7823 12538
rect 14176 12486 14228 12538
rect 14240 12486 14292 12538
rect 14304 12486 14356 12538
rect 14368 12486 14420 12538
rect 2780 12427 2832 12436
rect 2780 12393 2789 12427
rect 2789 12393 2823 12427
rect 2823 12393 2832 12427
rect 2780 12384 2832 12393
rect 4160 12384 4212 12436
rect 6920 12384 6972 12436
rect 7104 12384 7156 12436
rect 7288 12316 7340 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 3148 12248 3200 12300
rect 5356 12248 5408 12300
rect 5908 12248 5960 12300
rect 6368 12248 6420 12300
rect 8300 12384 8352 12436
rect 9036 12384 9088 12436
rect 10324 12384 10376 12436
rect 13268 12384 13320 12436
rect 13728 12384 13780 12436
rect 18604 12427 18656 12436
rect 10140 12316 10192 12368
rect 3516 12180 3568 12232
rect 4068 12180 4120 12232
rect 5540 12180 5592 12232
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 6276 12180 6328 12189
rect 2964 12112 3016 12164
rect 3976 12044 4028 12096
rect 6644 12044 6696 12096
rect 6920 12044 6972 12096
rect 7380 12044 7432 12096
rect 8116 12248 8168 12300
rect 8576 12248 8628 12300
rect 10600 12291 10652 12300
rect 10600 12257 10609 12291
rect 10609 12257 10643 12291
rect 10643 12257 10652 12291
rect 10600 12248 10652 12257
rect 9128 12180 9180 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10968 12248 11020 12300
rect 12624 12248 12676 12300
rect 13176 12248 13228 12300
rect 14740 12248 14792 12300
rect 15200 12316 15252 12368
rect 10232 12180 10284 12189
rect 11704 12180 11756 12232
rect 12440 12180 12492 12232
rect 12716 12180 12768 12232
rect 14648 12180 14700 12232
rect 15384 12248 15436 12300
rect 16028 12248 16080 12300
rect 16672 12248 16724 12300
rect 17776 12316 17828 12368
rect 18604 12393 18613 12427
rect 18613 12393 18647 12427
rect 18647 12393 18656 12427
rect 18604 12384 18656 12393
rect 19708 12384 19760 12436
rect 19156 12359 19208 12368
rect 19156 12325 19190 12359
rect 19190 12325 19208 12359
rect 19156 12316 19208 12325
rect 19432 12316 19484 12368
rect 20352 12316 20404 12368
rect 17132 12291 17184 12300
rect 15292 12223 15344 12232
rect 15292 12189 15301 12223
rect 15301 12189 15335 12223
rect 15335 12189 15344 12223
rect 15292 12180 15344 12189
rect 16304 12180 16356 12232
rect 11336 12044 11388 12096
rect 12900 12044 12952 12096
rect 13176 12044 13228 12096
rect 15200 12044 15252 12096
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17316 12248 17368 12300
rect 17224 12223 17276 12232
rect 17224 12189 17233 12223
rect 17233 12189 17267 12223
rect 17267 12189 17276 12223
rect 17224 12180 17276 12189
rect 17592 12180 17644 12232
rect 17868 12180 17920 12232
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 20168 12180 20220 12232
rect 20352 12044 20404 12096
rect 4280 11942 4332 11994
rect 4344 11942 4396 11994
rect 4408 11942 4460 11994
rect 4472 11942 4524 11994
rect 10878 11942 10930 11994
rect 10942 11942 10994 11994
rect 11006 11942 11058 11994
rect 11070 11942 11122 11994
rect 17475 11942 17527 11994
rect 17539 11942 17591 11994
rect 17603 11942 17655 11994
rect 17667 11942 17719 11994
rect 4896 11840 4948 11892
rect 5356 11883 5408 11892
rect 5356 11849 5365 11883
rect 5365 11849 5399 11883
rect 5399 11849 5408 11883
rect 5356 11840 5408 11849
rect 10508 11883 10560 11892
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 6828 11772 6880 11824
rect 6276 11704 6328 11756
rect 3976 11679 4028 11688
rect 3976 11645 3985 11679
rect 3985 11645 4019 11679
rect 4019 11645 4028 11679
rect 3976 11636 4028 11645
rect 6736 11636 6788 11688
rect 8484 11704 8536 11756
rect 7932 11636 7984 11688
rect 10508 11849 10517 11883
rect 10517 11849 10551 11883
rect 10551 11849 10560 11883
rect 10508 11840 10560 11849
rect 10692 11840 10744 11892
rect 14096 11840 14148 11892
rect 16672 11840 16724 11892
rect 17868 11883 17920 11892
rect 16028 11772 16080 11824
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 19800 11840 19852 11892
rect 10692 11747 10744 11756
rect 2320 11543 2372 11552
rect 2320 11509 2329 11543
rect 2329 11509 2363 11543
rect 2363 11509 2372 11543
rect 2320 11500 2372 11509
rect 4620 11568 4672 11620
rect 5448 11568 5500 11620
rect 7104 11611 7156 11620
rect 7104 11577 7138 11611
rect 7138 11577 7156 11611
rect 7104 11568 7156 11577
rect 7196 11568 7248 11620
rect 9128 11568 9180 11620
rect 9404 11568 9456 11620
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 12256 11704 12308 11756
rect 14556 11747 14608 11756
rect 14556 11713 14565 11747
rect 14565 11713 14599 11747
rect 14599 11713 14608 11747
rect 14556 11704 14608 11713
rect 11244 11636 11296 11688
rect 11336 11636 11388 11688
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3148 11500 3200 11509
rect 4160 11500 4212 11552
rect 7288 11500 7340 11552
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 8300 11500 8352 11552
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 11428 11568 11480 11620
rect 12532 11568 12584 11620
rect 13820 11568 13872 11620
rect 14832 11636 14884 11688
rect 14648 11568 14700 11620
rect 15292 11568 15344 11620
rect 16304 11568 16356 11620
rect 9772 11500 9824 11509
rect 11980 11500 12032 11552
rect 12164 11500 12216 11552
rect 13728 11500 13780 11552
rect 13912 11543 13964 11552
rect 13912 11509 13921 11543
rect 13921 11509 13955 11543
rect 13955 11509 13964 11543
rect 13912 11500 13964 11509
rect 14464 11543 14516 11552
rect 14464 11509 14473 11543
rect 14473 11509 14507 11543
rect 14507 11509 14516 11543
rect 14464 11500 14516 11509
rect 17776 11704 17828 11756
rect 20076 11704 20128 11756
rect 20352 11747 20404 11756
rect 20352 11713 20361 11747
rect 20361 11713 20395 11747
rect 20395 11713 20404 11747
rect 20352 11704 20404 11713
rect 20168 11679 20220 11688
rect 17132 11568 17184 11620
rect 17408 11568 17460 11620
rect 20168 11645 20177 11679
rect 20177 11645 20211 11679
rect 20211 11645 20220 11679
rect 20168 11636 20220 11645
rect 18880 11568 18932 11620
rect 16672 11500 16724 11552
rect 18420 11500 18472 11552
rect 19892 11500 19944 11552
rect 7579 11398 7631 11450
rect 7643 11398 7695 11450
rect 7707 11398 7759 11450
rect 7771 11398 7823 11450
rect 14176 11398 14228 11450
rect 14240 11398 14292 11450
rect 14304 11398 14356 11450
rect 14368 11398 14420 11450
rect 2320 11296 2372 11348
rect 5448 11339 5500 11348
rect 3332 11228 3384 11280
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 7196 11296 7248 11348
rect 8300 11339 8352 11348
rect 5540 11228 5592 11280
rect 1492 11160 1544 11212
rect 3240 11203 3292 11212
rect 3240 11169 3249 11203
rect 3249 11169 3283 11203
rect 3283 11169 3292 11203
rect 3240 11160 3292 11169
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 3792 11160 3844 11212
rect 4620 11160 4672 11212
rect 7656 11228 7708 11280
rect 6644 11160 6696 11212
rect 8300 11305 8309 11339
rect 8309 11305 8343 11339
rect 8343 11305 8352 11339
rect 8300 11296 8352 11305
rect 8116 11228 8168 11280
rect 9680 11228 9732 11280
rect 11244 11296 11296 11348
rect 13636 11296 13688 11348
rect 13728 11296 13780 11348
rect 14464 11296 14516 11348
rect 14832 11296 14884 11348
rect 15200 11296 15252 11348
rect 8852 11160 8904 11212
rect 9588 11160 9640 11212
rect 11980 11228 12032 11280
rect 13912 11228 13964 11280
rect 11520 11160 11572 11212
rect 12440 11160 12492 11212
rect 13820 11160 13872 11212
rect 16120 11228 16172 11280
rect 16764 11296 16816 11348
rect 18328 11296 18380 11348
rect 14648 11160 14700 11212
rect 15568 11203 15620 11212
rect 15568 11169 15602 11203
rect 15602 11169 15620 11203
rect 15568 11160 15620 11169
rect 16580 11160 16632 11212
rect 17040 11203 17092 11212
rect 17040 11169 17049 11203
rect 17049 11169 17083 11203
rect 17083 11169 17092 11203
rect 20076 11296 20128 11348
rect 20352 11228 20404 11280
rect 17040 11160 17092 11169
rect 19248 11160 19300 11212
rect 2780 11067 2832 11076
rect 2780 11033 2789 11067
rect 2789 11033 2823 11067
rect 2823 11033 2832 11067
rect 2780 11024 2832 11033
rect 7288 11092 7340 11144
rect 8116 11092 8168 11144
rect 8300 11092 8352 11144
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12808 11135 12860 11144
rect 4068 10956 4120 11008
rect 7104 11024 7156 11076
rect 7196 10956 7248 11008
rect 8576 11024 8628 11076
rect 8668 11024 8720 11076
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 12808 11092 12860 11101
rect 15292 11135 15344 11144
rect 7932 10956 7984 11008
rect 9312 10956 9364 11008
rect 12256 11024 12308 11076
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 17408 11135 17460 11144
rect 17408 11101 17417 11135
rect 17417 11101 17451 11135
rect 17451 11101 17460 11135
rect 17408 11092 17460 11101
rect 18880 11135 18932 11144
rect 18880 11101 18889 11135
rect 18889 11101 18923 11135
rect 18923 11101 18932 11135
rect 18880 11092 18932 11101
rect 18972 11092 19024 11144
rect 14464 11067 14516 11076
rect 14464 11033 14473 11067
rect 14473 11033 14507 11067
rect 14507 11033 14516 11067
rect 14464 11024 14516 11033
rect 11428 10999 11480 11008
rect 11428 10965 11437 10999
rect 11437 10965 11471 10999
rect 11471 10965 11480 10999
rect 11428 10956 11480 10965
rect 11612 10956 11664 11008
rect 12348 10956 12400 11008
rect 14924 10999 14976 11008
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 16304 11024 16356 11076
rect 17316 10956 17368 11008
rect 18696 10956 18748 11008
rect 4280 10854 4332 10906
rect 4344 10854 4396 10906
rect 4408 10854 4460 10906
rect 4472 10854 4524 10906
rect 10878 10854 10930 10906
rect 10942 10854 10994 10906
rect 11006 10854 11058 10906
rect 11070 10854 11122 10906
rect 17475 10854 17527 10906
rect 17539 10854 17591 10906
rect 17603 10854 17655 10906
rect 17667 10854 17719 10906
rect 3240 10752 3292 10804
rect 4160 10752 4212 10804
rect 4620 10752 4672 10804
rect 7104 10752 7156 10804
rect 7656 10795 7708 10804
rect 7656 10761 7665 10795
rect 7665 10761 7699 10795
rect 7699 10761 7708 10795
rect 7656 10752 7708 10761
rect 8024 10752 8076 10804
rect 6552 10684 6604 10736
rect 9772 10752 9824 10804
rect 10324 10752 10376 10804
rect 11336 10752 11388 10804
rect 11796 10752 11848 10804
rect 13176 10752 13228 10804
rect 13820 10795 13872 10804
rect 13820 10761 13829 10795
rect 13829 10761 13863 10795
rect 13863 10761 13872 10795
rect 13820 10752 13872 10761
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 2780 10548 2832 10600
rect 3148 10591 3200 10600
rect 3148 10557 3182 10591
rect 3182 10557 3200 10591
rect 3148 10548 3200 10557
rect 4068 10548 4120 10600
rect 5540 10616 5592 10668
rect 6460 10659 6512 10668
rect 6460 10625 6469 10659
rect 6469 10625 6503 10659
rect 6503 10625 6512 10659
rect 6460 10616 6512 10625
rect 5724 10548 5776 10600
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 4160 10480 4212 10532
rect 7012 10480 7064 10532
rect 7380 10480 7432 10532
rect 8300 10659 8352 10668
rect 8300 10625 8309 10659
rect 8309 10625 8343 10659
rect 8343 10625 8352 10659
rect 8300 10616 8352 10625
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 6000 10412 6052 10464
rect 6644 10412 6696 10464
rect 8208 10548 8260 10600
rect 7748 10480 7800 10532
rect 8024 10455 8076 10464
rect 8024 10421 8033 10455
rect 8033 10421 8067 10455
rect 8067 10421 8076 10455
rect 8024 10412 8076 10421
rect 12164 10684 12216 10736
rect 12256 10616 12308 10668
rect 15292 10752 15344 10804
rect 16028 10752 16080 10804
rect 16764 10795 16816 10804
rect 16764 10761 16773 10795
rect 16773 10761 16807 10795
rect 16807 10761 16816 10795
rect 16764 10752 16816 10761
rect 17224 10752 17276 10804
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 17500 10684 17552 10736
rect 17960 10684 18012 10736
rect 19340 10684 19392 10736
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 8576 10548 8628 10600
rect 8760 10548 8812 10600
rect 8852 10480 8904 10532
rect 10232 10480 10284 10532
rect 12256 10412 12308 10464
rect 12532 10548 12584 10600
rect 15108 10548 15160 10600
rect 15384 10591 15436 10600
rect 15384 10557 15393 10591
rect 15393 10557 15427 10591
rect 15427 10557 15436 10591
rect 15384 10548 15436 10557
rect 15936 10548 15988 10600
rect 17776 10548 17828 10600
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 15292 10455 15344 10464
rect 15292 10421 15301 10455
rect 15301 10421 15335 10455
rect 15335 10421 15344 10455
rect 15292 10412 15344 10421
rect 15568 10412 15620 10464
rect 18696 10480 18748 10532
rect 19708 10480 19760 10532
rect 20812 10480 20864 10532
rect 15844 10412 15896 10464
rect 16672 10412 16724 10464
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 17224 10412 17276 10464
rect 18052 10412 18104 10464
rect 18512 10412 18564 10464
rect 19524 10455 19576 10464
rect 19524 10421 19533 10455
rect 19533 10421 19567 10455
rect 19567 10421 19576 10455
rect 19524 10412 19576 10421
rect 19892 10455 19944 10464
rect 19892 10421 19901 10455
rect 19901 10421 19935 10455
rect 19935 10421 19944 10455
rect 19892 10412 19944 10421
rect 19984 10455 20036 10464
rect 19984 10421 19993 10455
rect 19993 10421 20027 10455
rect 20027 10421 20036 10455
rect 19984 10412 20036 10421
rect 7579 10310 7631 10362
rect 7643 10310 7695 10362
rect 7707 10310 7759 10362
rect 7771 10310 7823 10362
rect 14176 10310 14228 10362
rect 14240 10310 14292 10362
rect 14304 10310 14356 10362
rect 14368 10310 14420 10362
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 6920 10208 6972 10260
rect 7472 10208 7524 10260
rect 8024 10208 8076 10260
rect 8300 10208 8352 10260
rect 3240 10140 3292 10192
rect 5724 10140 5776 10192
rect 5816 10140 5868 10192
rect 4160 10072 4212 10124
rect 5908 10115 5960 10124
rect 5908 10081 5917 10115
rect 5917 10081 5951 10115
rect 5951 10081 5960 10115
rect 5908 10072 5960 10081
rect 7380 10115 7432 10124
rect 7380 10081 7389 10115
rect 7389 10081 7423 10115
rect 7423 10081 7432 10115
rect 7380 10072 7432 10081
rect 8116 10072 8168 10124
rect 8300 10115 8352 10124
rect 8300 10081 8309 10115
rect 8309 10081 8343 10115
rect 8343 10081 8352 10115
rect 9128 10115 9180 10124
rect 8300 10072 8352 10081
rect 9128 10081 9137 10115
rect 9137 10081 9171 10115
rect 9171 10081 9180 10115
rect 9128 10072 9180 10081
rect 9588 10140 9640 10192
rect 3792 10004 3844 10056
rect 5172 10004 5224 10056
rect 6276 10004 6328 10056
rect 7472 10047 7524 10056
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 8668 10004 8720 10056
rect 5172 9868 5224 9920
rect 6828 9936 6880 9988
rect 7932 9936 7984 9988
rect 7840 9868 7892 9920
rect 8392 9868 8444 9920
rect 9956 10072 10008 10124
rect 10324 10140 10376 10192
rect 11428 10208 11480 10260
rect 12164 10208 12216 10260
rect 17040 10208 17092 10260
rect 17132 10208 17184 10260
rect 17500 10208 17552 10260
rect 11796 10072 11848 10124
rect 9312 9936 9364 9988
rect 9496 10004 9548 10056
rect 12992 10140 13044 10192
rect 13360 10140 13412 10192
rect 15292 10140 15344 10192
rect 15660 10140 15712 10192
rect 12348 10072 12400 10124
rect 12716 10072 12768 10124
rect 14004 10072 14056 10124
rect 15476 10072 15528 10124
rect 16764 10072 16816 10124
rect 17776 10140 17828 10192
rect 19524 10208 19576 10260
rect 12808 10004 12860 10056
rect 13636 10004 13688 10056
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 15384 10004 15436 10056
rect 11520 9979 11572 9988
rect 11520 9945 11529 9979
rect 11529 9945 11563 9979
rect 11563 9945 11572 9979
rect 11520 9936 11572 9945
rect 12532 9936 12584 9988
rect 13176 9936 13228 9988
rect 11428 9868 11480 9920
rect 12992 9868 13044 9920
rect 13544 9868 13596 9920
rect 15108 9868 15160 9920
rect 15936 9868 15988 9920
rect 17040 10004 17092 10056
rect 17960 10072 18012 10124
rect 18880 10072 18932 10124
rect 20260 10072 20312 10124
rect 18052 10004 18104 10056
rect 18420 10004 18472 10056
rect 18604 10047 18656 10056
rect 18604 10013 18613 10047
rect 18613 10013 18647 10047
rect 18647 10013 18656 10047
rect 18604 10004 18656 10013
rect 18696 10004 18748 10056
rect 17224 9868 17276 9920
rect 17776 9868 17828 9920
rect 18604 9868 18656 9920
rect 19984 9936 20036 9988
rect 19708 9911 19760 9920
rect 19708 9877 19717 9911
rect 19717 9877 19751 9911
rect 19751 9877 19760 9911
rect 19708 9868 19760 9877
rect 20260 9868 20312 9920
rect 4280 9766 4332 9818
rect 4344 9766 4396 9818
rect 4408 9766 4460 9818
rect 4472 9766 4524 9818
rect 10878 9766 10930 9818
rect 10942 9766 10994 9818
rect 11006 9766 11058 9818
rect 11070 9766 11122 9818
rect 17475 9766 17527 9818
rect 17539 9766 17591 9818
rect 17603 9766 17655 9818
rect 17667 9766 17719 9818
rect 6000 9664 6052 9716
rect 7012 9664 7064 9716
rect 8760 9664 8812 9716
rect 8852 9664 8904 9716
rect 11428 9664 11480 9716
rect 12348 9664 12400 9716
rect 15108 9707 15160 9716
rect 1860 9596 1912 9648
rect 2964 9639 3016 9648
rect 2964 9605 2973 9639
rect 2973 9605 3007 9639
rect 3007 9605 3016 9639
rect 2964 9596 3016 9605
rect 6920 9596 6972 9648
rect 7472 9596 7524 9648
rect 9220 9639 9272 9648
rect 9220 9605 9229 9639
rect 9229 9605 9263 9639
rect 9263 9605 9272 9639
rect 9220 9596 9272 9605
rect 11888 9596 11940 9648
rect 12164 9596 12216 9648
rect 15108 9673 15117 9707
rect 15117 9673 15151 9707
rect 15151 9673 15160 9707
rect 15108 9664 15160 9673
rect 17868 9664 17920 9716
rect 2228 9435 2280 9444
rect 2228 9401 2237 9435
rect 2237 9401 2271 9435
rect 2271 9401 2280 9435
rect 2228 9392 2280 9401
rect 3332 9460 3384 9512
rect 3792 9503 3844 9512
rect 3792 9469 3801 9503
rect 3801 9469 3835 9503
rect 3835 9469 3844 9503
rect 3792 9460 3844 9469
rect 4988 9528 5040 9580
rect 6276 9528 6328 9580
rect 7656 9528 7708 9580
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 5172 9460 5224 9512
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 6276 9392 6328 9444
rect 3424 9324 3476 9333
rect 5080 9324 5132 9376
rect 5908 9324 5960 9376
rect 6000 9324 6052 9376
rect 8116 9435 8168 9444
rect 8116 9401 8150 9435
rect 8150 9401 8168 9435
rect 8116 9392 8168 9401
rect 8484 9392 8536 9444
rect 10692 9460 10744 9512
rect 11336 9460 11388 9512
rect 17684 9596 17736 9648
rect 18420 9639 18472 9648
rect 18420 9605 18429 9639
rect 18429 9605 18463 9639
rect 18463 9605 18472 9639
rect 18420 9596 18472 9605
rect 12164 9460 12216 9512
rect 9404 9392 9456 9444
rect 9680 9392 9732 9444
rect 12624 9460 12676 9512
rect 12808 9460 12860 9512
rect 13360 9528 13412 9580
rect 15108 9528 15160 9580
rect 15384 9571 15436 9580
rect 15384 9537 15393 9571
rect 15393 9537 15427 9571
rect 15427 9537 15436 9571
rect 15384 9528 15436 9537
rect 16488 9528 16540 9580
rect 17224 9528 17276 9580
rect 17776 9528 17828 9580
rect 18512 9528 18564 9580
rect 13176 9460 13228 9512
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 13544 9460 13596 9512
rect 14464 9460 14516 9512
rect 15660 9503 15712 9512
rect 15660 9469 15694 9503
rect 15694 9469 15712 9503
rect 15660 9460 15712 9469
rect 14556 9392 14608 9444
rect 16856 9460 16908 9512
rect 16948 9460 17000 9512
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 19248 9460 19300 9512
rect 10784 9324 10836 9376
rect 10876 9324 10928 9376
rect 11796 9324 11848 9376
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 12256 9324 12308 9376
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 15200 9324 15252 9376
rect 16672 9392 16724 9444
rect 18144 9392 18196 9444
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 17224 9367 17276 9376
rect 16856 9324 16908 9333
rect 17224 9333 17233 9367
rect 17233 9333 17267 9367
rect 17267 9333 17276 9367
rect 17224 9324 17276 9333
rect 17408 9324 17460 9376
rect 18604 9392 18656 9444
rect 18788 9392 18840 9444
rect 19156 9392 19208 9444
rect 18696 9324 18748 9376
rect 19432 9324 19484 9376
rect 7579 9222 7631 9274
rect 7643 9222 7695 9274
rect 7707 9222 7759 9274
rect 7771 9222 7823 9274
rect 14176 9222 14228 9274
rect 14240 9222 14292 9274
rect 14304 9222 14356 9274
rect 14368 9222 14420 9274
rect 2688 9163 2740 9172
rect 2688 9129 2697 9163
rect 2697 9129 2731 9163
rect 2731 9129 2740 9163
rect 2688 9120 2740 9129
rect 3792 9120 3844 9172
rect 3976 9052 4028 9104
rect 4252 9120 4304 9172
rect 5356 9120 5408 9172
rect 6000 9120 6052 9172
rect 7380 9120 7432 9172
rect 2964 8984 3016 9036
rect 2688 8848 2740 8900
rect 4160 8984 4212 9036
rect 5908 9052 5960 9104
rect 6920 9052 6972 9104
rect 7012 9052 7064 9104
rect 8024 9120 8076 9172
rect 8116 9120 8168 9172
rect 8208 9052 8260 9104
rect 4988 8984 5040 9036
rect 7840 8984 7892 9036
rect 9864 9120 9916 9172
rect 12440 9163 12492 9172
rect 4252 8848 4304 8900
rect 2872 8780 2924 8832
rect 3976 8780 4028 8832
rect 6920 8916 6972 8968
rect 10048 9052 10100 9104
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 12440 9120 12492 9129
rect 10508 8984 10560 9036
rect 11336 9027 11388 9036
rect 11336 8993 11370 9027
rect 11370 8993 11388 9027
rect 11336 8984 11388 8993
rect 12624 9052 12676 9104
rect 13176 9120 13228 9172
rect 13084 8984 13136 9036
rect 9312 8916 9364 8925
rect 10416 8916 10468 8968
rect 10692 8916 10744 8968
rect 10876 8959 10928 8968
rect 10876 8925 10885 8959
rect 10885 8925 10919 8959
rect 10919 8925 10928 8959
rect 10876 8916 10928 8925
rect 12256 8916 12308 8968
rect 14740 9027 14792 9036
rect 14740 8993 14749 9027
rect 14749 8993 14783 9027
rect 14783 8993 14792 9027
rect 14740 8984 14792 8993
rect 15384 8984 15436 9036
rect 16764 9052 16816 9104
rect 16856 9052 16908 9104
rect 17132 9027 17184 9036
rect 15016 8959 15068 8968
rect 4620 8780 4672 8832
rect 4712 8780 4764 8832
rect 10048 8848 10100 8900
rect 15016 8925 15025 8959
rect 15025 8925 15059 8959
rect 15059 8925 15068 8959
rect 15016 8916 15068 8925
rect 15108 8916 15160 8968
rect 9772 8780 9824 8832
rect 9956 8780 10008 8832
rect 12348 8780 12400 8832
rect 12532 8780 12584 8832
rect 14372 8823 14424 8832
rect 14372 8789 14381 8823
rect 14381 8789 14415 8823
rect 14415 8789 14424 8823
rect 14372 8780 14424 8789
rect 15200 8848 15252 8900
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 20536 9052 20588 9104
rect 19432 9027 19484 9036
rect 19432 8993 19466 9027
rect 19466 8993 19484 9027
rect 19432 8984 19484 8993
rect 16856 8916 16908 8968
rect 17316 8959 17368 8968
rect 17316 8925 17325 8959
rect 17325 8925 17359 8959
rect 17359 8925 17368 8959
rect 18144 8959 18196 8968
rect 17316 8916 17368 8925
rect 18144 8925 18153 8959
rect 18153 8925 18187 8959
rect 18187 8925 18196 8959
rect 18144 8916 18196 8925
rect 18512 8916 18564 8968
rect 17408 8848 17460 8900
rect 17500 8848 17552 8900
rect 18420 8848 18472 8900
rect 15936 8780 15988 8832
rect 16028 8780 16080 8832
rect 17316 8780 17368 8832
rect 18144 8780 18196 8832
rect 19524 8780 19576 8832
rect 4280 8678 4332 8730
rect 4344 8678 4396 8730
rect 4408 8678 4460 8730
rect 4472 8678 4524 8730
rect 10878 8678 10930 8730
rect 10942 8678 10994 8730
rect 11006 8678 11058 8730
rect 11070 8678 11122 8730
rect 17475 8678 17527 8730
rect 17539 8678 17591 8730
rect 17603 8678 17655 8730
rect 17667 8678 17719 8730
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 3884 8576 3936 8628
rect 4620 8576 4672 8628
rect 6276 8619 6328 8628
rect 4896 8508 4948 8560
rect 6276 8585 6285 8619
rect 6285 8585 6319 8619
rect 6319 8585 6328 8619
rect 6276 8576 6328 8585
rect 7840 8576 7892 8628
rect 8208 8576 8260 8628
rect 6460 8551 6512 8560
rect 6460 8517 6469 8551
rect 6469 8517 6503 8551
rect 6503 8517 6512 8551
rect 6460 8508 6512 8517
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3056 8483 3108 8492
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 3976 8440 4028 8492
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 4068 8372 4120 8424
rect 4804 8372 4856 8424
rect 4988 8372 5040 8424
rect 6000 8372 6052 8424
rect 6368 8372 6420 8424
rect 10508 8576 10560 8628
rect 12624 8576 12676 8628
rect 12808 8576 12860 8628
rect 13820 8576 13872 8628
rect 14464 8576 14516 8628
rect 14740 8576 14792 8628
rect 11428 8508 11480 8560
rect 11980 8508 12032 8560
rect 8484 8483 8536 8492
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 9496 8440 9548 8492
rect 7380 8304 7432 8356
rect 7472 8304 7524 8356
rect 9956 8372 10008 8424
rect 11980 8415 12032 8424
rect 10140 8304 10192 8356
rect 10416 8347 10468 8356
rect 10416 8313 10450 8347
rect 10450 8313 10468 8347
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 12900 8508 12952 8560
rect 13636 8508 13688 8560
rect 13360 8440 13412 8492
rect 13912 8508 13964 8560
rect 14188 8508 14240 8560
rect 16856 8576 16908 8628
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 19984 8576 20036 8628
rect 10416 8304 10468 8313
rect 12440 8304 12492 8356
rect 12808 8347 12860 8356
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 14556 8372 14608 8424
rect 16488 8508 16540 8560
rect 17040 8508 17092 8560
rect 15200 8440 15252 8492
rect 15476 8483 15528 8492
rect 15476 8449 15485 8483
rect 15485 8449 15519 8483
rect 15519 8449 15528 8483
rect 15476 8440 15528 8449
rect 16028 8372 16080 8424
rect 16212 8372 16264 8424
rect 18236 8440 18288 8492
rect 16672 8372 16724 8424
rect 18328 8372 18380 8424
rect 18788 8415 18840 8424
rect 18788 8381 18797 8415
rect 18797 8381 18831 8415
rect 18831 8381 18840 8415
rect 18788 8372 18840 8381
rect 17132 8304 17184 8356
rect 18052 8304 18104 8356
rect 20076 8304 20128 8356
rect 4988 8236 5040 8288
rect 9680 8236 9732 8288
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 12348 8236 12400 8288
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 13636 8279 13688 8288
rect 13636 8245 13645 8279
rect 13645 8245 13679 8279
rect 13679 8245 13688 8279
rect 13636 8236 13688 8245
rect 13728 8279 13780 8288
rect 13728 8245 13737 8279
rect 13737 8245 13771 8279
rect 13771 8245 13780 8279
rect 13728 8236 13780 8245
rect 14464 8236 14516 8288
rect 15844 8236 15896 8288
rect 16856 8279 16908 8288
rect 16856 8245 16865 8279
rect 16865 8245 16899 8279
rect 16899 8245 16908 8279
rect 16856 8236 16908 8245
rect 17224 8236 17276 8288
rect 7579 8134 7631 8186
rect 7643 8134 7695 8186
rect 7707 8134 7759 8186
rect 7771 8134 7823 8186
rect 14176 8134 14228 8186
rect 14240 8134 14292 8186
rect 14304 8134 14356 8186
rect 14368 8134 14420 8186
rect 4896 8032 4948 8084
rect 5632 7964 5684 8016
rect 5908 7964 5960 8016
rect 10416 8032 10468 8084
rect 11980 8032 12032 8084
rect 13360 8032 13412 8084
rect 13636 8075 13688 8084
rect 13636 8041 13645 8075
rect 13645 8041 13679 8075
rect 13679 8041 13688 8075
rect 13636 8032 13688 8041
rect 8852 7964 8904 8016
rect 9772 7964 9824 8016
rect 13728 7964 13780 8016
rect 15292 8032 15344 8084
rect 15752 8075 15804 8084
rect 15752 8041 15761 8075
rect 15761 8041 15795 8075
rect 15795 8041 15804 8075
rect 15752 8032 15804 8041
rect 17040 8032 17092 8084
rect 17132 8032 17184 8084
rect 15568 7964 15620 8016
rect 16212 7964 16264 8016
rect 18512 7964 18564 8016
rect 3608 7939 3660 7948
rect 3608 7905 3617 7939
rect 3617 7905 3651 7939
rect 3651 7905 3660 7939
rect 4988 7939 5040 7948
rect 3608 7896 3660 7905
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 5724 7896 5776 7948
rect 6644 7939 6696 7948
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 6000 7828 6052 7880
rect 5080 7760 5132 7812
rect 4068 7692 4120 7744
rect 5356 7692 5408 7744
rect 6000 7692 6052 7744
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 8024 7896 8076 7948
rect 8208 7896 8260 7948
rect 9864 7896 9916 7948
rect 10048 7939 10100 7948
rect 10048 7905 10082 7939
rect 10082 7905 10100 7939
rect 10048 7896 10100 7905
rect 13544 7896 13596 7948
rect 7472 7828 7524 7880
rect 7840 7760 7892 7812
rect 6736 7692 6788 7744
rect 7196 7692 7248 7744
rect 9496 7828 9548 7880
rect 11244 7828 11296 7880
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 14464 7896 14516 7948
rect 16028 7896 16080 7948
rect 16396 7939 16448 7948
rect 16396 7905 16405 7939
rect 16405 7905 16439 7939
rect 16439 7905 16448 7939
rect 16396 7896 16448 7905
rect 17040 7896 17092 7948
rect 17224 7896 17276 7948
rect 17776 7896 17828 7948
rect 19432 7939 19484 7948
rect 19432 7905 19466 7939
rect 19466 7905 19484 7939
rect 19432 7896 19484 7905
rect 18788 7871 18840 7880
rect 8392 7692 8444 7744
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 14924 7692 14976 7744
rect 15752 7692 15804 7744
rect 18052 7692 18104 7744
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 19892 7692 19944 7744
rect 4280 7590 4332 7642
rect 4344 7590 4396 7642
rect 4408 7590 4460 7642
rect 4472 7590 4524 7642
rect 10878 7590 10930 7642
rect 10942 7590 10994 7642
rect 11006 7590 11058 7642
rect 11070 7590 11122 7642
rect 17475 7590 17527 7642
rect 17539 7590 17591 7642
rect 17603 7590 17655 7642
rect 17667 7590 17719 7642
rect 6644 7488 6696 7540
rect 3608 7463 3660 7472
rect 3608 7429 3617 7463
rect 3617 7429 3651 7463
rect 3651 7429 3660 7463
rect 3608 7420 3660 7429
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 5080 7395 5132 7404
rect 5080 7361 5089 7395
rect 5089 7361 5123 7395
rect 5123 7361 5132 7395
rect 5080 7352 5132 7361
rect 5172 7352 5224 7404
rect 8300 7488 8352 7540
rect 11244 7488 11296 7540
rect 12808 7488 12860 7540
rect 13728 7488 13780 7540
rect 14924 7488 14976 7540
rect 17776 7531 17828 7540
rect 7840 7420 7892 7472
rect 9036 7420 9088 7472
rect 15476 7420 15528 7472
rect 17776 7497 17785 7531
rect 17785 7497 17819 7531
rect 17819 7497 17828 7531
rect 17776 7488 17828 7497
rect 18052 7420 18104 7472
rect 19064 7420 19116 7472
rect 9312 7352 9364 7404
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 13820 7352 13872 7404
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 16120 7395 16172 7404
rect 3976 7259 4028 7268
rect 3976 7225 3985 7259
rect 3985 7225 4019 7259
rect 4019 7225 4028 7259
rect 3976 7216 4028 7225
rect 6460 7284 6512 7336
rect 9496 7284 9548 7336
rect 10416 7284 10468 7336
rect 10692 7284 10744 7336
rect 12256 7284 12308 7336
rect 6276 7216 6328 7268
rect 5172 7148 5224 7200
rect 5356 7148 5408 7200
rect 11428 7216 11480 7268
rect 12808 7216 12860 7268
rect 12900 7216 12952 7268
rect 13820 7216 13872 7268
rect 15660 7284 15712 7336
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 16856 7284 16908 7336
rect 17868 7284 17920 7336
rect 18880 7284 18932 7336
rect 16948 7216 17000 7268
rect 17040 7216 17092 7268
rect 19892 7352 19944 7404
rect 8208 7191 8260 7200
rect 8208 7157 8217 7191
rect 8217 7157 8251 7191
rect 8251 7157 8260 7191
rect 8208 7148 8260 7157
rect 8760 7148 8812 7200
rect 9864 7148 9916 7200
rect 10048 7148 10100 7200
rect 14004 7148 14056 7200
rect 17224 7148 17276 7200
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 17868 7148 17920 7200
rect 18604 7148 18656 7200
rect 7579 7046 7631 7098
rect 7643 7046 7695 7098
rect 7707 7046 7759 7098
rect 7771 7046 7823 7098
rect 14176 7046 14228 7098
rect 14240 7046 14292 7098
rect 14304 7046 14356 7098
rect 14368 7046 14420 7098
rect 4252 6944 4304 6996
rect 6276 6987 6328 6996
rect 6276 6953 6285 6987
rect 6285 6953 6319 6987
rect 6319 6953 6328 6987
rect 6276 6944 6328 6953
rect 8300 6944 8352 6996
rect 11428 6987 11480 6996
rect 5724 6808 5776 6860
rect 6460 6808 6512 6860
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 8208 6876 8260 6928
rect 8576 6876 8628 6928
rect 8760 6876 8812 6928
rect 9036 6876 9088 6928
rect 11428 6953 11437 6987
rect 11437 6953 11471 6987
rect 11471 6953 11480 6987
rect 11428 6944 11480 6953
rect 10048 6876 10100 6928
rect 11244 6876 11296 6928
rect 13728 6944 13780 6996
rect 14464 6944 14516 6996
rect 15752 6987 15804 6996
rect 15752 6953 15761 6987
rect 15761 6953 15795 6987
rect 15795 6953 15804 6987
rect 15752 6944 15804 6953
rect 17224 6944 17276 6996
rect 18880 6944 18932 6996
rect 9864 6808 9916 6860
rect 4620 6740 4672 6792
rect 7104 6783 7156 6792
rect 7104 6749 7113 6783
rect 7113 6749 7147 6783
rect 7147 6749 7156 6783
rect 7104 6740 7156 6749
rect 8300 6740 8352 6792
rect 10140 6808 10192 6860
rect 10324 6851 10376 6860
rect 10324 6817 10358 6851
rect 10358 6817 10376 6851
rect 10324 6808 10376 6817
rect 10600 6808 10652 6860
rect 4160 6604 4212 6656
rect 9496 6604 9548 6656
rect 13268 6672 13320 6724
rect 11704 6604 11756 6656
rect 12624 6604 12676 6656
rect 13544 6851 13596 6860
rect 13544 6817 13553 6851
rect 13553 6817 13587 6851
rect 13587 6817 13596 6851
rect 13544 6808 13596 6817
rect 15660 6851 15712 6860
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 16120 6876 16172 6928
rect 17040 6876 17092 6928
rect 17316 6919 17368 6928
rect 17316 6885 17350 6919
rect 17350 6885 17368 6919
rect 17316 6876 17368 6885
rect 17500 6876 17552 6928
rect 19800 6876 19852 6928
rect 20996 6919 21048 6928
rect 20996 6885 21005 6919
rect 21005 6885 21039 6919
rect 21039 6885 21048 6919
rect 20996 6876 21048 6885
rect 18604 6808 18656 6860
rect 16856 6783 16908 6792
rect 13544 6672 13596 6724
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 18512 6740 18564 6792
rect 18788 6851 18840 6860
rect 18788 6817 18797 6851
rect 18797 6817 18831 6851
rect 18831 6817 18840 6851
rect 19984 6851 20036 6860
rect 18788 6808 18840 6817
rect 19984 6817 19993 6851
rect 19993 6817 20027 6851
rect 20027 6817 20036 6851
rect 19984 6808 20036 6817
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 16672 6672 16724 6724
rect 18052 6672 18104 6724
rect 13912 6604 13964 6656
rect 15660 6604 15712 6656
rect 16120 6604 16172 6656
rect 17040 6604 17092 6656
rect 17960 6604 18012 6656
rect 18604 6604 18656 6656
rect 18972 6647 19024 6656
rect 18972 6613 18981 6647
rect 18981 6613 19015 6647
rect 19015 6613 19024 6647
rect 18972 6604 19024 6613
rect 19432 6604 19484 6656
rect 4280 6502 4332 6554
rect 4344 6502 4396 6554
rect 4408 6502 4460 6554
rect 4472 6502 4524 6554
rect 10878 6502 10930 6554
rect 10942 6502 10994 6554
rect 11006 6502 11058 6554
rect 11070 6502 11122 6554
rect 17475 6502 17527 6554
rect 17539 6502 17591 6554
rect 17603 6502 17655 6554
rect 17667 6502 17719 6554
rect 5724 6400 5776 6452
rect 8300 6400 8352 6452
rect 9496 6400 9548 6452
rect 12532 6400 12584 6452
rect 13084 6400 13136 6452
rect 14648 6400 14700 6452
rect 18512 6400 18564 6452
rect 20536 6443 20588 6452
rect 20536 6409 20545 6443
rect 20545 6409 20579 6443
rect 20579 6409 20588 6443
rect 20536 6400 20588 6409
rect 6920 6332 6972 6384
rect 7656 6332 7708 6384
rect 11704 6332 11756 6384
rect 12900 6332 12952 6384
rect 13636 6332 13688 6384
rect 7472 6307 7524 6316
rect 4620 6196 4672 6248
rect 4252 6128 4304 6180
rect 5080 6196 5132 6248
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 6828 6196 6880 6248
rect 9128 6239 9180 6248
rect 5908 6128 5960 6180
rect 7104 6128 7156 6180
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 10140 6196 10192 6248
rect 10600 6239 10652 6248
rect 10600 6205 10609 6239
rect 10609 6205 10643 6239
rect 10643 6205 10652 6239
rect 10600 6196 10652 6205
rect 13544 6264 13596 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 16488 6264 16540 6316
rect 17316 6264 17368 6316
rect 17776 6264 17828 6316
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 7196 6103 7248 6112
rect 7196 6069 7205 6103
rect 7205 6069 7239 6103
rect 7239 6069 7248 6103
rect 7196 6060 7248 6069
rect 7380 6060 7432 6112
rect 8668 6128 8720 6180
rect 11796 6196 11848 6248
rect 12992 6196 13044 6248
rect 13360 6196 13412 6248
rect 13636 6239 13688 6248
rect 13636 6205 13645 6239
rect 13645 6205 13679 6239
rect 13679 6205 13688 6239
rect 13636 6196 13688 6205
rect 10876 6171 10928 6180
rect 10876 6137 10910 6171
rect 10910 6137 10928 6171
rect 10876 6128 10928 6137
rect 11612 6128 11664 6180
rect 18604 6239 18656 6248
rect 14556 6128 14608 6180
rect 8116 6060 8168 6112
rect 8392 6060 8444 6112
rect 9220 6060 9272 6112
rect 10140 6060 10192 6112
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 12992 6060 13044 6112
rect 13176 6103 13228 6112
rect 13176 6069 13185 6103
rect 13185 6069 13219 6103
rect 13219 6069 13228 6103
rect 13176 6060 13228 6069
rect 15016 6103 15068 6112
rect 15016 6069 15025 6103
rect 15025 6069 15059 6103
rect 15059 6069 15068 6103
rect 15016 6060 15068 6069
rect 15200 6103 15252 6112
rect 15200 6069 15209 6103
rect 15209 6069 15243 6103
rect 15243 6069 15252 6103
rect 15200 6060 15252 6069
rect 15476 6060 15528 6112
rect 15936 6060 15988 6112
rect 16120 6128 16172 6180
rect 18604 6205 18613 6239
rect 18613 6205 18647 6239
rect 18647 6205 18656 6239
rect 18604 6196 18656 6205
rect 19984 6196 20036 6248
rect 20168 6239 20220 6248
rect 20168 6205 20177 6239
rect 20177 6205 20211 6239
rect 20211 6205 20220 6239
rect 20168 6196 20220 6205
rect 19524 6128 19576 6180
rect 16304 6060 16356 6112
rect 16856 6103 16908 6112
rect 16856 6069 16865 6103
rect 16865 6069 16899 6103
rect 16899 6069 16908 6103
rect 16856 6060 16908 6069
rect 17040 6060 17092 6112
rect 18236 6103 18288 6112
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 19892 6060 19944 6112
rect 7579 5958 7631 6010
rect 7643 5958 7695 6010
rect 7707 5958 7759 6010
rect 7771 5958 7823 6010
rect 14176 5958 14228 6010
rect 14240 5958 14292 6010
rect 14304 5958 14356 6010
rect 14368 5958 14420 6010
rect 3608 5899 3660 5908
rect 3608 5865 3617 5899
rect 3617 5865 3651 5899
rect 3651 5865 3660 5899
rect 3608 5856 3660 5865
rect 4620 5856 4672 5908
rect 5908 5899 5960 5908
rect 5908 5865 5917 5899
rect 5917 5865 5951 5899
rect 5951 5865 5960 5899
rect 5908 5856 5960 5865
rect 6184 5856 6236 5908
rect 7472 5856 7524 5908
rect 10876 5856 10928 5908
rect 10968 5856 11020 5908
rect 13084 5856 13136 5908
rect 13268 5856 13320 5908
rect 16488 5856 16540 5908
rect 16764 5856 16816 5908
rect 19524 5899 19576 5908
rect 4160 5720 4212 5772
rect 4620 5720 4672 5772
rect 5816 5720 5868 5772
rect 4252 5652 4304 5704
rect 7288 5788 7340 5840
rect 6368 5720 6420 5772
rect 7564 5763 7616 5772
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 6552 5652 6604 5704
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 10048 5788 10100 5840
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 8392 5763 8444 5772
rect 8392 5729 8426 5763
rect 8426 5729 8444 5763
rect 8392 5720 8444 5729
rect 10784 5720 10836 5772
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 12808 5720 12860 5772
rect 13268 5763 13320 5772
rect 13268 5729 13302 5763
rect 13302 5729 13320 5763
rect 13268 5720 13320 5729
rect 13544 5720 13596 5772
rect 14648 5763 14700 5772
rect 6920 5652 6972 5661
rect 8116 5584 8168 5636
rect 6276 5516 6328 5568
rect 6368 5559 6420 5568
rect 6368 5525 6377 5559
rect 6377 5525 6411 5559
rect 6411 5525 6420 5559
rect 6368 5516 6420 5525
rect 6920 5516 6972 5568
rect 7380 5516 7432 5568
rect 10048 5584 10100 5636
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 11244 5652 11296 5704
rect 11428 5652 11480 5704
rect 11612 5652 11664 5704
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 12992 5695 13044 5704
rect 11796 5652 11848 5661
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 10140 5516 10192 5568
rect 10416 5516 10468 5568
rect 11336 5516 11388 5568
rect 12900 5559 12952 5568
rect 12900 5525 12909 5559
rect 12909 5525 12943 5559
rect 12943 5525 12952 5559
rect 12900 5516 12952 5525
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 15200 5720 15252 5772
rect 15568 5763 15620 5772
rect 15568 5729 15602 5763
rect 15602 5729 15620 5763
rect 15568 5720 15620 5729
rect 15936 5720 15988 5772
rect 15292 5695 15344 5704
rect 15292 5661 15301 5695
rect 15301 5661 15335 5695
rect 15335 5661 15344 5695
rect 15292 5652 15344 5661
rect 17960 5788 18012 5840
rect 18972 5788 19024 5840
rect 19524 5865 19533 5899
rect 19533 5865 19567 5899
rect 19567 5865 19576 5899
rect 19524 5856 19576 5865
rect 20720 5788 20772 5840
rect 19340 5720 19392 5772
rect 17776 5652 17828 5704
rect 18052 5652 18104 5704
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 15568 5516 15620 5568
rect 15936 5516 15988 5568
rect 17776 5559 17828 5568
rect 17776 5525 17785 5559
rect 17785 5525 17819 5559
rect 17819 5525 17828 5559
rect 17776 5516 17828 5525
rect 19616 5559 19668 5568
rect 19616 5525 19625 5559
rect 19625 5525 19659 5559
rect 19659 5525 19668 5559
rect 19616 5516 19668 5525
rect 4280 5414 4332 5466
rect 4344 5414 4396 5466
rect 4408 5414 4460 5466
rect 4472 5414 4524 5466
rect 10878 5414 10930 5466
rect 10942 5414 10994 5466
rect 11006 5414 11058 5466
rect 11070 5414 11122 5466
rect 17475 5414 17527 5466
rect 17539 5414 17591 5466
rect 17603 5414 17655 5466
rect 17667 5414 17719 5466
rect 5816 5312 5868 5364
rect 6276 5312 6328 5364
rect 6828 5312 6880 5364
rect 7288 5355 7340 5364
rect 7288 5321 7297 5355
rect 7297 5321 7331 5355
rect 7331 5321 7340 5355
rect 7288 5312 7340 5321
rect 8024 5312 8076 5364
rect 7196 5244 7248 5296
rect 10324 5312 10376 5364
rect 11336 5312 11388 5364
rect 13084 5312 13136 5364
rect 14372 5312 14424 5364
rect 15108 5312 15160 5364
rect 7012 5176 7064 5228
rect 8668 5219 8720 5228
rect 8668 5185 8677 5219
rect 8677 5185 8711 5219
rect 8711 5185 8720 5219
rect 8668 5176 8720 5185
rect 9128 5176 9180 5228
rect 11244 5244 11296 5296
rect 12164 5244 12216 5296
rect 19340 5312 19392 5364
rect 19984 5312 20036 5364
rect 10784 5219 10836 5228
rect 4620 5151 4672 5160
rect 4620 5117 4629 5151
rect 4629 5117 4663 5151
rect 4663 5117 4672 5151
rect 4620 5108 4672 5117
rect 6000 5108 6052 5160
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 7564 5108 7616 5160
rect 10508 5108 10560 5160
rect 10784 5185 10793 5219
rect 10793 5185 10827 5219
rect 10827 5185 10836 5219
rect 10784 5176 10836 5185
rect 11704 5176 11756 5228
rect 12256 5176 12308 5228
rect 13176 5176 13228 5228
rect 13544 5108 13596 5160
rect 19892 5244 19944 5296
rect 5816 5040 5868 5092
rect 7472 4972 7524 5024
rect 7932 4972 7984 5024
rect 8116 4972 8168 5024
rect 11520 5040 11572 5092
rect 12532 5040 12584 5092
rect 15292 5108 15344 5160
rect 15752 5108 15804 5160
rect 15936 5151 15988 5160
rect 15936 5117 15970 5151
rect 15970 5117 15988 5151
rect 15936 5108 15988 5117
rect 17776 5108 17828 5160
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 19432 5176 19484 5228
rect 18696 5108 18748 5160
rect 19616 5108 19668 5160
rect 16028 5040 16080 5092
rect 11428 5015 11480 5024
rect 11428 4981 11437 5015
rect 11437 4981 11471 5015
rect 11471 4981 11480 5015
rect 11428 4972 11480 4981
rect 11612 4972 11664 5024
rect 12072 4972 12124 5024
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 14648 4972 14700 5024
rect 15200 4972 15252 5024
rect 15660 4972 15712 5024
rect 16396 4972 16448 5024
rect 19340 5040 19392 5092
rect 17224 4972 17276 5024
rect 17592 4972 17644 5024
rect 18972 4972 19024 5024
rect 7579 4870 7631 4922
rect 7643 4870 7695 4922
rect 7707 4870 7759 4922
rect 7771 4870 7823 4922
rect 14176 4870 14228 4922
rect 14240 4870 14292 4922
rect 14304 4870 14356 4922
rect 14368 4870 14420 4922
rect 6000 4811 6052 4820
rect 6000 4777 6009 4811
rect 6009 4777 6043 4811
rect 6043 4777 6052 4811
rect 6000 4768 6052 4777
rect 7196 4811 7248 4820
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 7472 4768 7524 4820
rect 9772 4768 9824 4820
rect 10048 4768 10100 4820
rect 11336 4768 11388 4820
rect 11428 4768 11480 4820
rect 12624 4811 12676 4820
rect 12624 4777 12633 4811
rect 12633 4777 12667 4811
rect 12667 4777 12676 4811
rect 12624 4768 12676 4777
rect 15016 4768 15068 4820
rect 15660 4811 15712 4820
rect 15660 4777 15669 4811
rect 15669 4777 15703 4811
rect 15703 4777 15712 4811
rect 15660 4768 15712 4777
rect 15844 4768 15896 4820
rect 19340 4768 19392 4820
rect 19800 4768 19852 4820
rect 6092 4700 6144 4752
rect 9680 4700 9732 4752
rect 4620 4632 4672 4684
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 7656 4675 7708 4684
rect 7656 4641 7665 4675
rect 7665 4641 7699 4675
rect 7699 4641 7708 4675
rect 7656 4632 7708 4641
rect 8852 4675 8904 4684
rect 8852 4641 8861 4675
rect 8861 4641 8895 4675
rect 8895 4641 8904 4675
rect 8852 4632 8904 4641
rect 9036 4632 9088 4684
rect 9496 4632 9548 4684
rect 12808 4700 12860 4752
rect 14188 4700 14240 4752
rect 15568 4700 15620 4752
rect 19708 4700 19760 4752
rect 11980 4675 12032 4684
rect 11980 4641 11989 4675
rect 11989 4641 12023 4675
rect 12023 4641 12032 4675
rect 11980 4632 12032 4641
rect 12072 4632 12124 4684
rect 12992 4632 13044 4684
rect 6828 4564 6880 4616
rect 7472 4564 7524 4616
rect 9588 4564 9640 4616
rect 5908 4539 5960 4548
rect 5908 4505 5917 4539
rect 5917 4505 5951 4539
rect 5951 4505 5960 4539
rect 5908 4496 5960 4505
rect 7196 4496 7248 4548
rect 9128 4539 9180 4548
rect 9128 4505 9137 4539
rect 9137 4505 9171 4539
rect 9171 4505 9180 4539
rect 9128 4496 9180 4505
rect 8024 4471 8076 4480
rect 8024 4437 8033 4471
rect 8033 4437 8067 4471
rect 8067 4437 8076 4471
rect 8024 4428 8076 4437
rect 10140 4607 10192 4616
rect 10140 4573 10152 4607
rect 10152 4573 10186 4607
rect 10186 4573 10192 4607
rect 10140 4564 10192 4573
rect 11888 4564 11940 4616
rect 12440 4564 12492 4616
rect 13360 4564 13412 4616
rect 11336 4496 11388 4548
rect 11244 4428 11296 4480
rect 11428 4428 11480 4480
rect 11796 4428 11848 4480
rect 13544 4632 13596 4684
rect 15108 4675 15160 4684
rect 15108 4641 15117 4675
rect 15117 4641 15151 4675
rect 15151 4641 15160 4675
rect 15108 4632 15160 4641
rect 16396 4675 16448 4684
rect 15200 4564 15252 4616
rect 15384 4496 15436 4548
rect 16396 4641 16419 4675
rect 16419 4641 16448 4675
rect 16396 4632 16448 4641
rect 17316 4632 17368 4684
rect 18144 4632 18196 4684
rect 20536 4632 20588 4684
rect 17592 4607 17644 4616
rect 14832 4471 14884 4480
rect 14832 4437 14841 4471
rect 14841 4437 14875 4471
rect 14875 4437 14884 4471
rect 14832 4428 14884 4437
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 15752 4428 15804 4480
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 19156 4607 19208 4616
rect 19156 4573 19165 4607
rect 19165 4573 19199 4607
rect 19199 4573 19208 4607
rect 19156 4564 19208 4573
rect 17040 4428 17092 4480
rect 18604 4428 18656 4480
rect 4280 4326 4332 4378
rect 4344 4326 4396 4378
rect 4408 4326 4460 4378
rect 4472 4326 4524 4378
rect 10878 4326 10930 4378
rect 10942 4326 10994 4378
rect 11006 4326 11058 4378
rect 11070 4326 11122 4378
rect 17475 4326 17527 4378
rect 17539 4326 17591 4378
rect 17603 4326 17655 4378
rect 17667 4326 17719 4378
rect 5816 4267 5868 4276
rect 5816 4233 5825 4267
rect 5825 4233 5859 4267
rect 5859 4233 5868 4267
rect 5816 4224 5868 4233
rect 6368 4224 6420 4276
rect 7656 4224 7708 4276
rect 7932 4224 7984 4276
rect 9680 4224 9732 4276
rect 12624 4224 12676 4276
rect 14188 4267 14240 4276
rect 6736 4156 6788 4208
rect 7472 4156 7524 4208
rect 9404 4088 9456 4140
rect 10876 4156 10928 4208
rect 14188 4233 14197 4267
rect 14197 4233 14231 4267
rect 14231 4233 14240 4267
rect 14188 4224 14240 4233
rect 17224 4224 17276 4276
rect 19800 4224 19852 4276
rect 4436 4063 4488 4072
rect 4436 4029 4445 4063
rect 4445 4029 4479 4063
rect 4479 4029 4488 4063
rect 4436 4020 4488 4029
rect 5908 4020 5960 4072
rect 6276 4063 6328 4072
rect 6276 4029 6285 4063
rect 6285 4029 6319 4063
rect 6319 4029 6328 4063
rect 6276 4020 6328 4029
rect 8024 4020 8076 4072
rect 8116 4020 8168 4072
rect 9128 4020 9180 4072
rect 9864 4063 9916 4072
rect 9864 4029 9873 4063
rect 9873 4029 9907 4063
rect 9907 4029 9916 4063
rect 9864 4020 9916 4029
rect 11060 4088 11112 4140
rect 11796 4088 11848 4140
rect 14832 4156 14884 4208
rect 12348 4088 12400 4140
rect 15108 4088 15160 4140
rect 15292 4088 15344 4140
rect 17960 4156 18012 4208
rect 12072 4020 12124 4072
rect 14832 4020 14884 4072
rect 14924 4020 14976 4072
rect 18696 4156 18748 4208
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 8392 3884 8444 3936
rect 11060 3952 11112 4004
rect 15476 3952 15528 4004
rect 13268 3884 13320 3936
rect 14556 3927 14608 3936
rect 14556 3893 14565 3927
rect 14565 3893 14599 3927
rect 14599 3893 14608 3927
rect 14556 3884 14608 3893
rect 14648 3927 14700 3936
rect 14648 3893 14657 3927
rect 14657 3893 14691 3927
rect 14691 3893 14700 3927
rect 18236 4020 18288 4072
rect 19156 4063 19208 4072
rect 19156 4029 19165 4063
rect 19165 4029 19199 4063
rect 19199 4029 19208 4063
rect 19156 4020 19208 4029
rect 14648 3884 14700 3893
rect 16672 3927 16724 3936
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 16764 3927 16816 3936
rect 16764 3893 16773 3927
rect 16773 3893 16807 3927
rect 16807 3893 16816 3927
rect 17132 3927 17184 3936
rect 16764 3884 16816 3893
rect 17132 3893 17141 3927
rect 17141 3893 17175 3927
rect 17175 3893 17184 3927
rect 17132 3884 17184 3893
rect 17776 3884 17828 3936
rect 18696 3884 18748 3936
rect 20444 3952 20496 4004
rect 19800 3884 19852 3936
rect 7579 3782 7631 3834
rect 7643 3782 7695 3834
rect 7707 3782 7759 3834
rect 7771 3782 7823 3834
rect 14176 3782 14228 3834
rect 14240 3782 14292 3834
rect 14304 3782 14356 3834
rect 14368 3782 14420 3834
rect 4804 3680 4856 3732
rect 6368 3612 6420 3664
rect 4436 3587 4488 3596
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 6276 3544 6328 3596
rect 6460 3587 6512 3596
rect 6460 3553 6494 3587
rect 6494 3553 6512 3587
rect 6460 3544 6512 3553
rect 9680 3612 9732 3664
rect 12256 3680 12308 3732
rect 12348 3612 12400 3664
rect 14556 3680 14608 3732
rect 15660 3680 15712 3732
rect 18696 3723 18748 3732
rect 18696 3689 18705 3723
rect 18705 3689 18739 3723
rect 18739 3689 18748 3723
rect 18696 3680 18748 3689
rect 20444 3680 20496 3732
rect 16764 3612 16816 3664
rect 17132 3612 17184 3664
rect 8116 3587 8168 3596
rect 6092 3408 6144 3460
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 9312 3544 9364 3596
rect 9588 3476 9640 3528
rect 10324 3519 10376 3528
rect 10324 3485 10333 3519
rect 10333 3485 10367 3519
rect 10367 3485 10376 3519
rect 10324 3476 10376 3485
rect 10692 3476 10744 3528
rect 10784 3519 10836 3528
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 11152 3476 11204 3528
rect 11336 3476 11388 3528
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 12164 3544 12216 3596
rect 12992 3476 13044 3528
rect 13176 3519 13228 3528
rect 13176 3485 13188 3519
rect 13188 3485 13222 3519
rect 13222 3485 13228 3519
rect 13176 3476 13228 3485
rect 13544 3544 13596 3596
rect 14924 3544 14976 3596
rect 15016 3544 15068 3596
rect 15844 3587 15896 3596
rect 15844 3553 15878 3587
rect 15878 3553 15896 3587
rect 15844 3544 15896 3553
rect 17316 3587 17368 3596
rect 17316 3553 17350 3587
rect 17350 3553 17368 3587
rect 17316 3544 17368 3553
rect 19984 3544 20036 3596
rect 15476 3476 15528 3528
rect 15568 3519 15620 3528
rect 15568 3485 15577 3519
rect 15577 3485 15611 3519
rect 15611 3485 15620 3519
rect 17040 3519 17092 3528
rect 15568 3476 15620 3485
rect 9128 3408 9180 3460
rect 6552 3340 6604 3392
rect 9312 3340 9364 3392
rect 9772 3408 9824 3460
rect 14648 3408 14700 3460
rect 12256 3340 12308 3392
rect 12900 3340 12952 3392
rect 13544 3340 13596 3392
rect 15568 3340 15620 3392
rect 17040 3485 17049 3519
rect 17049 3485 17083 3519
rect 17083 3485 17092 3519
rect 17040 3476 17092 3485
rect 18696 3476 18748 3528
rect 19156 3519 19208 3528
rect 19156 3485 19165 3519
rect 19165 3485 19199 3519
rect 19199 3485 19208 3519
rect 19156 3476 19208 3485
rect 17224 3340 17276 3392
rect 4280 3238 4332 3290
rect 4344 3238 4396 3290
rect 4408 3238 4460 3290
rect 4472 3238 4524 3290
rect 10878 3238 10930 3290
rect 10942 3238 10994 3290
rect 11006 3238 11058 3290
rect 11070 3238 11122 3290
rect 17475 3238 17527 3290
rect 17539 3238 17591 3290
rect 17603 3238 17655 3290
rect 17667 3238 17719 3290
rect 4712 3136 4764 3188
rect 6460 3136 6512 3188
rect 9036 3136 9088 3188
rect 9496 3136 9548 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 11244 3136 11296 3188
rect 5080 3043 5132 3052
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 6276 3000 6328 3052
rect 4804 2975 4856 2984
rect 4804 2941 4813 2975
rect 4813 2941 4847 2975
rect 4847 2941 4856 2975
rect 4804 2932 4856 2941
rect 6552 2932 6604 2984
rect 6736 2932 6788 2984
rect 6920 2932 6972 2984
rect 6276 2864 6328 2916
rect 8208 2932 8260 2984
rect 7012 2796 7064 2848
rect 8300 2796 8352 2848
rect 9404 2932 9456 2984
rect 12440 3136 12492 3188
rect 12624 3136 12676 3188
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 11980 3000 12032 3052
rect 15108 3136 15160 3188
rect 15476 3136 15528 3188
rect 16672 3136 16724 3188
rect 19984 3136 20036 3188
rect 10692 2864 10744 2916
rect 12072 2932 12124 2984
rect 13268 2932 13320 2984
rect 13912 2975 13964 2984
rect 13912 2941 13921 2975
rect 13921 2941 13955 2975
rect 13955 2941 13964 2975
rect 13912 2932 13964 2941
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 17316 3000 17368 3052
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 16212 2932 16264 2984
rect 17040 2932 17092 2984
rect 17684 2932 17736 2984
rect 19248 2932 19300 2984
rect 20076 2932 20128 2984
rect 11520 2796 11572 2848
rect 13084 2796 13136 2848
rect 15660 2864 15712 2916
rect 17224 2864 17276 2916
rect 17592 2864 17644 2916
rect 18052 2864 18104 2916
rect 18972 2907 19024 2916
rect 18972 2873 19006 2907
rect 19006 2873 19024 2907
rect 18972 2864 19024 2873
rect 16212 2796 16264 2848
rect 7579 2694 7631 2746
rect 7643 2694 7695 2746
rect 7707 2694 7759 2746
rect 7771 2694 7823 2746
rect 14176 2694 14228 2746
rect 14240 2694 14292 2746
rect 14304 2694 14356 2746
rect 14368 2694 14420 2746
rect 6460 2635 6512 2644
rect 6460 2601 6469 2635
rect 6469 2601 6503 2635
rect 6503 2601 6512 2635
rect 6460 2592 6512 2601
rect 6828 2592 6880 2644
rect 8300 2635 8352 2644
rect 6368 2567 6420 2576
rect 6368 2533 6377 2567
rect 6377 2533 6411 2567
rect 6411 2533 6420 2567
rect 6368 2524 6420 2533
rect 7012 2524 7064 2576
rect 6736 2456 6788 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 11888 2592 11940 2644
rect 12900 2592 12952 2644
rect 13360 2592 13412 2644
rect 17316 2635 17368 2644
rect 17316 2601 17325 2635
rect 17325 2601 17359 2635
rect 17359 2601 17368 2635
rect 17316 2592 17368 2601
rect 17776 2592 17828 2644
rect 18972 2592 19024 2644
rect 19800 2635 19852 2644
rect 19800 2601 19809 2635
rect 19809 2601 19843 2635
rect 19843 2601 19852 2635
rect 19800 2592 19852 2601
rect 19984 2592 20036 2644
rect 11704 2524 11756 2576
rect 15108 2524 15160 2576
rect 16212 2567 16264 2576
rect 16212 2533 16246 2567
rect 16246 2533 16264 2567
rect 16212 2524 16264 2533
rect 9864 2456 9916 2508
rect 10324 2456 10376 2508
rect 12532 2456 12584 2508
rect 13912 2499 13964 2508
rect 13912 2465 13921 2499
rect 13921 2465 13955 2499
rect 13955 2465 13964 2499
rect 13912 2456 13964 2465
rect 15476 2456 15528 2508
rect 20444 2524 20496 2576
rect 18604 2499 18656 2508
rect 18604 2465 18638 2499
rect 18638 2465 18656 2499
rect 18604 2456 18656 2465
rect 13084 2388 13136 2440
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 18052 2431 18104 2440
rect 18052 2397 18061 2431
rect 18061 2397 18095 2431
rect 18095 2397 18104 2431
rect 18052 2388 18104 2397
rect 8392 2363 8444 2372
rect 8392 2329 8401 2363
rect 8401 2329 8435 2363
rect 8435 2329 8444 2363
rect 8392 2320 8444 2329
rect 17684 2320 17736 2372
rect 5356 2252 5408 2304
rect 7196 2252 7248 2304
rect 11704 2295 11756 2304
rect 11704 2261 11713 2295
rect 11713 2261 11747 2295
rect 11747 2261 11756 2295
rect 11704 2252 11756 2261
rect 18052 2252 18104 2304
rect 4280 2150 4332 2202
rect 4344 2150 4396 2202
rect 4408 2150 4460 2202
rect 4472 2150 4524 2202
rect 10878 2150 10930 2202
rect 10942 2150 10994 2202
rect 11006 2150 11058 2202
rect 11070 2150 11122 2202
rect 17475 2150 17527 2202
rect 17539 2150 17591 2202
rect 17603 2150 17655 2202
rect 17667 2150 17719 2202
rect 1768 1232 1820 1284
rect 9588 1232 9640 1284
<< metal2 >>
rect 294 21520 350 22000
rect 846 21520 902 22000
rect 1490 21520 1546 22000
rect 2042 21520 2098 22000
rect 2686 21520 2742 22000
rect 3330 21520 3386 22000
rect 3882 21520 3938 22000
rect 4526 21520 4582 22000
rect 5170 21520 5226 22000
rect 5722 21520 5778 22000
rect 6366 21520 6422 22000
rect 7010 21520 7066 22000
rect 7562 21520 7618 22000
rect 8206 21520 8262 22000
rect 8758 21520 8814 22000
rect 9402 21520 9458 22000
rect 10046 21520 10102 22000
rect 10598 21520 10654 22000
rect 11242 21520 11298 22000
rect 11886 21520 11942 22000
rect 12438 21520 12494 22000
rect 13082 21520 13138 22000
rect 13726 21520 13782 22000
rect 14278 21520 14334 22000
rect 14922 21520 14978 22000
rect 15474 21520 15530 22000
rect 16118 21520 16174 22000
rect 16394 21720 16450 21729
rect 16394 21655 16450 21664
rect 308 18630 336 21520
rect 860 18970 888 21520
rect 1504 19242 1532 21520
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1492 19236 1544 19242
rect 1492 19178 1544 19184
rect 848 18964 900 18970
rect 848 18906 900 18912
rect 296 18624 348 18630
rect 296 18566 348 18572
rect 1596 18408 1624 19246
rect 1676 19168 1728 19174
rect 2056 19156 2084 21520
rect 1676 19110 1728 19116
rect 1780 19128 2084 19156
rect 2136 19168 2188 19174
rect 1688 18970 1716 19110
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1596 18380 1716 18408
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1306 17776 1362 17785
rect 1412 17746 1440 18158
rect 1688 17746 1716 18380
rect 1306 17711 1362 17720
rect 1400 17740 1452 17746
rect 1320 17134 1348 17711
rect 1400 17682 1452 17688
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1412 17218 1440 17682
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1412 17190 1532 17218
rect 1504 17134 1532 17190
rect 1308 17128 1360 17134
rect 1308 17070 1360 17076
rect 1492 17128 1544 17134
rect 1492 17070 1544 17076
rect 1504 16658 1532 17070
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1596 16590 1624 17478
rect 1688 16998 1716 17682
rect 1780 17270 1808 19128
rect 2136 19110 2188 19116
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 1768 17264 1820 17270
rect 1768 17206 1820 17212
rect 2148 17066 2176 19110
rect 2410 19000 2466 19009
rect 2410 18935 2466 18944
rect 2424 18834 2452 18935
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2240 18222 2268 18770
rect 2424 18426 2452 18770
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2412 17604 2464 17610
rect 2412 17546 2464 17552
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 2148 16726 2176 17002
rect 2424 16810 2452 17546
rect 2332 16794 2452 16810
rect 2320 16788 2452 16794
rect 2372 16782 2452 16788
rect 2320 16730 2372 16736
rect 2044 16720 2096 16726
rect 2042 16688 2044 16697
rect 2136 16720 2188 16726
rect 2096 16688 2098 16697
rect 1860 16652 1912 16658
rect 2136 16662 2188 16668
rect 2042 16623 2098 16632
rect 1860 16594 1912 16600
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1872 16114 1900 16594
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1872 15570 1900 16050
rect 2608 15978 2636 19110
rect 2700 17066 2728 21520
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2792 17882 2820 18090
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 2596 15972 2648 15978
rect 2596 15914 2648 15920
rect 2884 15638 2912 19110
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2976 15910 3004 16390
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1872 15162 1900 15506
rect 2884 15162 2912 15574
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1412 14482 1440 14962
rect 2964 14952 3016 14958
rect 3068 14940 3096 19110
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3160 17134 3188 18906
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3252 15570 3280 16934
rect 3344 16522 3372 21520
rect 3896 19394 3924 21520
rect 4540 19802 4568 21520
rect 4540 19774 4660 19802
rect 4254 19612 4550 19632
rect 4310 19610 4334 19612
rect 4390 19610 4414 19612
rect 4470 19610 4494 19612
rect 4332 19558 4334 19610
rect 4396 19558 4408 19610
rect 4470 19558 4472 19610
rect 4310 19556 4334 19558
rect 4390 19556 4414 19558
rect 4470 19556 4494 19558
rect 4254 19536 4550 19556
rect 3896 19366 4016 19394
rect 3988 19292 4016 19366
rect 4160 19304 4212 19310
rect 3988 19264 4160 19292
rect 4160 19246 4212 19252
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3620 18986 3648 19178
rect 4068 19168 4120 19174
rect 3974 19136 4030 19145
rect 4068 19110 4120 19116
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 3974 19071 4030 19080
rect 3528 18970 3648 18986
rect 3528 18964 3660 18970
rect 3528 18958 3608 18964
rect 3528 18222 3556 18958
rect 3608 18906 3660 18912
rect 3606 18864 3662 18873
rect 3606 18799 3608 18808
rect 3660 18799 3662 18808
rect 3608 18770 3660 18776
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3896 18426 3924 18566
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 3422 17912 3478 17921
rect 3422 17847 3478 17856
rect 3436 16697 3464 17847
rect 3516 17060 3568 17066
rect 3516 17002 3568 17008
rect 3528 16794 3556 17002
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3422 16688 3478 16697
rect 3422 16623 3478 16632
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 3436 16182 3464 16623
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 3620 16114 3648 18158
rect 3988 17814 4016 19071
rect 4080 17882 4108 19110
rect 4172 18816 4200 19110
rect 4632 18970 4660 19774
rect 4896 19440 4948 19446
rect 4896 19382 4948 19388
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4712 19168 4764 19174
rect 4816 19145 4844 19178
rect 4712 19110 4764 19116
rect 4802 19136 4858 19145
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4335 18828 4387 18834
rect 4172 18788 4335 18816
rect 4172 18426 4200 18788
rect 4335 18770 4387 18776
rect 4254 18524 4550 18544
rect 4310 18522 4334 18524
rect 4390 18522 4414 18524
rect 4470 18522 4494 18524
rect 4332 18470 4334 18522
rect 4396 18470 4408 18522
rect 4470 18470 4472 18522
rect 4310 18468 4334 18470
rect 4390 18468 4414 18470
rect 4470 18468 4494 18470
rect 4254 18448 4550 18468
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 3976 17808 4028 17814
rect 3976 17750 4028 17756
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3896 17202 3924 17614
rect 3974 17232 4030 17241
rect 3884 17196 3936 17202
rect 3974 17167 4030 17176
rect 3884 17138 3936 17144
rect 3698 17096 3754 17105
rect 3698 17031 3754 17040
rect 3712 16658 3740 17031
rect 3700 16652 3752 16658
rect 3752 16612 3832 16640
rect 3700 16594 3752 16600
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3620 15434 3648 16050
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3608 15428 3660 15434
rect 3608 15370 3660 15376
rect 3016 14912 3096 14940
rect 2964 14894 3016 14900
rect 3068 14550 3096 14912
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3344 14550 3372 14894
rect 3056 14544 3108 14550
rect 3056 14486 3108 14492
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1412 13938 1440 14418
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3068 14074 3096 14350
rect 3056 14068 3108 14074
rect 3108 14028 3280 14056
rect 3056 14010 3108 14016
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12782 1440 13262
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 12306 1440 12718
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1400 11144 1452 11150
rect 1504 11121 1532 11154
rect 1400 11086 1452 11092
rect 1490 11112 1546 11121
rect 1412 10606 1440 11086
rect 1490 11047 1546 11056
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1872 9654 1900 12582
rect 2516 11762 2544 13398
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2884 12986 2912 13330
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2976 12782 3004 13874
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 12442 2820 12650
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2976 12170 3004 12718
rect 3160 12306 3188 13466
rect 3252 12782 3280 14028
rect 3344 13734 3372 14350
rect 3528 14074 3556 14894
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3620 13802 3648 14282
rect 3608 13796 3660 13802
rect 3608 13738 3660 13744
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3344 13410 3372 13670
rect 3712 13530 3740 15982
rect 3804 15450 3832 16612
rect 3896 16046 3924 17138
rect 3988 16726 4016 17167
rect 4172 17134 4200 18022
rect 4620 17672 4672 17678
rect 4724 17660 4752 19110
rect 4802 19071 4858 19080
rect 4908 18970 4936 19382
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 5092 18290 5120 19314
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 4816 17921 4844 18022
rect 4802 17912 4858 17921
rect 4802 17847 4858 17856
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 4672 17632 4752 17660
rect 4804 17672 4856 17678
rect 4620 17614 4672 17620
rect 4804 17614 4856 17620
rect 4254 17436 4550 17456
rect 4310 17434 4334 17436
rect 4390 17434 4414 17436
rect 4470 17434 4494 17436
rect 4332 17382 4334 17434
rect 4396 17382 4408 17434
rect 4470 17382 4472 17434
rect 4310 17380 4334 17382
rect 4390 17380 4414 17382
rect 4470 17380 4494 17382
rect 4254 17360 4550 17380
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 4080 16114 4108 16934
rect 4356 16794 4384 17002
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4172 16250 4200 16594
rect 4254 16348 4550 16368
rect 4310 16346 4334 16348
rect 4390 16346 4414 16348
rect 4470 16346 4494 16348
rect 4332 16294 4334 16346
rect 4396 16294 4408 16346
rect 4470 16294 4472 16346
rect 4310 16292 4334 16294
rect 4390 16292 4414 16294
rect 4470 16292 4494 16294
rect 4254 16272 4550 16292
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 3884 16040 3936 16046
rect 4264 15994 4292 16050
rect 3884 15982 3936 15988
rect 4080 15966 4292 15994
rect 4080 15910 4108 15966
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4080 15502 4108 15846
rect 4632 15638 4660 16934
rect 4724 16590 4752 17138
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4620 15632 4672 15638
rect 4620 15574 4672 15580
rect 4068 15496 4120 15502
rect 3804 15422 3924 15450
rect 4068 15438 4120 15444
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 14482 3832 15302
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 3344 13382 3464 13410
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3344 12714 3372 13262
rect 3436 13190 3464 13382
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3528 12238 3556 13262
rect 3516 12232 3568 12238
rect 3344 12192 3516 12220
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 3344 11762 3372 12192
rect 3516 12174 3568 12180
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 2332 11354 2360 11494
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 10606 2820 11018
rect 2870 10704 2926 10713
rect 2870 10639 2926 10648
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2884 10146 2912 10639
rect 3160 10606 3188 11494
rect 3344 11286 3372 11698
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3804 11218 3832 14214
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3252 10810 3280 11154
rect 3330 11112 3386 11121
rect 3330 11047 3386 11056
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3160 10266 3188 10542
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3252 10198 3280 10746
rect 2792 10118 2912 10146
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 2226 9480 2282 9489
rect 2226 9415 2228 9424
rect 2280 9415 2282 9424
rect 2228 9386 2280 9392
rect 2410 9344 2466 9353
rect 2410 9279 2466 9288
rect 2424 8634 2452 9279
rect 2686 9208 2742 9217
rect 2686 9143 2688 9152
rect 2740 9143 2742 9152
rect 2688 9114 2740 9120
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2700 8401 2728 8842
rect 2792 8430 2820 10118
rect 2964 9648 3016 9654
rect 2962 9616 2964 9625
rect 3016 9616 3018 9625
rect 2962 9551 3018 9560
rect 3344 9518 3372 11047
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 9518 3832 9998
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8498 2912 8774
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2780 8424 2832 8430
rect 2686 8392 2742 8401
rect 2780 8366 2832 8372
rect 2686 8327 2742 8336
rect 2976 8129 3004 8978
rect 3344 8809 3372 9318
rect 3436 9081 3464 9318
rect 3804 9178 3832 9454
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3422 9072 3478 9081
rect 3422 9007 3478 9016
rect 3330 8800 3386 8809
rect 3330 8735 3386 8744
rect 3896 8634 3924 15422
rect 4080 15162 4108 15438
rect 4254 15260 4550 15280
rect 4310 15258 4334 15260
rect 4390 15258 4414 15260
rect 4470 15258 4494 15260
rect 4332 15206 4334 15258
rect 4396 15206 4408 15258
rect 4470 15206 4472 15258
rect 4310 15204 4334 15206
rect 4390 15204 4414 15206
rect 4470 15204 4494 15206
rect 4254 15184 4550 15204
rect 4632 15162 4660 15574
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3988 13394 4016 14418
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 3988 12102 4016 13330
rect 4080 12918 4108 15098
rect 4172 14890 4200 15098
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4620 14408 4672 14414
rect 4724 14396 4752 15846
rect 4816 15706 4844 17614
rect 4908 17082 4936 17818
rect 5000 17814 5028 18022
rect 4988 17808 5040 17814
rect 4988 17750 5040 17756
rect 5092 17218 5120 18226
rect 5000 17202 5120 17218
rect 4988 17196 5120 17202
rect 5040 17190 5120 17196
rect 4988 17138 5040 17144
rect 5080 17128 5132 17134
rect 4908 17054 5028 17082
rect 5080 17070 5132 17076
rect 5000 16998 5028 17054
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4896 16720 4948 16726
rect 4896 16662 4948 16668
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4672 14368 4752 14396
rect 4620 14350 4672 14356
rect 4172 13954 4200 14350
rect 4254 14172 4550 14192
rect 4310 14170 4334 14172
rect 4390 14170 4414 14172
rect 4470 14170 4494 14172
rect 4332 14118 4334 14170
rect 4396 14118 4408 14170
rect 4470 14118 4472 14170
rect 4310 14116 4334 14118
rect 4390 14116 4414 14118
rect 4470 14116 4494 14118
rect 4254 14096 4550 14116
rect 4172 13926 4292 13954
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 12986 4200 13806
rect 4264 13326 4292 13926
rect 4632 13530 4660 14350
rect 4816 13954 4844 15302
rect 4908 15094 4936 16662
rect 5000 16250 5028 16934
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5092 15366 5120 17070
rect 5184 15570 5212 21520
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5460 19281 5488 19314
rect 5446 19272 5502 19281
rect 5446 19207 5502 19216
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5276 19009 5304 19110
rect 5262 19000 5318 19009
rect 5262 18935 5318 18944
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5276 18290 5304 18566
rect 5736 18306 5764 21520
rect 6380 19292 6408 21520
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6460 19304 6512 19310
rect 6380 19264 6460 19292
rect 6460 19246 6512 19252
rect 6276 19168 6328 19174
rect 6328 19128 6408 19156
rect 6276 19110 6328 19116
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5644 18278 5764 18306
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5552 17202 5580 17614
rect 5356 17196 5408 17202
rect 5540 17196 5592 17202
rect 5408 17156 5488 17184
rect 5356 17138 5408 17144
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 4896 15088 4948 15094
rect 4896 15030 4948 15036
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 5000 14074 5028 14486
rect 5092 14482 5120 15302
rect 5460 15042 5488 17156
rect 5540 17138 5592 17144
rect 5644 17082 5672 18278
rect 5724 18148 5776 18154
rect 5724 18090 5776 18096
rect 5736 17338 5764 18090
rect 6288 17814 6316 18770
rect 6380 18290 6408 19128
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6472 18222 6500 18566
rect 6460 18216 6512 18222
rect 6460 18158 6512 18164
rect 6276 17808 6328 17814
rect 6276 17750 6328 17756
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 5816 17672 5868 17678
rect 5920 17649 5948 17682
rect 5816 17614 5868 17620
rect 5906 17640 5962 17649
rect 5828 17338 5856 17614
rect 5906 17575 5962 17584
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 6472 17202 6500 18158
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 5552 17054 5672 17082
rect 5552 16046 5580 17054
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5644 16794 5672 16934
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5736 16250 5764 17138
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5828 15162 5856 16594
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 6012 15910 6040 16526
rect 6104 16454 6132 16934
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6564 16153 6592 19314
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18193 6868 19110
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6826 18184 6882 18193
rect 6826 18119 6882 18128
rect 6932 17814 6960 18226
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6656 17134 6684 17614
rect 6748 17202 6776 17750
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6932 16794 6960 17070
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6550 16144 6606 16153
rect 6550 16079 6606 16088
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 15638 6224 15846
rect 6840 15638 6868 15914
rect 6932 15706 6960 16730
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5460 15026 5580 15042
rect 6196 15026 6224 15574
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 5460 15020 5592 15026
rect 5460 15014 5540 15020
rect 5540 14962 5592 14968
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6840 14958 6868 15370
rect 6932 15366 6960 15506
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6932 14890 6960 15302
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 5276 14074 5304 14418
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 4816 13938 5028 13954
rect 4816 13932 5040 13938
rect 4816 13926 4988 13932
rect 4988 13874 5040 13880
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4254 13084 4550 13104
rect 4310 13082 4334 13084
rect 4390 13082 4414 13084
rect 4470 13082 4494 13084
rect 4332 13030 4334 13082
rect 4396 13030 4408 13082
rect 4470 13030 4472 13082
rect 4310 13028 4334 13030
rect 4390 13028 4414 13030
rect 4470 13028 4494 13030
rect 4254 13008 4550 13028
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 4172 12442 4200 12650
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3976 11688 4028 11694
rect 4080 11676 4108 12174
rect 4254 11996 4550 12016
rect 4310 11994 4334 11996
rect 4390 11994 4414 11996
rect 4470 11994 4494 11996
rect 4332 11942 4334 11994
rect 4396 11942 4408 11994
rect 4470 11942 4472 11994
rect 4310 11940 4334 11942
rect 4390 11940 4414 11942
rect 4470 11940 4494 11942
rect 4254 11920 4550 11940
rect 4028 11648 4108 11676
rect 3976 11630 4028 11636
rect 4080 11014 4108 11648
rect 4632 11626 4660 13330
rect 4724 12782 4752 13670
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10606 4108 10950
rect 4172 10810 4200 11494
rect 4620 11212 4672 11218
rect 4816 11200 4844 13398
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4908 11898 4936 13330
rect 5000 13326 5028 13874
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5092 12986 5120 13262
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5552 12918 5580 14350
rect 6104 13870 6132 14418
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6104 13530 6132 13806
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6288 13462 6316 13670
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 5828 12986 5856 13398
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5920 12306 5948 12922
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5368 11898 5396 12242
rect 6288 12238 6316 12922
rect 6380 12850 6408 13126
rect 6840 12986 6868 14486
rect 7024 13938 7052 21520
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7104 19168 7156 19174
rect 7156 19128 7420 19156
rect 7104 19110 7156 19116
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7116 16794 7144 18702
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7300 17746 7328 18294
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7300 16794 7328 17682
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7116 16046 7144 16594
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7208 15706 7236 16458
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7300 16114 7328 16390
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7208 14890 7236 15642
rect 7392 14958 7420 19128
rect 7484 17785 7512 19450
rect 7576 19310 7604 21520
rect 8220 19530 8248 21520
rect 7944 19502 8248 19530
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7553 19068 7849 19088
rect 7609 19066 7633 19068
rect 7689 19066 7713 19068
rect 7769 19066 7793 19068
rect 7631 19014 7633 19066
rect 7695 19014 7707 19066
rect 7769 19014 7771 19066
rect 7609 19012 7633 19014
rect 7689 19012 7713 19014
rect 7769 19012 7793 19014
rect 7553 18992 7849 19012
rect 7553 17980 7849 18000
rect 7609 17978 7633 17980
rect 7689 17978 7713 17980
rect 7769 17978 7793 17980
rect 7631 17926 7633 17978
rect 7695 17926 7707 17978
rect 7769 17926 7771 17978
rect 7609 17924 7633 17926
rect 7689 17924 7713 17926
rect 7769 17924 7793 17926
rect 7553 17904 7849 17924
rect 7944 17814 7972 19502
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8024 19168 8076 19174
rect 8024 19110 8076 19116
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 8036 18970 8064 19110
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 7932 17808 7984 17814
rect 7470 17776 7526 17785
rect 7932 17750 7984 17756
rect 7470 17711 7526 17720
rect 8036 17610 8064 18770
rect 8128 17610 8156 19110
rect 8220 18630 8248 19314
rect 8298 19272 8354 19281
rect 8298 19207 8354 19216
rect 8312 19174 8340 19207
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18154 8248 18566
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8208 18148 8260 18154
rect 8208 18090 8260 18096
rect 8024 17604 8076 17610
rect 8024 17546 8076 17552
rect 8116 17604 8168 17610
rect 8116 17546 8168 17552
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7484 16590 7512 17002
rect 7944 16998 7972 17138
rect 8496 17134 8524 18158
rect 8666 17640 8722 17649
rect 8666 17575 8722 17584
rect 8680 17338 8708 17575
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8484 17128 8536 17134
rect 8220 17076 8484 17082
rect 8220 17070 8536 17076
rect 8220 17054 8524 17070
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 7553 16892 7849 16912
rect 7609 16890 7633 16892
rect 7689 16890 7713 16892
rect 7769 16890 7793 16892
rect 7631 16838 7633 16890
rect 7695 16838 7707 16890
rect 7769 16838 7771 16890
rect 7609 16836 7633 16838
rect 7689 16836 7713 16838
rect 7769 16836 7793 16838
rect 7553 16816 7849 16836
rect 8036 16776 8064 16934
rect 7852 16748 8064 16776
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7852 16114 7880 16748
rect 7944 16646 8156 16674
rect 7944 16250 7972 16646
rect 8128 16590 8156 16646
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7840 16108 7892 16114
rect 7484 16068 7840 16096
rect 7380 14952 7432 14958
rect 7300 14912 7380 14940
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7116 13870 7144 14486
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6840 12850 6868 12922
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6932 12442 6960 13330
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5354 11656 5410 11665
rect 5354 11591 5410 11600
rect 5448 11620 5500 11626
rect 4672 11172 4844 11200
rect 4620 11154 4672 11160
rect 4254 10908 4550 10928
rect 4310 10906 4334 10908
rect 4390 10906 4414 10908
rect 4470 10906 4494 10908
rect 4332 10854 4334 10906
rect 4396 10854 4408 10906
rect 4470 10854 4472 10906
rect 4310 10852 4334 10854
rect 4390 10852 4414 10854
rect 4470 10852 4494 10854
rect 4254 10832 4550 10852
rect 4632 10810 4660 11154
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 3974 10160 4030 10169
rect 4172 10130 4200 10474
rect 3974 10095 4030 10104
rect 4160 10124 4212 10130
rect 3988 9110 4016 10095
rect 4160 10066 4212 10072
rect 5172 10056 5224 10062
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 5078 10024 5134 10033
rect 5172 9998 5224 10004
rect 5078 9959 5134 9968
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3054 8528 3110 8537
rect 3988 8498 4016 8774
rect 3054 8463 3056 8472
rect 3108 8463 3110 8472
rect 3884 8492 3936 8498
rect 3056 8434 3108 8440
rect 3884 8434 3936 8440
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3896 8265 3924 8434
rect 4080 8430 4108 9959
rect 4254 9820 4550 9840
rect 4310 9818 4334 9820
rect 4390 9818 4414 9820
rect 4470 9818 4494 9820
rect 4332 9766 4334 9818
rect 4396 9766 4408 9818
rect 4470 9766 4472 9818
rect 4310 9764 4334 9766
rect 4390 9764 4414 9766
rect 4470 9764 4494 9766
rect 4254 9744 4550 9764
rect 4802 9752 4858 9761
rect 4802 9687 4858 9696
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3882 8256 3938 8265
rect 3882 8191 3938 8200
rect 2962 8120 3018 8129
rect 2962 8055 3018 8064
rect 3606 7984 3662 7993
rect 3606 7919 3608 7928
rect 3660 7919 3662 7928
rect 3608 7890 3660 7896
rect 3792 7880 3844 7886
rect 3790 7848 3792 7857
rect 3844 7848 3846 7857
rect 3790 7783 3846 7792
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 3608 7472 3660 7478
rect 3606 7440 3608 7449
rect 3660 7440 3662 7449
rect 4080 7410 4108 7686
rect 3606 7375 3662 7384
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3974 7304 4030 7313
rect 3974 7239 3976 7248
rect 4028 7239 4030 7248
rect 3976 7210 4028 7216
rect 4172 6662 4200 8978
rect 4264 8906 4292 9114
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4254 8732 4550 8752
rect 4310 8730 4334 8732
rect 4390 8730 4414 8732
rect 4470 8730 4494 8732
rect 4332 8678 4334 8730
rect 4396 8678 4408 8730
rect 4470 8678 4472 8730
rect 4310 8676 4334 8678
rect 4390 8676 4414 8678
rect 4470 8676 4494 8678
rect 4254 8656 4550 8676
rect 4632 8634 4660 8774
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4724 8498 4752 8774
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4816 8430 4844 9687
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5000 9042 5028 9522
rect 5092 9382 5120 9959
rect 5184 9926 5212 9998
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5184 9518 5212 9862
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5368 9178 5396 11591
rect 5448 11562 5500 11568
rect 5460 11354 5488 11562
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5552 11286 5580 12174
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5552 10266 5580 10610
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5736 10198 5764 10542
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 6000 10464 6052 10470
rect 6288 10441 6316 11698
rect 6000 10406 6052 10412
rect 6274 10432 6330 10441
rect 5828 10198 5856 10406
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5920 9382 5948 10066
rect 6012 9722 6040 10406
rect 6274 10367 6330 10376
rect 6288 10062 6316 10367
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6288 9586 6316 9998
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6276 9444 6328 9450
rect 6276 9386 6328 9392
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4908 8090 4936 8502
rect 5000 8430 5028 8978
rect 4988 8424 5040 8430
rect 5040 8372 5212 8378
rect 4988 8366 5212 8372
rect 5000 8350 5212 8366
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 5000 7954 5028 8230
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 4254 7644 4550 7664
rect 4310 7642 4334 7644
rect 4390 7642 4414 7644
rect 4470 7642 4494 7644
rect 4332 7590 4334 7642
rect 4396 7590 4408 7642
rect 4470 7590 4472 7642
rect 4310 7588 4334 7590
rect 4390 7588 4414 7590
rect 4470 7588 4494 7590
rect 4254 7568 4550 7588
rect 5092 7410 5120 7754
rect 5184 7410 5212 8350
rect 5368 7750 5396 9114
rect 5920 9110 5948 9318
rect 6012 9178 6040 9318
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 6012 8430 6040 9114
rect 6288 8634 6316 9386
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6380 8430 6408 12242
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6656 11778 6684 12038
rect 6828 11824 6880 11830
rect 6656 11750 6776 11778
rect 6932 11778 6960 12038
rect 6880 11772 6960 11778
rect 6828 11766 6960 11772
rect 6840 11750 6960 11766
rect 6748 11694 6776 11750
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6458 10840 6514 10849
rect 6458 10775 6514 10784
rect 6472 10674 6500 10775
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 5644 8078 5948 8106
rect 5644 8022 5672 8078
rect 5920 8022 5948 8078
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 4264 7002 4292 7346
rect 5172 7200 5224 7206
rect 5356 7200 5408 7206
rect 5224 7160 5356 7188
rect 5172 7142 5224 7148
rect 5356 7142 5408 7148
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 5736 6866 5764 7890
rect 6000 7880 6052 7886
rect 5920 7828 6000 7834
rect 5920 7822 6052 7828
rect 5920 7806 6040 7822
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 3606 6216 3662 6225
rect 3606 6151 3662 6160
rect 3620 5914 3648 6151
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 4172 5778 4200 6598
rect 4254 6556 4550 6576
rect 4310 6554 4334 6556
rect 4390 6554 4414 6556
rect 4470 6554 4494 6556
rect 4332 6502 4334 6554
rect 4396 6502 4408 6554
rect 4470 6502 4472 6554
rect 4310 6500 4334 6502
rect 4390 6500 4414 6502
rect 4470 6500 4494 6502
rect 4254 6480 4550 6500
rect 4632 6254 4660 6734
rect 5736 6458 5764 6802
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4264 5710 4292 6122
rect 4632 5914 4660 6190
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4632 5778 4660 5850
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4254 5468 4550 5488
rect 4310 5466 4334 5468
rect 4390 5466 4414 5468
rect 4470 5466 4494 5468
rect 4332 5414 4334 5466
rect 4396 5414 4408 5466
rect 4470 5414 4472 5466
rect 4310 5412 4334 5414
rect 4390 5412 4414 5414
rect 4470 5412 4494 5414
rect 4254 5392 4550 5412
rect 4632 5166 4660 5714
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4632 4690 4660 5102
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4254 4380 4550 4400
rect 4310 4378 4334 4380
rect 4390 4378 4414 4380
rect 4470 4378 4494 4380
rect 4332 4326 4334 4378
rect 4396 4326 4408 4378
rect 4470 4326 4472 4378
rect 4310 4324 4334 4326
rect 4390 4324 4414 4326
rect 4470 4324 4494 4326
rect 4254 4304 4550 4324
rect 4632 4264 4660 4626
rect 4448 4236 4660 4264
rect 4448 4078 4476 4236
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4448 3602 4476 4014
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4254 3292 4550 3312
rect 4310 3290 4334 3292
rect 4390 3290 4414 3292
rect 4470 3290 4494 3292
rect 4332 3238 4334 3290
rect 4396 3238 4408 3290
rect 4470 3238 4472 3290
rect 4310 3236 4334 3238
rect 4390 3236 4414 3238
rect 4470 3236 4494 3238
rect 4254 3216 4550 3236
rect 4710 3224 4766 3233
rect 4710 3159 4712 3168
rect 4764 3159 4766 3168
rect 4712 3130 4764 3136
rect 4816 2990 4844 3674
rect 5092 3058 5120 6190
rect 5920 6186 5948 7806
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 6254 6040 7686
rect 6472 7342 6500 8502
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6288 7002 6316 7210
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6472 6866 6500 7278
rect 6564 6882 6592 10678
rect 6656 10470 6684 11154
rect 7024 10656 7052 13398
rect 7300 13326 7328 14912
rect 7380 14894 7432 14900
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7116 11626 7144 12378
rect 7300 12374 7328 12582
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7208 11354 7236 11562
rect 7300 11558 7328 12310
rect 7392 12102 7420 13262
rect 7484 12782 7512 16068
rect 7840 16050 7892 16056
rect 8036 16046 8064 16526
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7553 15804 7849 15824
rect 7609 15802 7633 15804
rect 7689 15802 7713 15804
rect 7769 15802 7793 15804
rect 7631 15750 7633 15802
rect 7695 15750 7707 15802
rect 7769 15750 7771 15802
rect 7609 15748 7633 15750
rect 7689 15748 7713 15750
rect 7769 15748 7793 15750
rect 7553 15728 7849 15748
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7668 14958 7696 15302
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7944 14822 7972 15914
rect 8036 15366 8064 15982
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 8220 14958 8248 17054
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8312 15892 8340 16526
rect 8404 16046 8432 16730
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8680 15910 8708 16730
rect 8772 16250 8800 21520
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8864 18154 8892 19110
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 18426 9076 18566
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 8864 16794 8892 17682
rect 9048 17610 9076 18158
rect 9140 17882 9168 18906
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9324 18086 9352 18702
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8864 16114 8892 16730
rect 9140 16454 9168 17478
rect 9232 16561 9260 18022
rect 9324 17134 9352 18022
rect 9416 17814 9444 21520
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9508 19378 9536 19654
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9600 16590 9628 17682
rect 9692 17678 9720 19246
rect 9876 19174 9904 19450
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 9968 18986 9996 19110
rect 9876 18958 9996 18986
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9876 17066 9904 18958
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9968 17202 9996 18770
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 9588 16584 9640 16590
rect 9218 16552 9274 16561
rect 9588 16526 9640 16532
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9218 16487 9274 16496
rect 9128 16448 9180 16454
rect 9876 16436 9904 16526
rect 9128 16390 9180 16396
rect 9600 16408 9904 16436
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 9600 15910 9628 16408
rect 8392 15904 8444 15910
rect 8312 15864 8392 15892
rect 8392 15846 8444 15852
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7553 14716 7849 14736
rect 7609 14714 7633 14716
rect 7689 14714 7713 14716
rect 7769 14714 7793 14716
rect 7631 14662 7633 14714
rect 7695 14662 7707 14714
rect 7769 14662 7771 14714
rect 7609 14660 7633 14662
rect 7689 14660 7713 14662
rect 7769 14660 7793 14662
rect 7553 14640 7849 14660
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7852 14074 7880 14418
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7553 13628 7849 13648
rect 7609 13626 7633 13628
rect 7689 13626 7713 13628
rect 7769 13626 7793 13628
rect 7631 13574 7633 13626
rect 7695 13574 7707 13626
rect 7769 13574 7771 13626
rect 7609 13572 7633 13574
rect 7689 13572 7713 13574
rect 7769 13572 7793 13574
rect 7553 13552 7849 13572
rect 7944 13462 7972 14758
rect 8312 14482 8340 15438
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8404 13530 8432 14418
rect 8680 14278 8708 14826
rect 9324 14346 9352 15030
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 8680 13938 8708 14214
rect 9232 13938 9260 14214
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8680 13530 8708 13738
rect 9600 13734 9628 15846
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9692 15026 9720 15438
rect 9784 15162 9812 15506
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 8772 13326 8800 13670
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 8128 12986 8340 13002
rect 8116 12980 8340 12986
rect 8168 12974 8340 12980
rect 8116 12922 8168 12928
rect 8312 12850 8340 12974
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 8312 12646 8340 12786
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 7553 12540 7849 12560
rect 7609 12538 7633 12540
rect 7689 12538 7713 12540
rect 7769 12538 7793 12540
rect 7631 12486 7633 12538
rect 7695 12486 7707 12538
rect 7769 12486 7771 12538
rect 7609 12484 7633 12486
rect 7689 12484 7713 12486
rect 7769 12484 7793 12486
rect 7553 12464 7849 12484
rect 8312 12442 8340 12582
rect 9048 12442 9076 12650
rect 9600 12646 9628 13262
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7553 11452 7849 11472
rect 7609 11450 7633 11452
rect 7689 11450 7713 11452
rect 7769 11450 7793 11452
rect 7631 11398 7633 11450
rect 7695 11398 7707 11450
rect 7769 11398 7771 11450
rect 7609 11396 7633 11398
rect 7689 11396 7713 11398
rect 7769 11396 7793 11398
rect 7553 11376 7849 11396
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7116 10810 7144 11018
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6932 10628 7052 10656
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6932 10266 6960 10628
rect 7208 10606 7236 10950
rect 7196 10600 7248 10606
rect 7102 10568 7158 10577
rect 7012 10532 7064 10538
rect 7196 10542 7248 10548
rect 7102 10503 7158 10512
rect 7012 10474 7064 10480
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6656 7546 6684 7890
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6564 6866 6684 6882
rect 6460 6860 6512 6866
rect 6564 6860 6696 6866
rect 6564 6854 6644 6860
rect 6460 6802 6512 6808
rect 6644 6802 6696 6808
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5920 5914 5948 6122
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5914 6224 6054
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6274 5808 6330 5817
rect 5816 5772 5868 5778
rect 6274 5743 6330 5752
rect 6368 5772 6420 5778
rect 5816 5714 5868 5720
rect 5828 5370 5856 5714
rect 6288 5574 6316 5743
rect 6368 5714 6420 5720
rect 6380 5574 6408 5714
rect 6552 5704 6604 5710
rect 6550 5672 6552 5681
rect 6604 5672 6606 5681
rect 6550 5607 6606 5616
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5828 4282 5856 5034
rect 6012 4826 6040 5102
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 5908 4548 5960 4554
rect 5908 4490 5960 4496
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5920 4078 5948 4490
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 6104 3466 6132 4694
rect 6288 4078 6316 5306
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6380 4282 6408 4626
rect 6748 4604 6776 7686
rect 6840 6254 6868 9930
rect 7024 9722 7052 10474
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6932 9110 6960 9590
rect 7116 9489 7144 10503
rect 7102 9480 7158 9489
rect 7102 9415 7158 9424
rect 7102 9344 7158 9353
rect 7102 9279 7158 9288
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 8498 6960 8910
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7024 8129 7052 9046
rect 7116 8673 7144 9279
rect 7102 8664 7158 8673
rect 7102 8599 7158 8608
rect 7300 8265 7328 11086
rect 7668 10810 7696 11222
rect 7944 11014 7972 11630
rect 8128 11286 8156 12242
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8128 11150 8156 11222
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8036 10588 8064 10746
rect 8220 10606 8248 11494
rect 8312 11354 8340 11494
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8496 11150 8524 11698
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8312 10849 8340 11086
rect 8588 11082 8616 12242
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8298 10840 8354 10849
rect 8298 10775 8354 10784
rect 8312 10674 8340 10775
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 7944 10560 8064 10588
rect 8208 10600 8260 10606
rect 7380 10532 7432 10538
rect 7748 10532 7800 10538
rect 7380 10474 7432 10480
rect 7484 10492 7748 10520
rect 7392 10441 7420 10474
rect 7378 10432 7434 10441
rect 7378 10367 7434 10376
rect 7484 10266 7512 10492
rect 7748 10474 7800 10480
rect 7553 10364 7849 10384
rect 7609 10362 7633 10364
rect 7689 10362 7713 10364
rect 7769 10362 7793 10364
rect 7631 10310 7633 10362
rect 7695 10310 7707 10362
rect 7769 10310 7771 10362
rect 7609 10308 7633 10310
rect 7689 10308 7713 10310
rect 7769 10308 7793 10310
rect 7553 10288 7849 10308
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7392 9178 7420 10066
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7484 9654 7512 9998
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7668 9586 7696 9998
rect 7944 9994 7972 10560
rect 8208 10542 8260 10548
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 10266 8064 10406
rect 8312 10266 8340 10610
rect 8576 10600 8628 10606
rect 8404 10560 8576 10588
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8116 10124 8168 10130
rect 8300 10124 8352 10130
rect 8116 10066 8168 10072
rect 8220 10084 8300 10112
rect 7932 9988 7984 9994
rect 7932 9930 7984 9936
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9586 7880 9862
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 8128 9450 8156 10066
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8022 9344 8078 9353
rect 7553 9276 7849 9296
rect 8022 9279 8078 9288
rect 7609 9274 7633 9276
rect 7689 9274 7713 9276
rect 7769 9274 7793 9276
rect 7631 9222 7633 9274
rect 7695 9222 7707 9274
rect 7769 9222 7771 9274
rect 7609 9220 7633 9222
rect 7689 9220 7713 9222
rect 7769 9220 7793 9222
rect 7553 9200 7849 9220
rect 7930 9208 7986 9217
rect 7380 9172 7432 9178
rect 8036 9178 8064 9279
rect 8128 9178 8156 9386
rect 7930 9143 7986 9152
rect 8024 9172 8076 9178
rect 7380 9114 7432 9120
rect 7392 8362 7420 9114
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7852 8634 7880 8978
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7944 8401 7972 9143
rect 8024 9114 8076 9120
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8220 9110 8248 10084
rect 8300 10066 8352 10072
rect 8404 9926 8432 10560
rect 8576 10542 8628 10548
rect 8482 10296 8538 10305
rect 8482 10231 8538 10240
rect 8392 9920 8444 9926
rect 8496 9897 8524 10231
rect 8680 10062 8708 11018
rect 8758 10704 8814 10713
rect 8758 10639 8814 10648
rect 8772 10606 8800 10639
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8864 10538 8892 11154
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8392 9862 8444 9868
rect 8482 9888 8538 9897
rect 8404 9432 8432 9862
rect 8482 9823 8538 9832
rect 8864 9722 8892 10474
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8484 9444 8536 9450
rect 8404 9404 8484 9432
rect 8484 9386 8536 9392
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8220 8634 8248 9046
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8496 8498 8524 9386
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 7930 8392 7986 8401
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7472 8356 7524 8362
rect 7930 8327 7986 8336
rect 7472 8298 7524 8304
rect 7286 8256 7342 8265
rect 7286 8191 7342 8200
rect 7010 8120 7066 8129
rect 7010 8055 7066 8064
rect 7484 7886 7512 8298
rect 7553 8188 7849 8208
rect 7609 8186 7633 8188
rect 7689 8186 7713 8188
rect 7769 8186 7793 8188
rect 7631 8134 7633 8186
rect 7695 8134 7707 8186
rect 7769 8134 7771 8186
rect 7609 8132 7633 8134
rect 7689 8132 7713 8134
rect 7769 8132 7793 8134
rect 7553 8112 7849 8132
rect 8496 7970 8524 8434
rect 8220 7954 8524 7970
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8208 7948 8524 7954
rect 8260 7942 8524 7948
rect 8208 7890 8260 7896
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6932 5710 6960 6326
rect 7116 6186 7144 6734
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 7208 6118 7236 7686
rect 7852 7478 7880 7754
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7553 7100 7849 7120
rect 7609 7098 7633 7100
rect 7689 7098 7713 7100
rect 7769 7098 7793 7100
rect 7631 7046 7633 7098
rect 7695 7046 7707 7098
rect 7769 7046 7771 7098
rect 7609 7044 7633 7046
rect 7689 7044 7713 7046
rect 7769 7044 7793 7046
rect 7553 7024 7849 7044
rect 7654 6760 7710 6769
rect 7654 6695 7710 6704
rect 7668 6390 7696 6695
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6920 5704 6972 5710
rect 6972 5652 7052 5658
rect 6920 5646 7052 5652
rect 6840 5370 6868 5646
rect 6932 5630 7052 5646
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6932 5166 6960 5510
rect 7024 5234 7052 5630
rect 7208 5302 7236 6054
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7300 5370 7328 5782
rect 7392 5574 7420 6054
rect 7484 5914 7512 6258
rect 7553 6012 7849 6032
rect 7609 6010 7633 6012
rect 7689 6010 7713 6012
rect 7769 6010 7793 6012
rect 7631 5958 7633 6010
rect 7695 5958 7707 6010
rect 7769 5958 7771 6010
rect 7609 5956 7633 5958
rect 7689 5956 7713 5958
rect 7769 5956 7793 5958
rect 7553 5936 7849 5956
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7576 5166 7604 5714
rect 8036 5370 8064 7890
rect 8312 7546 8340 7942
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8298 7168 8354 7177
rect 8220 6934 8248 7142
rect 8298 7103 8354 7112
rect 8312 7002 8340 7103
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8312 6458 8340 6734
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8404 6118 8432 7686
rect 8772 7206 8800 9658
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8772 6934 8800 7142
rect 8576 6928 8628 6934
rect 8760 6928 8812 6934
rect 8628 6888 8708 6916
rect 8576 6870 8628 6876
rect 8680 6186 8708 6888
rect 8760 6870 8812 6876
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8128 5778 8156 6054
rect 8404 5778 8432 6054
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 8128 5030 8156 5578
rect 8680 5234 8708 6122
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 7484 4826 7512 4966
rect 7553 4924 7849 4944
rect 7609 4922 7633 4924
rect 7689 4922 7713 4924
rect 7769 4922 7793 4924
rect 7631 4870 7633 4922
rect 7695 4870 7707 4922
rect 7769 4870 7771 4922
rect 7609 4868 7633 4870
rect 7689 4868 7713 4870
rect 7769 4868 7793 4870
rect 7553 4848 7849 4868
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 6828 4616 6880 4622
rect 6748 4576 6828 4604
rect 6828 4558 6880 4564
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6736 4208 6788 4214
rect 6840 4162 6868 4558
rect 7208 4554 7236 4762
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7484 4214 7512 4558
rect 7668 4282 7696 4626
rect 7944 4282 7972 4966
rect 8864 4690 8892 7958
rect 9048 7478 9076 12378
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 11626 9168 12174
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9416 11150 9444 11562
rect 9600 11218 9628 12582
rect 9692 11665 9720 14826
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9784 14618 9812 14758
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 14074 9904 14214
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9784 12646 9812 13330
rect 9968 13274 9996 17002
rect 10060 13530 10088 21520
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10336 19009 10364 19110
rect 10322 19000 10378 19009
rect 10322 18935 10324 18944
rect 10376 18935 10378 18944
rect 10324 18906 10376 18912
rect 10336 18875 10364 18906
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10152 16250 10180 18702
rect 10244 18426 10272 18702
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10336 18306 10364 18770
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10244 18278 10364 18306
rect 10428 18290 10456 18634
rect 10416 18284 10468 18290
rect 10244 16998 10272 18278
rect 10416 18226 10468 18232
rect 10414 18048 10470 18057
rect 10414 17983 10470 17992
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10152 14958 10180 16186
rect 10244 16046 10272 16934
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 16046 10364 16390
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10152 13938 10180 14894
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10244 13462 10272 15506
rect 10336 15366 10364 15982
rect 10428 15570 10456 17983
rect 10520 16114 10548 19110
rect 10612 17066 10640 21520
rect 10852 19612 11148 19632
rect 10908 19610 10932 19612
rect 10988 19610 11012 19612
rect 11068 19610 11092 19612
rect 10930 19558 10932 19610
rect 10994 19558 11006 19610
rect 11068 19558 11070 19610
rect 10908 19556 10932 19558
rect 10988 19556 11012 19558
rect 11068 19556 11092 19558
rect 10852 19536 11148 19556
rect 11256 19530 11284 21520
rect 11256 19502 11376 19530
rect 10874 19408 10930 19417
rect 10874 19343 10930 19352
rect 11244 19372 11296 19378
rect 10888 18970 10916 19343
rect 11244 19314 11296 19320
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11072 18970 11100 19110
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10888 18850 10916 18906
rect 11164 18850 11192 19110
rect 10784 18828 10836 18834
rect 10888 18822 11192 18850
rect 10784 18770 10836 18776
rect 10796 18222 10824 18770
rect 10852 18524 11148 18544
rect 10908 18522 10932 18524
rect 10988 18522 11012 18524
rect 11068 18522 11092 18524
rect 10930 18470 10932 18522
rect 10994 18470 11006 18522
rect 11068 18470 11070 18522
rect 10908 18468 10932 18470
rect 10988 18468 11012 18470
rect 11068 18468 11092 18470
rect 10852 18448 11148 18468
rect 10874 18320 10930 18329
rect 10874 18255 10930 18264
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10796 17270 10824 18158
rect 10888 18154 10916 18255
rect 11256 18154 11284 19314
rect 11348 18834 11376 19502
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11532 18902 11560 19110
rect 11612 18964 11664 18970
rect 11612 18906 11664 18912
rect 11428 18896 11480 18902
rect 11428 18838 11480 18844
rect 11520 18896 11572 18902
rect 11520 18838 11572 18844
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11440 18426 11468 18838
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 11256 17882 11284 18090
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 10852 17436 11148 17456
rect 10908 17434 10932 17436
rect 10988 17434 11012 17436
rect 11068 17434 11092 17436
rect 10930 17382 10932 17434
rect 10994 17382 11006 17434
rect 11068 17382 11070 17434
rect 10908 17380 10932 17382
rect 10988 17380 11012 17382
rect 11068 17380 11092 17382
rect 10852 17360 11148 17380
rect 11256 17338 11284 17614
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 10784 17264 10836 17270
rect 10784 17206 10836 17212
rect 11242 17232 11298 17241
rect 11242 17167 11298 17176
rect 10600 17060 10652 17066
rect 10600 17002 10652 17008
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10704 15706 10732 16934
rect 10852 16348 11148 16368
rect 10908 16346 10932 16348
rect 10988 16346 11012 16348
rect 11068 16346 11092 16348
rect 10930 16294 10932 16346
rect 10994 16294 11006 16346
rect 11068 16294 11070 16346
rect 10908 16292 10932 16294
rect 10988 16292 11012 16294
rect 11068 16292 11092 16294
rect 10852 16272 11148 16292
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10336 13870 10364 15302
rect 10796 15094 10824 16050
rect 11256 15586 11284 17167
rect 11348 16522 11376 17750
rect 11428 17060 11480 17066
rect 11428 17002 11480 17008
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11440 16969 11468 17002
rect 11426 16960 11482 16969
rect 11426 16895 11482 16904
rect 11532 16726 11560 17002
rect 11624 16794 11652 18906
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11520 16720 11572 16726
rect 11520 16662 11572 16668
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 11348 15706 11376 16458
rect 11532 16454 11560 16662
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11428 15632 11480 15638
rect 11256 15558 11376 15586
rect 11428 15574 11480 15580
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 10852 15260 11148 15280
rect 10908 15258 10932 15260
rect 10988 15258 11012 15260
rect 11068 15258 11092 15260
rect 10930 15206 10932 15258
rect 10994 15206 11006 15258
rect 11068 15206 11070 15258
rect 10908 15204 10932 15206
rect 10988 15204 11012 15206
rect 11068 15204 11092 15206
rect 10852 15184 11148 15204
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 9876 13246 9996 13274
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9876 12594 9904 13246
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9968 12714 9996 13126
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9784 12458 9812 12582
rect 9876 12566 9996 12594
rect 9784 12430 9904 12458
rect 9678 11656 9734 11665
rect 9678 11591 9734 11600
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9692 11286 9720 11494
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9140 9897 9168 10066
rect 9232 9976 9260 11086
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 9994 9352 10950
rect 9586 10296 9642 10305
rect 9692 10282 9720 11086
rect 9784 10810 9812 11494
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9692 10254 9812 10282
rect 9586 10231 9642 10240
rect 9600 10198 9628 10231
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9312 9988 9364 9994
rect 9232 9948 9263 9976
rect 9126 9888 9182 9897
rect 9235 9874 9263 9948
rect 9312 9930 9364 9936
rect 9126 9823 9182 9832
rect 9232 9846 9263 9874
rect 9232 9654 9260 9846
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9324 8974 9352 9930
rect 9404 9444 9456 9450
rect 9508 9432 9536 9998
rect 9678 9888 9734 9897
rect 9678 9823 9734 9832
rect 9692 9450 9720 9823
rect 9456 9404 9536 9432
rect 9404 9386 9456 9392
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 9324 7410 9352 8910
rect 9508 8498 9536 9404
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9784 8922 9812 10254
rect 9876 9178 9904 12430
rect 9968 10130 9996 12566
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 10060 9110 10088 13126
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 10152 10033 10180 12310
rect 10244 12238 10272 13398
rect 10336 12986 10364 13806
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10336 12442 10364 12582
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10138 10024 10194 10033
rect 10138 9959 10194 9968
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9692 8894 9812 8922
rect 10048 8900 10100 8906
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9508 7886 9536 8434
rect 9692 8294 9720 8894
rect 10048 8842 10100 8848
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9784 8022 9812 8774
rect 9968 8430 9996 8774
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9876 7954 9904 8230
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9496 7880 9548 7886
rect 9416 7828 9496 7834
rect 9416 7822 9548 7828
rect 9416 7806 9536 7822
rect 9416 7410 9444 7806
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9508 7342 9536 7686
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9876 7206 9904 7890
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9862 7032 9918 7041
rect 9862 6967 9918 6976
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 9048 4690 9076 6870
rect 9876 6866 9904 6967
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9496 6656 9548 6662
rect 9968 6644 9996 8366
rect 10060 7954 10088 8842
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10152 8265 10180 8298
rect 10138 8256 10194 8265
rect 10138 8191 10194 8200
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 10060 7206 10088 7890
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 9496 6598 9548 6604
rect 9692 6616 9996 6644
rect 9508 6458 9536 6598
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9218 6216 9274 6225
rect 9140 5234 9168 6190
rect 9218 6151 9274 6160
rect 9232 6118 9260 6151
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 9140 4554 9168 5170
rect 9692 4842 9720 6616
rect 10060 5846 10088 6870
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10152 6254 10180 6802
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10140 6112 10192 6118
rect 10138 6080 10140 6089
rect 10192 6080 10194 6089
rect 10138 6015 10194 6024
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 9600 4814 9720 4842
rect 10060 4826 10088 5578
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 9772 4820 9824 4826
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9128 4548 9180 4554
rect 9128 4490 9180 4496
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 6788 4156 6868 4162
rect 6736 4150 6868 4156
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 6748 4134 6868 4150
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 6288 3058 6316 3538
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 6288 2922 6316 2994
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6380 2582 6408 3606
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6472 3194 6500 3538
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6472 2650 6500 3130
rect 6564 2990 6592 3334
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 6748 2514 6776 2926
rect 6840 2650 6868 4134
rect 8036 4078 8064 4422
rect 9140 4078 9168 4490
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6932 2514 6960 2926
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7024 2582 7052 2790
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7208 2310 7236 3878
rect 7553 3836 7849 3856
rect 7609 3834 7633 3836
rect 7689 3834 7713 3836
rect 7769 3834 7793 3836
rect 7631 3782 7633 3834
rect 7695 3782 7707 3834
rect 7769 3782 7771 3834
rect 7609 3780 7633 3782
rect 7689 3780 7713 3782
rect 7769 3780 7793 3782
rect 7553 3760 7849 3780
rect 8128 3602 8156 4014
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8128 2972 8156 3538
rect 8208 2984 8260 2990
rect 8128 2944 8208 2972
rect 8208 2926 8260 2932
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 7553 2748 7849 2768
rect 7609 2746 7633 2748
rect 7689 2746 7713 2748
rect 7769 2746 7793 2748
rect 7631 2694 7633 2746
rect 7695 2694 7707 2746
rect 7769 2694 7771 2746
rect 7609 2692 7633 2694
rect 7689 2692 7713 2694
rect 7769 2692 7793 2694
rect 7553 2672 7849 2692
rect 8312 2650 8340 2790
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 2378 8432 3878
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 9140 3233 9168 3402
rect 9324 3398 9352 3538
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9126 3224 9182 3233
rect 9036 3188 9088 3194
rect 9126 3159 9182 3168
rect 9036 3130 9088 3136
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 4254 2204 4550 2224
rect 4310 2202 4334 2204
rect 4390 2202 4414 2204
rect 4470 2202 4494 2204
rect 4332 2150 4334 2202
rect 4396 2150 4408 2202
rect 4470 2150 4472 2202
rect 4310 2148 4334 2150
rect 4390 2148 4414 2150
rect 4470 2148 4494 2150
rect 4254 2128 4550 2148
rect 1768 1284 1820 1290
rect 1768 1226 1820 1232
rect 1780 480 1808 1226
rect 5368 480 5396 2246
rect 9048 480 9076 3130
rect 9416 2990 9444 4082
rect 9508 3194 9536 4626
rect 9600 4622 9628 4814
rect 9772 4762 9824 4768
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9692 4282 9720 4694
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9600 1290 9628 3470
rect 9692 3194 9720 3606
rect 9784 3466 9812 4762
rect 10152 4622 10180 5510
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10244 4185 10272 10474
rect 10336 10198 10364 10746
rect 10324 10192 10376 10198
rect 10324 10134 10376 10140
rect 10428 9761 10456 14758
rect 10612 14550 10640 14962
rect 11256 14958 11284 15438
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10888 14482 10916 14758
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10852 14172 11148 14192
rect 10908 14170 10932 14172
rect 10988 14170 11012 14172
rect 11068 14170 11092 14172
rect 10930 14118 10932 14170
rect 10994 14118 11006 14170
rect 11068 14118 11070 14170
rect 10908 14116 10932 14118
rect 10988 14116 11012 14118
rect 11068 14116 11092 14118
rect 10852 14096 11148 14116
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10704 13394 10732 13806
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10520 11898 10548 12786
rect 10612 12306 10640 12922
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10612 12209 10640 12242
rect 10598 12200 10654 12209
rect 10598 12135 10654 12144
rect 10704 11898 10732 13330
rect 10980 13258 11008 13806
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10852 13084 11148 13104
rect 10908 13082 10932 13084
rect 10988 13082 11012 13084
rect 11068 13082 11092 13084
rect 10930 13030 10932 13082
rect 10994 13030 11006 13082
rect 11068 13030 11070 13082
rect 10908 13028 10932 13030
rect 10988 13028 11012 13030
rect 11068 13028 11092 13030
rect 10852 13008 11148 13028
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11256 12866 11284 12922
rect 11072 12838 11284 12866
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 12481 11008 12718
rect 11072 12714 11100 12838
rect 11348 12714 11376 15558
rect 11440 15026 11468 15574
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11716 14482 11744 14554
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11532 13462 11560 13670
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11152 12640 11204 12646
rect 11150 12608 11152 12617
rect 11204 12608 11206 12617
rect 11150 12543 11206 12552
rect 10966 12472 11022 12481
rect 10966 12407 11022 12416
rect 10966 12336 11022 12345
rect 10966 12271 10968 12280
rect 11020 12271 11022 12280
rect 10968 12242 11020 12248
rect 10852 11996 11148 12016
rect 10908 11994 10932 11996
rect 10988 11994 11012 11996
rect 11068 11994 11092 11996
rect 10930 11942 10932 11994
rect 10994 11942 11006 11994
rect 11068 11942 11070 11994
rect 10908 11940 10932 11942
rect 10988 11940 11012 11942
rect 11068 11940 11092 11942
rect 10852 11920 11148 11940
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10704 11762 10732 11834
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 11256 11694 11284 12650
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11348 11694 11376 12038
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11256 11354 11284 11630
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 10852 10908 11148 10928
rect 10908 10906 10932 10908
rect 10988 10906 11012 10908
rect 11068 10906 11092 10908
rect 10930 10854 10932 10906
rect 10994 10854 11006 10906
rect 11068 10854 11070 10906
rect 10908 10852 10932 10854
rect 10988 10852 11012 10854
rect 11068 10852 11092 10854
rect 10852 10832 11148 10852
rect 11348 10810 11376 11630
rect 11440 11626 11468 12582
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11532 11336 11560 13398
rect 11624 13308 11652 14010
rect 11716 13462 11744 14418
rect 11808 14278 11836 15506
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11624 13280 11744 13308
rect 11610 12608 11666 12617
rect 11610 12543 11666 12552
rect 11440 11308 11560 11336
rect 11440 11121 11468 11308
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11426 11112 11482 11121
rect 11426 11047 11482 11056
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 10782 10704 10838 10713
rect 10782 10639 10838 10648
rect 10414 9752 10470 9761
rect 10414 9687 10470 9696
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10428 8362 10456 8910
rect 10520 8634 10548 8978
rect 10704 8974 10732 9454
rect 10796 9382 10824 10639
rect 11440 10266 11468 10950
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11532 9994 11560 11154
rect 11624 11014 11652 12543
rect 11716 12238 11744 13280
rect 11900 12986 11928 21520
rect 12254 19408 12310 19417
rect 12072 19372 12124 19378
rect 12254 19343 12256 19352
rect 12072 19314 12124 19320
rect 12308 19343 12310 19352
rect 12256 19314 12308 19320
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 11992 19145 12020 19246
rect 11978 19136 12034 19145
rect 11978 19071 12034 19080
rect 12084 18630 12112 19314
rect 12452 19310 12480 21520
rect 12544 19366 12848 19394
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12544 19174 12572 19366
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12820 19258 12848 19366
rect 12256 19168 12308 19174
rect 12532 19168 12584 19174
rect 12308 19128 12480 19156
rect 12256 19110 12308 19116
rect 12254 18728 12310 18737
rect 12254 18663 12310 18672
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12084 17814 12112 18566
rect 12176 18057 12204 18566
rect 12162 18048 12218 18057
rect 12162 17983 12218 17992
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 12268 17241 12296 18663
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12360 17814 12388 18362
rect 12452 17882 12480 19128
rect 12532 19110 12584 19116
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12544 18222 12572 18770
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12348 17808 12400 17814
rect 12348 17750 12400 17756
rect 12544 17338 12572 18158
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12254 17232 12310 17241
rect 12254 17167 12310 17176
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 11992 16794 12020 16934
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12084 16250 12112 16526
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 12268 15706 12296 16934
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12360 14890 12388 16934
rect 12544 16658 12572 17274
rect 12636 16658 12664 19110
rect 12728 18834 12756 19246
rect 12820 19230 12940 19258
rect 12806 19136 12862 19145
rect 12806 19071 12862 19080
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12728 16969 12756 17546
rect 12714 16960 12770 16969
rect 12714 16895 12770 16904
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12544 15978 12572 16594
rect 12622 16144 12678 16153
rect 12622 16079 12624 16088
rect 12676 16079 12678 16088
rect 12624 16050 12676 16056
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12440 15632 12492 15638
rect 12728 15586 12756 15914
rect 12492 15580 12756 15586
rect 12440 15574 12756 15580
rect 12452 15558 12756 15574
rect 12452 15162 12480 15558
rect 12820 15366 12848 19071
rect 12912 18086 12940 19230
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 13004 18970 13032 19178
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13004 17066 13032 17614
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16794 12940 16934
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 13096 16250 13124 21520
rect 13266 19000 13322 19009
rect 13266 18935 13322 18944
rect 13280 18630 13308 18935
rect 13636 18760 13688 18766
rect 13464 18720 13636 18748
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13266 18456 13322 18465
rect 13266 18391 13322 18400
rect 13280 17338 13308 18391
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13188 16969 13216 17138
rect 13174 16960 13230 16969
rect 13174 16895 13230 16904
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 13004 15502 13032 15914
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 13004 15026 13032 15438
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 12084 14618 12112 14758
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12084 13530 12112 14418
rect 12636 14074 12664 14894
rect 13464 14074 13492 18720
rect 13636 18702 13688 18708
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 16794 13584 18022
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13648 17134 13676 17614
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13740 15638 13768 21520
rect 14292 19938 14320 21520
rect 14292 19910 14596 19938
rect 13910 19408 13966 19417
rect 13910 19343 13966 19352
rect 13924 19174 13952 19343
rect 14188 19304 14240 19310
rect 14186 19272 14188 19281
rect 14240 19272 14242 19281
rect 14186 19207 14242 19216
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13832 18698 13860 18906
rect 14016 18850 14044 19110
rect 14150 19068 14446 19088
rect 14206 19066 14230 19068
rect 14286 19066 14310 19068
rect 14366 19066 14390 19068
rect 14228 19014 14230 19066
rect 14292 19014 14304 19066
rect 14366 19014 14368 19066
rect 14206 19012 14230 19014
rect 14286 19012 14310 19014
rect 14366 19012 14390 19014
rect 14150 18992 14446 19012
rect 14016 18822 14136 18850
rect 13820 18692 13872 18698
rect 13820 18634 13872 18640
rect 14108 18290 14136 18822
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14292 18601 14320 18770
rect 14278 18592 14334 18601
rect 14278 18527 14334 18536
rect 14384 18465 14412 18770
rect 14370 18456 14426 18465
rect 14280 18420 14332 18426
rect 14370 18391 14426 18400
rect 14280 18362 14332 18368
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13832 17202 13860 18022
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13832 16726 13860 17138
rect 13924 17134 13952 18022
rect 14016 17882 14044 18158
rect 14292 18154 14320 18362
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 14150 17980 14446 18000
rect 14206 17978 14230 17980
rect 14286 17978 14310 17980
rect 14366 17978 14390 17980
rect 14228 17926 14230 17978
rect 14292 17926 14304 17978
rect 14366 17926 14368 17978
rect 14206 17924 14230 17926
rect 14286 17924 14310 17926
rect 14366 17924 14390 17926
rect 14150 17904 14446 17924
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 14096 17808 14148 17814
rect 14096 17750 14148 17756
rect 14476 17762 14504 19110
rect 14568 18850 14596 19910
rect 14936 19530 14964 21520
rect 15934 20360 15990 20369
rect 15934 20295 15990 20304
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 14844 19502 14964 19530
rect 15200 19508 15252 19514
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14660 18970 14688 19110
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14568 18834 14780 18850
rect 14568 18828 14792 18834
rect 14568 18822 14740 18828
rect 14740 18770 14792 18776
rect 14738 18320 14794 18329
rect 14738 18255 14794 18264
rect 14752 18222 14780 18255
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14844 17814 14872 19502
rect 15200 19450 15252 19456
rect 14924 19372 14976 19378
rect 14976 19332 15056 19360
rect 14924 19314 14976 19320
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14832 17808 14884 17814
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 14108 17066 14136 17750
rect 14476 17734 14688 17762
rect 14832 17750 14884 17756
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14096 17060 14148 17066
rect 14096 17002 14148 17008
rect 14464 17060 14516 17066
rect 14464 17002 14516 17008
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13832 15570 13860 16526
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 13924 16046 13952 16458
rect 14016 16402 14044 16934
rect 14150 16892 14446 16912
rect 14206 16890 14230 16892
rect 14286 16890 14310 16892
rect 14366 16890 14390 16892
rect 14228 16838 14230 16890
rect 14292 16838 14304 16890
rect 14366 16838 14368 16890
rect 14206 16836 14230 16838
rect 14286 16836 14310 16838
rect 14366 16836 14390 16838
rect 14150 16816 14446 16836
rect 14476 16726 14504 17002
rect 14568 16794 14596 17614
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14464 16720 14516 16726
rect 14464 16662 14516 16668
rect 14016 16374 14136 16402
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 14016 14958 14044 16186
rect 14108 15978 14136 16374
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 14150 15804 14446 15824
rect 14206 15802 14230 15804
rect 14286 15802 14310 15804
rect 14366 15802 14390 15804
rect 14228 15750 14230 15802
rect 14292 15750 14304 15802
rect 14366 15750 14368 15802
rect 14206 15748 14230 15750
rect 14286 15748 14310 15750
rect 14366 15748 14390 15750
rect 14150 15728 14446 15748
rect 14476 15706 14504 16662
rect 14554 16416 14610 16425
rect 14554 16351 14610 16360
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 14568 14906 14596 16351
rect 14660 15978 14688 17734
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14752 16794 14780 17682
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14844 16658 14872 17478
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14830 16552 14886 16561
rect 14936 16522 14964 18702
rect 14830 16487 14886 16496
rect 14924 16516 14976 16522
rect 14738 16008 14794 16017
rect 14648 15972 14700 15978
rect 14738 15943 14794 15952
rect 14648 15914 14700 15920
rect 14752 15706 14780 15943
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14844 15026 14872 16487
rect 14924 16458 14976 16464
rect 14924 16244 14976 16250
rect 15028 16232 15056 19332
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 14976 16204 15056 16232
rect 14924 16186 14976 16192
rect 14924 15972 14976 15978
rect 14924 15914 14976 15920
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14568 14878 14688 14906
rect 14936 14890 14964 15914
rect 15016 15632 15068 15638
rect 15016 15574 15068 15580
rect 15028 14958 15056 15574
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 13556 14414 13584 14758
rect 14150 14716 14446 14736
rect 14206 14714 14230 14716
rect 14286 14714 14310 14716
rect 14366 14714 14390 14716
rect 14228 14662 14230 14714
rect 14292 14662 14304 14714
rect 14366 14662 14368 14714
rect 14206 14660 14230 14662
rect 14286 14660 14310 14662
rect 14366 14660 14390 14662
rect 14150 14640 14446 14660
rect 14568 14482 14596 14758
rect 14556 14476 14608 14482
rect 14660 14464 14688 14878
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14660 14436 14780 14464
rect 14556 14418 14608 14424
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 12084 12850 12112 13466
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11704 12232 11756 12238
rect 12360 12220 12388 13806
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12452 12782 12480 13670
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12440 12232 12492 12238
rect 12360 12200 12440 12220
rect 12492 12200 12494 12209
rect 12360 12192 12438 12200
rect 11704 12174 11756 12180
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11716 10169 11744 12174
rect 12438 12135 12494 12144
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 11980 11552 12032 11558
rect 12164 11552 12216 11558
rect 11980 11494 12032 11500
rect 12084 11512 12164 11540
rect 11992 11286 12020 11494
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11702 10160 11758 10169
rect 11808 10130 11836 10746
rect 11702 10095 11758 10104
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 10852 9820 11148 9840
rect 10908 9818 10932 9820
rect 10988 9818 11012 9820
rect 11068 9818 11092 9820
rect 10930 9766 10932 9818
rect 10994 9766 11006 9818
rect 11068 9766 11070 9818
rect 10908 9764 10932 9766
rect 10988 9764 11012 9766
rect 11068 9764 11092 9766
rect 10852 9744 11148 9764
rect 11440 9722 11468 9862
rect 11794 9752 11850 9761
rect 11428 9716 11480 9722
rect 11794 9687 11850 9696
rect 11428 9658 11480 9664
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 8974 10916 9318
rect 11348 9042 11376 9454
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 8090 10456 8298
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10704 7342 10732 8910
rect 10852 8732 11148 8752
rect 10908 8730 10932 8732
rect 10988 8730 11012 8732
rect 11068 8730 11092 8732
rect 10930 8678 10932 8730
rect 10994 8678 11006 8730
rect 11068 8678 11070 8730
rect 10908 8676 10932 8678
rect 10988 8676 11012 8678
rect 11068 8676 11092 8678
rect 10852 8656 11148 8676
rect 11440 8566 11468 9658
rect 11808 9382 11836 9687
rect 11900 9654 11928 11086
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11992 9432 12020 10095
rect 11900 9404 12020 9432
rect 11796 9376 11848 9382
rect 11702 9344 11758 9353
rect 11796 9318 11848 9324
rect 11702 9279 11758 9288
rect 11716 8673 11744 9279
rect 11702 8664 11758 8673
rect 11702 8599 11758 8608
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 10852 7644 11148 7664
rect 10908 7642 10932 7644
rect 10988 7642 11012 7644
rect 11068 7642 11092 7644
rect 10930 7590 10932 7642
rect 10994 7590 11006 7642
rect 11068 7590 11070 7642
rect 10908 7588 10932 7590
rect 10988 7588 11012 7590
rect 11068 7588 11092 7590
rect 10852 7568 11148 7588
rect 11256 7546 11284 7822
rect 11334 7576 11390 7585
rect 11244 7540 11296 7546
rect 11334 7511 11390 7520
rect 11244 7482 11296 7488
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10428 6848 10456 7278
rect 11348 7177 11376 7511
rect 11428 7268 11480 7274
rect 11428 7210 11480 7216
rect 11334 7168 11390 7177
rect 11334 7103 11390 7112
rect 11440 7002 11468 7210
rect 11794 7032 11850 7041
rect 11428 6996 11480 7002
rect 11794 6967 11850 6976
rect 11428 6938 11480 6944
rect 11244 6928 11296 6934
rect 11244 6870 11296 6876
rect 10600 6860 10652 6866
rect 10428 6820 10600 6848
rect 10336 5710 10364 6802
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10336 5370 10364 5646
rect 10428 5574 10456 6820
rect 10600 6802 10652 6808
rect 10852 6556 11148 6576
rect 10908 6554 10932 6556
rect 10988 6554 11012 6556
rect 11068 6554 11092 6556
rect 10930 6502 10932 6554
rect 10994 6502 11006 6554
rect 11068 6502 11070 6554
rect 10908 6500 10932 6502
rect 10988 6500 11012 6502
rect 11068 6500 11092 6502
rect 10852 6480 11148 6500
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5953 10548 6054
rect 10506 5944 10562 5953
rect 10506 5879 10562 5888
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10520 5166 10548 5879
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10230 4176 10286 4185
rect 10230 4111 10286 4120
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9876 2514 9904 4014
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10336 2514 10364 3470
rect 10612 2904 10640 6190
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10888 5914 10916 6122
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10980 5778 11008 5850
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10796 5234 10824 5714
rect 11256 5710 11284 6870
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11716 6390 11744 6598
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11808 6254 11836 6967
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11624 5710 11652 6122
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11428 5704 11480 5710
rect 11612 5704 11664 5710
rect 11428 5646 11480 5652
rect 11532 5664 11612 5692
rect 10852 5468 11148 5488
rect 10908 5466 10932 5468
rect 10988 5466 11012 5468
rect 11068 5466 11092 5468
rect 10930 5414 10932 5466
rect 10994 5414 11006 5466
rect 11068 5414 11070 5466
rect 10908 5412 10932 5414
rect 10988 5412 11012 5414
rect 11068 5412 11092 5414
rect 10852 5392 11148 5412
rect 11256 5302 11284 5646
rect 11336 5568 11388 5574
rect 11440 5545 11468 5646
rect 11336 5510 11388 5516
rect 11426 5536 11482 5545
rect 11348 5370 11376 5510
rect 11426 5471 11482 5480
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 11256 4486 11284 5238
rect 11532 5098 11560 5664
rect 11612 5646 11664 5652
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11428 5024 11480 5030
rect 11612 5024 11664 5030
rect 11428 4966 11480 4972
rect 11532 4972 11612 4978
rect 11532 4966 11664 4972
rect 11440 4826 11468 4966
rect 11532 4950 11652 4966
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11348 4706 11376 4762
rect 11348 4678 11468 4706
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 10852 4380 11148 4400
rect 10908 4378 10932 4380
rect 10988 4378 11012 4380
rect 11068 4378 11092 4380
rect 10930 4326 10932 4378
rect 10994 4326 11006 4378
rect 11068 4326 11070 4378
rect 10908 4324 10932 4326
rect 10988 4324 11012 4326
rect 11068 4324 11092 4326
rect 10852 4304 11148 4324
rect 10876 4208 10928 4214
rect 10704 4168 10876 4196
rect 10704 3534 10732 4168
rect 10876 4150 10928 4156
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11072 4010 11100 4082
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10782 3632 10838 3641
rect 10782 3567 10838 3576
rect 10796 3534 10824 3567
rect 11348 3534 11376 4490
rect 11440 4486 11468 4678
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11532 3534 11560 4950
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 11152 3528 11204 3534
rect 11336 3528 11388 3534
rect 11204 3505 11284 3516
rect 11204 3496 11298 3505
rect 11204 3488 11242 3496
rect 11152 3470 11204 3476
rect 11336 3470 11388 3476
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11242 3431 11298 3440
rect 10852 3292 11148 3312
rect 10908 3290 10932 3292
rect 10988 3290 11012 3292
rect 11068 3290 11092 3292
rect 10930 3238 10932 3290
rect 10994 3238 11006 3290
rect 11068 3238 11070 3290
rect 10908 3236 10932 3238
rect 10988 3236 11012 3238
rect 11068 3236 11092 3238
rect 10852 3216 11148 3236
rect 11256 3194 11284 3431
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11716 3126 11744 5170
rect 11808 4486 11836 5646
rect 11900 5545 11928 9404
rect 11978 9344 12034 9353
rect 11978 9279 12034 9288
rect 11992 8566 12020 9279
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11992 8090 12020 8366
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11886 5536 11942 5545
rect 11886 5471 11942 5480
rect 12084 5030 12112 11512
rect 12164 11494 12216 11500
rect 12268 11082 12296 11698
rect 12544 11626 12572 13126
rect 12636 12345 12664 13670
rect 13556 13394 13584 14350
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 13924 13870 13952 14010
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13832 13530 13860 13806
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12622 12336 12678 12345
rect 12622 12271 12624 12280
rect 12676 12271 12678 12280
rect 12624 12242 12676 12248
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12176 10266 12204 10678
rect 12268 10674 12296 11018
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12162 10024 12218 10033
rect 12162 9959 12218 9968
rect 12176 9654 12204 9959
rect 12268 9874 12296 10406
rect 12360 10130 12388 10950
rect 12452 10554 12480 11154
rect 12532 10600 12584 10606
rect 12452 10548 12532 10554
rect 12452 10542 12584 10548
rect 12452 10526 12572 10542
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12268 9846 12388 9874
rect 12360 9722 12388 9846
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12176 9382 12204 9454
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 9058 12296 9318
rect 12452 9178 12480 10526
rect 12636 10441 12664 12242
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12622 10432 12678 10441
rect 12622 10367 12678 10376
rect 12728 10248 12756 12174
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12806 11248 12862 11257
rect 12806 11183 12862 11192
rect 12820 11150 12848 11183
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12636 10220 12756 10248
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12544 9353 12572 9930
rect 12636 9897 12664 10220
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12622 9888 12678 9897
rect 12622 9823 12678 9832
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12530 9344 12586 9353
rect 12530 9279 12586 9288
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12636 9110 12664 9454
rect 12176 9030 12296 9058
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12176 8809 12204 9030
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12360 8945 12572 8956
rect 12360 8936 12586 8945
rect 12360 8928 12530 8936
rect 12162 8800 12218 8809
rect 12162 8735 12218 8744
rect 12162 8392 12218 8401
rect 12162 8327 12218 8336
rect 12176 6905 12204 8327
rect 12268 7886 12296 8910
rect 12360 8838 12388 8928
rect 12530 8871 12586 8880
rect 12348 8832 12400 8838
rect 12532 8832 12584 8838
rect 12348 8774 12400 8780
rect 12452 8780 12532 8786
rect 12452 8774 12584 8780
rect 12452 8758 12572 8774
rect 12452 8362 12480 8758
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12348 8288 12400 8294
rect 12348 8230 12400 8236
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7342 12296 7822
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12162 6896 12218 6905
rect 12162 6831 12218 6840
rect 12254 5944 12310 5953
rect 12254 5879 12310 5888
rect 12164 5296 12216 5302
rect 12164 5238 12216 5244
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11900 4162 11928 4558
rect 11808 4146 11928 4162
rect 11796 4140 11928 4146
rect 11848 4134 11928 4140
rect 11796 4082 11848 4088
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11518 2952 11574 2961
rect 10692 2916 10744 2922
rect 10612 2876 10692 2904
rect 11518 2887 11574 2896
rect 10692 2858 10744 2864
rect 11532 2854 11560 2887
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11716 2582 11744 3062
rect 11900 2650 11928 4134
rect 11992 3058 12020 4626
rect 12084 4078 12112 4626
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12084 2990 12112 4014
rect 12176 3641 12204 5238
rect 12268 5234 12296 5879
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12360 4146 12388 8230
rect 12636 6662 12664 8570
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12544 6361 12572 6394
rect 12530 6352 12586 6361
rect 12530 6287 12586 6296
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12162 3632 12218 3641
rect 12162 3567 12164 3576
rect 12216 3567 12218 3576
rect 12164 3538 12216 3544
rect 12176 3507 12204 3538
rect 12268 3398 12296 3674
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12360 3097 12388 3606
rect 12452 3194 12480 4558
rect 12544 4264 12572 5034
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12636 4729 12664 4762
rect 12622 4720 12678 4729
rect 12622 4655 12678 4664
rect 12624 4276 12676 4282
rect 12544 4236 12624 4264
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12346 3088 12402 3097
rect 12346 3023 12402 3032
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 12544 2514 12572 4236
rect 12624 4218 12676 4224
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12636 3097 12664 3130
rect 12622 3088 12678 3097
rect 12622 3023 12678 3032
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 10852 2204 11148 2224
rect 10908 2202 10932 2204
rect 10988 2202 11012 2204
rect 11068 2202 11092 2204
rect 10930 2150 10932 2202
rect 10994 2150 11006 2202
rect 11068 2150 11070 2202
rect 10908 2148 10932 2150
rect 10988 2148 11012 2150
rect 11068 2148 11092 2150
rect 10852 2128 11148 2148
rect 9588 1284 9640 1290
rect 9588 1226 9640 1232
rect 11716 921 11744 2246
rect 11702 912 11758 921
rect 11702 847 11758 856
rect 12728 480 12756 10066
rect 12820 10062 12848 11086
rect 12912 10577 12940 12038
rect 12898 10568 12954 10577
rect 12898 10503 12954 10512
rect 13004 10198 13032 13126
rect 13556 12986 13584 13330
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13924 12730 13952 13806
rect 14384 13784 14412 14010
rect 14384 13756 14504 13784
rect 14150 13628 14446 13648
rect 14206 13626 14230 13628
rect 14286 13626 14310 13628
rect 14366 13626 14390 13628
rect 14228 13574 14230 13626
rect 14292 13574 14304 13626
rect 14366 13574 14368 13626
rect 14206 13572 14230 13574
rect 14286 13572 14310 13574
rect 14366 13572 14390 13574
rect 14150 13552 14446 13572
rect 13740 12702 13952 12730
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 12808 9512 12860 9518
rect 12860 9472 12940 9500
rect 12808 9454 12860 9460
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 8634 12848 9318
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12912 8566 12940 9472
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12820 7546 12848 8298
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12820 7274 12848 7482
rect 12912 7274 12940 8230
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12806 5808 12862 5817
rect 12806 5743 12808 5752
rect 12860 5743 12862 5752
rect 12808 5714 12860 5720
rect 12912 5574 12940 6326
rect 13004 6254 13032 9862
rect 13096 9625 13124 12582
rect 13542 12472 13598 12481
rect 13268 12436 13320 12442
rect 13740 12442 13768 12702
rect 13542 12407 13598 12416
rect 13728 12436 13780 12442
rect 13268 12378 13320 12384
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13188 12102 13216 12242
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13188 9994 13216 10746
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 13082 9616 13138 9625
rect 13082 9551 13138 9560
rect 13280 9518 13308 12378
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 13372 9586 13400 10134
rect 13556 9926 13584 12407
rect 13728 12378 13780 12384
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11354 13768 11494
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13648 10690 13676 11290
rect 13832 11218 13860 11562
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13924 11286 13952 11494
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13832 10810 13860 11154
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13648 10662 13860 10690
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13544 9920 13596 9926
rect 13464 9880 13544 9908
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13188 9178 13216 9454
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13096 6458 13124 8978
rect 13372 8498 13400 9522
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13372 8090 13400 8434
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13464 7698 13492 9880
rect 13544 9862 13596 9868
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13556 7954 13584 9454
rect 13648 8566 13676 9998
rect 13832 8634 13860 10662
rect 14016 10130 14044 12718
rect 14150 12540 14446 12560
rect 14206 12538 14230 12540
rect 14286 12538 14310 12540
rect 14366 12538 14390 12540
rect 14228 12486 14230 12538
rect 14292 12486 14304 12538
rect 14366 12486 14368 12538
rect 14206 12484 14230 12486
rect 14286 12484 14310 12486
rect 14366 12484 14390 12486
rect 14150 12464 14446 12484
rect 14094 11928 14150 11937
rect 14094 11863 14096 11872
rect 14148 11863 14150 11872
rect 14096 11834 14148 11840
rect 14476 11558 14504 13756
rect 14568 11762 14596 14418
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14660 13394 14688 14282
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14752 13258 14780 14436
rect 14844 13938 14872 14758
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14646 12744 14702 12753
rect 14752 12714 14780 13194
rect 14646 12679 14702 12688
rect 14740 12708 14792 12714
rect 14660 12238 14688 12679
rect 14740 12650 14792 12656
rect 14738 12608 14794 12617
rect 14738 12543 14794 12552
rect 14752 12306 14780 12543
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14844 11694 14872 13874
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14150 11452 14446 11472
rect 14206 11450 14230 11452
rect 14286 11450 14310 11452
rect 14366 11450 14390 11452
rect 14228 11398 14230 11450
rect 14292 11398 14304 11450
rect 14366 11398 14368 11450
rect 14206 11396 14230 11398
rect 14286 11396 14310 11398
rect 14366 11396 14390 11398
rect 14150 11376 14446 11396
rect 14476 11354 14504 11494
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14660 11218 14688 11562
rect 14936 11506 14964 12854
rect 14752 11478 14964 11506
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14150 10364 14446 10384
rect 14206 10362 14230 10364
rect 14286 10362 14310 10364
rect 14366 10362 14390 10364
rect 14228 10310 14230 10362
rect 14292 10310 14304 10362
rect 14366 10310 14368 10362
rect 14206 10308 14230 10310
rect 14286 10308 14310 10310
rect 14366 10308 14390 10310
rect 14150 10288 14446 10308
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14476 9518 14504 11018
rect 14646 10704 14702 10713
rect 14752 10656 14780 11478
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14702 10648 14780 10656
rect 14646 10639 14780 10648
rect 14660 10628 14780 10639
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14150 9276 14446 9296
rect 14206 9274 14230 9276
rect 14286 9274 14310 9276
rect 14366 9274 14390 9276
rect 14228 9222 14230 9274
rect 14292 9222 14304 9274
rect 14366 9222 14368 9274
rect 14206 9220 14230 9222
rect 14286 9220 14310 9222
rect 14366 9220 14390 9222
rect 14150 9200 14446 9220
rect 14372 8832 14424 8838
rect 14186 8800 14242 8809
rect 14186 8735 14242 8744
rect 14370 8800 14372 8809
rect 14424 8800 14426 8809
rect 14370 8735 14426 8744
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 14200 8566 14228 8735
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 13636 8288 13688 8294
rect 13634 8256 13636 8265
rect 13728 8288 13780 8294
rect 13688 8256 13690 8265
rect 13728 8230 13780 8236
rect 13634 8191 13690 8200
rect 13648 8090 13676 8191
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13740 8022 13768 8230
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13464 7670 13584 7698
rect 13556 6866 13584 7670
rect 13740 7546 13768 7958
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13820 7404 13872 7410
rect 13740 7364 13820 7392
rect 13740 7002 13768 7364
rect 13820 7346 13872 7352
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13268 6724 13320 6730
rect 13544 6724 13596 6730
rect 13268 6666 13320 6672
rect 13464 6684 13544 6712
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13004 5817 13032 6054
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 12990 5808 13046 5817
rect 12990 5743 13046 5752
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12820 4758 12848 4966
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 13004 4690 13032 5646
rect 13096 5370 13124 5850
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13188 5234 13216 6054
rect 13280 5914 13308 6666
rect 13360 6248 13412 6254
rect 13464 6236 13492 6684
rect 13544 6666 13596 6672
rect 13832 6474 13860 7210
rect 13924 6662 13952 8502
rect 14476 8294 14504 8570
rect 14568 8430 14596 9386
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14464 8288 14516 8294
rect 14660 8242 14688 10628
rect 14844 9761 14872 11290
rect 14922 11112 14978 11121
rect 15028 11098 15056 13330
rect 14978 11070 15056 11098
rect 14922 11047 14978 11056
rect 14936 11014 14964 11047
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 15120 10826 15148 19246
rect 15212 18222 15240 19450
rect 15290 18456 15346 18465
rect 15290 18391 15346 18400
rect 15304 18358 15332 18391
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15200 18216 15252 18222
rect 15200 18158 15252 18164
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15212 14346 15240 17138
rect 15304 15570 15332 17206
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15396 15450 15424 19654
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15580 18850 15608 19246
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15856 18970 15884 19178
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15580 18822 15700 18850
rect 15672 18766 15700 18822
rect 15660 18760 15712 18766
rect 15712 18708 15884 18714
rect 15660 18702 15884 18708
rect 15672 18686 15884 18702
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15488 17134 15516 17818
rect 15476 17128 15528 17134
rect 15672 17082 15700 18566
rect 15764 18222 15792 18566
rect 15856 18358 15884 18686
rect 15844 18352 15896 18358
rect 15844 18294 15896 18300
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15856 17762 15884 18294
rect 15948 17882 15976 20295
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 16040 18222 16068 19654
rect 16132 19394 16160 21520
rect 16132 19366 16252 19394
rect 16224 19310 16252 19366
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16132 18902 16160 19110
rect 16120 18896 16172 18902
rect 16120 18838 16172 18844
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15856 17734 15976 17762
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15476 17070 15528 17076
rect 15488 16998 15516 17070
rect 15580 17054 15700 17082
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15488 16425 15516 16730
rect 15474 16416 15530 16425
rect 15474 16351 15530 16360
rect 15580 15978 15608 17054
rect 15660 16992 15712 16998
rect 15712 16952 15792 16980
rect 15660 16934 15712 16940
rect 15764 16658 15792 16952
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15672 16250 15700 16594
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 15706 15516 15846
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15488 15502 15516 15642
rect 15672 15638 15700 16186
rect 15764 16046 15792 16594
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15750 15872 15806 15881
rect 15750 15807 15806 15816
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 15304 15422 15424 15450
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15304 15162 15332 15422
rect 15488 15314 15516 15438
rect 15488 15286 15608 15314
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15304 13938 15332 14894
rect 15580 14482 15608 15286
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15304 12782 15332 13874
rect 15566 13696 15622 13705
rect 15566 13631 15622 13640
rect 15580 13410 15608 13631
rect 15488 13382 15608 13410
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15212 12374 15240 12650
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15304 12238 15332 12718
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15212 11354 15240 12038
rect 15304 11626 15332 12174
rect 15396 11801 15424 12242
rect 15382 11792 15438 11801
rect 15382 11727 15438 11736
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15304 11150 15332 11562
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 14936 10798 15148 10826
rect 15304 10810 15332 11086
rect 15292 10804 15344 10810
rect 14830 9752 14886 9761
rect 14830 9687 14886 9696
rect 14844 9217 14872 9687
rect 14830 9208 14886 9217
rect 14830 9143 14886 9152
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14752 8634 14780 8978
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14936 8514 14964 10798
rect 15292 10746 15344 10752
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15120 9926 15148 10542
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15304 10198 15332 10406
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15396 10062 15424 10542
rect 15488 10130 15516 13382
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15580 12209 15608 13262
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15672 13025 15700 13126
rect 15658 13016 15714 13025
rect 15658 12951 15714 12960
rect 15658 12472 15714 12481
rect 15658 12407 15714 12416
rect 15566 12200 15622 12209
rect 15566 12135 15622 12144
rect 15568 11212 15620 11218
rect 15672 11200 15700 12407
rect 15620 11172 15700 11200
rect 15568 11154 15620 11160
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15120 9722 15148 9862
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15120 8974 15148 9522
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 14464 8230 14516 8236
rect 14568 8214 14688 8242
rect 14752 8486 14964 8514
rect 14150 8188 14446 8208
rect 14206 8186 14230 8188
rect 14286 8186 14310 8188
rect 14366 8186 14390 8188
rect 14228 8134 14230 8186
rect 14292 8134 14304 8186
rect 14366 8134 14368 8186
rect 14206 8132 14230 8134
rect 14286 8132 14310 8134
rect 14366 8132 14390 8134
rect 14150 8112 14446 8132
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14002 7712 14058 7721
rect 14002 7647 14058 7656
rect 14016 7410 14044 7647
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13648 6446 13860 6474
rect 13648 6390 13676 6446
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13412 6208 13492 6236
rect 13360 6190 13412 6196
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13280 5778 13308 5850
rect 13556 5778 13584 6258
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13544 5160 13596 5166
rect 13648 5148 13676 6190
rect 14016 5545 14044 7142
rect 14150 7100 14446 7120
rect 14206 7098 14230 7100
rect 14286 7098 14310 7100
rect 14366 7098 14390 7100
rect 14228 7046 14230 7098
rect 14292 7046 14304 7098
rect 14366 7046 14368 7098
rect 14206 7044 14230 7046
rect 14286 7044 14310 7046
rect 14366 7044 14390 7046
rect 14150 7024 14446 7044
rect 14476 7002 14504 7890
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14568 6186 14596 8214
rect 14752 6905 14780 8486
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14936 7546 14964 7686
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14738 6896 14794 6905
rect 14738 6831 14794 6840
rect 15028 6769 15056 8910
rect 15120 8514 15148 8910
rect 15212 8906 15240 9318
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15120 8498 15240 8514
rect 15120 8492 15252 8498
rect 15120 8486 15200 8492
rect 15200 8434 15252 8440
rect 15304 8090 15332 9998
rect 15396 9586 15424 9998
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15014 6760 15070 6769
rect 15014 6695 15070 6704
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14150 6012 14446 6032
rect 14206 6010 14230 6012
rect 14286 6010 14310 6012
rect 14366 6010 14390 6012
rect 14228 5958 14230 6010
rect 14292 5958 14304 6010
rect 14366 5958 14368 6010
rect 14206 5956 14230 5958
rect 14286 5956 14310 5958
rect 14366 5956 14390 5958
rect 14150 5936 14446 5956
rect 14660 5778 14688 6394
rect 15014 6216 15070 6225
rect 15014 6151 15070 6160
rect 15028 6118 15056 6151
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5778 15240 6054
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 14464 5568 14516 5574
rect 14002 5536 14058 5545
rect 14002 5471 14058 5480
rect 14384 5528 14464 5556
rect 14384 5370 14412 5528
rect 14464 5510 14516 5516
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 13596 5120 13676 5148
rect 13544 5102 13596 5108
rect 13556 4690 13584 5102
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14150 4924 14446 4944
rect 14206 4922 14230 4924
rect 14286 4922 14310 4924
rect 14366 4922 14390 4924
rect 14228 4870 14230 4922
rect 14292 4870 14304 4922
rect 14366 4870 14368 4922
rect 14206 4868 14230 4870
rect 14286 4868 14310 4870
rect 14366 4868 14390 4870
rect 14150 4848 14446 4868
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13174 3632 13230 3641
rect 13174 3567 13230 3576
rect 13188 3534 13216 3567
rect 12992 3528 13044 3534
rect 12990 3496 12992 3505
rect 13176 3528 13228 3534
rect 13044 3496 13046 3505
rect 13176 3470 13228 3476
rect 12990 3431 13046 3440
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 2650 12940 3334
rect 13280 2990 13308 3878
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13096 2446 13124 2790
rect 13280 2446 13308 2926
rect 13372 2650 13400 4558
rect 14200 4282 14228 4694
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14660 3942 14688 4966
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14844 4214 14872 4422
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 14844 4078 14872 4150
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14150 3836 14446 3856
rect 14206 3834 14230 3836
rect 14286 3834 14310 3836
rect 14366 3834 14390 3836
rect 14228 3782 14230 3834
rect 14292 3782 14304 3834
rect 14366 3782 14368 3834
rect 14206 3780 14230 3782
rect 14286 3780 14310 3782
rect 14366 3780 14390 3782
rect 14150 3760 14446 3780
rect 14568 3738 14596 3878
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14568 3641 14596 3674
rect 14554 3632 14610 3641
rect 13544 3596 13596 3602
rect 14554 3567 14610 3576
rect 13544 3538 13596 3544
rect 13556 3398 13584 3538
rect 14660 3466 14688 3878
rect 14936 3602 14964 4014
rect 15028 3602 15056 4762
rect 15120 4690 15148 5306
rect 15304 5166 15332 5646
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15212 4622 15240 4966
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15396 4554 15424 8978
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15488 7478 15516 8434
rect 15580 8022 15608 10406
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15672 9518 15700 10134
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15658 9344 15714 9353
rect 15658 9279 15714 9288
rect 15672 8945 15700 9279
rect 15658 8936 15714 8945
rect 15658 8871 15714 8880
rect 15764 8378 15792 15807
rect 15856 10470 15884 17614
rect 15948 16658 15976 17734
rect 16040 17202 16068 18158
rect 16132 17882 16160 18838
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 16132 17134 16160 17478
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15948 16114 15976 16594
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15948 15706 15976 16050
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 16040 14278 16068 14962
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 16040 13977 16068 14214
rect 16026 13968 16082 13977
rect 16026 13903 16082 13912
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16132 13433 16160 13738
rect 16118 13424 16174 13433
rect 16118 13359 16174 13368
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15948 11257 15976 13194
rect 16118 12880 16174 12889
rect 16118 12815 16174 12824
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 16040 11830 16068 12242
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 16132 11286 16160 12815
rect 16120 11280 16172 11286
rect 15934 11248 15990 11257
rect 16120 11222 16172 11228
rect 15934 11183 15990 11192
rect 15948 10792 15976 11183
rect 16028 10804 16080 10810
rect 15948 10764 16028 10792
rect 16028 10746 16080 10752
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15948 9926 15976 10542
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15934 8936 15990 8945
rect 15934 8871 15990 8880
rect 15948 8838 15976 8871
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16040 8430 16068 8774
rect 16224 8514 16252 17682
rect 16408 17678 16436 21655
rect 16762 21520 16818 22000
rect 17314 21520 17370 22000
rect 17958 21520 18014 22000
rect 18602 21520 18658 22000
rect 19154 21520 19210 22000
rect 19798 21520 19854 22000
rect 20442 21520 20498 22000
rect 20994 21520 21050 22000
rect 21638 21520 21694 22000
rect 16578 21040 16634 21049
rect 16578 20975 16634 20984
rect 16592 19242 16620 20975
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 16500 17882 16528 18838
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16592 17678 16620 18906
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16592 17202 16620 17614
rect 16684 17610 16712 19246
rect 16776 18834 16804 21520
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16960 18970 16988 19314
rect 17328 19258 17356 21520
rect 17866 19680 17922 19689
rect 17449 19612 17745 19632
rect 17866 19615 17922 19624
rect 17505 19610 17529 19612
rect 17585 19610 17609 19612
rect 17665 19610 17689 19612
rect 17527 19558 17529 19610
rect 17591 19558 17603 19610
rect 17665 19558 17667 19610
rect 17505 19556 17529 19558
rect 17585 19556 17609 19558
rect 17665 19556 17689 19558
rect 17449 19536 17745 19556
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17236 19230 17356 19258
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16592 16454 16620 17138
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16658 16712 16934
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16684 16250 16712 16594
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16500 14278 16528 14826
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16592 14385 16620 14486
rect 16578 14376 16634 14385
rect 16578 14311 16634 14320
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16776 14090 16804 17070
rect 16868 15570 16896 18702
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16592 14062 16804 14090
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16316 13326 16344 13738
rect 16592 13512 16620 14062
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16408 13484 16620 13512
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16316 12782 16344 13262
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16316 12238 16344 12582
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16304 11620 16356 11626
rect 16304 11562 16356 11568
rect 16316 11082 16344 11562
rect 16408 11098 16436 13484
rect 16486 13424 16542 13433
rect 16486 13359 16542 13368
rect 16580 13388 16632 13394
rect 16500 13326 16528 13359
rect 16580 13330 16632 13336
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16500 12594 16528 13126
rect 16592 12782 16620 13330
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16684 12594 16712 13874
rect 16868 13394 16896 15098
rect 16960 13818 16988 18770
rect 17144 18222 17172 18906
rect 17236 18465 17264 19230
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17328 18601 17356 19110
rect 17604 18970 17632 19110
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17696 18834 17724 19314
rect 17774 19000 17830 19009
rect 17774 18935 17830 18944
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17314 18592 17370 18601
rect 17314 18527 17370 18536
rect 17222 18456 17278 18465
rect 17222 18391 17278 18400
rect 17328 18358 17356 18527
rect 17449 18524 17745 18544
rect 17505 18522 17529 18524
rect 17585 18522 17609 18524
rect 17665 18522 17689 18524
rect 17527 18470 17529 18522
rect 17591 18470 17603 18522
rect 17665 18470 17667 18522
rect 17505 18468 17529 18470
rect 17585 18468 17609 18470
rect 17665 18468 17689 18470
rect 17449 18448 17745 18468
rect 17788 18358 17816 18935
rect 17880 18630 17908 19615
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17316 18352 17368 18358
rect 17316 18294 17368 18300
rect 17776 18352 17828 18358
rect 17776 18294 17828 18300
rect 17132 18216 17184 18222
rect 17038 18184 17094 18193
rect 17132 18158 17184 18164
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17038 18119 17094 18128
rect 17052 18034 17080 18119
rect 17224 18080 17276 18086
rect 17052 18006 17172 18034
rect 17224 18022 17276 18028
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17052 16046 17080 16934
rect 17144 16182 17172 18006
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 17236 16046 17264 18022
rect 17696 17678 17724 18022
rect 17774 17776 17830 17785
rect 17774 17711 17776 17720
rect 17828 17711 17830 17720
rect 17776 17682 17828 17688
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17774 17640 17830 17649
rect 17774 17575 17830 17584
rect 17449 17436 17745 17456
rect 17505 17434 17529 17436
rect 17585 17434 17609 17436
rect 17665 17434 17689 17436
rect 17527 17382 17529 17434
rect 17591 17382 17603 17434
rect 17665 17382 17667 17434
rect 17505 17380 17529 17382
rect 17585 17380 17609 17382
rect 17665 17380 17689 17382
rect 17449 17360 17745 17380
rect 17788 17338 17816 17575
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17328 16794 17356 16934
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17449 16348 17745 16368
rect 17505 16346 17529 16348
rect 17585 16346 17609 16348
rect 17665 16346 17689 16348
rect 17527 16294 17529 16346
rect 17591 16294 17603 16346
rect 17665 16294 17667 16346
rect 17505 16292 17529 16294
rect 17585 16292 17609 16294
rect 17665 16292 17689 16294
rect 17449 16272 17745 16292
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17052 15706 17080 15982
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 17316 15632 17368 15638
rect 17316 15574 17368 15580
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 17052 13938 17080 14894
rect 17328 14822 17356 15574
rect 17449 15260 17745 15280
rect 17505 15258 17529 15260
rect 17585 15258 17609 15260
rect 17665 15258 17689 15260
rect 17527 15206 17529 15258
rect 17591 15206 17603 15258
rect 17665 15206 17667 15258
rect 17505 15204 17529 15206
rect 17585 15204 17609 15206
rect 17665 15204 17689 15206
rect 17449 15184 17745 15204
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17500 14476 17552 14482
rect 17328 14436 17500 14464
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17132 13864 17184 13870
rect 16960 13790 17080 13818
rect 17132 13806 17184 13812
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 16960 13530 16988 13670
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16776 12986 16804 13194
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16960 12714 16988 13262
rect 17052 12986 17080 13790
rect 17144 13462 17172 13806
rect 17236 13802 17264 14214
rect 17328 13938 17356 14436
rect 17500 14418 17552 14424
rect 17449 14172 17745 14192
rect 17505 14170 17529 14172
rect 17585 14170 17609 14172
rect 17665 14170 17689 14172
rect 17527 14118 17529 14170
rect 17591 14118 17603 14170
rect 17665 14118 17667 14170
rect 17505 14116 17529 14118
rect 17585 14116 17609 14118
rect 17665 14116 17689 14118
rect 17449 14096 17745 14116
rect 17498 13968 17554 13977
rect 17316 13932 17368 13938
rect 17498 13903 17500 13912
rect 17316 13874 17368 13880
rect 17552 13903 17554 13912
rect 17500 13874 17552 13880
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17144 12918 17172 13398
rect 17512 13326 17540 13874
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17222 13016 17278 13025
rect 17222 12951 17278 12960
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16500 12566 16712 12594
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16592 11218 16620 12566
rect 16776 12458 16804 12582
rect 16684 12430 16804 12458
rect 16684 12306 16712 12430
rect 16762 12336 16818 12345
rect 16672 12300 16724 12306
rect 16762 12271 16818 12280
rect 16672 12242 16724 12248
rect 16672 12096 16724 12102
rect 16670 12064 16672 12073
rect 16724 12064 16726 12073
rect 16670 11999 16726 12008
rect 16670 11928 16726 11937
rect 16670 11863 16672 11872
rect 16724 11863 16726 11872
rect 16672 11834 16724 11840
rect 16672 11552 16724 11558
rect 16776 11540 16804 12271
rect 16960 12073 16988 12650
rect 16946 12064 17002 12073
rect 16946 11999 17002 12008
rect 16724 11512 16804 11540
rect 16672 11494 16724 11500
rect 16776 11354 16804 11512
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 17052 11218 17080 12786
rect 17236 12730 17264 12951
rect 17328 12850 17356 13262
rect 17449 13084 17745 13104
rect 17505 13082 17529 13084
rect 17585 13082 17609 13084
rect 17665 13082 17689 13084
rect 17527 13030 17529 13082
rect 17591 13030 17603 13082
rect 17665 13030 17667 13082
rect 17505 13028 17529 13030
rect 17585 13028 17609 13030
rect 17665 13028 17689 13030
rect 17449 13008 17745 13028
rect 17316 12844 17368 12850
rect 17368 12804 17632 12832
rect 17316 12786 17368 12792
rect 17236 12702 17356 12730
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 12345 17264 12582
rect 17222 12336 17278 12345
rect 17132 12300 17184 12306
rect 17328 12306 17356 12702
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17222 12271 17278 12280
rect 17316 12300 17368 12306
rect 17132 12242 17184 12248
rect 17316 12242 17368 12248
rect 17144 11626 17172 12242
rect 17224 12232 17276 12238
rect 17512 12209 17540 12582
rect 17604 12238 17632 12804
rect 17788 12782 17816 14758
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17774 12472 17830 12481
rect 17774 12407 17830 12416
rect 17788 12374 17816 12407
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17880 12322 17908 18158
rect 17972 17921 18000 21520
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17958 17912 18014 17921
rect 18064 17882 18092 19110
rect 18328 18828 18380 18834
rect 18328 18770 18380 18776
rect 18236 18760 18288 18766
rect 18156 18708 18236 18714
rect 18156 18702 18288 18708
rect 18156 18686 18276 18702
rect 18156 18222 18184 18686
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 17958 17847 18014 17856
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18156 17814 18184 18158
rect 18340 18154 18368 18770
rect 18616 18737 18644 21520
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18602 18728 18658 18737
rect 18602 18663 18658 18672
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18340 17882 18368 18090
rect 18708 18057 18736 19110
rect 18694 18048 18750 18057
rect 18694 17983 18750 17992
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 17960 17808 18012 17814
rect 18144 17808 18196 17814
rect 17960 17750 18012 17756
rect 18050 17776 18106 17785
rect 17972 16794 18000 17750
rect 18144 17750 18196 17756
rect 18050 17711 18106 17720
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17972 15978 18000 16730
rect 18064 16726 18092 17711
rect 18156 17134 18184 17750
rect 18144 17128 18196 17134
rect 18196 17076 18276 17082
rect 18144 17070 18276 17076
rect 18156 17054 18276 17070
rect 18248 16726 18276 17054
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 18236 16720 18288 16726
rect 18236 16662 18288 16668
rect 18064 16250 18092 16662
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18248 16130 18276 16662
rect 18880 16516 18932 16522
rect 18880 16458 18932 16464
rect 18892 16153 18920 16458
rect 18156 16102 18276 16130
rect 18878 16144 18934 16153
rect 18156 16046 18184 16102
rect 18878 16079 18934 16088
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 18156 15570 18184 15982
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18156 15162 18184 15506
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18156 14550 18184 15098
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 18432 13802 18460 14962
rect 18616 13938 18644 15982
rect 18696 15972 18748 15978
rect 18696 15914 18748 15920
rect 18708 14958 18736 15914
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18892 13938 18920 15302
rect 18984 14822 19012 19314
rect 19168 19258 19196 21520
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19720 19378 19748 19654
rect 19812 19417 19840 21520
rect 19798 19408 19854 19417
rect 19708 19372 19760 19378
rect 19798 19343 19854 19352
rect 19708 19314 19760 19320
rect 19076 19230 19196 19258
rect 19076 17105 19104 19230
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19168 18630 19196 19110
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19444 18358 19472 18770
rect 19432 18352 19484 18358
rect 19154 18320 19210 18329
rect 19432 18294 19484 18300
rect 19154 18255 19210 18264
rect 19168 17678 19196 18255
rect 19248 18148 19300 18154
rect 19248 18090 19300 18096
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19062 17096 19118 17105
rect 19062 17031 19118 17040
rect 19168 15042 19196 17478
rect 19260 17134 19288 18090
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19444 17746 19472 18022
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19444 17338 19472 17682
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19260 16794 19288 17070
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19076 15026 19196 15042
rect 19064 15020 19196 15026
rect 19116 15014 19196 15020
rect 19064 14962 19116 14968
rect 19352 14890 19380 16390
rect 19444 15706 19472 16526
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 19444 14550 19472 15642
rect 19536 14618 19564 17070
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19628 15570 19656 16594
rect 19720 16522 19748 18770
rect 19812 17338 19840 19343
rect 20456 19281 20484 21520
rect 20720 19304 20772 19310
rect 20442 19272 20498 19281
rect 20720 19246 20772 19252
rect 20442 19207 20498 19216
rect 19892 17808 19944 17814
rect 19892 17750 19944 17756
rect 19800 17332 19852 17338
rect 19800 17274 19852 17280
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19628 14618 19656 15506
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18892 13818 18920 13874
rect 19064 13864 19116 13870
rect 18420 13796 18472 13802
rect 18892 13790 19012 13818
rect 19064 13806 19116 13812
rect 18420 13738 18472 13744
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18248 12782 18276 13670
rect 18432 13394 18460 13738
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18236 12776 18288 12782
rect 18142 12744 18198 12753
rect 18236 12718 18288 12724
rect 18142 12679 18198 12688
rect 18156 12646 18184 12679
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 17880 12294 18000 12322
rect 17592 12232 17644 12238
rect 17224 12174 17276 12180
rect 17498 12200 17554 12209
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 16946 11112 17002 11121
rect 16304 11076 16356 11082
rect 16408 11070 16620 11098
rect 16304 11018 16356 11024
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16500 9353 16528 9522
rect 16486 9344 16542 9353
rect 16486 9279 16542 9288
rect 16488 8560 16540 8566
rect 16408 8520 16488 8548
rect 16224 8486 16344 8514
rect 16028 8424 16080 8430
rect 15764 8350 15976 8378
rect 16028 8366 16080 8372
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 15844 8288 15896 8294
rect 15750 8256 15806 8265
rect 15844 8230 15896 8236
rect 15750 8191 15806 8200
rect 15764 8090 15792 8191
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15568 8016 15620 8022
rect 15568 7958 15620 7964
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15672 6866 15700 7278
rect 15764 7002 15792 7686
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15672 6662 15700 6802
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15764 6225 15792 6258
rect 15566 6216 15622 6225
rect 15566 6151 15622 6160
rect 15750 6216 15806 6225
rect 15750 6151 15806 6160
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15304 4146 15332 4422
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 15120 3194 15148 4082
rect 15488 4010 15516 6054
rect 15580 5778 15608 6151
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15580 4758 15608 5510
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15672 4826 15700 4966
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15764 4486 15792 5102
rect 15856 4826 15884 8230
rect 15948 6746 15976 8350
rect 16040 7954 16068 8366
rect 16224 8022 16252 8366
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16132 6934 16160 7346
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 15948 6718 16252 6746
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 6186 16160 6598
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 15936 6112 15988 6118
rect 15988 6072 16068 6100
rect 15936 6054 15988 6060
rect 15934 5808 15990 5817
rect 15934 5743 15936 5752
rect 15988 5743 15990 5752
rect 15936 5714 15988 5720
rect 15934 5672 15990 5681
rect 15934 5607 15990 5616
rect 15948 5574 15976 5607
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15948 5166 15976 5510
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 16040 5098 16068 6072
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15488 3194 15516 3470
rect 15580 3398 15608 3470
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13924 2514 13952 2926
rect 14150 2748 14446 2768
rect 14206 2746 14230 2748
rect 14286 2746 14310 2748
rect 14366 2746 14390 2748
rect 14228 2694 14230 2746
rect 14292 2694 14304 2746
rect 14366 2694 14368 2746
rect 14206 2692 14230 2694
rect 14286 2692 14310 2694
rect 14366 2692 14390 2694
rect 14150 2672 14446 2692
rect 15120 2582 15148 3130
rect 15580 3074 15608 3334
rect 15488 3046 15608 3074
rect 15488 2990 15516 3046
rect 15476 2984 15528 2990
rect 15672 2961 15700 3674
rect 15856 3602 15884 4762
rect 16224 3754 16252 6718
rect 16316 6118 16344 8486
rect 16408 7954 16436 8520
rect 16488 8502 16540 8508
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16408 7721 16436 7890
rect 16394 7712 16450 7721
rect 16394 7647 16450 7656
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16500 5914 16528 6258
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16408 4690 16436 4966
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16224 3726 16436 3754
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 16212 2984 16264 2990
rect 15476 2926 15528 2932
rect 15658 2952 15714 2961
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15488 2514 15516 2926
rect 16212 2926 16264 2932
rect 15658 2887 15660 2896
rect 15712 2887 15714 2896
rect 15660 2858 15712 2864
rect 16224 2854 16252 2926
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16224 2582 16252 2790
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 16408 480 16436 3726
rect 16592 921 16620 11070
rect 16946 11047 17002 11056
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16672 10464 16724 10470
rect 16670 10432 16672 10441
rect 16724 10432 16726 10441
rect 16670 10367 16726 10376
rect 16776 10130 16804 10746
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16670 9616 16726 9625
rect 16670 9551 16726 9560
rect 16684 9450 16712 9551
rect 16868 9518 16896 10406
rect 16960 9518 16988 11047
rect 17038 10296 17094 10305
rect 17144 10266 17172 11562
rect 17236 10810 17264 12174
rect 17592 12174 17644 12180
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17498 12135 17554 12144
rect 17449 11996 17745 12016
rect 17505 11994 17529 11996
rect 17585 11994 17609 11996
rect 17665 11994 17689 11996
rect 17527 11942 17529 11994
rect 17591 11942 17603 11994
rect 17665 11942 17667 11994
rect 17505 11940 17529 11942
rect 17585 11940 17609 11942
rect 17665 11940 17689 11942
rect 17449 11920 17745 11940
rect 17880 11898 17908 12174
rect 17868 11892 17920 11898
rect 17788 11852 17868 11880
rect 17788 11762 17816 11852
rect 17868 11834 17920 11840
rect 17972 11778 18000 12294
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17880 11750 18000 11778
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17420 11150 17448 11562
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17880 11064 17908 11750
rect 17880 11036 18000 11064
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17866 10976 17922 10985
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17328 10674 17356 10950
rect 17449 10908 17745 10928
rect 17866 10911 17922 10920
rect 17505 10906 17529 10908
rect 17585 10906 17609 10908
rect 17665 10906 17689 10908
rect 17527 10854 17529 10906
rect 17591 10854 17603 10906
rect 17665 10854 17667 10906
rect 17505 10852 17529 10854
rect 17585 10852 17609 10854
rect 17665 10852 17689 10854
rect 17449 10832 17745 10852
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17512 10554 17540 10678
rect 17328 10526 17540 10554
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17038 10231 17040 10240
rect 17092 10231 17094 10240
rect 17132 10260 17184 10266
rect 17040 10202 17092 10208
rect 17132 10202 17184 10208
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16764 9376 16816 9382
rect 16670 9344 16726 9353
rect 16764 9318 16816 9324
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16670 9279 16726 9288
rect 16684 8673 16712 9279
rect 16776 9110 16804 9318
rect 16868 9110 16896 9318
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16762 8800 16818 8809
rect 16762 8735 16818 8744
rect 16670 8664 16726 8673
rect 16670 8599 16726 8608
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16684 6730 16712 8366
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 16776 5914 16804 8735
rect 16868 8634 16896 8910
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16868 7342 16896 8230
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16868 6798 16896 7278
rect 16960 7274 16988 8570
rect 17052 8566 17080 9998
rect 17236 9926 17264 10406
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17236 9382 17264 9522
rect 17328 9466 17356 10526
rect 17498 10432 17554 10441
rect 17498 10367 17554 10376
rect 17512 10266 17540 10367
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17788 10198 17816 10542
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17449 9820 17745 9840
rect 17505 9818 17529 9820
rect 17585 9818 17609 9820
rect 17665 9818 17689 9820
rect 17527 9766 17529 9818
rect 17591 9766 17603 9818
rect 17665 9766 17667 9818
rect 17505 9764 17529 9766
rect 17585 9764 17609 9766
rect 17665 9764 17689 9766
rect 17449 9744 17745 9764
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17328 9438 17540 9466
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17314 9208 17370 9217
rect 17314 9143 17370 9152
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 17144 8362 17172 8978
rect 17328 8974 17356 9143
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17420 8906 17448 9318
rect 17512 8906 17540 9438
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17316 8832 17368 8838
rect 17696 8820 17724 9590
rect 17788 9586 17816 9862
rect 17880 9722 17908 10911
rect 17972 10742 18000 11036
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18064 10470 18092 10542
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18050 10160 18106 10169
rect 17960 10124 18012 10130
rect 18050 10095 18106 10104
rect 17960 10066 18012 10072
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17696 8792 17908 8820
rect 17316 8774 17368 8780
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17224 8288 17276 8294
rect 17052 8236 17224 8242
rect 17328 8265 17356 8774
rect 17449 8732 17745 8752
rect 17505 8730 17529 8732
rect 17585 8730 17609 8732
rect 17665 8730 17689 8732
rect 17527 8678 17529 8730
rect 17591 8678 17603 8730
rect 17665 8678 17667 8730
rect 17505 8676 17529 8678
rect 17585 8676 17609 8678
rect 17665 8676 17689 8678
rect 17449 8656 17745 8676
rect 17052 8230 17276 8236
rect 17314 8256 17370 8265
rect 17052 8214 17264 8230
rect 17052 8090 17080 8214
rect 17314 8191 17370 8200
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17038 7984 17094 7993
rect 17038 7919 17040 7928
rect 17092 7919 17094 7928
rect 17040 7890 17092 7896
rect 17144 7585 17172 8026
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17130 7576 17186 7585
rect 17130 7511 17186 7520
rect 16948 7268 17000 7274
rect 16948 7210 17000 7216
rect 17040 7268 17092 7274
rect 17040 7210 17092 7216
rect 17052 6934 17080 7210
rect 17236 7206 17264 7890
rect 17449 7644 17745 7664
rect 17505 7642 17529 7644
rect 17585 7642 17609 7644
rect 17665 7642 17689 7644
rect 17527 7590 17529 7642
rect 17591 7590 17603 7642
rect 17665 7590 17667 7642
rect 17505 7588 17529 7590
rect 17585 7588 17609 7590
rect 17665 7588 17689 7590
rect 17449 7568 17745 7588
rect 17788 7546 17816 7890
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17880 7342 17908 8792
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17236 7002 17264 7142
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17512 6934 17540 7142
rect 17040 6928 17092 6934
rect 16946 6896 17002 6905
rect 17040 6870 17092 6876
rect 17316 6928 17368 6934
rect 17316 6870 17368 6876
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 16946 6831 17002 6840
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16684 3194 16712 3878
rect 16776 3670 16804 3878
rect 16764 3664 16816 3670
rect 16868 3641 16896 6054
rect 16960 4593 16988 6831
rect 17052 6798 17080 6870
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17052 6118 17080 6598
rect 17328 6322 17356 6870
rect 17449 6556 17745 6576
rect 17505 6554 17529 6556
rect 17585 6554 17609 6556
rect 17665 6554 17689 6556
rect 17527 6502 17529 6554
rect 17591 6502 17603 6554
rect 17665 6502 17667 6554
rect 17505 6500 17529 6502
rect 17585 6500 17609 6502
rect 17665 6500 17689 6502
rect 17449 6480 17745 6500
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 17788 5710 17816 6258
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17449 5468 17745 5488
rect 17505 5466 17529 5468
rect 17585 5466 17609 5468
rect 17665 5466 17689 5468
rect 17527 5414 17529 5466
rect 17591 5414 17603 5466
rect 17665 5414 17667 5466
rect 17505 5412 17529 5414
rect 17585 5412 17609 5414
rect 17665 5412 17689 5414
rect 17449 5392 17745 5412
rect 17788 5166 17816 5510
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 16946 4584 17002 4593
rect 16946 4519 17002 4528
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16764 3606 16816 3612
rect 16854 3632 16910 3641
rect 16854 3567 16910 3576
rect 17052 3534 17080 4422
rect 17236 4282 17264 4966
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17328 4162 17356 4626
rect 17604 4622 17632 4966
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17449 4380 17745 4400
rect 17505 4378 17529 4380
rect 17585 4378 17609 4380
rect 17665 4378 17689 4380
rect 17527 4326 17529 4378
rect 17591 4326 17603 4378
rect 17665 4326 17667 4378
rect 17505 4324 17529 4326
rect 17585 4324 17609 4326
rect 17665 4324 17689 4326
rect 17449 4304 17745 4324
rect 17236 4134 17356 4162
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17144 3670 17172 3878
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 17052 2990 17080 3470
rect 17236 3398 17264 4134
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17236 2922 17264 3334
rect 17328 3058 17356 3538
rect 17449 3292 17745 3312
rect 17505 3290 17529 3292
rect 17585 3290 17609 3292
rect 17665 3290 17689 3292
rect 17527 3238 17529 3290
rect 17591 3238 17603 3290
rect 17665 3238 17667 3290
rect 17505 3236 17529 3238
rect 17585 3236 17609 3238
rect 17665 3236 17689 3238
rect 17449 3216 17745 3236
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 17328 2650 17356 2994
rect 17604 2922 17632 2994
rect 17684 2984 17736 2990
rect 17684 2926 17736 2932
rect 17592 2916 17644 2922
rect 17592 2858 17644 2864
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17696 2378 17724 2926
rect 17788 2650 17816 3878
rect 17880 2961 17908 7142
rect 17972 6662 18000 10066
rect 18064 10062 18092 10095
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18064 8362 18092 9998
rect 18248 9518 18276 12718
rect 18340 11354 18368 13262
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18432 12628 18460 13126
rect 18524 12986 18552 13670
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18512 12640 18564 12646
rect 18432 12608 18512 12628
rect 18564 12608 18566 12617
rect 18432 12600 18510 12608
rect 18510 12543 18566 12552
rect 18418 12472 18474 12481
rect 18616 12442 18644 13330
rect 18984 13326 19012 13790
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18800 12850 18828 13194
rect 19076 12850 19104 13806
rect 19156 13456 19208 13462
rect 19156 13398 19208 13404
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 18418 12407 18474 12416
rect 18604 12436 18656 12442
rect 18432 11558 18460 12407
rect 18604 12378 18656 12384
rect 18892 12238 18920 12786
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18892 11626 18920 12174
rect 18880 11620 18932 11626
rect 18932 11580 19012 11608
rect 18880 11562 18932 11568
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18984 11150 19012 11580
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18708 10538 18736 10950
rect 18696 10532 18748 10538
rect 18696 10474 18748 10480
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18432 9654 18460 9998
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18236 9512 18288 9518
rect 18432 9489 18460 9590
rect 18524 9586 18552 10406
rect 18708 10062 18736 10474
rect 18892 10130 18920 11086
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18616 9926 18644 9998
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18236 9454 18288 9460
rect 18418 9480 18474 9489
rect 18144 9444 18196 9450
rect 18418 9415 18474 9424
rect 18144 9386 18196 9392
rect 18156 8974 18184 9386
rect 18524 8974 18552 9522
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18064 7478 18092 7686
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 18050 6760 18106 6769
rect 18050 6695 18052 6704
rect 18104 6695 18106 6704
rect 18052 6666 18104 6672
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 18064 5794 18092 6666
rect 18156 6225 18184 8774
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18248 7449 18276 8434
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18340 7993 18368 8366
rect 18326 7984 18382 7993
rect 18326 7919 18382 7928
rect 18234 7440 18290 7449
rect 18234 7375 18290 7384
rect 18432 6361 18460 8842
rect 18524 8022 18552 8910
rect 18512 8016 18564 8022
rect 18512 7958 18564 7964
rect 18616 7868 18644 9386
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18524 7840 18644 7868
rect 18524 6798 18552 7840
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18616 6866 18644 7142
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18524 6458 18552 6734
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18418 6352 18474 6361
rect 18418 6287 18474 6296
rect 18142 6216 18198 6225
rect 18142 6151 18198 6160
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 17972 4214 18000 5782
rect 18064 5766 18184 5794
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 18064 5166 18092 5646
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18156 4808 18184 5766
rect 18064 4780 18184 4808
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17866 2952 17922 2961
rect 18064 2922 18092 4780
rect 18142 4720 18198 4729
rect 18142 4655 18144 4664
rect 18196 4655 18198 4664
rect 18144 4626 18196 4632
rect 18248 4078 18276 6054
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 17866 2887 17922 2896
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 18064 2446 18092 2858
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 17684 2372 17736 2378
rect 17684 2314 17736 2320
rect 18064 2310 18092 2382
rect 18052 2304 18104 2310
rect 18432 2281 18460 6287
rect 18616 6254 18644 6598
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18708 5166 18736 9318
rect 18800 9081 18828 9386
rect 18786 9072 18842 9081
rect 18786 9007 18842 9016
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18800 7886 18828 8366
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18892 7342 18920 7822
rect 19076 7478 19104 12650
rect 19168 12646 19196 13398
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 12374 19196 12582
rect 19156 12368 19208 12374
rect 19156 12310 19208 12316
rect 19352 11234 19380 13330
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19720 12442 19748 13262
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19444 11801 19472 12310
rect 19812 11898 19840 17002
rect 19904 13682 19932 17750
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20088 16998 20116 17614
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 20088 16114 20116 16526
rect 20166 16280 20222 16289
rect 20166 16215 20222 16224
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19996 15706 20024 15846
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19996 14958 20024 15642
rect 20074 15600 20130 15609
rect 20074 15535 20076 15544
rect 20128 15535 20130 15544
rect 20076 15506 20128 15512
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 20180 14550 20208 16215
rect 20272 15065 20300 17682
rect 20350 16960 20406 16969
rect 20350 16895 20406 16904
rect 20364 16794 20392 16895
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20258 15056 20314 15065
rect 20258 14991 20314 15000
rect 20364 14822 20392 15914
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 20364 13870 20392 14758
rect 20444 14476 20496 14482
rect 20444 14418 20496 14424
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20456 13734 20484 14418
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20444 13728 20496 13734
rect 19904 13654 20392 13682
rect 20444 13670 20496 13676
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19430 11792 19486 11801
rect 20088 11762 20116 13126
rect 20364 12374 20392 13654
rect 20456 12782 20484 13670
rect 20548 13394 20576 14214
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20352 12368 20404 12374
rect 20352 12310 20404 12316
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 19430 11727 19486 11736
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 20180 11694 20208 12174
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20364 11762 20392 12038
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19260 11218 19380 11234
rect 19248 11212 19380 11218
rect 19300 11206 19380 11212
rect 19248 11154 19300 11160
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19352 9602 19380 10678
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19536 10266 19564 10406
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19720 9926 19748 10474
rect 19904 10470 19932 11494
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20088 10674 20116 11290
rect 20364 11286 20392 11698
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19168 9574 19380 9602
rect 19168 9450 19196 9574
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19156 9444 19208 9450
rect 19156 9386 19208 9392
rect 19154 9344 19210 9353
rect 19154 9279 19210 9288
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18786 7032 18842 7041
rect 18892 7002 18920 7278
rect 18786 6967 18842 6976
rect 18880 6996 18932 7002
rect 18800 6866 18828 6967
rect 18880 6938 18932 6944
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18984 5846 19012 6598
rect 18972 5840 19024 5846
rect 18972 5782 19024 5788
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18616 2514 18644 4422
rect 18708 4214 18736 5102
rect 18984 5030 19012 5782
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 19168 4740 19196 9279
rect 19260 7721 19288 9454
rect 19432 9376 19484 9382
rect 19720 9353 19748 9862
rect 19432 9318 19484 9324
rect 19706 9344 19762 9353
rect 19444 9042 19472 9318
rect 19706 9279 19762 9288
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19444 8537 19472 8978
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19430 8528 19486 8537
rect 19430 8463 19486 8472
rect 19432 7948 19484 7954
rect 19536 7936 19564 8774
rect 19904 8129 19932 10406
rect 19996 9994 20024 10406
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 19996 8634 20024 9930
rect 20272 9926 20300 10066
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 19890 8120 19946 8129
rect 19890 8055 19946 8064
rect 19484 7908 19564 7936
rect 19432 7890 19484 7896
rect 19444 7857 19472 7890
rect 19430 7848 19486 7857
rect 19430 7783 19486 7792
rect 19892 7744 19944 7750
rect 19246 7712 19302 7721
rect 19892 7686 19944 7692
rect 19246 7647 19302 7656
rect 19904 7410 19932 7686
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 20088 7313 20116 8298
rect 20166 8256 20222 8265
rect 20166 8191 20222 8200
rect 20074 7304 20130 7313
rect 20074 7239 20130 7248
rect 19800 6928 19852 6934
rect 19800 6870 19852 6876
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19352 5370 19380 5714
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 5234 19472 6598
rect 19628 6202 19656 6734
rect 19524 6180 19576 6186
rect 19628 6174 19748 6202
rect 19524 6122 19576 6128
rect 19536 5914 19564 6122
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19616 5568 19668 5574
rect 19616 5510 19668 5516
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19628 5166 19656 5510
rect 19616 5160 19668 5166
rect 19616 5102 19668 5108
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 19352 4826 19380 5034
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19720 4758 19748 6174
rect 19812 4826 19840 6870
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 19996 6361 20024 6802
rect 19982 6352 20038 6361
rect 19982 6287 20038 6296
rect 20180 6254 20208 8191
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 19892 6112 19944 6118
rect 19892 6054 19944 6060
rect 19904 5302 19932 6054
rect 19996 5370 20024 6190
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19892 5296 19944 5302
rect 19892 5238 19944 5244
rect 20272 5001 20300 9862
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20548 6458 20576 9046
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20640 6338 20668 16594
rect 20548 6310 20668 6338
rect 20258 4992 20314 5001
rect 20258 4927 20314 4936
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19708 4752 19760 4758
rect 19168 4712 19288 4740
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 19168 4078 19196 4558
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18708 3738 18736 3878
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 19168 3534 19196 4014
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 19156 3528 19208 3534
rect 19156 3470 19208 3476
rect 18708 3058 18736 3470
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 19260 2990 19288 4712
rect 19708 4694 19760 4700
rect 19720 4298 19748 4694
rect 20548 4690 20576 6310
rect 20732 5846 20760 19246
rect 21008 18970 21036 21520
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20812 18828 20864 18834
rect 20812 18770 20864 18776
rect 20824 10538 20852 18770
rect 21652 18698 21680 21520
rect 21640 18692 21692 18698
rect 21640 18634 21692 18640
rect 20996 18352 21048 18358
rect 20994 18320 20996 18329
rect 21048 18320 21050 18329
rect 20994 18255 21050 18264
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 21008 8401 21036 17546
rect 20994 8392 21050 8401
rect 20994 8327 21050 8336
rect 20996 6928 21048 6934
rect 20996 6870 21048 6876
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 19720 4282 19840 4298
rect 19720 4276 19852 4282
rect 19720 4270 19800 4276
rect 19800 4218 19852 4224
rect 20444 4004 20496 4010
rect 20444 3946 20496 3952
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 18972 2916 19024 2922
rect 18972 2858 19024 2864
rect 18984 2650 19012 2858
rect 19812 2650 19840 3878
rect 20456 3738 20484 3946
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19996 3194 20024 3538
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19996 2650 20024 3130
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 19800 2644 19852 2650
rect 19800 2586 19852 2592
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 18052 2246 18104 2252
rect 18418 2272 18474 2281
rect 17449 2204 17745 2224
rect 18418 2207 18474 2216
rect 17505 2202 17529 2204
rect 17585 2202 17609 2204
rect 17665 2202 17689 2204
rect 17527 2150 17529 2202
rect 17591 2150 17603 2202
rect 17665 2150 17667 2202
rect 17505 2148 17529 2150
rect 17585 2148 17609 2150
rect 17665 2148 17689 2150
rect 17449 2128 17745 2148
rect 16578 912 16634 921
rect 16578 847 16634 856
rect 20088 480 20116 2926
rect 20456 2582 20484 3674
rect 20444 2576 20496 2582
rect 20444 2518 20496 2524
rect 1766 0 1822 480
rect 5354 0 5410 480
rect 9034 0 9090 480
rect 12714 0 12770 480
rect 16394 0 16450 480
rect 20074 0 20130 480
rect 20548 377 20576 4626
rect 20732 1601 20760 5782
rect 21008 5681 21036 6870
rect 20994 5672 21050 5681
rect 20994 5607 21050 5616
rect 20718 1592 20774 1601
rect 20718 1527 20774 1536
rect 20534 368 20590 377
rect 20534 303 20590 312
<< via2 >>
rect 16394 21664 16450 21720
rect 1306 17720 1362 17776
rect 2410 18944 2466 19000
rect 2042 16668 2044 16688
rect 2044 16668 2096 16688
rect 2096 16668 2098 16688
rect 2042 16632 2098 16668
rect 4254 19610 4310 19612
rect 4334 19610 4390 19612
rect 4414 19610 4470 19612
rect 4494 19610 4550 19612
rect 4254 19558 4280 19610
rect 4280 19558 4310 19610
rect 4334 19558 4344 19610
rect 4344 19558 4390 19610
rect 4414 19558 4460 19610
rect 4460 19558 4470 19610
rect 4494 19558 4524 19610
rect 4524 19558 4550 19610
rect 4254 19556 4310 19558
rect 4334 19556 4390 19558
rect 4414 19556 4470 19558
rect 4494 19556 4550 19558
rect 3974 19080 4030 19136
rect 3606 18828 3662 18864
rect 3606 18808 3608 18828
rect 3608 18808 3660 18828
rect 3660 18808 3662 18828
rect 3422 17856 3478 17912
rect 3422 16632 3478 16688
rect 4254 18522 4310 18524
rect 4334 18522 4390 18524
rect 4414 18522 4470 18524
rect 4494 18522 4550 18524
rect 4254 18470 4280 18522
rect 4280 18470 4310 18522
rect 4334 18470 4344 18522
rect 4344 18470 4390 18522
rect 4414 18470 4460 18522
rect 4460 18470 4470 18522
rect 4494 18470 4524 18522
rect 4524 18470 4550 18522
rect 4254 18468 4310 18470
rect 4334 18468 4390 18470
rect 4414 18468 4470 18470
rect 4494 18468 4550 18470
rect 3974 17176 4030 17232
rect 3698 17040 3754 17096
rect 1490 11056 1546 11112
rect 4802 19080 4858 19136
rect 4802 17856 4858 17912
rect 4254 17434 4310 17436
rect 4334 17434 4390 17436
rect 4414 17434 4470 17436
rect 4494 17434 4550 17436
rect 4254 17382 4280 17434
rect 4280 17382 4310 17434
rect 4334 17382 4344 17434
rect 4344 17382 4390 17434
rect 4414 17382 4460 17434
rect 4460 17382 4470 17434
rect 4494 17382 4524 17434
rect 4524 17382 4550 17434
rect 4254 17380 4310 17382
rect 4334 17380 4390 17382
rect 4414 17380 4470 17382
rect 4494 17380 4550 17382
rect 4254 16346 4310 16348
rect 4334 16346 4390 16348
rect 4414 16346 4470 16348
rect 4494 16346 4550 16348
rect 4254 16294 4280 16346
rect 4280 16294 4310 16346
rect 4334 16294 4344 16346
rect 4344 16294 4390 16346
rect 4414 16294 4460 16346
rect 4460 16294 4470 16346
rect 4494 16294 4524 16346
rect 4524 16294 4550 16346
rect 4254 16292 4310 16294
rect 4334 16292 4390 16294
rect 4414 16292 4470 16294
rect 4494 16292 4550 16294
rect 2870 10648 2926 10704
rect 3330 11056 3386 11112
rect 2226 9444 2282 9480
rect 2226 9424 2228 9444
rect 2228 9424 2280 9444
rect 2280 9424 2282 9444
rect 2410 9288 2466 9344
rect 2686 9172 2742 9208
rect 2686 9152 2688 9172
rect 2688 9152 2740 9172
rect 2740 9152 2742 9172
rect 2962 9596 2964 9616
rect 2964 9596 3016 9616
rect 3016 9596 3018 9616
rect 2962 9560 3018 9596
rect 2686 8336 2742 8392
rect 3422 9016 3478 9072
rect 3330 8744 3386 8800
rect 4254 15258 4310 15260
rect 4334 15258 4390 15260
rect 4414 15258 4470 15260
rect 4494 15258 4550 15260
rect 4254 15206 4280 15258
rect 4280 15206 4310 15258
rect 4334 15206 4344 15258
rect 4344 15206 4390 15258
rect 4414 15206 4460 15258
rect 4460 15206 4470 15258
rect 4494 15206 4524 15258
rect 4524 15206 4550 15258
rect 4254 15204 4310 15206
rect 4334 15204 4390 15206
rect 4414 15204 4470 15206
rect 4494 15204 4550 15206
rect 4254 14170 4310 14172
rect 4334 14170 4390 14172
rect 4414 14170 4470 14172
rect 4494 14170 4550 14172
rect 4254 14118 4280 14170
rect 4280 14118 4310 14170
rect 4334 14118 4344 14170
rect 4344 14118 4390 14170
rect 4414 14118 4460 14170
rect 4460 14118 4470 14170
rect 4494 14118 4524 14170
rect 4524 14118 4550 14170
rect 4254 14116 4310 14118
rect 4334 14116 4390 14118
rect 4414 14116 4470 14118
rect 4494 14116 4550 14118
rect 5446 19216 5502 19272
rect 5262 18944 5318 19000
rect 5906 17584 5962 17640
rect 6826 18128 6882 18184
rect 6550 16088 6606 16144
rect 4254 13082 4310 13084
rect 4334 13082 4390 13084
rect 4414 13082 4470 13084
rect 4494 13082 4550 13084
rect 4254 13030 4280 13082
rect 4280 13030 4310 13082
rect 4334 13030 4344 13082
rect 4344 13030 4390 13082
rect 4414 13030 4460 13082
rect 4460 13030 4470 13082
rect 4494 13030 4524 13082
rect 4524 13030 4550 13082
rect 4254 13028 4310 13030
rect 4334 13028 4390 13030
rect 4414 13028 4470 13030
rect 4494 13028 4550 13030
rect 4254 11994 4310 11996
rect 4334 11994 4390 11996
rect 4414 11994 4470 11996
rect 4494 11994 4550 11996
rect 4254 11942 4280 11994
rect 4280 11942 4310 11994
rect 4334 11942 4344 11994
rect 4344 11942 4390 11994
rect 4414 11942 4460 11994
rect 4460 11942 4470 11994
rect 4494 11942 4524 11994
rect 4524 11942 4550 11994
rect 4254 11940 4310 11942
rect 4334 11940 4390 11942
rect 4414 11940 4470 11942
rect 4494 11940 4550 11942
rect 7553 19066 7609 19068
rect 7633 19066 7689 19068
rect 7713 19066 7769 19068
rect 7793 19066 7849 19068
rect 7553 19014 7579 19066
rect 7579 19014 7609 19066
rect 7633 19014 7643 19066
rect 7643 19014 7689 19066
rect 7713 19014 7759 19066
rect 7759 19014 7769 19066
rect 7793 19014 7823 19066
rect 7823 19014 7849 19066
rect 7553 19012 7609 19014
rect 7633 19012 7689 19014
rect 7713 19012 7769 19014
rect 7793 19012 7849 19014
rect 7553 17978 7609 17980
rect 7633 17978 7689 17980
rect 7713 17978 7769 17980
rect 7793 17978 7849 17980
rect 7553 17926 7579 17978
rect 7579 17926 7609 17978
rect 7633 17926 7643 17978
rect 7643 17926 7689 17978
rect 7713 17926 7759 17978
rect 7759 17926 7769 17978
rect 7793 17926 7823 17978
rect 7823 17926 7849 17978
rect 7553 17924 7609 17926
rect 7633 17924 7689 17926
rect 7713 17924 7769 17926
rect 7793 17924 7849 17926
rect 7470 17720 7526 17776
rect 8298 19216 8354 19272
rect 8666 17584 8722 17640
rect 7553 16890 7609 16892
rect 7633 16890 7689 16892
rect 7713 16890 7769 16892
rect 7793 16890 7849 16892
rect 7553 16838 7579 16890
rect 7579 16838 7609 16890
rect 7633 16838 7643 16890
rect 7643 16838 7689 16890
rect 7713 16838 7759 16890
rect 7759 16838 7769 16890
rect 7793 16838 7823 16890
rect 7823 16838 7849 16890
rect 7553 16836 7609 16838
rect 7633 16836 7689 16838
rect 7713 16836 7769 16838
rect 7793 16836 7849 16838
rect 5354 11600 5410 11656
rect 4254 10906 4310 10908
rect 4334 10906 4390 10908
rect 4414 10906 4470 10908
rect 4494 10906 4550 10908
rect 4254 10854 4280 10906
rect 4280 10854 4310 10906
rect 4334 10854 4344 10906
rect 4344 10854 4390 10906
rect 4414 10854 4460 10906
rect 4460 10854 4470 10906
rect 4494 10854 4524 10906
rect 4524 10854 4550 10906
rect 4254 10852 4310 10854
rect 4334 10852 4390 10854
rect 4414 10852 4470 10854
rect 4494 10852 4550 10854
rect 3974 10104 4030 10160
rect 4066 9968 4122 10024
rect 5078 9968 5134 10024
rect 3054 8492 3110 8528
rect 3054 8472 3056 8492
rect 3056 8472 3108 8492
rect 3108 8472 3110 8492
rect 4254 9818 4310 9820
rect 4334 9818 4390 9820
rect 4414 9818 4470 9820
rect 4494 9818 4550 9820
rect 4254 9766 4280 9818
rect 4280 9766 4310 9818
rect 4334 9766 4344 9818
rect 4344 9766 4390 9818
rect 4414 9766 4460 9818
rect 4460 9766 4470 9818
rect 4494 9766 4524 9818
rect 4524 9766 4550 9818
rect 4254 9764 4310 9766
rect 4334 9764 4390 9766
rect 4414 9764 4470 9766
rect 4494 9764 4550 9766
rect 4802 9696 4858 9752
rect 3882 8200 3938 8256
rect 2962 8064 3018 8120
rect 3606 7948 3662 7984
rect 3606 7928 3608 7948
rect 3608 7928 3660 7948
rect 3660 7928 3662 7948
rect 3790 7828 3792 7848
rect 3792 7828 3844 7848
rect 3844 7828 3846 7848
rect 3790 7792 3846 7828
rect 3606 7420 3608 7440
rect 3608 7420 3660 7440
rect 3660 7420 3662 7440
rect 3606 7384 3662 7420
rect 3974 7268 4030 7304
rect 3974 7248 3976 7268
rect 3976 7248 4028 7268
rect 4028 7248 4030 7268
rect 4254 8730 4310 8732
rect 4334 8730 4390 8732
rect 4414 8730 4470 8732
rect 4494 8730 4550 8732
rect 4254 8678 4280 8730
rect 4280 8678 4310 8730
rect 4334 8678 4344 8730
rect 4344 8678 4390 8730
rect 4414 8678 4460 8730
rect 4460 8678 4470 8730
rect 4494 8678 4524 8730
rect 4524 8678 4550 8730
rect 4254 8676 4310 8678
rect 4334 8676 4390 8678
rect 4414 8676 4470 8678
rect 4494 8676 4550 8678
rect 6274 10376 6330 10432
rect 4254 7642 4310 7644
rect 4334 7642 4390 7644
rect 4414 7642 4470 7644
rect 4494 7642 4550 7644
rect 4254 7590 4280 7642
rect 4280 7590 4310 7642
rect 4334 7590 4344 7642
rect 4344 7590 4390 7642
rect 4414 7590 4460 7642
rect 4460 7590 4470 7642
rect 4494 7590 4524 7642
rect 4524 7590 4550 7642
rect 4254 7588 4310 7590
rect 4334 7588 4390 7590
rect 4414 7588 4470 7590
rect 4494 7588 4550 7590
rect 6458 10784 6514 10840
rect 3606 6160 3662 6216
rect 4254 6554 4310 6556
rect 4334 6554 4390 6556
rect 4414 6554 4470 6556
rect 4494 6554 4550 6556
rect 4254 6502 4280 6554
rect 4280 6502 4310 6554
rect 4334 6502 4344 6554
rect 4344 6502 4390 6554
rect 4414 6502 4460 6554
rect 4460 6502 4470 6554
rect 4494 6502 4524 6554
rect 4524 6502 4550 6554
rect 4254 6500 4310 6502
rect 4334 6500 4390 6502
rect 4414 6500 4470 6502
rect 4494 6500 4550 6502
rect 4254 5466 4310 5468
rect 4334 5466 4390 5468
rect 4414 5466 4470 5468
rect 4494 5466 4550 5468
rect 4254 5414 4280 5466
rect 4280 5414 4310 5466
rect 4334 5414 4344 5466
rect 4344 5414 4390 5466
rect 4414 5414 4460 5466
rect 4460 5414 4470 5466
rect 4494 5414 4524 5466
rect 4524 5414 4550 5466
rect 4254 5412 4310 5414
rect 4334 5412 4390 5414
rect 4414 5412 4470 5414
rect 4494 5412 4550 5414
rect 4254 4378 4310 4380
rect 4334 4378 4390 4380
rect 4414 4378 4470 4380
rect 4494 4378 4550 4380
rect 4254 4326 4280 4378
rect 4280 4326 4310 4378
rect 4334 4326 4344 4378
rect 4344 4326 4390 4378
rect 4414 4326 4460 4378
rect 4460 4326 4470 4378
rect 4494 4326 4524 4378
rect 4524 4326 4550 4378
rect 4254 4324 4310 4326
rect 4334 4324 4390 4326
rect 4414 4324 4470 4326
rect 4494 4324 4550 4326
rect 4254 3290 4310 3292
rect 4334 3290 4390 3292
rect 4414 3290 4470 3292
rect 4494 3290 4550 3292
rect 4254 3238 4280 3290
rect 4280 3238 4310 3290
rect 4334 3238 4344 3290
rect 4344 3238 4390 3290
rect 4414 3238 4460 3290
rect 4460 3238 4470 3290
rect 4494 3238 4524 3290
rect 4524 3238 4550 3290
rect 4254 3236 4310 3238
rect 4334 3236 4390 3238
rect 4414 3236 4470 3238
rect 4494 3236 4550 3238
rect 4710 3188 4766 3224
rect 4710 3168 4712 3188
rect 4712 3168 4764 3188
rect 4764 3168 4766 3188
rect 7553 15802 7609 15804
rect 7633 15802 7689 15804
rect 7713 15802 7769 15804
rect 7793 15802 7849 15804
rect 7553 15750 7579 15802
rect 7579 15750 7609 15802
rect 7633 15750 7643 15802
rect 7643 15750 7689 15802
rect 7713 15750 7759 15802
rect 7759 15750 7769 15802
rect 7793 15750 7823 15802
rect 7823 15750 7849 15802
rect 7553 15748 7609 15750
rect 7633 15748 7689 15750
rect 7713 15748 7769 15750
rect 7793 15748 7849 15750
rect 9218 16496 9274 16552
rect 7553 14714 7609 14716
rect 7633 14714 7689 14716
rect 7713 14714 7769 14716
rect 7793 14714 7849 14716
rect 7553 14662 7579 14714
rect 7579 14662 7609 14714
rect 7633 14662 7643 14714
rect 7643 14662 7689 14714
rect 7713 14662 7759 14714
rect 7759 14662 7769 14714
rect 7793 14662 7823 14714
rect 7823 14662 7849 14714
rect 7553 14660 7609 14662
rect 7633 14660 7689 14662
rect 7713 14660 7769 14662
rect 7793 14660 7849 14662
rect 7553 13626 7609 13628
rect 7633 13626 7689 13628
rect 7713 13626 7769 13628
rect 7793 13626 7849 13628
rect 7553 13574 7579 13626
rect 7579 13574 7609 13626
rect 7633 13574 7643 13626
rect 7643 13574 7689 13626
rect 7713 13574 7759 13626
rect 7759 13574 7769 13626
rect 7793 13574 7823 13626
rect 7823 13574 7849 13626
rect 7553 13572 7609 13574
rect 7633 13572 7689 13574
rect 7713 13572 7769 13574
rect 7793 13572 7849 13574
rect 7553 12538 7609 12540
rect 7633 12538 7689 12540
rect 7713 12538 7769 12540
rect 7793 12538 7849 12540
rect 7553 12486 7579 12538
rect 7579 12486 7609 12538
rect 7633 12486 7643 12538
rect 7643 12486 7689 12538
rect 7713 12486 7759 12538
rect 7759 12486 7769 12538
rect 7793 12486 7823 12538
rect 7823 12486 7849 12538
rect 7553 12484 7609 12486
rect 7633 12484 7689 12486
rect 7713 12484 7769 12486
rect 7793 12484 7849 12486
rect 7553 11450 7609 11452
rect 7633 11450 7689 11452
rect 7713 11450 7769 11452
rect 7793 11450 7849 11452
rect 7553 11398 7579 11450
rect 7579 11398 7609 11450
rect 7633 11398 7643 11450
rect 7643 11398 7689 11450
rect 7713 11398 7759 11450
rect 7759 11398 7769 11450
rect 7793 11398 7823 11450
rect 7823 11398 7849 11450
rect 7553 11396 7609 11398
rect 7633 11396 7689 11398
rect 7713 11396 7769 11398
rect 7793 11396 7849 11398
rect 7102 10512 7158 10568
rect 6274 5752 6330 5808
rect 6550 5652 6552 5672
rect 6552 5652 6604 5672
rect 6604 5652 6606 5672
rect 6550 5616 6606 5652
rect 7102 9424 7158 9480
rect 7102 9288 7158 9344
rect 7102 8608 7158 8664
rect 8298 10784 8354 10840
rect 7378 10376 7434 10432
rect 7553 10362 7609 10364
rect 7633 10362 7689 10364
rect 7713 10362 7769 10364
rect 7793 10362 7849 10364
rect 7553 10310 7579 10362
rect 7579 10310 7609 10362
rect 7633 10310 7643 10362
rect 7643 10310 7689 10362
rect 7713 10310 7759 10362
rect 7759 10310 7769 10362
rect 7793 10310 7823 10362
rect 7823 10310 7849 10362
rect 7553 10308 7609 10310
rect 7633 10308 7689 10310
rect 7713 10308 7769 10310
rect 7793 10308 7849 10310
rect 8022 9288 8078 9344
rect 7553 9274 7609 9276
rect 7633 9274 7689 9276
rect 7713 9274 7769 9276
rect 7793 9274 7849 9276
rect 7553 9222 7579 9274
rect 7579 9222 7609 9274
rect 7633 9222 7643 9274
rect 7643 9222 7689 9274
rect 7713 9222 7759 9274
rect 7759 9222 7769 9274
rect 7793 9222 7823 9274
rect 7823 9222 7849 9274
rect 7553 9220 7609 9222
rect 7633 9220 7689 9222
rect 7713 9220 7769 9222
rect 7793 9220 7849 9222
rect 7930 9152 7986 9208
rect 8482 10240 8538 10296
rect 8758 10648 8814 10704
rect 8482 9832 8538 9888
rect 7930 8336 7986 8392
rect 7286 8200 7342 8256
rect 7010 8064 7066 8120
rect 7553 8186 7609 8188
rect 7633 8186 7689 8188
rect 7713 8186 7769 8188
rect 7793 8186 7849 8188
rect 7553 8134 7579 8186
rect 7579 8134 7609 8186
rect 7633 8134 7643 8186
rect 7643 8134 7689 8186
rect 7713 8134 7759 8186
rect 7759 8134 7769 8186
rect 7793 8134 7823 8186
rect 7823 8134 7849 8186
rect 7553 8132 7609 8134
rect 7633 8132 7689 8134
rect 7713 8132 7769 8134
rect 7793 8132 7849 8134
rect 7553 7098 7609 7100
rect 7633 7098 7689 7100
rect 7713 7098 7769 7100
rect 7793 7098 7849 7100
rect 7553 7046 7579 7098
rect 7579 7046 7609 7098
rect 7633 7046 7643 7098
rect 7643 7046 7689 7098
rect 7713 7046 7759 7098
rect 7759 7046 7769 7098
rect 7793 7046 7823 7098
rect 7823 7046 7849 7098
rect 7553 7044 7609 7046
rect 7633 7044 7689 7046
rect 7713 7044 7769 7046
rect 7793 7044 7849 7046
rect 7654 6704 7710 6760
rect 7553 6010 7609 6012
rect 7633 6010 7689 6012
rect 7713 6010 7769 6012
rect 7793 6010 7849 6012
rect 7553 5958 7579 6010
rect 7579 5958 7609 6010
rect 7633 5958 7643 6010
rect 7643 5958 7689 6010
rect 7713 5958 7759 6010
rect 7759 5958 7769 6010
rect 7793 5958 7823 6010
rect 7823 5958 7849 6010
rect 7553 5956 7609 5958
rect 7633 5956 7689 5958
rect 7713 5956 7769 5958
rect 7793 5956 7849 5958
rect 8298 7112 8354 7168
rect 7553 4922 7609 4924
rect 7633 4922 7689 4924
rect 7713 4922 7769 4924
rect 7793 4922 7849 4924
rect 7553 4870 7579 4922
rect 7579 4870 7609 4922
rect 7633 4870 7643 4922
rect 7643 4870 7689 4922
rect 7713 4870 7759 4922
rect 7759 4870 7769 4922
rect 7793 4870 7823 4922
rect 7823 4870 7849 4922
rect 7553 4868 7609 4870
rect 7633 4868 7689 4870
rect 7713 4868 7769 4870
rect 7793 4868 7849 4870
rect 10322 18964 10378 19000
rect 10322 18944 10324 18964
rect 10324 18944 10376 18964
rect 10376 18944 10378 18964
rect 10414 17992 10470 18048
rect 10852 19610 10908 19612
rect 10932 19610 10988 19612
rect 11012 19610 11068 19612
rect 11092 19610 11148 19612
rect 10852 19558 10878 19610
rect 10878 19558 10908 19610
rect 10932 19558 10942 19610
rect 10942 19558 10988 19610
rect 11012 19558 11058 19610
rect 11058 19558 11068 19610
rect 11092 19558 11122 19610
rect 11122 19558 11148 19610
rect 10852 19556 10908 19558
rect 10932 19556 10988 19558
rect 11012 19556 11068 19558
rect 11092 19556 11148 19558
rect 10874 19352 10930 19408
rect 10852 18522 10908 18524
rect 10932 18522 10988 18524
rect 11012 18522 11068 18524
rect 11092 18522 11148 18524
rect 10852 18470 10878 18522
rect 10878 18470 10908 18522
rect 10932 18470 10942 18522
rect 10942 18470 10988 18522
rect 11012 18470 11058 18522
rect 11058 18470 11068 18522
rect 11092 18470 11122 18522
rect 11122 18470 11148 18522
rect 10852 18468 10908 18470
rect 10932 18468 10988 18470
rect 11012 18468 11068 18470
rect 11092 18468 11148 18470
rect 10874 18264 10930 18320
rect 10852 17434 10908 17436
rect 10932 17434 10988 17436
rect 11012 17434 11068 17436
rect 11092 17434 11148 17436
rect 10852 17382 10878 17434
rect 10878 17382 10908 17434
rect 10932 17382 10942 17434
rect 10942 17382 10988 17434
rect 11012 17382 11058 17434
rect 11058 17382 11068 17434
rect 11092 17382 11122 17434
rect 11122 17382 11148 17434
rect 10852 17380 10908 17382
rect 10932 17380 10988 17382
rect 11012 17380 11068 17382
rect 11092 17380 11148 17382
rect 11242 17176 11298 17232
rect 10852 16346 10908 16348
rect 10932 16346 10988 16348
rect 11012 16346 11068 16348
rect 11092 16346 11148 16348
rect 10852 16294 10878 16346
rect 10878 16294 10908 16346
rect 10932 16294 10942 16346
rect 10942 16294 10988 16346
rect 11012 16294 11058 16346
rect 11058 16294 11068 16346
rect 11092 16294 11122 16346
rect 11122 16294 11148 16346
rect 10852 16292 10908 16294
rect 10932 16292 10988 16294
rect 11012 16292 11068 16294
rect 11092 16292 11148 16294
rect 11426 16904 11482 16960
rect 10852 15258 10908 15260
rect 10932 15258 10988 15260
rect 11012 15258 11068 15260
rect 11092 15258 11148 15260
rect 10852 15206 10878 15258
rect 10878 15206 10908 15258
rect 10932 15206 10942 15258
rect 10942 15206 10988 15258
rect 11012 15206 11058 15258
rect 11058 15206 11068 15258
rect 11092 15206 11122 15258
rect 11122 15206 11148 15258
rect 10852 15204 10908 15206
rect 10932 15204 10988 15206
rect 11012 15204 11068 15206
rect 11092 15204 11148 15206
rect 9678 11600 9734 11656
rect 9586 10240 9642 10296
rect 9126 9832 9182 9888
rect 9678 9832 9734 9888
rect 10138 9968 10194 10024
rect 9862 6976 9918 7032
rect 10138 8200 10194 8256
rect 9218 6160 9274 6216
rect 10138 6060 10140 6080
rect 10140 6060 10192 6080
rect 10192 6060 10194 6080
rect 10138 6024 10194 6060
rect 7553 3834 7609 3836
rect 7633 3834 7689 3836
rect 7713 3834 7769 3836
rect 7793 3834 7849 3836
rect 7553 3782 7579 3834
rect 7579 3782 7609 3834
rect 7633 3782 7643 3834
rect 7643 3782 7689 3834
rect 7713 3782 7759 3834
rect 7759 3782 7769 3834
rect 7793 3782 7823 3834
rect 7823 3782 7849 3834
rect 7553 3780 7609 3782
rect 7633 3780 7689 3782
rect 7713 3780 7769 3782
rect 7793 3780 7849 3782
rect 7553 2746 7609 2748
rect 7633 2746 7689 2748
rect 7713 2746 7769 2748
rect 7793 2746 7849 2748
rect 7553 2694 7579 2746
rect 7579 2694 7609 2746
rect 7633 2694 7643 2746
rect 7643 2694 7689 2746
rect 7713 2694 7759 2746
rect 7759 2694 7769 2746
rect 7793 2694 7823 2746
rect 7823 2694 7849 2746
rect 7553 2692 7609 2694
rect 7633 2692 7689 2694
rect 7713 2692 7769 2694
rect 7793 2692 7849 2694
rect 9126 3168 9182 3224
rect 4254 2202 4310 2204
rect 4334 2202 4390 2204
rect 4414 2202 4470 2204
rect 4494 2202 4550 2204
rect 4254 2150 4280 2202
rect 4280 2150 4310 2202
rect 4334 2150 4344 2202
rect 4344 2150 4390 2202
rect 4414 2150 4460 2202
rect 4460 2150 4470 2202
rect 4494 2150 4524 2202
rect 4524 2150 4550 2202
rect 4254 2148 4310 2150
rect 4334 2148 4390 2150
rect 4414 2148 4470 2150
rect 4494 2148 4550 2150
rect 10852 14170 10908 14172
rect 10932 14170 10988 14172
rect 11012 14170 11068 14172
rect 11092 14170 11148 14172
rect 10852 14118 10878 14170
rect 10878 14118 10908 14170
rect 10932 14118 10942 14170
rect 10942 14118 10988 14170
rect 11012 14118 11058 14170
rect 11058 14118 11068 14170
rect 11092 14118 11122 14170
rect 11122 14118 11148 14170
rect 10852 14116 10908 14118
rect 10932 14116 10988 14118
rect 11012 14116 11068 14118
rect 11092 14116 11148 14118
rect 10598 12144 10654 12200
rect 10852 13082 10908 13084
rect 10932 13082 10988 13084
rect 11012 13082 11068 13084
rect 11092 13082 11148 13084
rect 10852 13030 10878 13082
rect 10878 13030 10908 13082
rect 10932 13030 10942 13082
rect 10942 13030 10988 13082
rect 11012 13030 11058 13082
rect 11058 13030 11068 13082
rect 11092 13030 11122 13082
rect 11122 13030 11148 13082
rect 10852 13028 10908 13030
rect 10932 13028 10988 13030
rect 11012 13028 11068 13030
rect 11092 13028 11148 13030
rect 11150 12588 11152 12608
rect 11152 12588 11204 12608
rect 11204 12588 11206 12608
rect 11150 12552 11206 12588
rect 10966 12416 11022 12472
rect 10966 12300 11022 12336
rect 10966 12280 10968 12300
rect 10968 12280 11020 12300
rect 11020 12280 11022 12300
rect 10852 11994 10908 11996
rect 10932 11994 10988 11996
rect 11012 11994 11068 11996
rect 11092 11994 11148 11996
rect 10852 11942 10878 11994
rect 10878 11942 10908 11994
rect 10932 11942 10942 11994
rect 10942 11942 10988 11994
rect 11012 11942 11058 11994
rect 11058 11942 11068 11994
rect 11092 11942 11122 11994
rect 11122 11942 11148 11994
rect 10852 11940 10908 11942
rect 10932 11940 10988 11942
rect 11012 11940 11068 11942
rect 11092 11940 11148 11942
rect 10852 10906 10908 10908
rect 10932 10906 10988 10908
rect 11012 10906 11068 10908
rect 11092 10906 11148 10908
rect 10852 10854 10878 10906
rect 10878 10854 10908 10906
rect 10932 10854 10942 10906
rect 10942 10854 10988 10906
rect 11012 10854 11058 10906
rect 11058 10854 11068 10906
rect 11092 10854 11122 10906
rect 11122 10854 11148 10906
rect 10852 10852 10908 10854
rect 10932 10852 10988 10854
rect 11012 10852 11068 10854
rect 11092 10852 11148 10854
rect 11610 12552 11666 12608
rect 11426 11056 11482 11112
rect 10782 10648 10838 10704
rect 10414 9696 10470 9752
rect 12254 19372 12310 19408
rect 12254 19352 12256 19372
rect 12256 19352 12308 19372
rect 12308 19352 12310 19372
rect 11978 19080 12034 19136
rect 12254 18672 12310 18728
rect 12162 17992 12218 18048
rect 12254 17176 12310 17232
rect 12806 19080 12862 19136
rect 12714 16904 12770 16960
rect 12622 16108 12678 16144
rect 12622 16088 12624 16108
rect 12624 16088 12676 16108
rect 12676 16088 12678 16108
rect 13266 18944 13322 19000
rect 13266 18400 13322 18456
rect 13174 16904 13230 16960
rect 13910 19352 13966 19408
rect 14186 19252 14188 19272
rect 14188 19252 14240 19272
rect 14240 19252 14242 19272
rect 14186 19216 14242 19252
rect 14150 19066 14206 19068
rect 14230 19066 14286 19068
rect 14310 19066 14366 19068
rect 14390 19066 14446 19068
rect 14150 19014 14176 19066
rect 14176 19014 14206 19066
rect 14230 19014 14240 19066
rect 14240 19014 14286 19066
rect 14310 19014 14356 19066
rect 14356 19014 14366 19066
rect 14390 19014 14420 19066
rect 14420 19014 14446 19066
rect 14150 19012 14206 19014
rect 14230 19012 14286 19014
rect 14310 19012 14366 19014
rect 14390 19012 14446 19014
rect 14278 18536 14334 18592
rect 14370 18400 14426 18456
rect 14150 17978 14206 17980
rect 14230 17978 14286 17980
rect 14310 17978 14366 17980
rect 14390 17978 14446 17980
rect 14150 17926 14176 17978
rect 14176 17926 14206 17978
rect 14230 17926 14240 17978
rect 14240 17926 14286 17978
rect 14310 17926 14356 17978
rect 14356 17926 14366 17978
rect 14390 17926 14420 17978
rect 14420 17926 14446 17978
rect 14150 17924 14206 17926
rect 14230 17924 14286 17926
rect 14310 17924 14366 17926
rect 14390 17924 14446 17926
rect 15934 20304 15990 20360
rect 14738 18264 14794 18320
rect 14150 16890 14206 16892
rect 14230 16890 14286 16892
rect 14310 16890 14366 16892
rect 14390 16890 14446 16892
rect 14150 16838 14176 16890
rect 14176 16838 14206 16890
rect 14230 16838 14240 16890
rect 14240 16838 14286 16890
rect 14310 16838 14356 16890
rect 14356 16838 14366 16890
rect 14390 16838 14420 16890
rect 14420 16838 14446 16890
rect 14150 16836 14206 16838
rect 14230 16836 14286 16838
rect 14310 16836 14366 16838
rect 14390 16836 14446 16838
rect 14150 15802 14206 15804
rect 14230 15802 14286 15804
rect 14310 15802 14366 15804
rect 14390 15802 14446 15804
rect 14150 15750 14176 15802
rect 14176 15750 14206 15802
rect 14230 15750 14240 15802
rect 14240 15750 14286 15802
rect 14310 15750 14356 15802
rect 14356 15750 14366 15802
rect 14390 15750 14420 15802
rect 14420 15750 14446 15802
rect 14150 15748 14206 15750
rect 14230 15748 14286 15750
rect 14310 15748 14366 15750
rect 14390 15748 14446 15750
rect 14554 16360 14610 16416
rect 14830 16496 14886 16552
rect 14738 15952 14794 16008
rect 14150 14714 14206 14716
rect 14230 14714 14286 14716
rect 14310 14714 14366 14716
rect 14390 14714 14446 14716
rect 14150 14662 14176 14714
rect 14176 14662 14206 14714
rect 14230 14662 14240 14714
rect 14240 14662 14286 14714
rect 14310 14662 14356 14714
rect 14356 14662 14366 14714
rect 14390 14662 14420 14714
rect 14420 14662 14446 14714
rect 14150 14660 14206 14662
rect 14230 14660 14286 14662
rect 14310 14660 14366 14662
rect 14390 14660 14446 14662
rect 12438 12180 12440 12200
rect 12440 12180 12492 12200
rect 12492 12180 12494 12200
rect 12438 12144 12494 12180
rect 11702 10104 11758 10160
rect 10852 9818 10908 9820
rect 10932 9818 10988 9820
rect 11012 9818 11068 9820
rect 11092 9818 11148 9820
rect 10852 9766 10878 9818
rect 10878 9766 10908 9818
rect 10932 9766 10942 9818
rect 10942 9766 10988 9818
rect 11012 9766 11058 9818
rect 11058 9766 11068 9818
rect 11092 9766 11122 9818
rect 11122 9766 11148 9818
rect 10852 9764 10908 9766
rect 10932 9764 10988 9766
rect 11012 9764 11068 9766
rect 11092 9764 11148 9766
rect 11794 9696 11850 9752
rect 10852 8730 10908 8732
rect 10932 8730 10988 8732
rect 11012 8730 11068 8732
rect 11092 8730 11148 8732
rect 10852 8678 10878 8730
rect 10878 8678 10908 8730
rect 10932 8678 10942 8730
rect 10942 8678 10988 8730
rect 11012 8678 11058 8730
rect 11058 8678 11068 8730
rect 11092 8678 11122 8730
rect 11122 8678 11148 8730
rect 10852 8676 10908 8678
rect 10932 8676 10988 8678
rect 11012 8676 11068 8678
rect 11092 8676 11148 8678
rect 11978 10104 12034 10160
rect 11702 9288 11758 9344
rect 11702 8608 11758 8664
rect 10852 7642 10908 7644
rect 10932 7642 10988 7644
rect 11012 7642 11068 7644
rect 11092 7642 11148 7644
rect 10852 7590 10878 7642
rect 10878 7590 10908 7642
rect 10932 7590 10942 7642
rect 10942 7590 10988 7642
rect 11012 7590 11058 7642
rect 11058 7590 11068 7642
rect 11092 7590 11122 7642
rect 11122 7590 11148 7642
rect 10852 7588 10908 7590
rect 10932 7588 10988 7590
rect 11012 7588 11068 7590
rect 11092 7588 11148 7590
rect 11334 7520 11390 7576
rect 11334 7112 11390 7168
rect 11794 6976 11850 7032
rect 10852 6554 10908 6556
rect 10932 6554 10988 6556
rect 11012 6554 11068 6556
rect 11092 6554 11148 6556
rect 10852 6502 10878 6554
rect 10878 6502 10908 6554
rect 10932 6502 10942 6554
rect 10942 6502 10988 6554
rect 11012 6502 11058 6554
rect 11058 6502 11068 6554
rect 11092 6502 11122 6554
rect 11122 6502 11148 6554
rect 10852 6500 10908 6502
rect 10932 6500 10988 6502
rect 11012 6500 11068 6502
rect 11092 6500 11148 6502
rect 10506 5888 10562 5944
rect 10230 4120 10286 4176
rect 10852 5466 10908 5468
rect 10932 5466 10988 5468
rect 11012 5466 11068 5468
rect 11092 5466 11148 5468
rect 10852 5414 10878 5466
rect 10878 5414 10908 5466
rect 10932 5414 10942 5466
rect 10942 5414 10988 5466
rect 11012 5414 11058 5466
rect 11058 5414 11068 5466
rect 11092 5414 11122 5466
rect 11122 5414 11148 5466
rect 10852 5412 10908 5414
rect 10932 5412 10988 5414
rect 11012 5412 11068 5414
rect 11092 5412 11148 5414
rect 11426 5480 11482 5536
rect 10852 4378 10908 4380
rect 10932 4378 10988 4380
rect 11012 4378 11068 4380
rect 11092 4378 11148 4380
rect 10852 4326 10878 4378
rect 10878 4326 10908 4378
rect 10932 4326 10942 4378
rect 10942 4326 10988 4378
rect 11012 4326 11058 4378
rect 11058 4326 11068 4378
rect 11092 4326 11122 4378
rect 11122 4326 11148 4378
rect 10852 4324 10908 4326
rect 10932 4324 10988 4326
rect 11012 4324 11068 4326
rect 11092 4324 11148 4326
rect 10782 3576 10838 3632
rect 11242 3440 11298 3496
rect 10852 3290 10908 3292
rect 10932 3290 10988 3292
rect 11012 3290 11068 3292
rect 11092 3290 11148 3292
rect 10852 3238 10878 3290
rect 10878 3238 10908 3290
rect 10932 3238 10942 3290
rect 10942 3238 10988 3290
rect 11012 3238 11058 3290
rect 11058 3238 11068 3290
rect 11092 3238 11122 3290
rect 11122 3238 11148 3290
rect 10852 3236 10908 3238
rect 10932 3236 10988 3238
rect 11012 3236 11068 3238
rect 11092 3236 11148 3238
rect 11978 9288 12034 9344
rect 11886 5480 11942 5536
rect 12622 12300 12678 12336
rect 12622 12280 12624 12300
rect 12624 12280 12676 12300
rect 12676 12280 12678 12300
rect 12162 9968 12218 10024
rect 12622 10376 12678 10432
rect 12806 11192 12862 11248
rect 12622 9832 12678 9888
rect 12530 9288 12586 9344
rect 12162 8744 12218 8800
rect 12162 8336 12218 8392
rect 12530 8880 12586 8936
rect 12162 6840 12218 6896
rect 12254 5888 12310 5944
rect 11518 2896 11574 2952
rect 12530 6296 12586 6352
rect 12162 3596 12218 3632
rect 12162 3576 12164 3596
rect 12164 3576 12216 3596
rect 12216 3576 12218 3596
rect 12622 4664 12678 4720
rect 12346 3032 12402 3088
rect 12622 3032 12678 3088
rect 10852 2202 10908 2204
rect 10932 2202 10988 2204
rect 11012 2202 11068 2204
rect 11092 2202 11148 2204
rect 10852 2150 10878 2202
rect 10878 2150 10908 2202
rect 10932 2150 10942 2202
rect 10942 2150 10988 2202
rect 11012 2150 11058 2202
rect 11058 2150 11068 2202
rect 11092 2150 11122 2202
rect 11122 2150 11148 2202
rect 10852 2148 10908 2150
rect 10932 2148 10988 2150
rect 11012 2148 11068 2150
rect 11092 2148 11148 2150
rect 11702 856 11758 912
rect 12898 10512 12954 10568
rect 14150 13626 14206 13628
rect 14230 13626 14286 13628
rect 14310 13626 14366 13628
rect 14390 13626 14446 13628
rect 14150 13574 14176 13626
rect 14176 13574 14206 13626
rect 14230 13574 14240 13626
rect 14240 13574 14286 13626
rect 14310 13574 14356 13626
rect 14356 13574 14366 13626
rect 14390 13574 14420 13626
rect 14420 13574 14446 13626
rect 14150 13572 14206 13574
rect 14230 13572 14286 13574
rect 14310 13572 14366 13574
rect 14390 13572 14446 13574
rect 12806 5772 12862 5808
rect 12806 5752 12808 5772
rect 12808 5752 12860 5772
rect 12860 5752 12862 5772
rect 13542 12416 13598 12472
rect 13082 9560 13138 9616
rect 14150 12538 14206 12540
rect 14230 12538 14286 12540
rect 14310 12538 14366 12540
rect 14390 12538 14446 12540
rect 14150 12486 14176 12538
rect 14176 12486 14206 12538
rect 14230 12486 14240 12538
rect 14240 12486 14286 12538
rect 14310 12486 14356 12538
rect 14356 12486 14366 12538
rect 14390 12486 14420 12538
rect 14420 12486 14446 12538
rect 14150 12484 14206 12486
rect 14230 12484 14286 12486
rect 14310 12484 14366 12486
rect 14390 12484 14446 12486
rect 14094 11892 14150 11928
rect 14094 11872 14096 11892
rect 14096 11872 14148 11892
rect 14148 11872 14150 11892
rect 14646 12688 14702 12744
rect 14738 12552 14794 12608
rect 14150 11450 14206 11452
rect 14230 11450 14286 11452
rect 14310 11450 14366 11452
rect 14390 11450 14446 11452
rect 14150 11398 14176 11450
rect 14176 11398 14206 11450
rect 14230 11398 14240 11450
rect 14240 11398 14286 11450
rect 14310 11398 14356 11450
rect 14356 11398 14366 11450
rect 14390 11398 14420 11450
rect 14420 11398 14446 11450
rect 14150 11396 14206 11398
rect 14230 11396 14286 11398
rect 14310 11396 14366 11398
rect 14390 11396 14446 11398
rect 14150 10362 14206 10364
rect 14230 10362 14286 10364
rect 14310 10362 14366 10364
rect 14390 10362 14446 10364
rect 14150 10310 14176 10362
rect 14176 10310 14206 10362
rect 14230 10310 14240 10362
rect 14240 10310 14286 10362
rect 14310 10310 14356 10362
rect 14356 10310 14366 10362
rect 14390 10310 14420 10362
rect 14420 10310 14446 10362
rect 14150 10308 14206 10310
rect 14230 10308 14286 10310
rect 14310 10308 14366 10310
rect 14390 10308 14446 10310
rect 14646 10648 14702 10704
rect 14150 9274 14206 9276
rect 14230 9274 14286 9276
rect 14310 9274 14366 9276
rect 14390 9274 14446 9276
rect 14150 9222 14176 9274
rect 14176 9222 14206 9274
rect 14230 9222 14240 9274
rect 14240 9222 14286 9274
rect 14310 9222 14356 9274
rect 14356 9222 14366 9274
rect 14390 9222 14420 9274
rect 14420 9222 14446 9274
rect 14150 9220 14206 9222
rect 14230 9220 14286 9222
rect 14310 9220 14366 9222
rect 14390 9220 14446 9222
rect 14186 8744 14242 8800
rect 14370 8780 14372 8800
rect 14372 8780 14424 8800
rect 14424 8780 14426 8800
rect 14370 8744 14426 8780
rect 13634 8236 13636 8256
rect 13636 8236 13688 8256
rect 13688 8236 13690 8256
rect 13634 8200 13690 8236
rect 12990 5752 13046 5808
rect 14922 11056 14978 11112
rect 15290 18400 15346 18456
rect 15474 16360 15530 16416
rect 15750 15816 15806 15872
rect 15566 13640 15622 13696
rect 15382 11736 15438 11792
rect 14830 9696 14886 9752
rect 14830 9152 14886 9208
rect 15658 12960 15714 13016
rect 15658 12416 15714 12472
rect 15566 12144 15622 12200
rect 14150 8186 14206 8188
rect 14230 8186 14286 8188
rect 14310 8186 14366 8188
rect 14390 8186 14446 8188
rect 14150 8134 14176 8186
rect 14176 8134 14206 8186
rect 14230 8134 14240 8186
rect 14240 8134 14286 8186
rect 14310 8134 14356 8186
rect 14356 8134 14366 8186
rect 14390 8134 14420 8186
rect 14420 8134 14446 8186
rect 14150 8132 14206 8134
rect 14230 8132 14286 8134
rect 14310 8132 14366 8134
rect 14390 8132 14446 8134
rect 14002 7656 14058 7712
rect 14150 7098 14206 7100
rect 14230 7098 14286 7100
rect 14310 7098 14366 7100
rect 14390 7098 14446 7100
rect 14150 7046 14176 7098
rect 14176 7046 14206 7098
rect 14230 7046 14240 7098
rect 14240 7046 14286 7098
rect 14310 7046 14356 7098
rect 14356 7046 14366 7098
rect 14390 7046 14420 7098
rect 14420 7046 14446 7098
rect 14150 7044 14206 7046
rect 14230 7044 14286 7046
rect 14310 7044 14366 7046
rect 14390 7044 14446 7046
rect 14738 6840 14794 6896
rect 15014 6704 15070 6760
rect 14150 6010 14206 6012
rect 14230 6010 14286 6012
rect 14310 6010 14366 6012
rect 14390 6010 14446 6012
rect 14150 5958 14176 6010
rect 14176 5958 14206 6010
rect 14230 5958 14240 6010
rect 14240 5958 14286 6010
rect 14310 5958 14356 6010
rect 14356 5958 14366 6010
rect 14390 5958 14420 6010
rect 14420 5958 14446 6010
rect 14150 5956 14206 5958
rect 14230 5956 14286 5958
rect 14310 5956 14366 5958
rect 14390 5956 14446 5958
rect 15014 6160 15070 6216
rect 14002 5480 14058 5536
rect 14150 4922 14206 4924
rect 14230 4922 14286 4924
rect 14310 4922 14366 4924
rect 14390 4922 14446 4924
rect 14150 4870 14176 4922
rect 14176 4870 14206 4922
rect 14230 4870 14240 4922
rect 14240 4870 14286 4922
rect 14310 4870 14356 4922
rect 14356 4870 14366 4922
rect 14390 4870 14420 4922
rect 14420 4870 14446 4922
rect 14150 4868 14206 4870
rect 14230 4868 14286 4870
rect 14310 4868 14366 4870
rect 14390 4868 14446 4870
rect 13174 3576 13230 3632
rect 12990 3476 12992 3496
rect 12992 3476 13044 3496
rect 13044 3476 13046 3496
rect 12990 3440 13046 3476
rect 14150 3834 14206 3836
rect 14230 3834 14286 3836
rect 14310 3834 14366 3836
rect 14390 3834 14446 3836
rect 14150 3782 14176 3834
rect 14176 3782 14206 3834
rect 14230 3782 14240 3834
rect 14240 3782 14286 3834
rect 14310 3782 14356 3834
rect 14356 3782 14366 3834
rect 14390 3782 14420 3834
rect 14420 3782 14446 3834
rect 14150 3780 14206 3782
rect 14230 3780 14286 3782
rect 14310 3780 14366 3782
rect 14390 3780 14446 3782
rect 14554 3576 14610 3632
rect 15658 9288 15714 9344
rect 15658 8880 15714 8936
rect 16026 13912 16082 13968
rect 16118 13368 16174 13424
rect 16118 12824 16174 12880
rect 15934 11192 15990 11248
rect 15934 8880 15990 8936
rect 16578 20984 16634 21040
rect 17866 19624 17922 19680
rect 17449 19610 17505 19612
rect 17529 19610 17585 19612
rect 17609 19610 17665 19612
rect 17689 19610 17745 19612
rect 17449 19558 17475 19610
rect 17475 19558 17505 19610
rect 17529 19558 17539 19610
rect 17539 19558 17585 19610
rect 17609 19558 17655 19610
rect 17655 19558 17665 19610
rect 17689 19558 17719 19610
rect 17719 19558 17745 19610
rect 17449 19556 17505 19558
rect 17529 19556 17585 19558
rect 17609 19556 17665 19558
rect 17689 19556 17745 19558
rect 16578 14320 16634 14376
rect 16486 13368 16542 13424
rect 17774 18944 17830 19000
rect 17314 18536 17370 18592
rect 17222 18400 17278 18456
rect 17449 18522 17505 18524
rect 17529 18522 17585 18524
rect 17609 18522 17665 18524
rect 17689 18522 17745 18524
rect 17449 18470 17475 18522
rect 17475 18470 17505 18522
rect 17529 18470 17539 18522
rect 17539 18470 17585 18522
rect 17609 18470 17655 18522
rect 17655 18470 17665 18522
rect 17689 18470 17719 18522
rect 17719 18470 17745 18522
rect 17449 18468 17505 18470
rect 17529 18468 17585 18470
rect 17609 18468 17665 18470
rect 17689 18468 17745 18470
rect 17038 18128 17094 18184
rect 17774 17740 17830 17776
rect 17774 17720 17776 17740
rect 17776 17720 17828 17740
rect 17828 17720 17830 17740
rect 17774 17584 17830 17640
rect 17449 17434 17505 17436
rect 17529 17434 17585 17436
rect 17609 17434 17665 17436
rect 17689 17434 17745 17436
rect 17449 17382 17475 17434
rect 17475 17382 17505 17434
rect 17529 17382 17539 17434
rect 17539 17382 17585 17434
rect 17609 17382 17655 17434
rect 17655 17382 17665 17434
rect 17689 17382 17719 17434
rect 17719 17382 17745 17434
rect 17449 17380 17505 17382
rect 17529 17380 17585 17382
rect 17609 17380 17665 17382
rect 17689 17380 17745 17382
rect 17449 16346 17505 16348
rect 17529 16346 17585 16348
rect 17609 16346 17665 16348
rect 17689 16346 17745 16348
rect 17449 16294 17475 16346
rect 17475 16294 17505 16346
rect 17529 16294 17539 16346
rect 17539 16294 17585 16346
rect 17609 16294 17655 16346
rect 17655 16294 17665 16346
rect 17689 16294 17719 16346
rect 17719 16294 17745 16346
rect 17449 16292 17505 16294
rect 17529 16292 17585 16294
rect 17609 16292 17665 16294
rect 17689 16292 17745 16294
rect 17449 15258 17505 15260
rect 17529 15258 17585 15260
rect 17609 15258 17665 15260
rect 17689 15258 17745 15260
rect 17449 15206 17475 15258
rect 17475 15206 17505 15258
rect 17529 15206 17539 15258
rect 17539 15206 17585 15258
rect 17609 15206 17655 15258
rect 17655 15206 17665 15258
rect 17689 15206 17719 15258
rect 17719 15206 17745 15258
rect 17449 15204 17505 15206
rect 17529 15204 17585 15206
rect 17609 15204 17665 15206
rect 17689 15204 17745 15206
rect 17449 14170 17505 14172
rect 17529 14170 17585 14172
rect 17609 14170 17665 14172
rect 17689 14170 17745 14172
rect 17449 14118 17475 14170
rect 17475 14118 17505 14170
rect 17529 14118 17539 14170
rect 17539 14118 17585 14170
rect 17609 14118 17655 14170
rect 17655 14118 17665 14170
rect 17689 14118 17719 14170
rect 17719 14118 17745 14170
rect 17449 14116 17505 14118
rect 17529 14116 17585 14118
rect 17609 14116 17665 14118
rect 17689 14116 17745 14118
rect 17498 13932 17554 13968
rect 17498 13912 17500 13932
rect 17500 13912 17552 13932
rect 17552 13912 17554 13932
rect 17222 12960 17278 13016
rect 16762 12280 16818 12336
rect 16670 12044 16672 12064
rect 16672 12044 16724 12064
rect 16724 12044 16726 12064
rect 16670 12008 16726 12044
rect 16670 11892 16726 11928
rect 16670 11872 16672 11892
rect 16672 11872 16724 11892
rect 16724 11872 16726 11892
rect 16946 12008 17002 12064
rect 17449 13082 17505 13084
rect 17529 13082 17585 13084
rect 17609 13082 17665 13084
rect 17689 13082 17745 13084
rect 17449 13030 17475 13082
rect 17475 13030 17505 13082
rect 17529 13030 17539 13082
rect 17539 13030 17585 13082
rect 17609 13030 17655 13082
rect 17655 13030 17665 13082
rect 17689 13030 17719 13082
rect 17719 13030 17745 13082
rect 17449 13028 17505 13030
rect 17529 13028 17585 13030
rect 17609 13028 17665 13030
rect 17689 13028 17745 13030
rect 17222 12280 17278 12336
rect 17774 12416 17830 12472
rect 17958 17856 18014 17912
rect 18602 18672 18658 18728
rect 18694 17992 18750 18048
rect 18050 17720 18106 17776
rect 18878 16088 18934 16144
rect 19798 19352 19854 19408
rect 19154 18264 19210 18320
rect 19062 17040 19118 17096
rect 20442 19216 20498 19272
rect 18142 12688 18198 12744
rect 16486 9288 16542 9344
rect 15750 8200 15806 8256
rect 15566 6160 15622 6216
rect 15750 6160 15806 6216
rect 15934 5772 15990 5808
rect 15934 5752 15936 5772
rect 15936 5752 15988 5772
rect 15988 5752 15990 5772
rect 15934 5616 15990 5672
rect 14150 2746 14206 2748
rect 14230 2746 14286 2748
rect 14310 2746 14366 2748
rect 14390 2746 14446 2748
rect 14150 2694 14176 2746
rect 14176 2694 14206 2746
rect 14230 2694 14240 2746
rect 14240 2694 14286 2746
rect 14310 2694 14356 2746
rect 14356 2694 14366 2746
rect 14390 2694 14420 2746
rect 14420 2694 14446 2746
rect 14150 2692 14206 2694
rect 14230 2692 14286 2694
rect 14310 2692 14366 2694
rect 14390 2692 14446 2694
rect 16394 7656 16450 7712
rect 15658 2916 15714 2952
rect 15658 2896 15660 2916
rect 15660 2896 15712 2916
rect 15712 2896 15714 2916
rect 16946 11056 17002 11112
rect 16670 10412 16672 10432
rect 16672 10412 16724 10432
rect 16724 10412 16726 10432
rect 16670 10376 16726 10412
rect 16670 9560 16726 9616
rect 17038 10260 17094 10296
rect 17498 12144 17554 12200
rect 17449 11994 17505 11996
rect 17529 11994 17585 11996
rect 17609 11994 17665 11996
rect 17689 11994 17745 11996
rect 17449 11942 17475 11994
rect 17475 11942 17505 11994
rect 17529 11942 17539 11994
rect 17539 11942 17585 11994
rect 17609 11942 17655 11994
rect 17655 11942 17665 11994
rect 17689 11942 17719 11994
rect 17719 11942 17745 11994
rect 17449 11940 17505 11942
rect 17529 11940 17585 11942
rect 17609 11940 17665 11942
rect 17689 11940 17745 11942
rect 17866 10920 17922 10976
rect 17449 10906 17505 10908
rect 17529 10906 17585 10908
rect 17609 10906 17665 10908
rect 17689 10906 17745 10908
rect 17449 10854 17475 10906
rect 17475 10854 17505 10906
rect 17529 10854 17539 10906
rect 17539 10854 17585 10906
rect 17609 10854 17655 10906
rect 17655 10854 17665 10906
rect 17689 10854 17719 10906
rect 17719 10854 17745 10906
rect 17449 10852 17505 10854
rect 17529 10852 17585 10854
rect 17609 10852 17665 10854
rect 17689 10852 17745 10854
rect 17038 10240 17040 10260
rect 17040 10240 17092 10260
rect 17092 10240 17094 10260
rect 16670 9288 16726 9344
rect 16762 8744 16818 8800
rect 16670 8608 16726 8664
rect 17498 10376 17554 10432
rect 17449 9818 17505 9820
rect 17529 9818 17585 9820
rect 17609 9818 17665 9820
rect 17689 9818 17745 9820
rect 17449 9766 17475 9818
rect 17475 9766 17505 9818
rect 17529 9766 17539 9818
rect 17539 9766 17585 9818
rect 17609 9766 17655 9818
rect 17655 9766 17665 9818
rect 17689 9766 17719 9818
rect 17719 9766 17745 9818
rect 17449 9764 17505 9766
rect 17529 9764 17585 9766
rect 17609 9764 17665 9766
rect 17689 9764 17745 9766
rect 17314 9152 17370 9208
rect 18050 10104 18106 10160
rect 17449 8730 17505 8732
rect 17529 8730 17585 8732
rect 17609 8730 17665 8732
rect 17689 8730 17745 8732
rect 17449 8678 17475 8730
rect 17475 8678 17505 8730
rect 17529 8678 17539 8730
rect 17539 8678 17585 8730
rect 17609 8678 17655 8730
rect 17655 8678 17665 8730
rect 17689 8678 17719 8730
rect 17719 8678 17745 8730
rect 17449 8676 17505 8678
rect 17529 8676 17585 8678
rect 17609 8676 17665 8678
rect 17689 8676 17745 8678
rect 17314 8200 17370 8256
rect 17038 7948 17094 7984
rect 17038 7928 17040 7948
rect 17040 7928 17092 7948
rect 17092 7928 17094 7948
rect 17130 7520 17186 7576
rect 17449 7642 17505 7644
rect 17529 7642 17585 7644
rect 17609 7642 17665 7644
rect 17689 7642 17745 7644
rect 17449 7590 17475 7642
rect 17475 7590 17505 7642
rect 17529 7590 17539 7642
rect 17539 7590 17585 7642
rect 17609 7590 17655 7642
rect 17655 7590 17665 7642
rect 17689 7590 17719 7642
rect 17719 7590 17745 7642
rect 17449 7588 17505 7590
rect 17529 7588 17585 7590
rect 17609 7588 17665 7590
rect 17689 7588 17745 7590
rect 16946 6840 17002 6896
rect 17449 6554 17505 6556
rect 17529 6554 17585 6556
rect 17609 6554 17665 6556
rect 17689 6554 17745 6556
rect 17449 6502 17475 6554
rect 17475 6502 17505 6554
rect 17529 6502 17539 6554
rect 17539 6502 17585 6554
rect 17609 6502 17655 6554
rect 17655 6502 17665 6554
rect 17689 6502 17719 6554
rect 17719 6502 17745 6554
rect 17449 6500 17505 6502
rect 17529 6500 17585 6502
rect 17609 6500 17665 6502
rect 17689 6500 17745 6502
rect 17449 5466 17505 5468
rect 17529 5466 17585 5468
rect 17609 5466 17665 5468
rect 17689 5466 17745 5468
rect 17449 5414 17475 5466
rect 17475 5414 17505 5466
rect 17529 5414 17539 5466
rect 17539 5414 17585 5466
rect 17609 5414 17655 5466
rect 17655 5414 17665 5466
rect 17689 5414 17719 5466
rect 17719 5414 17745 5466
rect 17449 5412 17505 5414
rect 17529 5412 17585 5414
rect 17609 5412 17665 5414
rect 17689 5412 17745 5414
rect 16946 4528 17002 4584
rect 16854 3576 16910 3632
rect 17449 4378 17505 4380
rect 17529 4378 17585 4380
rect 17609 4378 17665 4380
rect 17689 4378 17745 4380
rect 17449 4326 17475 4378
rect 17475 4326 17505 4378
rect 17529 4326 17539 4378
rect 17539 4326 17585 4378
rect 17609 4326 17655 4378
rect 17655 4326 17665 4378
rect 17689 4326 17719 4378
rect 17719 4326 17745 4378
rect 17449 4324 17505 4326
rect 17529 4324 17585 4326
rect 17609 4324 17665 4326
rect 17689 4324 17745 4326
rect 17449 3290 17505 3292
rect 17529 3290 17585 3292
rect 17609 3290 17665 3292
rect 17689 3290 17745 3292
rect 17449 3238 17475 3290
rect 17475 3238 17505 3290
rect 17529 3238 17539 3290
rect 17539 3238 17585 3290
rect 17609 3238 17655 3290
rect 17655 3238 17665 3290
rect 17689 3238 17719 3290
rect 17719 3238 17745 3290
rect 17449 3236 17505 3238
rect 17529 3236 17585 3238
rect 17609 3236 17665 3238
rect 17689 3236 17745 3238
rect 18510 12588 18512 12608
rect 18512 12588 18564 12608
rect 18564 12588 18566 12608
rect 18510 12552 18566 12588
rect 18418 12416 18474 12472
rect 18418 9424 18474 9480
rect 18050 6724 18106 6760
rect 18050 6704 18052 6724
rect 18052 6704 18104 6724
rect 18104 6704 18106 6724
rect 18326 7928 18382 7984
rect 18234 7384 18290 7440
rect 18418 6296 18474 6352
rect 18142 6160 18198 6216
rect 17866 2896 17922 2952
rect 18142 4684 18198 4720
rect 18142 4664 18144 4684
rect 18144 4664 18196 4684
rect 18196 4664 18198 4684
rect 18786 9016 18842 9072
rect 20166 16224 20222 16280
rect 20074 15564 20130 15600
rect 20074 15544 20076 15564
rect 20076 15544 20128 15564
rect 20128 15544 20130 15564
rect 20350 16904 20406 16960
rect 20258 15000 20314 15056
rect 19430 11736 19486 11792
rect 19154 9288 19210 9344
rect 18786 6976 18842 7032
rect 19706 9288 19762 9344
rect 19430 8472 19486 8528
rect 19890 8064 19946 8120
rect 19430 7792 19486 7848
rect 19246 7656 19302 7712
rect 20166 8200 20222 8256
rect 20074 7248 20130 7304
rect 19982 6296 20038 6352
rect 20258 4936 20314 4992
rect 20994 18300 20996 18320
rect 20996 18300 21048 18320
rect 21048 18300 21050 18320
rect 20994 18264 21050 18300
rect 20994 8336 21050 8392
rect 18418 2216 18474 2272
rect 17449 2202 17505 2204
rect 17529 2202 17585 2204
rect 17609 2202 17665 2204
rect 17689 2202 17745 2204
rect 17449 2150 17475 2202
rect 17475 2150 17505 2202
rect 17529 2150 17539 2202
rect 17539 2150 17585 2202
rect 17609 2150 17655 2202
rect 17655 2150 17665 2202
rect 17689 2150 17719 2202
rect 17719 2150 17745 2202
rect 17449 2148 17505 2150
rect 17529 2148 17585 2150
rect 17609 2148 17665 2150
rect 17689 2148 17745 2150
rect 16578 856 16634 912
rect 20994 5616 21050 5672
rect 20718 1536 20774 1592
rect 20534 312 20590 368
<< metal3 >>
rect 16389 21722 16455 21725
rect 21520 21722 22000 21752
rect 16389 21720 22000 21722
rect 16389 21664 16394 21720
rect 16450 21664 22000 21720
rect 16389 21662 22000 21664
rect 16389 21659 16455 21662
rect 21520 21632 22000 21662
rect 16573 21042 16639 21045
rect 21520 21042 22000 21072
rect 16573 21040 22000 21042
rect 16573 20984 16578 21040
rect 16634 20984 22000 21040
rect 16573 20982 22000 20984
rect 16573 20979 16639 20982
rect 21520 20952 22000 20982
rect 15929 20362 15995 20365
rect 21520 20362 22000 20392
rect 15929 20360 22000 20362
rect 15929 20304 15934 20360
rect 15990 20304 22000 20360
rect 15929 20302 22000 20304
rect 15929 20299 15995 20302
rect 21520 20272 22000 20302
rect 17861 19682 17927 19685
rect 21520 19682 22000 19712
rect 17861 19680 22000 19682
rect 17861 19624 17866 19680
rect 17922 19624 22000 19680
rect 17861 19622 22000 19624
rect 17861 19619 17927 19622
rect 4242 19616 4562 19617
rect 4242 19552 4250 19616
rect 4314 19552 4330 19616
rect 4394 19552 4410 19616
rect 4474 19552 4490 19616
rect 4554 19552 4562 19616
rect 4242 19551 4562 19552
rect 10840 19616 11160 19617
rect 10840 19552 10848 19616
rect 10912 19552 10928 19616
rect 10992 19552 11008 19616
rect 11072 19552 11088 19616
rect 11152 19552 11160 19616
rect 10840 19551 11160 19552
rect 17437 19616 17757 19617
rect 17437 19552 17445 19616
rect 17509 19552 17525 19616
rect 17589 19552 17605 19616
rect 17669 19552 17685 19616
rect 17749 19552 17757 19616
rect 21520 19592 22000 19622
rect 17437 19551 17757 19552
rect 10869 19410 10935 19413
rect 12249 19410 12315 19413
rect 10869 19408 12315 19410
rect 10869 19352 10874 19408
rect 10930 19352 12254 19408
rect 12310 19352 12315 19408
rect 10869 19350 12315 19352
rect 10869 19347 10935 19350
rect 12249 19347 12315 19350
rect 13905 19410 13971 19413
rect 19793 19410 19859 19413
rect 13905 19408 19859 19410
rect 13905 19352 13910 19408
rect 13966 19352 19798 19408
rect 19854 19352 19859 19408
rect 13905 19350 19859 19352
rect 13905 19347 13971 19350
rect 19793 19347 19859 19350
rect 5441 19274 5507 19277
rect 8293 19274 8359 19277
rect 14181 19274 14247 19277
rect 20437 19274 20503 19277
rect 5441 19272 8359 19274
rect 5441 19216 5446 19272
rect 5502 19216 8298 19272
rect 8354 19216 8359 19272
rect 5441 19214 8359 19216
rect 5441 19211 5507 19214
rect 8293 19211 8359 19214
rect 13862 19272 20503 19274
rect 13862 19216 14186 19272
rect 14242 19216 20442 19272
rect 20498 19216 20503 19272
rect 13862 19214 20503 19216
rect 3969 19138 4035 19141
rect 4797 19138 4863 19141
rect 3969 19136 4863 19138
rect 3969 19080 3974 19136
rect 4030 19080 4802 19136
rect 4858 19080 4863 19136
rect 3969 19078 4863 19080
rect 3969 19075 4035 19078
rect 4797 19075 4863 19078
rect 11973 19138 12039 19141
rect 12801 19138 12867 19141
rect 11973 19136 12867 19138
rect 11973 19080 11978 19136
rect 12034 19080 12806 19136
rect 12862 19080 12867 19136
rect 11973 19078 12867 19080
rect 11973 19075 12039 19078
rect 12801 19075 12867 19078
rect 7541 19072 7861 19073
rect 7541 19008 7549 19072
rect 7613 19008 7629 19072
rect 7693 19008 7709 19072
rect 7773 19008 7789 19072
rect 7853 19008 7861 19072
rect 7541 19007 7861 19008
rect 2405 19002 2471 19005
rect 5257 19002 5323 19005
rect 2405 19000 5323 19002
rect 2405 18944 2410 19000
rect 2466 18944 5262 19000
rect 5318 18944 5323 19000
rect 2405 18942 5323 18944
rect 2405 18939 2471 18942
rect 5257 18939 5323 18942
rect 10317 19002 10383 19005
rect 13261 19002 13327 19005
rect 10317 19000 13327 19002
rect 10317 18944 10322 19000
rect 10378 18944 13266 19000
rect 13322 18944 13327 19000
rect 10317 18942 13327 18944
rect 10317 18939 10383 18942
rect 13261 18939 13327 18942
rect 3601 18866 3667 18869
rect 13862 18866 13922 19214
rect 14181 19211 14247 19214
rect 20437 19211 20503 19214
rect 14138 19072 14458 19073
rect 14138 19008 14146 19072
rect 14210 19008 14226 19072
rect 14290 19008 14306 19072
rect 14370 19008 14386 19072
rect 14450 19008 14458 19072
rect 14138 19007 14458 19008
rect 17769 19002 17835 19005
rect 21520 19002 22000 19032
rect 17769 19000 22000 19002
rect 17769 18944 17774 19000
rect 17830 18944 22000 19000
rect 17769 18942 22000 18944
rect 17769 18939 17835 18942
rect 21520 18912 22000 18942
rect 3601 18864 13922 18866
rect 3601 18808 3606 18864
rect 3662 18808 13922 18864
rect 3601 18806 13922 18808
rect 3601 18803 3667 18806
rect 12249 18730 12315 18733
rect 18597 18730 18663 18733
rect 12249 18728 18663 18730
rect 12249 18672 12254 18728
rect 12310 18672 18602 18728
rect 18658 18672 18663 18728
rect 12249 18670 18663 18672
rect 12249 18667 12315 18670
rect 18597 18667 18663 18670
rect 14273 18594 14339 18597
rect 17309 18594 17375 18597
rect 14273 18592 17375 18594
rect 14273 18536 14278 18592
rect 14334 18536 17314 18592
rect 17370 18536 17375 18592
rect 14273 18534 17375 18536
rect 14273 18531 14339 18534
rect 17309 18531 17375 18534
rect 4242 18528 4562 18529
rect 0 18368 480 18488
rect 4242 18464 4250 18528
rect 4314 18464 4330 18528
rect 4394 18464 4410 18528
rect 4474 18464 4490 18528
rect 4554 18464 4562 18528
rect 4242 18463 4562 18464
rect 10840 18528 11160 18529
rect 10840 18464 10848 18528
rect 10912 18464 10928 18528
rect 10992 18464 11008 18528
rect 11072 18464 11088 18528
rect 11152 18464 11160 18528
rect 10840 18463 11160 18464
rect 17437 18528 17757 18529
rect 17437 18464 17445 18528
rect 17509 18464 17525 18528
rect 17589 18464 17605 18528
rect 17669 18464 17685 18528
rect 17749 18464 17757 18528
rect 17437 18463 17757 18464
rect 13261 18458 13327 18461
rect 14365 18458 14431 18461
rect 15285 18458 15351 18461
rect 17217 18458 17283 18461
rect 13261 18456 14980 18458
rect 13261 18400 13266 18456
rect 13322 18400 14370 18456
rect 14426 18400 14980 18456
rect 13261 18398 14980 18400
rect 13261 18395 13327 18398
rect 14365 18395 14431 18398
rect 10869 18322 10935 18325
rect 14733 18322 14799 18325
rect 10869 18320 14799 18322
rect 10869 18264 10874 18320
rect 10930 18264 14738 18320
rect 14794 18264 14799 18320
rect 10869 18262 14799 18264
rect 14920 18322 14980 18398
rect 15285 18456 17283 18458
rect 15285 18400 15290 18456
rect 15346 18400 17222 18456
rect 17278 18400 17283 18456
rect 15285 18398 17283 18400
rect 15285 18395 15351 18398
rect 17217 18395 17283 18398
rect 19149 18322 19215 18325
rect 14920 18320 19215 18322
rect 14920 18264 19154 18320
rect 19210 18264 19215 18320
rect 14920 18262 19215 18264
rect 10869 18259 10935 18262
rect 14733 18259 14799 18262
rect 19149 18259 19215 18262
rect 20989 18322 21055 18325
rect 21520 18322 22000 18352
rect 20989 18320 22000 18322
rect 20989 18264 20994 18320
rect 21050 18264 22000 18320
rect 20989 18262 22000 18264
rect 20989 18259 21055 18262
rect 21520 18232 22000 18262
rect 6821 18186 6887 18189
rect 17033 18186 17099 18189
rect 6821 18184 17099 18186
rect 6821 18128 6826 18184
rect 6882 18128 17038 18184
rect 17094 18128 17099 18184
rect 6821 18126 17099 18128
rect 6821 18123 6887 18126
rect 17033 18123 17099 18126
rect 10409 18050 10475 18053
rect 12157 18050 12223 18053
rect 10409 18048 12223 18050
rect 10409 17992 10414 18048
rect 10470 17992 12162 18048
rect 12218 17992 12223 18048
rect 10409 17990 12223 17992
rect 10409 17987 10475 17990
rect 12157 17987 12223 17990
rect 14958 17988 14964 18052
rect 15028 18050 15034 18052
rect 18689 18050 18755 18053
rect 15028 18048 18755 18050
rect 15028 17992 18694 18048
rect 18750 17992 18755 18048
rect 15028 17990 18755 17992
rect 15028 17988 15034 17990
rect 18689 17987 18755 17990
rect 7541 17984 7861 17985
rect 7541 17920 7549 17984
rect 7613 17920 7629 17984
rect 7693 17920 7709 17984
rect 7773 17920 7789 17984
rect 7853 17920 7861 17984
rect 7541 17919 7861 17920
rect 14138 17984 14458 17985
rect 14138 17920 14146 17984
rect 14210 17920 14226 17984
rect 14290 17920 14306 17984
rect 14370 17920 14386 17984
rect 14450 17920 14458 17984
rect 14138 17919 14458 17920
rect 3417 17914 3483 17917
rect 4797 17914 4863 17917
rect 17953 17914 18019 17917
rect 3417 17912 4863 17914
rect 3417 17856 3422 17912
rect 3478 17856 4802 17912
rect 4858 17856 4863 17912
rect 3417 17854 4863 17856
rect 3417 17851 3483 17854
rect 4797 17851 4863 17854
rect 15150 17912 18019 17914
rect 15150 17856 17958 17912
rect 18014 17856 18019 17912
rect 15150 17854 18019 17856
rect 1301 17778 1367 17781
rect 7465 17778 7531 17781
rect 1301 17776 8954 17778
rect 1301 17720 1306 17776
rect 1362 17720 7470 17776
rect 7526 17720 8954 17776
rect 1301 17718 8954 17720
rect 1301 17715 1367 17718
rect 7465 17715 7531 17718
rect 5901 17642 5967 17645
rect 8661 17642 8727 17645
rect 5901 17640 8727 17642
rect 5901 17584 5906 17640
rect 5962 17584 8666 17640
rect 8722 17584 8727 17640
rect 5901 17582 8727 17584
rect 8894 17642 8954 17718
rect 15150 17642 15210 17854
rect 17953 17851 18019 17854
rect 17769 17778 17835 17781
rect 18045 17778 18111 17781
rect 17769 17776 18111 17778
rect 17769 17720 17774 17776
rect 17830 17720 18050 17776
rect 18106 17720 18111 17776
rect 17769 17718 18111 17720
rect 17769 17715 17835 17718
rect 18045 17715 18111 17718
rect 8894 17582 15210 17642
rect 17769 17642 17835 17645
rect 21520 17642 22000 17672
rect 17769 17640 22000 17642
rect 17769 17584 17774 17640
rect 17830 17584 22000 17640
rect 17769 17582 22000 17584
rect 5901 17579 5967 17582
rect 8661 17579 8727 17582
rect 17769 17579 17835 17582
rect 21520 17552 22000 17582
rect 4242 17440 4562 17441
rect 4242 17376 4250 17440
rect 4314 17376 4330 17440
rect 4394 17376 4410 17440
rect 4474 17376 4490 17440
rect 4554 17376 4562 17440
rect 4242 17375 4562 17376
rect 10840 17440 11160 17441
rect 10840 17376 10848 17440
rect 10912 17376 10928 17440
rect 10992 17376 11008 17440
rect 11072 17376 11088 17440
rect 11152 17376 11160 17440
rect 10840 17375 11160 17376
rect 17437 17440 17757 17441
rect 17437 17376 17445 17440
rect 17509 17376 17525 17440
rect 17589 17376 17605 17440
rect 17669 17376 17685 17440
rect 17749 17376 17757 17440
rect 17437 17375 17757 17376
rect 3969 17234 4035 17237
rect 11237 17234 11303 17237
rect 12249 17234 12315 17237
rect 3969 17232 12315 17234
rect 3969 17176 3974 17232
rect 4030 17176 11242 17232
rect 11298 17176 12254 17232
rect 12310 17176 12315 17232
rect 3969 17174 12315 17176
rect 3969 17171 4035 17174
rect 11237 17171 11303 17174
rect 12249 17171 12315 17174
rect 3693 17098 3759 17101
rect 19057 17098 19123 17101
rect 3693 17096 19123 17098
rect 3693 17040 3698 17096
rect 3754 17040 19062 17096
rect 19118 17040 19123 17096
rect 3693 17038 19123 17040
rect 3693 17035 3759 17038
rect 19057 17035 19123 17038
rect 11421 16962 11487 16965
rect 12709 16962 12775 16965
rect 13169 16962 13235 16965
rect 11421 16960 13235 16962
rect 11421 16904 11426 16960
rect 11482 16904 12714 16960
rect 12770 16904 13174 16960
rect 13230 16904 13235 16960
rect 11421 16902 13235 16904
rect 11421 16899 11487 16902
rect 12709 16899 12775 16902
rect 13169 16899 13235 16902
rect 20345 16962 20411 16965
rect 21520 16962 22000 16992
rect 20345 16960 22000 16962
rect 20345 16904 20350 16960
rect 20406 16904 22000 16960
rect 20345 16902 22000 16904
rect 20345 16899 20411 16902
rect 7541 16896 7861 16897
rect 7541 16832 7549 16896
rect 7613 16832 7629 16896
rect 7693 16832 7709 16896
rect 7773 16832 7789 16896
rect 7853 16832 7861 16896
rect 7541 16831 7861 16832
rect 14138 16896 14458 16897
rect 14138 16832 14146 16896
rect 14210 16832 14226 16896
rect 14290 16832 14306 16896
rect 14370 16832 14386 16896
rect 14450 16832 14458 16896
rect 21520 16872 22000 16902
rect 14138 16831 14458 16832
rect 2037 16690 2103 16693
rect 3417 16690 3483 16693
rect 2037 16688 3483 16690
rect 2037 16632 2042 16688
rect 2098 16632 3422 16688
rect 3478 16632 3483 16688
rect 2037 16630 3483 16632
rect 2037 16627 2103 16630
rect 3417 16627 3483 16630
rect 9213 16554 9279 16557
rect 14825 16554 14891 16557
rect 14958 16554 14964 16556
rect 9213 16552 14964 16554
rect 9213 16496 9218 16552
rect 9274 16496 14830 16552
rect 14886 16496 14964 16552
rect 9213 16494 14964 16496
rect 9213 16491 9279 16494
rect 14825 16491 14891 16494
rect 14958 16492 14964 16494
rect 15028 16492 15034 16556
rect 14549 16418 14615 16421
rect 15469 16418 15535 16421
rect 14549 16416 15535 16418
rect 14549 16360 14554 16416
rect 14610 16360 15474 16416
rect 15530 16360 15535 16416
rect 14549 16358 15535 16360
rect 14549 16355 14615 16358
rect 15469 16355 15535 16358
rect 4242 16352 4562 16353
rect 4242 16288 4250 16352
rect 4314 16288 4330 16352
rect 4394 16288 4410 16352
rect 4474 16288 4490 16352
rect 4554 16288 4562 16352
rect 4242 16287 4562 16288
rect 10840 16352 11160 16353
rect 10840 16288 10848 16352
rect 10912 16288 10928 16352
rect 10992 16288 11008 16352
rect 11072 16288 11088 16352
rect 11152 16288 11160 16352
rect 10840 16287 11160 16288
rect 17437 16352 17757 16353
rect 17437 16288 17445 16352
rect 17509 16288 17525 16352
rect 17589 16288 17605 16352
rect 17669 16288 17685 16352
rect 17749 16288 17757 16352
rect 17437 16287 17757 16288
rect 20161 16282 20227 16285
rect 21520 16282 22000 16312
rect 20161 16280 22000 16282
rect 20161 16224 20166 16280
rect 20222 16224 22000 16280
rect 20161 16222 22000 16224
rect 20161 16219 20227 16222
rect 21520 16192 22000 16222
rect 6545 16146 6611 16149
rect 12617 16146 12683 16149
rect 18873 16146 18939 16149
rect 6545 16144 12220 16146
rect 6545 16088 6550 16144
rect 6606 16088 12220 16144
rect 6545 16086 12220 16088
rect 6545 16083 6611 16086
rect 12160 16010 12220 16086
rect 12617 16144 18939 16146
rect 12617 16088 12622 16144
rect 12678 16088 18878 16144
rect 18934 16088 18939 16144
rect 12617 16086 18939 16088
rect 12617 16083 12683 16086
rect 14733 16010 14799 16013
rect 12160 16008 14799 16010
rect 12160 15952 14738 16008
rect 14794 15952 14799 16008
rect 12160 15950 14799 15952
rect 14733 15947 14799 15950
rect 15702 15877 15762 16086
rect 18873 16083 18939 16086
rect 15702 15872 15811 15877
rect 15702 15816 15750 15872
rect 15806 15816 15811 15872
rect 15702 15814 15811 15816
rect 15745 15811 15811 15814
rect 7541 15808 7861 15809
rect 7541 15744 7549 15808
rect 7613 15744 7629 15808
rect 7693 15744 7709 15808
rect 7773 15744 7789 15808
rect 7853 15744 7861 15808
rect 7541 15743 7861 15744
rect 14138 15808 14458 15809
rect 14138 15744 14146 15808
rect 14210 15744 14226 15808
rect 14290 15744 14306 15808
rect 14370 15744 14386 15808
rect 14450 15744 14458 15808
rect 14138 15743 14458 15744
rect 20069 15602 20135 15605
rect 21520 15602 22000 15632
rect 20069 15600 22000 15602
rect 20069 15544 20074 15600
rect 20130 15544 22000 15600
rect 20069 15542 22000 15544
rect 20069 15539 20135 15542
rect 21520 15512 22000 15542
rect 4242 15264 4562 15265
rect 4242 15200 4250 15264
rect 4314 15200 4330 15264
rect 4394 15200 4410 15264
rect 4474 15200 4490 15264
rect 4554 15200 4562 15264
rect 4242 15199 4562 15200
rect 10840 15264 11160 15265
rect 10840 15200 10848 15264
rect 10912 15200 10928 15264
rect 10992 15200 11008 15264
rect 11072 15200 11088 15264
rect 11152 15200 11160 15264
rect 10840 15199 11160 15200
rect 17437 15264 17757 15265
rect 17437 15200 17445 15264
rect 17509 15200 17525 15264
rect 17589 15200 17605 15264
rect 17669 15200 17685 15264
rect 17749 15200 17757 15264
rect 17437 15199 17757 15200
rect 20253 15058 20319 15061
rect 21520 15058 22000 15088
rect 20253 15056 22000 15058
rect 20253 15000 20258 15056
rect 20314 15000 22000 15056
rect 20253 14998 22000 15000
rect 20253 14995 20319 14998
rect 21520 14968 22000 14998
rect 7541 14720 7861 14721
rect 7541 14656 7549 14720
rect 7613 14656 7629 14720
rect 7693 14656 7709 14720
rect 7773 14656 7789 14720
rect 7853 14656 7861 14720
rect 7541 14655 7861 14656
rect 14138 14720 14458 14721
rect 14138 14656 14146 14720
rect 14210 14656 14226 14720
rect 14290 14656 14306 14720
rect 14370 14656 14386 14720
rect 14450 14656 14458 14720
rect 14138 14655 14458 14656
rect 16573 14378 16639 14381
rect 21520 14378 22000 14408
rect 16573 14376 22000 14378
rect 16573 14320 16578 14376
rect 16634 14320 22000 14376
rect 16573 14318 22000 14320
rect 16573 14315 16639 14318
rect 21520 14288 22000 14318
rect 4242 14176 4562 14177
rect 4242 14112 4250 14176
rect 4314 14112 4330 14176
rect 4394 14112 4410 14176
rect 4474 14112 4490 14176
rect 4554 14112 4562 14176
rect 4242 14111 4562 14112
rect 10840 14176 11160 14177
rect 10840 14112 10848 14176
rect 10912 14112 10928 14176
rect 10992 14112 11008 14176
rect 11072 14112 11088 14176
rect 11152 14112 11160 14176
rect 10840 14111 11160 14112
rect 17437 14176 17757 14177
rect 17437 14112 17445 14176
rect 17509 14112 17525 14176
rect 17589 14112 17605 14176
rect 17669 14112 17685 14176
rect 17749 14112 17757 14176
rect 17437 14111 17757 14112
rect 16021 13970 16087 13973
rect 17493 13970 17559 13973
rect 16021 13968 17559 13970
rect 16021 13912 16026 13968
rect 16082 13912 17498 13968
rect 17554 13912 17559 13968
rect 16021 13910 17559 13912
rect 16021 13907 16087 13910
rect 17493 13907 17559 13910
rect 15561 13698 15627 13701
rect 21520 13698 22000 13728
rect 15561 13696 22000 13698
rect 15561 13640 15566 13696
rect 15622 13640 22000 13696
rect 15561 13638 22000 13640
rect 15561 13635 15627 13638
rect 7541 13632 7861 13633
rect 7541 13568 7549 13632
rect 7613 13568 7629 13632
rect 7693 13568 7709 13632
rect 7773 13568 7789 13632
rect 7853 13568 7861 13632
rect 7541 13567 7861 13568
rect 14138 13632 14458 13633
rect 14138 13568 14146 13632
rect 14210 13568 14226 13632
rect 14290 13568 14306 13632
rect 14370 13568 14386 13632
rect 14450 13568 14458 13632
rect 21520 13608 22000 13638
rect 14138 13567 14458 13568
rect 16113 13426 16179 13429
rect 16481 13426 16547 13429
rect 16113 13424 16547 13426
rect 16113 13368 16118 13424
rect 16174 13368 16486 13424
rect 16542 13368 16547 13424
rect 16113 13366 16547 13368
rect 16113 13363 16179 13366
rect 16481 13363 16547 13366
rect 4242 13088 4562 13089
rect 4242 13024 4250 13088
rect 4314 13024 4330 13088
rect 4394 13024 4410 13088
rect 4474 13024 4490 13088
rect 4554 13024 4562 13088
rect 4242 13023 4562 13024
rect 10840 13088 11160 13089
rect 10840 13024 10848 13088
rect 10912 13024 10928 13088
rect 10992 13024 11008 13088
rect 11072 13024 11088 13088
rect 11152 13024 11160 13088
rect 10840 13023 11160 13024
rect 17437 13088 17757 13089
rect 17437 13024 17445 13088
rect 17509 13024 17525 13088
rect 17589 13024 17605 13088
rect 17669 13024 17685 13088
rect 17749 13024 17757 13088
rect 17437 13023 17757 13024
rect 15653 13018 15719 13021
rect 17217 13018 17283 13021
rect 21520 13018 22000 13048
rect 15653 13016 17283 13018
rect 15653 12960 15658 13016
rect 15714 12960 17222 13016
rect 17278 12960 17283 13016
rect 15653 12958 17283 12960
rect 15653 12955 15719 12958
rect 17217 12955 17283 12958
rect 17910 12958 22000 13018
rect 16113 12882 16179 12885
rect 17910 12882 17970 12958
rect 21520 12928 22000 12958
rect 16113 12880 17970 12882
rect 16113 12824 16118 12880
rect 16174 12824 17970 12880
rect 16113 12822 17970 12824
rect 16113 12819 16179 12822
rect 14641 12746 14707 12749
rect 18137 12746 18203 12749
rect 14641 12744 18203 12746
rect 14641 12688 14646 12744
rect 14702 12688 18142 12744
rect 18198 12688 18203 12744
rect 14641 12686 18203 12688
rect 14641 12683 14707 12686
rect 18137 12683 18203 12686
rect 11145 12610 11211 12613
rect 11605 12610 11671 12613
rect 11145 12608 11671 12610
rect 11145 12552 11150 12608
rect 11206 12552 11610 12608
rect 11666 12552 11671 12608
rect 11145 12550 11671 12552
rect 11145 12547 11211 12550
rect 11605 12547 11671 12550
rect 14733 12610 14799 12613
rect 18505 12610 18571 12613
rect 14733 12608 18571 12610
rect 14733 12552 14738 12608
rect 14794 12552 18510 12608
rect 18566 12552 18571 12608
rect 14733 12550 18571 12552
rect 14733 12547 14799 12550
rect 18505 12547 18571 12550
rect 7541 12544 7861 12545
rect 7541 12480 7549 12544
rect 7613 12480 7629 12544
rect 7693 12480 7709 12544
rect 7773 12480 7789 12544
rect 7853 12480 7861 12544
rect 7541 12479 7861 12480
rect 14138 12544 14458 12545
rect 14138 12480 14146 12544
rect 14210 12480 14226 12544
rect 14290 12480 14306 12544
rect 14370 12480 14386 12544
rect 14450 12480 14458 12544
rect 14138 12479 14458 12480
rect 10961 12474 11027 12477
rect 13537 12474 13603 12477
rect 10961 12472 13603 12474
rect 10961 12416 10966 12472
rect 11022 12416 13542 12472
rect 13598 12416 13603 12472
rect 10961 12414 13603 12416
rect 10961 12411 11027 12414
rect 13537 12411 13603 12414
rect 15653 12474 15719 12477
rect 17769 12474 17835 12477
rect 18413 12474 18479 12477
rect 15653 12472 18479 12474
rect 15653 12416 15658 12472
rect 15714 12416 17774 12472
rect 17830 12416 18418 12472
rect 18474 12416 18479 12472
rect 15653 12414 18479 12416
rect 15653 12411 15719 12414
rect 17769 12411 17835 12414
rect 18413 12411 18479 12414
rect 10961 12338 11027 12341
rect 12617 12338 12683 12341
rect 10961 12336 12683 12338
rect 10961 12280 10966 12336
rect 11022 12280 12622 12336
rect 12678 12280 12683 12336
rect 10961 12278 12683 12280
rect 10961 12275 11027 12278
rect 12617 12275 12683 12278
rect 16757 12338 16823 12341
rect 17217 12338 17283 12341
rect 21520 12338 22000 12368
rect 16757 12336 17283 12338
rect 16757 12280 16762 12336
rect 16818 12280 17222 12336
rect 17278 12280 17283 12336
rect 16757 12278 17283 12280
rect 16757 12275 16823 12278
rect 17217 12275 17283 12278
rect 17358 12278 22000 12338
rect 10593 12202 10659 12205
rect 12433 12202 12499 12205
rect 10593 12200 12499 12202
rect 10593 12144 10598 12200
rect 10654 12144 12438 12200
rect 12494 12144 12499 12200
rect 10593 12142 12499 12144
rect 10593 12139 10659 12142
rect 12433 12139 12499 12142
rect 15561 12202 15627 12205
rect 17358 12202 17418 12278
rect 21520 12248 22000 12278
rect 15561 12200 17418 12202
rect 15561 12144 15566 12200
rect 15622 12144 17418 12200
rect 15561 12142 17418 12144
rect 17493 12202 17559 12205
rect 17493 12200 19626 12202
rect 17493 12144 17498 12200
rect 17554 12144 19626 12200
rect 17493 12142 19626 12144
rect 15561 12139 15627 12142
rect 17493 12139 17559 12142
rect 16665 12066 16731 12069
rect 16941 12066 17007 12069
rect 16665 12064 17007 12066
rect 16665 12008 16670 12064
rect 16726 12008 16946 12064
rect 17002 12008 17007 12064
rect 16665 12006 17007 12008
rect 16665 12003 16731 12006
rect 16941 12003 17007 12006
rect 4242 12000 4562 12001
rect 4242 11936 4250 12000
rect 4314 11936 4330 12000
rect 4394 11936 4410 12000
rect 4474 11936 4490 12000
rect 4554 11936 4562 12000
rect 4242 11935 4562 11936
rect 10840 12000 11160 12001
rect 10840 11936 10848 12000
rect 10912 11936 10928 12000
rect 10992 11936 11008 12000
rect 11072 11936 11088 12000
rect 11152 11936 11160 12000
rect 10840 11935 11160 11936
rect 17437 12000 17757 12001
rect 17437 11936 17445 12000
rect 17509 11936 17525 12000
rect 17589 11936 17605 12000
rect 17669 11936 17685 12000
rect 17749 11936 17757 12000
rect 17437 11935 17757 11936
rect 14089 11930 14155 11933
rect 16665 11930 16731 11933
rect 14089 11928 16731 11930
rect 14089 11872 14094 11928
rect 14150 11872 16670 11928
rect 16726 11872 16731 11928
rect 14089 11870 16731 11872
rect 14089 11867 14155 11870
rect 16665 11867 16731 11870
rect 15377 11794 15443 11797
rect 19425 11794 19491 11797
rect 15377 11792 19491 11794
rect 15377 11736 15382 11792
rect 15438 11736 19430 11792
rect 19486 11736 19491 11792
rect 15377 11734 19491 11736
rect 15377 11731 15443 11734
rect 19425 11731 19491 11734
rect 5349 11658 5415 11661
rect 9673 11658 9739 11661
rect 5349 11656 9739 11658
rect 5349 11600 5354 11656
rect 5410 11600 9678 11656
rect 9734 11600 9739 11656
rect 5349 11598 9739 11600
rect 19566 11658 19626 12142
rect 21520 11658 22000 11688
rect 19566 11598 22000 11658
rect 5349 11595 5415 11598
rect 9673 11595 9739 11598
rect 21520 11568 22000 11598
rect 7541 11456 7861 11457
rect 7541 11392 7549 11456
rect 7613 11392 7629 11456
rect 7693 11392 7709 11456
rect 7773 11392 7789 11456
rect 7853 11392 7861 11456
rect 7541 11391 7861 11392
rect 14138 11456 14458 11457
rect 14138 11392 14146 11456
rect 14210 11392 14226 11456
rect 14290 11392 14306 11456
rect 14370 11392 14386 11456
rect 14450 11392 14458 11456
rect 14138 11391 14458 11392
rect 12801 11250 12867 11253
rect 15929 11250 15995 11253
rect 12801 11248 15995 11250
rect 12801 11192 12806 11248
rect 12862 11192 15934 11248
rect 15990 11192 15995 11248
rect 12801 11190 15995 11192
rect 12801 11187 12867 11190
rect 15929 11187 15995 11190
rect 0 11114 480 11144
rect 1485 11114 1551 11117
rect 0 11112 1551 11114
rect 0 11056 1490 11112
rect 1546 11056 1551 11112
rect 0 11054 1551 11056
rect 0 11024 480 11054
rect 1485 11051 1551 11054
rect 3325 11114 3391 11117
rect 11421 11114 11487 11117
rect 3325 11112 11487 11114
rect 3325 11056 3330 11112
rect 3386 11056 11426 11112
rect 11482 11056 11487 11112
rect 3325 11054 11487 11056
rect 3325 11051 3391 11054
rect 11421 11051 11487 11054
rect 14917 11114 14983 11117
rect 16941 11114 17007 11117
rect 14917 11112 17007 11114
rect 14917 11056 14922 11112
rect 14978 11056 16946 11112
rect 17002 11056 17007 11112
rect 14917 11054 17007 11056
rect 14917 11051 14983 11054
rect 16941 11051 17007 11054
rect 17861 10978 17927 10981
rect 21520 10978 22000 11008
rect 17861 10976 22000 10978
rect 17861 10920 17866 10976
rect 17922 10920 22000 10976
rect 17861 10918 22000 10920
rect 17861 10915 17927 10918
rect 4242 10912 4562 10913
rect 4242 10848 4250 10912
rect 4314 10848 4330 10912
rect 4394 10848 4410 10912
rect 4474 10848 4490 10912
rect 4554 10848 4562 10912
rect 4242 10847 4562 10848
rect 10840 10912 11160 10913
rect 10840 10848 10848 10912
rect 10912 10848 10928 10912
rect 10992 10848 11008 10912
rect 11072 10848 11088 10912
rect 11152 10848 11160 10912
rect 10840 10847 11160 10848
rect 17437 10912 17757 10913
rect 17437 10848 17445 10912
rect 17509 10848 17525 10912
rect 17589 10848 17605 10912
rect 17669 10848 17685 10912
rect 17749 10848 17757 10912
rect 21520 10888 22000 10918
rect 17437 10847 17757 10848
rect 6453 10842 6519 10845
rect 8293 10842 8359 10845
rect 6453 10840 8359 10842
rect 6453 10784 6458 10840
rect 6514 10784 8298 10840
rect 8354 10784 8359 10840
rect 6453 10782 8359 10784
rect 6453 10779 6519 10782
rect 8293 10779 8359 10782
rect 2865 10706 2931 10709
rect 8753 10706 8819 10709
rect 2865 10704 8819 10706
rect 2865 10648 2870 10704
rect 2926 10648 8758 10704
rect 8814 10648 8819 10704
rect 2865 10646 8819 10648
rect 2865 10643 2931 10646
rect 8753 10643 8819 10646
rect 10777 10706 10843 10709
rect 14641 10706 14707 10709
rect 10777 10704 14707 10706
rect 10777 10648 10782 10704
rect 10838 10648 14646 10704
rect 14702 10648 14707 10704
rect 10777 10646 14707 10648
rect 10777 10643 10843 10646
rect 14641 10643 14707 10646
rect 7097 10570 7163 10573
rect 12893 10570 12959 10573
rect 7097 10568 12959 10570
rect 7097 10512 7102 10568
rect 7158 10512 12898 10568
rect 12954 10512 12959 10568
rect 7097 10510 12959 10512
rect 7097 10507 7163 10510
rect 12893 10507 12959 10510
rect 6269 10434 6335 10437
rect 7373 10434 7439 10437
rect 6269 10432 7439 10434
rect 6269 10376 6274 10432
rect 6330 10376 7378 10432
rect 7434 10376 7439 10432
rect 6269 10374 7439 10376
rect 6269 10371 6335 10374
rect 7373 10371 7439 10374
rect 12617 10432 12683 10437
rect 12617 10376 12622 10432
rect 12678 10376 12683 10432
rect 12617 10371 12683 10376
rect 16665 10434 16731 10437
rect 17493 10434 17559 10437
rect 16665 10432 17559 10434
rect 16665 10376 16670 10432
rect 16726 10376 17498 10432
rect 17554 10376 17559 10432
rect 16665 10374 17559 10376
rect 16665 10371 16731 10374
rect 17493 10371 17559 10374
rect 7541 10368 7861 10369
rect 7541 10304 7549 10368
rect 7613 10304 7629 10368
rect 7693 10304 7709 10368
rect 7773 10304 7789 10368
rect 7853 10304 7861 10368
rect 7541 10303 7861 10304
rect 8477 10298 8543 10301
rect 9581 10298 9647 10301
rect 8477 10296 9647 10298
rect 8477 10240 8482 10296
rect 8538 10240 9586 10296
rect 9642 10240 9647 10296
rect 8477 10238 9647 10240
rect 8477 10235 8543 10238
rect 9581 10235 9647 10238
rect 3969 10162 4035 10165
rect 11697 10162 11763 10165
rect 3969 10160 11763 10162
rect 3969 10104 3974 10160
rect 4030 10104 11702 10160
rect 11758 10104 11763 10160
rect 3969 10102 11763 10104
rect 3969 10099 4035 10102
rect 11697 10099 11763 10102
rect 11973 10162 12039 10165
rect 12620 10162 12680 10371
rect 14138 10368 14458 10369
rect 14138 10304 14146 10368
rect 14210 10304 14226 10368
rect 14290 10304 14306 10368
rect 14370 10304 14386 10368
rect 14450 10304 14458 10368
rect 14138 10303 14458 10304
rect 17033 10298 17099 10301
rect 21520 10298 22000 10328
rect 17033 10296 22000 10298
rect 17033 10240 17038 10296
rect 17094 10240 22000 10296
rect 17033 10238 22000 10240
rect 17033 10235 17099 10238
rect 21520 10208 22000 10238
rect 18045 10162 18111 10165
rect 11973 10160 18111 10162
rect 11973 10104 11978 10160
rect 12034 10104 18050 10160
rect 18106 10104 18111 10160
rect 11973 10102 18111 10104
rect 11973 10099 12039 10102
rect 18045 10099 18111 10102
rect 4061 10026 4127 10029
rect 5073 10026 5139 10029
rect 10133 10026 10199 10029
rect 12157 10026 12223 10029
rect 4061 10024 4722 10026
rect 4061 9968 4066 10024
rect 4122 9968 4722 10024
rect 4061 9966 4722 9968
rect 4061 9963 4127 9966
rect 4662 9890 4722 9966
rect 5073 10024 12223 10026
rect 5073 9968 5078 10024
rect 5134 9968 10138 10024
rect 10194 9968 12162 10024
rect 12218 9968 12223 10024
rect 5073 9966 12223 9968
rect 5073 9963 5139 9966
rect 10133 9963 10199 9966
rect 12157 9963 12223 9966
rect 8477 9890 8543 9893
rect 4662 9888 8543 9890
rect 4662 9832 8482 9888
rect 8538 9832 8543 9888
rect 4662 9830 8543 9832
rect 8477 9827 8543 9830
rect 9121 9890 9187 9893
rect 9673 9890 9739 9893
rect 12617 9890 12683 9893
rect 9121 9888 9739 9890
rect 9121 9832 9126 9888
rect 9182 9832 9678 9888
rect 9734 9832 9739 9888
rect 9121 9830 9739 9832
rect 9121 9827 9187 9830
rect 9673 9827 9739 9830
rect 11654 9888 12683 9890
rect 11654 9832 12622 9888
rect 12678 9832 12683 9888
rect 11654 9830 12683 9832
rect 4242 9824 4562 9825
rect 4242 9760 4250 9824
rect 4314 9760 4330 9824
rect 4394 9760 4410 9824
rect 4474 9760 4490 9824
rect 4554 9760 4562 9824
rect 4242 9759 4562 9760
rect 10840 9824 11160 9825
rect 10840 9760 10848 9824
rect 10912 9760 10928 9824
rect 10992 9760 11008 9824
rect 11072 9760 11088 9824
rect 11152 9760 11160 9824
rect 10840 9759 11160 9760
rect 4797 9754 4863 9757
rect 10409 9754 10475 9757
rect 4797 9752 10475 9754
rect 4797 9696 4802 9752
rect 4858 9696 10414 9752
rect 10470 9696 10475 9752
rect 4797 9694 10475 9696
rect 4797 9691 4863 9694
rect 10409 9691 10475 9694
rect 2957 9618 3023 9621
rect 11654 9618 11714 9830
rect 12617 9827 12683 9830
rect 17437 9824 17757 9825
rect 17437 9760 17445 9824
rect 17509 9760 17525 9824
rect 17589 9760 17605 9824
rect 17669 9760 17685 9824
rect 17749 9760 17757 9824
rect 17437 9759 17757 9760
rect 11789 9754 11855 9757
rect 14825 9754 14891 9757
rect 11789 9752 14891 9754
rect 11789 9696 11794 9752
rect 11850 9696 14830 9752
rect 14886 9696 14891 9752
rect 11789 9694 14891 9696
rect 11789 9691 11855 9694
rect 14825 9691 14891 9694
rect 2957 9616 11714 9618
rect 2957 9560 2962 9616
rect 3018 9560 11714 9616
rect 2957 9558 11714 9560
rect 2957 9555 3023 9558
rect 11830 9556 11836 9620
rect 11900 9618 11906 9620
rect 13077 9618 13143 9621
rect 11900 9616 13143 9618
rect 11900 9560 13082 9616
rect 13138 9560 13143 9616
rect 11900 9558 13143 9560
rect 11900 9556 11906 9558
rect 13077 9555 13143 9558
rect 16665 9618 16731 9621
rect 21520 9618 22000 9648
rect 16665 9616 22000 9618
rect 16665 9560 16670 9616
rect 16726 9560 22000 9616
rect 16665 9558 22000 9560
rect 16665 9555 16731 9558
rect 21520 9528 22000 9558
rect 2221 9482 2287 9485
rect 7097 9482 7163 9485
rect 18413 9482 18479 9485
rect 2221 9480 7163 9482
rect 2221 9424 2226 9480
rect 2282 9424 7102 9480
rect 7158 9424 7163 9480
rect 2221 9422 7163 9424
rect 2221 9419 2287 9422
rect 7097 9419 7163 9422
rect 7238 9480 18479 9482
rect 7238 9424 18418 9480
rect 18474 9424 18479 9480
rect 7238 9422 18479 9424
rect 2405 9346 2471 9349
rect 7097 9346 7163 9349
rect 2405 9344 7163 9346
rect 2405 9288 2410 9344
rect 2466 9288 7102 9344
rect 7158 9288 7163 9344
rect 2405 9286 7163 9288
rect 2405 9283 2471 9286
rect 7097 9283 7163 9286
rect 2681 9210 2747 9213
rect 7238 9210 7298 9422
rect 18413 9419 18479 9422
rect 8017 9346 8083 9349
rect 11697 9346 11763 9349
rect 8017 9344 11763 9346
rect 8017 9288 8022 9344
rect 8078 9288 11702 9344
rect 11758 9288 11763 9344
rect 8017 9286 11763 9288
rect 8017 9283 8083 9286
rect 11697 9283 11763 9286
rect 11973 9346 12039 9349
rect 12525 9346 12591 9349
rect 11973 9344 12591 9346
rect 11973 9288 11978 9344
rect 12034 9288 12530 9344
rect 12586 9288 12591 9344
rect 11973 9286 12591 9288
rect 11973 9283 12039 9286
rect 12525 9283 12591 9286
rect 15653 9346 15719 9349
rect 16481 9346 16547 9349
rect 15653 9344 16547 9346
rect 15653 9288 15658 9344
rect 15714 9288 16486 9344
rect 16542 9288 16547 9344
rect 15653 9286 16547 9288
rect 15653 9283 15719 9286
rect 16481 9283 16547 9286
rect 16665 9346 16731 9349
rect 19149 9346 19215 9349
rect 19701 9346 19767 9349
rect 16665 9344 19767 9346
rect 16665 9288 16670 9344
rect 16726 9288 19154 9344
rect 19210 9288 19706 9344
rect 19762 9288 19767 9344
rect 16665 9286 19767 9288
rect 16665 9283 16731 9286
rect 19149 9283 19215 9286
rect 19701 9283 19767 9286
rect 7541 9280 7861 9281
rect 7541 9216 7549 9280
rect 7613 9216 7629 9280
rect 7693 9216 7709 9280
rect 7773 9216 7789 9280
rect 7853 9216 7861 9280
rect 7541 9215 7861 9216
rect 14138 9280 14458 9281
rect 14138 9216 14146 9280
rect 14210 9216 14226 9280
rect 14290 9216 14306 9280
rect 14370 9216 14386 9280
rect 14450 9216 14458 9280
rect 14138 9215 14458 9216
rect 2681 9208 7298 9210
rect 2681 9152 2686 9208
rect 2742 9152 7298 9208
rect 2681 9150 7298 9152
rect 7925 9210 7991 9213
rect 14825 9210 14891 9213
rect 17309 9210 17375 9213
rect 7925 9208 13002 9210
rect 7925 9152 7930 9208
rect 7986 9152 13002 9208
rect 7925 9150 13002 9152
rect 2681 9147 2747 9150
rect 7925 9147 7991 9150
rect 3417 9074 3483 9077
rect 12382 9074 12388 9076
rect 3417 9072 12388 9074
rect 3417 9016 3422 9072
rect 3478 9016 12388 9072
rect 3417 9014 12388 9016
rect 3417 9011 3483 9014
rect 12382 9012 12388 9014
rect 12452 9012 12458 9076
rect 12942 9074 13002 9150
rect 14825 9208 17375 9210
rect 14825 9152 14830 9208
rect 14886 9152 17314 9208
rect 17370 9152 17375 9208
rect 14825 9150 17375 9152
rect 14825 9147 14891 9150
rect 17309 9147 17375 9150
rect 18781 9074 18847 9077
rect 12942 9072 18847 9074
rect 12942 9016 18786 9072
rect 18842 9016 18847 9072
rect 12942 9014 18847 9016
rect 18781 9011 18847 9014
rect 11830 8938 11836 8940
rect 4110 8844 4722 8904
rect 3325 8802 3391 8805
rect 4110 8802 4170 8844
rect 3325 8800 4170 8802
rect 3325 8744 3330 8800
rect 3386 8744 4170 8800
rect 3325 8742 4170 8744
rect 4662 8802 4722 8844
rect 10550 8878 11836 8938
rect 4662 8742 8218 8802
rect 3325 8739 3391 8742
rect 4242 8736 4562 8737
rect 4242 8672 4250 8736
rect 4314 8672 4330 8736
rect 4394 8672 4410 8736
rect 4474 8672 4490 8736
rect 4554 8672 4562 8736
rect 4242 8671 4562 8672
rect 7097 8666 7163 8669
rect 7966 8666 7972 8668
rect 7097 8664 7972 8666
rect 7097 8608 7102 8664
rect 7158 8608 7972 8664
rect 7097 8606 7972 8608
rect 7097 8603 7163 8606
rect 7966 8604 7972 8606
rect 8036 8604 8042 8668
rect 8158 8666 8218 8742
rect 10550 8666 10610 8878
rect 11830 8876 11836 8878
rect 11900 8876 11906 8940
rect 12525 8938 12591 8941
rect 15653 8938 15719 8941
rect 12525 8936 15719 8938
rect 12525 8880 12530 8936
rect 12586 8880 15658 8936
rect 15714 8880 15719 8936
rect 12525 8878 15719 8880
rect 12525 8875 12591 8878
rect 15653 8875 15719 8878
rect 15929 8938 15995 8941
rect 21520 8938 22000 8968
rect 15929 8936 22000 8938
rect 15929 8880 15934 8936
rect 15990 8880 22000 8936
rect 15929 8878 22000 8880
rect 15929 8875 15995 8878
rect 21520 8848 22000 8878
rect 12157 8802 12223 8805
rect 14181 8802 14247 8805
rect 12157 8800 14247 8802
rect 12157 8744 12162 8800
rect 12218 8744 14186 8800
rect 14242 8744 14247 8800
rect 12157 8742 14247 8744
rect 12157 8739 12223 8742
rect 14181 8739 14247 8742
rect 14365 8802 14431 8805
rect 16757 8802 16823 8805
rect 14365 8800 16823 8802
rect 14365 8744 14370 8800
rect 14426 8744 16762 8800
rect 16818 8744 16823 8800
rect 14365 8742 16823 8744
rect 14365 8739 14431 8742
rect 16757 8739 16823 8742
rect 10840 8736 11160 8737
rect 10840 8672 10848 8736
rect 10912 8672 10928 8736
rect 10992 8672 11008 8736
rect 11072 8672 11088 8736
rect 11152 8672 11160 8736
rect 10840 8671 11160 8672
rect 17437 8736 17757 8737
rect 17437 8672 17445 8736
rect 17509 8672 17525 8736
rect 17589 8672 17605 8736
rect 17669 8672 17685 8736
rect 17749 8672 17757 8736
rect 17437 8671 17757 8672
rect 8158 8606 10610 8666
rect 11697 8666 11763 8669
rect 16665 8666 16731 8669
rect 11697 8664 16731 8666
rect 11697 8608 11702 8664
rect 11758 8608 16670 8664
rect 16726 8608 16731 8664
rect 11697 8606 16731 8608
rect 11697 8603 11763 8606
rect 16665 8603 16731 8606
rect 3049 8530 3115 8533
rect 19425 8530 19491 8533
rect 3049 8528 19491 8530
rect 3049 8472 3054 8528
rect 3110 8472 19430 8528
rect 19486 8472 19491 8528
rect 3049 8470 19491 8472
rect 3049 8467 3115 8470
rect 19425 8467 19491 8470
rect 2681 8394 2747 8397
rect 7925 8394 7991 8397
rect 2681 8392 7991 8394
rect 2681 8336 2686 8392
rect 2742 8336 7930 8392
rect 7986 8336 7991 8392
rect 2681 8334 7991 8336
rect 2681 8331 2747 8334
rect 7925 8331 7991 8334
rect 8150 8332 8156 8396
rect 8220 8394 8226 8396
rect 12157 8394 12223 8397
rect 8220 8392 12223 8394
rect 8220 8336 12162 8392
rect 12218 8336 12223 8392
rect 8220 8334 12223 8336
rect 8220 8332 8226 8334
rect 12157 8331 12223 8334
rect 12382 8332 12388 8396
rect 12452 8394 12458 8396
rect 20989 8394 21055 8397
rect 12452 8392 21055 8394
rect 12452 8336 20994 8392
rect 21050 8336 21055 8392
rect 12452 8334 21055 8336
rect 12452 8332 12458 8334
rect 20989 8331 21055 8334
rect 3877 8258 3943 8261
rect 7281 8258 7347 8261
rect 3877 8256 7347 8258
rect 3877 8200 3882 8256
rect 3938 8200 7286 8256
rect 7342 8200 7347 8256
rect 3877 8198 7347 8200
rect 3877 8195 3943 8198
rect 7281 8195 7347 8198
rect 10133 8258 10199 8261
rect 13629 8258 13695 8261
rect 10133 8256 13695 8258
rect 10133 8200 10138 8256
rect 10194 8200 13634 8256
rect 13690 8200 13695 8256
rect 10133 8198 13695 8200
rect 10133 8195 10199 8198
rect 13629 8195 13695 8198
rect 15745 8258 15811 8261
rect 17309 8258 17375 8261
rect 15745 8256 17375 8258
rect 15745 8200 15750 8256
rect 15806 8200 17314 8256
rect 17370 8200 17375 8256
rect 15745 8198 17375 8200
rect 15745 8195 15811 8198
rect 17309 8195 17375 8198
rect 20161 8258 20227 8261
rect 21520 8258 22000 8288
rect 20161 8256 22000 8258
rect 20161 8200 20166 8256
rect 20222 8200 22000 8256
rect 20161 8198 22000 8200
rect 20161 8195 20227 8198
rect 7541 8192 7861 8193
rect 7541 8128 7549 8192
rect 7613 8128 7629 8192
rect 7693 8128 7709 8192
rect 7773 8128 7789 8192
rect 7853 8128 7861 8192
rect 7541 8127 7861 8128
rect 14138 8192 14458 8193
rect 14138 8128 14146 8192
rect 14210 8128 14226 8192
rect 14290 8128 14306 8192
rect 14370 8128 14386 8192
rect 14450 8128 14458 8192
rect 21520 8168 22000 8198
rect 14138 8127 14458 8128
rect 2957 8122 3023 8125
rect 7005 8122 7071 8125
rect 19885 8122 19951 8125
rect 2957 8120 7071 8122
rect 2957 8064 2962 8120
rect 3018 8064 7010 8120
rect 7066 8064 7071 8120
rect 2957 8062 7071 8064
rect 2957 8059 3023 8062
rect 7005 8059 7071 8062
rect 16254 8120 19951 8122
rect 16254 8064 19890 8120
rect 19946 8064 19951 8120
rect 16254 8062 19951 8064
rect 3601 7986 3667 7989
rect 16254 7986 16314 8062
rect 19885 8059 19951 8062
rect 3601 7984 16314 7986
rect 3601 7928 3606 7984
rect 3662 7928 16314 7984
rect 3601 7926 16314 7928
rect 17033 7986 17099 7989
rect 18321 7986 18387 7989
rect 17033 7984 18387 7986
rect 17033 7928 17038 7984
rect 17094 7928 18326 7984
rect 18382 7928 18387 7984
rect 17033 7926 18387 7928
rect 3601 7923 3667 7926
rect 17033 7923 17099 7926
rect 18321 7923 18387 7926
rect 3785 7850 3851 7853
rect 19425 7850 19491 7853
rect 3785 7848 19491 7850
rect 3785 7792 3790 7848
rect 3846 7792 19430 7848
rect 19486 7792 19491 7848
rect 3785 7790 19491 7792
rect 3785 7787 3851 7790
rect 19425 7787 19491 7790
rect 13997 7714 14063 7717
rect 16389 7714 16455 7717
rect 13997 7712 16455 7714
rect 13997 7656 14002 7712
rect 14058 7656 16394 7712
rect 16450 7656 16455 7712
rect 13997 7654 16455 7656
rect 13997 7651 14063 7654
rect 16389 7651 16455 7654
rect 19241 7714 19307 7717
rect 21520 7714 22000 7744
rect 19241 7712 22000 7714
rect 19241 7656 19246 7712
rect 19302 7656 22000 7712
rect 19241 7654 22000 7656
rect 19241 7651 19307 7654
rect 4242 7648 4562 7649
rect 4242 7584 4250 7648
rect 4314 7584 4330 7648
rect 4394 7584 4410 7648
rect 4474 7584 4490 7648
rect 4554 7584 4562 7648
rect 4242 7583 4562 7584
rect 10840 7648 11160 7649
rect 10840 7584 10848 7648
rect 10912 7584 10928 7648
rect 10992 7584 11008 7648
rect 11072 7584 11088 7648
rect 11152 7584 11160 7648
rect 10840 7583 11160 7584
rect 17437 7648 17757 7649
rect 17437 7584 17445 7648
rect 17509 7584 17525 7648
rect 17589 7584 17605 7648
rect 17669 7584 17685 7648
rect 17749 7584 17757 7648
rect 21520 7624 22000 7654
rect 17437 7583 17757 7584
rect 11329 7578 11395 7581
rect 17125 7578 17191 7581
rect 11329 7576 17191 7578
rect 11329 7520 11334 7576
rect 11390 7520 17130 7576
rect 17186 7520 17191 7576
rect 11329 7518 17191 7520
rect 11329 7515 11395 7518
rect 17125 7515 17191 7518
rect 3601 7442 3667 7445
rect 18229 7442 18295 7445
rect 3601 7440 18295 7442
rect 3601 7384 3606 7440
rect 3662 7384 18234 7440
rect 18290 7384 18295 7440
rect 3601 7382 18295 7384
rect 3601 7379 3667 7382
rect 18229 7379 18295 7382
rect 3969 7306 4035 7309
rect 20069 7306 20135 7309
rect 3969 7304 20135 7306
rect 3969 7248 3974 7304
rect 4030 7248 20074 7304
rect 20130 7248 20135 7304
rect 3969 7246 20135 7248
rect 3969 7243 4035 7246
rect 20069 7243 20135 7246
rect 8293 7170 8359 7173
rect 11329 7170 11395 7173
rect 8293 7168 11395 7170
rect 8293 7112 8298 7168
rect 8354 7112 11334 7168
rect 11390 7112 11395 7168
rect 8293 7110 11395 7112
rect 8293 7107 8359 7110
rect 11329 7107 11395 7110
rect 7541 7104 7861 7105
rect 7541 7040 7549 7104
rect 7613 7040 7629 7104
rect 7693 7040 7709 7104
rect 7773 7040 7789 7104
rect 7853 7040 7861 7104
rect 7541 7039 7861 7040
rect 14138 7104 14458 7105
rect 14138 7040 14146 7104
rect 14210 7040 14226 7104
rect 14290 7040 14306 7104
rect 14370 7040 14386 7104
rect 14450 7040 14458 7104
rect 14138 7039 14458 7040
rect 9857 7034 9923 7037
rect 11789 7034 11855 7037
rect 9857 7032 11855 7034
rect 9857 6976 9862 7032
rect 9918 6976 11794 7032
rect 11850 6976 11855 7032
rect 9857 6974 11855 6976
rect 9857 6971 9923 6974
rect 11789 6971 11855 6974
rect 18781 7034 18847 7037
rect 21520 7034 22000 7064
rect 18781 7032 22000 7034
rect 18781 6976 18786 7032
rect 18842 6976 22000 7032
rect 18781 6974 22000 6976
rect 18781 6971 18847 6974
rect 21520 6944 22000 6974
rect 12157 6898 12223 6901
rect 14733 6898 14799 6901
rect 16941 6898 17007 6901
rect 12157 6896 17007 6898
rect 12157 6840 12162 6896
rect 12218 6840 14738 6896
rect 14794 6840 16946 6896
rect 17002 6840 17007 6896
rect 12157 6838 17007 6840
rect 12157 6835 12223 6838
rect 14733 6835 14799 6838
rect 16941 6835 17007 6838
rect 7649 6762 7715 6765
rect 15009 6762 15075 6765
rect 18045 6762 18111 6765
rect 7649 6760 18111 6762
rect 7649 6704 7654 6760
rect 7710 6704 15014 6760
rect 15070 6704 18050 6760
rect 18106 6704 18111 6760
rect 7649 6702 18111 6704
rect 7649 6699 7715 6702
rect 15009 6699 15075 6702
rect 18045 6699 18111 6702
rect 4242 6560 4562 6561
rect 4242 6496 4250 6560
rect 4314 6496 4330 6560
rect 4394 6496 4410 6560
rect 4474 6496 4490 6560
rect 4554 6496 4562 6560
rect 4242 6495 4562 6496
rect 10840 6560 11160 6561
rect 10840 6496 10848 6560
rect 10912 6496 10928 6560
rect 10992 6496 11008 6560
rect 11072 6496 11088 6560
rect 11152 6496 11160 6560
rect 10840 6495 11160 6496
rect 17437 6560 17757 6561
rect 17437 6496 17445 6560
rect 17509 6496 17525 6560
rect 17589 6496 17605 6560
rect 17669 6496 17685 6560
rect 17749 6496 17757 6560
rect 17437 6495 17757 6496
rect 12525 6354 12591 6357
rect 18413 6354 18479 6357
rect 12525 6352 18479 6354
rect 12525 6296 12530 6352
rect 12586 6296 18418 6352
rect 18474 6296 18479 6352
rect 12525 6294 18479 6296
rect 12525 6291 12591 6294
rect 18413 6291 18479 6294
rect 19977 6354 20043 6357
rect 21520 6354 22000 6384
rect 19977 6352 22000 6354
rect 19977 6296 19982 6352
rect 20038 6296 22000 6352
rect 19977 6294 22000 6296
rect 19977 6291 20043 6294
rect 21520 6264 22000 6294
rect 3601 6218 3667 6221
rect 9213 6218 9279 6221
rect 15009 6218 15075 6221
rect 15561 6218 15627 6221
rect 3601 6216 9279 6218
rect 3601 6160 3606 6216
rect 3662 6160 9218 6216
rect 9274 6160 9279 6216
rect 3601 6158 9279 6160
rect 3601 6155 3667 6158
rect 9213 6155 9279 6158
rect 13310 6216 15627 6218
rect 13310 6160 15014 6216
rect 15070 6160 15566 6216
rect 15622 6160 15627 6216
rect 13310 6158 15627 6160
rect 10133 6082 10199 6085
rect 13310 6082 13370 6158
rect 15009 6155 15075 6158
rect 15561 6155 15627 6158
rect 15745 6218 15811 6221
rect 18137 6218 18203 6221
rect 15745 6216 18203 6218
rect 15745 6160 15750 6216
rect 15806 6160 18142 6216
rect 18198 6160 18203 6216
rect 15745 6158 18203 6160
rect 15745 6155 15811 6158
rect 18137 6155 18203 6158
rect 10133 6080 13370 6082
rect 10133 6024 10138 6080
rect 10194 6024 13370 6080
rect 10133 6022 13370 6024
rect 10133 6019 10199 6022
rect 7541 6016 7861 6017
rect 7541 5952 7549 6016
rect 7613 5952 7629 6016
rect 7693 5952 7709 6016
rect 7773 5952 7789 6016
rect 7853 5952 7861 6016
rect 7541 5951 7861 5952
rect 14138 6016 14458 6017
rect 14138 5952 14146 6016
rect 14210 5952 14226 6016
rect 14290 5952 14306 6016
rect 14370 5952 14386 6016
rect 14450 5952 14458 6016
rect 14138 5951 14458 5952
rect 10501 5946 10567 5949
rect 12249 5946 12315 5949
rect 10501 5944 12315 5946
rect 10501 5888 10506 5944
rect 10562 5888 12254 5944
rect 12310 5888 12315 5944
rect 10501 5886 12315 5888
rect 10501 5883 10567 5886
rect 12249 5883 12315 5886
rect 6269 5810 6335 5813
rect 12801 5810 12867 5813
rect 6269 5808 12867 5810
rect 6269 5752 6274 5808
rect 6330 5752 12806 5808
rect 12862 5752 12867 5808
rect 6269 5750 12867 5752
rect 6269 5747 6335 5750
rect 12801 5747 12867 5750
rect 12985 5810 13051 5813
rect 15929 5810 15995 5813
rect 12985 5808 15995 5810
rect 12985 5752 12990 5808
rect 13046 5752 15934 5808
rect 15990 5752 15995 5808
rect 12985 5750 15995 5752
rect 12985 5747 13051 5750
rect 15929 5747 15995 5750
rect 6545 5674 6611 5677
rect 15929 5674 15995 5677
rect 6545 5672 15995 5674
rect 6545 5616 6550 5672
rect 6606 5616 15934 5672
rect 15990 5616 15995 5672
rect 6545 5614 15995 5616
rect 6545 5611 6611 5614
rect 15929 5611 15995 5614
rect 20989 5674 21055 5677
rect 21520 5674 22000 5704
rect 20989 5672 22000 5674
rect 20989 5616 20994 5672
rect 21050 5616 22000 5672
rect 20989 5614 22000 5616
rect 20989 5611 21055 5614
rect 21520 5584 22000 5614
rect 11421 5540 11487 5541
rect 11421 5538 11468 5540
rect 11376 5536 11468 5538
rect 11532 5538 11538 5540
rect 11881 5538 11947 5541
rect 13997 5538 14063 5541
rect 11532 5536 14063 5538
rect 11376 5480 11426 5536
rect 11532 5480 11886 5536
rect 11942 5480 14002 5536
rect 14058 5480 14063 5536
rect 11376 5478 11468 5480
rect 11421 5476 11468 5478
rect 11532 5478 14063 5480
rect 11532 5476 11538 5478
rect 11421 5475 11487 5476
rect 11881 5475 11947 5478
rect 13997 5475 14063 5478
rect 4242 5472 4562 5473
rect 4242 5408 4250 5472
rect 4314 5408 4330 5472
rect 4394 5408 4410 5472
rect 4474 5408 4490 5472
rect 4554 5408 4562 5472
rect 4242 5407 4562 5408
rect 10840 5472 11160 5473
rect 10840 5408 10848 5472
rect 10912 5408 10928 5472
rect 10992 5408 11008 5472
rect 11072 5408 11088 5472
rect 11152 5408 11160 5472
rect 10840 5407 11160 5408
rect 17437 5472 17757 5473
rect 17437 5408 17445 5472
rect 17509 5408 17525 5472
rect 17589 5408 17605 5472
rect 17669 5408 17685 5472
rect 17749 5408 17757 5472
rect 17437 5407 17757 5408
rect 20253 4994 20319 4997
rect 21520 4994 22000 5024
rect 20253 4992 22000 4994
rect 20253 4936 20258 4992
rect 20314 4936 22000 4992
rect 20253 4934 22000 4936
rect 20253 4931 20319 4934
rect 7541 4928 7861 4929
rect 7541 4864 7549 4928
rect 7613 4864 7629 4928
rect 7693 4864 7709 4928
rect 7773 4864 7789 4928
rect 7853 4864 7861 4928
rect 7541 4863 7861 4864
rect 14138 4928 14458 4929
rect 14138 4864 14146 4928
rect 14210 4864 14226 4928
rect 14290 4864 14306 4928
rect 14370 4864 14386 4928
rect 14450 4864 14458 4928
rect 21520 4904 22000 4934
rect 14138 4863 14458 4864
rect 12617 4722 12683 4725
rect 18137 4722 18203 4725
rect 12617 4720 18203 4722
rect 12617 4664 12622 4720
rect 12678 4664 18142 4720
rect 18198 4664 18203 4720
rect 12617 4662 18203 4664
rect 12617 4659 12683 4662
rect 18137 4659 18203 4662
rect 16941 4586 17007 4589
rect 16941 4584 17970 4586
rect 16941 4528 16946 4584
rect 17002 4528 17970 4584
rect 16941 4526 17970 4528
rect 16941 4523 17007 4526
rect 4242 4384 4562 4385
rect 4242 4320 4250 4384
rect 4314 4320 4330 4384
rect 4394 4320 4410 4384
rect 4474 4320 4490 4384
rect 4554 4320 4562 4384
rect 4242 4319 4562 4320
rect 10840 4384 11160 4385
rect 10840 4320 10848 4384
rect 10912 4320 10928 4384
rect 10992 4320 11008 4384
rect 11072 4320 11088 4384
rect 11152 4320 11160 4384
rect 10840 4319 11160 4320
rect 17437 4384 17757 4385
rect 17437 4320 17445 4384
rect 17509 4320 17525 4384
rect 17589 4320 17605 4384
rect 17669 4320 17685 4384
rect 17749 4320 17757 4384
rect 17437 4319 17757 4320
rect 17910 4314 17970 4526
rect 21520 4314 22000 4344
rect 17910 4254 22000 4314
rect 21520 4224 22000 4254
rect 10225 4178 10291 4181
rect 4800 4176 10291 4178
rect 4800 4120 10230 4176
rect 10286 4120 10291 4176
rect 4800 4118 10291 4120
rect 0 3770 480 3800
rect 4800 3770 4860 4118
rect 10225 4115 10291 4118
rect 7541 3840 7861 3841
rect 7541 3776 7549 3840
rect 7613 3776 7629 3840
rect 7693 3776 7709 3840
rect 7773 3776 7789 3840
rect 7853 3776 7861 3840
rect 7541 3775 7861 3776
rect 14138 3840 14458 3841
rect 14138 3776 14146 3840
rect 14210 3776 14226 3840
rect 14290 3776 14306 3840
rect 14370 3776 14386 3840
rect 14450 3776 14458 3840
rect 14138 3775 14458 3776
rect 0 3710 4860 3770
rect 0 3680 480 3710
rect 10777 3634 10843 3637
rect 12157 3634 12223 3637
rect 10777 3632 12223 3634
rect 10777 3576 10782 3632
rect 10838 3576 12162 3632
rect 12218 3576 12223 3632
rect 10777 3574 12223 3576
rect 10777 3571 10843 3574
rect 12157 3571 12223 3574
rect 13169 3634 13235 3637
rect 14549 3634 14615 3637
rect 13169 3632 14615 3634
rect 13169 3576 13174 3632
rect 13230 3576 14554 3632
rect 14610 3576 14615 3632
rect 13169 3574 14615 3576
rect 13169 3571 13235 3574
rect 14549 3571 14615 3574
rect 16849 3634 16915 3637
rect 21520 3634 22000 3664
rect 16849 3632 22000 3634
rect 16849 3576 16854 3632
rect 16910 3576 22000 3632
rect 16849 3574 22000 3576
rect 16849 3571 16915 3574
rect 21520 3544 22000 3574
rect 11237 3498 11303 3501
rect 11462 3498 11468 3500
rect 11237 3496 11468 3498
rect 11237 3440 11242 3496
rect 11298 3440 11468 3496
rect 11237 3438 11468 3440
rect 11237 3435 11303 3438
rect 11462 3436 11468 3438
rect 11532 3498 11538 3500
rect 12985 3498 13051 3501
rect 11532 3496 13051 3498
rect 11532 3440 12990 3496
rect 13046 3440 13051 3496
rect 11532 3438 13051 3440
rect 11532 3436 11538 3438
rect 12985 3435 13051 3438
rect 4242 3296 4562 3297
rect 4242 3232 4250 3296
rect 4314 3232 4330 3296
rect 4394 3232 4410 3296
rect 4474 3232 4490 3296
rect 4554 3232 4562 3296
rect 4242 3231 4562 3232
rect 10840 3296 11160 3297
rect 10840 3232 10848 3296
rect 10912 3232 10928 3296
rect 10992 3232 11008 3296
rect 11072 3232 11088 3296
rect 11152 3232 11160 3296
rect 10840 3231 11160 3232
rect 17437 3296 17757 3297
rect 17437 3232 17445 3296
rect 17509 3232 17525 3296
rect 17589 3232 17605 3296
rect 17669 3232 17685 3296
rect 17749 3232 17757 3296
rect 17437 3231 17757 3232
rect 4705 3226 4771 3229
rect 9121 3226 9187 3229
rect 4705 3224 9187 3226
rect 4705 3168 4710 3224
rect 4766 3168 9126 3224
rect 9182 3168 9187 3224
rect 4705 3166 9187 3168
rect 4705 3163 4771 3166
rect 9121 3163 9187 3166
rect 12341 3090 12407 3093
rect 12617 3090 12683 3093
rect 12341 3088 12683 3090
rect 12341 3032 12346 3088
rect 12402 3032 12622 3088
rect 12678 3032 12683 3088
rect 12341 3030 12683 3032
rect 12341 3027 12407 3030
rect 12617 3027 12683 3030
rect 11513 2954 11579 2957
rect 15653 2954 15719 2957
rect 11513 2952 15719 2954
rect 11513 2896 11518 2952
rect 11574 2896 15658 2952
rect 15714 2896 15719 2952
rect 11513 2894 15719 2896
rect 11513 2891 11579 2894
rect 15653 2891 15719 2894
rect 17861 2954 17927 2957
rect 21520 2954 22000 2984
rect 17861 2952 22000 2954
rect 17861 2896 17866 2952
rect 17922 2896 22000 2952
rect 17861 2894 22000 2896
rect 17861 2891 17927 2894
rect 21520 2864 22000 2894
rect 7541 2752 7861 2753
rect 7541 2688 7549 2752
rect 7613 2688 7629 2752
rect 7693 2688 7709 2752
rect 7773 2688 7789 2752
rect 7853 2688 7861 2752
rect 7541 2687 7861 2688
rect 14138 2752 14458 2753
rect 14138 2688 14146 2752
rect 14210 2688 14226 2752
rect 14290 2688 14306 2752
rect 14370 2688 14386 2752
rect 14450 2688 14458 2752
rect 14138 2687 14458 2688
rect 18413 2274 18479 2277
rect 21520 2274 22000 2304
rect 18413 2272 22000 2274
rect 18413 2216 18418 2272
rect 18474 2216 22000 2272
rect 18413 2214 22000 2216
rect 18413 2211 18479 2214
rect 4242 2208 4562 2209
rect 4242 2144 4250 2208
rect 4314 2144 4330 2208
rect 4394 2144 4410 2208
rect 4474 2144 4490 2208
rect 4554 2144 4562 2208
rect 4242 2143 4562 2144
rect 10840 2208 11160 2209
rect 10840 2144 10848 2208
rect 10912 2144 10928 2208
rect 10992 2144 11008 2208
rect 11072 2144 11088 2208
rect 11152 2144 11160 2208
rect 10840 2143 11160 2144
rect 17437 2208 17757 2209
rect 17437 2144 17445 2208
rect 17509 2144 17525 2208
rect 17589 2144 17605 2208
rect 17669 2144 17685 2208
rect 17749 2144 17757 2208
rect 21520 2184 22000 2214
rect 17437 2143 17757 2144
rect 20713 1594 20779 1597
rect 21520 1594 22000 1624
rect 20713 1592 22000 1594
rect 20713 1536 20718 1592
rect 20774 1536 22000 1592
rect 20713 1534 22000 1536
rect 20713 1531 20779 1534
rect 21520 1504 22000 1534
rect 11697 914 11763 917
rect 16573 914 16639 917
rect 21520 914 22000 944
rect 11697 912 22000 914
rect 11697 856 11702 912
rect 11758 856 16578 912
rect 16634 856 22000 912
rect 11697 854 22000 856
rect 11697 851 11763 854
rect 16573 851 16639 854
rect 21520 824 22000 854
rect 20529 370 20595 373
rect 21520 370 22000 400
rect 20529 368 22000 370
rect 20529 312 20534 368
rect 20590 312 22000 368
rect 20529 310 22000 312
rect 20529 307 20595 310
rect 21520 280 22000 310
<< via3 >>
rect 4250 19612 4314 19616
rect 4250 19556 4254 19612
rect 4254 19556 4310 19612
rect 4310 19556 4314 19612
rect 4250 19552 4314 19556
rect 4330 19612 4394 19616
rect 4330 19556 4334 19612
rect 4334 19556 4390 19612
rect 4390 19556 4394 19612
rect 4330 19552 4394 19556
rect 4410 19612 4474 19616
rect 4410 19556 4414 19612
rect 4414 19556 4470 19612
rect 4470 19556 4474 19612
rect 4410 19552 4474 19556
rect 4490 19612 4554 19616
rect 4490 19556 4494 19612
rect 4494 19556 4550 19612
rect 4550 19556 4554 19612
rect 4490 19552 4554 19556
rect 10848 19612 10912 19616
rect 10848 19556 10852 19612
rect 10852 19556 10908 19612
rect 10908 19556 10912 19612
rect 10848 19552 10912 19556
rect 10928 19612 10992 19616
rect 10928 19556 10932 19612
rect 10932 19556 10988 19612
rect 10988 19556 10992 19612
rect 10928 19552 10992 19556
rect 11008 19612 11072 19616
rect 11008 19556 11012 19612
rect 11012 19556 11068 19612
rect 11068 19556 11072 19612
rect 11008 19552 11072 19556
rect 11088 19612 11152 19616
rect 11088 19556 11092 19612
rect 11092 19556 11148 19612
rect 11148 19556 11152 19612
rect 11088 19552 11152 19556
rect 17445 19612 17509 19616
rect 17445 19556 17449 19612
rect 17449 19556 17505 19612
rect 17505 19556 17509 19612
rect 17445 19552 17509 19556
rect 17525 19612 17589 19616
rect 17525 19556 17529 19612
rect 17529 19556 17585 19612
rect 17585 19556 17589 19612
rect 17525 19552 17589 19556
rect 17605 19612 17669 19616
rect 17605 19556 17609 19612
rect 17609 19556 17665 19612
rect 17665 19556 17669 19612
rect 17605 19552 17669 19556
rect 17685 19612 17749 19616
rect 17685 19556 17689 19612
rect 17689 19556 17745 19612
rect 17745 19556 17749 19612
rect 17685 19552 17749 19556
rect 7549 19068 7613 19072
rect 7549 19012 7553 19068
rect 7553 19012 7609 19068
rect 7609 19012 7613 19068
rect 7549 19008 7613 19012
rect 7629 19068 7693 19072
rect 7629 19012 7633 19068
rect 7633 19012 7689 19068
rect 7689 19012 7693 19068
rect 7629 19008 7693 19012
rect 7709 19068 7773 19072
rect 7709 19012 7713 19068
rect 7713 19012 7769 19068
rect 7769 19012 7773 19068
rect 7709 19008 7773 19012
rect 7789 19068 7853 19072
rect 7789 19012 7793 19068
rect 7793 19012 7849 19068
rect 7849 19012 7853 19068
rect 7789 19008 7853 19012
rect 14146 19068 14210 19072
rect 14146 19012 14150 19068
rect 14150 19012 14206 19068
rect 14206 19012 14210 19068
rect 14146 19008 14210 19012
rect 14226 19068 14290 19072
rect 14226 19012 14230 19068
rect 14230 19012 14286 19068
rect 14286 19012 14290 19068
rect 14226 19008 14290 19012
rect 14306 19068 14370 19072
rect 14306 19012 14310 19068
rect 14310 19012 14366 19068
rect 14366 19012 14370 19068
rect 14306 19008 14370 19012
rect 14386 19068 14450 19072
rect 14386 19012 14390 19068
rect 14390 19012 14446 19068
rect 14446 19012 14450 19068
rect 14386 19008 14450 19012
rect 4250 18524 4314 18528
rect 4250 18468 4254 18524
rect 4254 18468 4310 18524
rect 4310 18468 4314 18524
rect 4250 18464 4314 18468
rect 4330 18524 4394 18528
rect 4330 18468 4334 18524
rect 4334 18468 4390 18524
rect 4390 18468 4394 18524
rect 4330 18464 4394 18468
rect 4410 18524 4474 18528
rect 4410 18468 4414 18524
rect 4414 18468 4470 18524
rect 4470 18468 4474 18524
rect 4410 18464 4474 18468
rect 4490 18524 4554 18528
rect 4490 18468 4494 18524
rect 4494 18468 4550 18524
rect 4550 18468 4554 18524
rect 4490 18464 4554 18468
rect 10848 18524 10912 18528
rect 10848 18468 10852 18524
rect 10852 18468 10908 18524
rect 10908 18468 10912 18524
rect 10848 18464 10912 18468
rect 10928 18524 10992 18528
rect 10928 18468 10932 18524
rect 10932 18468 10988 18524
rect 10988 18468 10992 18524
rect 10928 18464 10992 18468
rect 11008 18524 11072 18528
rect 11008 18468 11012 18524
rect 11012 18468 11068 18524
rect 11068 18468 11072 18524
rect 11008 18464 11072 18468
rect 11088 18524 11152 18528
rect 11088 18468 11092 18524
rect 11092 18468 11148 18524
rect 11148 18468 11152 18524
rect 11088 18464 11152 18468
rect 17445 18524 17509 18528
rect 17445 18468 17449 18524
rect 17449 18468 17505 18524
rect 17505 18468 17509 18524
rect 17445 18464 17509 18468
rect 17525 18524 17589 18528
rect 17525 18468 17529 18524
rect 17529 18468 17585 18524
rect 17585 18468 17589 18524
rect 17525 18464 17589 18468
rect 17605 18524 17669 18528
rect 17605 18468 17609 18524
rect 17609 18468 17665 18524
rect 17665 18468 17669 18524
rect 17605 18464 17669 18468
rect 17685 18524 17749 18528
rect 17685 18468 17689 18524
rect 17689 18468 17745 18524
rect 17745 18468 17749 18524
rect 17685 18464 17749 18468
rect 14964 17988 15028 18052
rect 7549 17980 7613 17984
rect 7549 17924 7553 17980
rect 7553 17924 7609 17980
rect 7609 17924 7613 17980
rect 7549 17920 7613 17924
rect 7629 17980 7693 17984
rect 7629 17924 7633 17980
rect 7633 17924 7689 17980
rect 7689 17924 7693 17980
rect 7629 17920 7693 17924
rect 7709 17980 7773 17984
rect 7709 17924 7713 17980
rect 7713 17924 7769 17980
rect 7769 17924 7773 17980
rect 7709 17920 7773 17924
rect 7789 17980 7853 17984
rect 7789 17924 7793 17980
rect 7793 17924 7849 17980
rect 7849 17924 7853 17980
rect 7789 17920 7853 17924
rect 14146 17980 14210 17984
rect 14146 17924 14150 17980
rect 14150 17924 14206 17980
rect 14206 17924 14210 17980
rect 14146 17920 14210 17924
rect 14226 17980 14290 17984
rect 14226 17924 14230 17980
rect 14230 17924 14286 17980
rect 14286 17924 14290 17980
rect 14226 17920 14290 17924
rect 14306 17980 14370 17984
rect 14306 17924 14310 17980
rect 14310 17924 14366 17980
rect 14366 17924 14370 17980
rect 14306 17920 14370 17924
rect 14386 17980 14450 17984
rect 14386 17924 14390 17980
rect 14390 17924 14446 17980
rect 14446 17924 14450 17980
rect 14386 17920 14450 17924
rect 4250 17436 4314 17440
rect 4250 17380 4254 17436
rect 4254 17380 4310 17436
rect 4310 17380 4314 17436
rect 4250 17376 4314 17380
rect 4330 17436 4394 17440
rect 4330 17380 4334 17436
rect 4334 17380 4390 17436
rect 4390 17380 4394 17436
rect 4330 17376 4394 17380
rect 4410 17436 4474 17440
rect 4410 17380 4414 17436
rect 4414 17380 4470 17436
rect 4470 17380 4474 17436
rect 4410 17376 4474 17380
rect 4490 17436 4554 17440
rect 4490 17380 4494 17436
rect 4494 17380 4550 17436
rect 4550 17380 4554 17436
rect 4490 17376 4554 17380
rect 10848 17436 10912 17440
rect 10848 17380 10852 17436
rect 10852 17380 10908 17436
rect 10908 17380 10912 17436
rect 10848 17376 10912 17380
rect 10928 17436 10992 17440
rect 10928 17380 10932 17436
rect 10932 17380 10988 17436
rect 10988 17380 10992 17436
rect 10928 17376 10992 17380
rect 11008 17436 11072 17440
rect 11008 17380 11012 17436
rect 11012 17380 11068 17436
rect 11068 17380 11072 17436
rect 11008 17376 11072 17380
rect 11088 17436 11152 17440
rect 11088 17380 11092 17436
rect 11092 17380 11148 17436
rect 11148 17380 11152 17436
rect 11088 17376 11152 17380
rect 17445 17436 17509 17440
rect 17445 17380 17449 17436
rect 17449 17380 17505 17436
rect 17505 17380 17509 17436
rect 17445 17376 17509 17380
rect 17525 17436 17589 17440
rect 17525 17380 17529 17436
rect 17529 17380 17585 17436
rect 17585 17380 17589 17436
rect 17525 17376 17589 17380
rect 17605 17436 17669 17440
rect 17605 17380 17609 17436
rect 17609 17380 17665 17436
rect 17665 17380 17669 17436
rect 17605 17376 17669 17380
rect 17685 17436 17749 17440
rect 17685 17380 17689 17436
rect 17689 17380 17745 17436
rect 17745 17380 17749 17436
rect 17685 17376 17749 17380
rect 7549 16892 7613 16896
rect 7549 16836 7553 16892
rect 7553 16836 7609 16892
rect 7609 16836 7613 16892
rect 7549 16832 7613 16836
rect 7629 16892 7693 16896
rect 7629 16836 7633 16892
rect 7633 16836 7689 16892
rect 7689 16836 7693 16892
rect 7629 16832 7693 16836
rect 7709 16892 7773 16896
rect 7709 16836 7713 16892
rect 7713 16836 7769 16892
rect 7769 16836 7773 16892
rect 7709 16832 7773 16836
rect 7789 16892 7853 16896
rect 7789 16836 7793 16892
rect 7793 16836 7849 16892
rect 7849 16836 7853 16892
rect 7789 16832 7853 16836
rect 14146 16892 14210 16896
rect 14146 16836 14150 16892
rect 14150 16836 14206 16892
rect 14206 16836 14210 16892
rect 14146 16832 14210 16836
rect 14226 16892 14290 16896
rect 14226 16836 14230 16892
rect 14230 16836 14286 16892
rect 14286 16836 14290 16892
rect 14226 16832 14290 16836
rect 14306 16892 14370 16896
rect 14306 16836 14310 16892
rect 14310 16836 14366 16892
rect 14366 16836 14370 16892
rect 14306 16832 14370 16836
rect 14386 16892 14450 16896
rect 14386 16836 14390 16892
rect 14390 16836 14446 16892
rect 14446 16836 14450 16892
rect 14386 16832 14450 16836
rect 14964 16492 15028 16556
rect 4250 16348 4314 16352
rect 4250 16292 4254 16348
rect 4254 16292 4310 16348
rect 4310 16292 4314 16348
rect 4250 16288 4314 16292
rect 4330 16348 4394 16352
rect 4330 16292 4334 16348
rect 4334 16292 4390 16348
rect 4390 16292 4394 16348
rect 4330 16288 4394 16292
rect 4410 16348 4474 16352
rect 4410 16292 4414 16348
rect 4414 16292 4470 16348
rect 4470 16292 4474 16348
rect 4410 16288 4474 16292
rect 4490 16348 4554 16352
rect 4490 16292 4494 16348
rect 4494 16292 4550 16348
rect 4550 16292 4554 16348
rect 4490 16288 4554 16292
rect 10848 16348 10912 16352
rect 10848 16292 10852 16348
rect 10852 16292 10908 16348
rect 10908 16292 10912 16348
rect 10848 16288 10912 16292
rect 10928 16348 10992 16352
rect 10928 16292 10932 16348
rect 10932 16292 10988 16348
rect 10988 16292 10992 16348
rect 10928 16288 10992 16292
rect 11008 16348 11072 16352
rect 11008 16292 11012 16348
rect 11012 16292 11068 16348
rect 11068 16292 11072 16348
rect 11008 16288 11072 16292
rect 11088 16348 11152 16352
rect 11088 16292 11092 16348
rect 11092 16292 11148 16348
rect 11148 16292 11152 16348
rect 11088 16288 11152 16292
rect 17445 16348 17509 16352
rect 17445 16292 17449 16348
rect 17449 16292 17505 16348
rect 17505 16292 17509 16348
rect 17445 16288 17509 16292
rect 17525 16348 17589 16352
rect 17525 16292 17529 16348
rect 17529 16292 17585 16348
rect 17585 16292 17589 16348
rect 17525 16288 17589 16292
rect 17605 16348 17669 16352
rect 17605 16292 17609 16348
rect 17609 16292 17665 16348
rect 17665 16292 17669 16348
rect 17605 16288 17669 16292
rect 17685 16348 17749 16352
rect 17685 16292 17689 16348
rect 17689 16292 17745 16348
rect 17745 16292 17749 16348
rect 17685 16288 17749 16292
rect 7549 15804 7613 15808
rect 7549 15748 7553 15804
rect 7553 15748 7609 15804
rect 7609 15748 7613 15804
rect 7549 15744 7613 15748
rect 7629 15804 7693 15808
rect 7629 15748 7633 15804
rect 7633 15748 7689 15804
rect 7689 15748 7693 15804
rect 7629 15744 7693 15748
rect 7709 15804 7773 15808
rect 7709 15748 7713 15804
rect 7713 15748 7769 15804
rect 7769 15748 7773 15804
rect 7709 15744 7773 15748
rect 7789 15804 7853 15808
rect 7789 15748 7793 15804
rect 7793 15748 7849 15804
rect 7849 15748 7853 15804
rect 7789 15744 7853 15748
rect 14146 15804 14210 15808
rect 14146 15748 14150 15804
rect 14150 15748 14206 15804
rect 14206 15748 14210 15804
rect 14146 15744 14210 15748
rect 14226 15804 14290 15808
rect 14226 15748 14230 15804
rect 14230 15748 14286 15804
rect 14286 15748 14290 15804
rect 14226 15744 14290 15748
rect 14306 15804 14370 15808
rect 14306 15748 14310 15804
rect 14310 15748 14366 15804
rect 14366 15748 14370 15804
rect 14306 15744 14370 15748
rect 14386 15804 14450 15808
rect 14386 15748 14390 15804
rect 14390 15748 14446 15804
rect 14446 15748 14450 15804
rect 14386 15744 14450 15748
rect 4250 15260 4314 15264
rect 4250 15204 4254 15260
rect 4254 15204 4310 15260
rect 4310 15204 4314 15260
rect 4250 15200 4314 15204
rect 4330 15260 4394 15264
rect 4330 15204 4334 15260
rect 4334 15204 4390 15260
rect 4390 15204 4394 15260
rect 4330 15200 4394 15204
rect 4410 15260 4474 15264
rect 4410 15204 4414 15260
rect 4414 15204 4470 15260
rect 4470 15204 4474 15260
rect 4410 15200 4474 15204
rect 4490 15260 4554 15264
rect 4490 15204 4494 15260
rect 4494 15204 4550 15260
rect 4550 15204 4554 15260
rect 4490 15200 4554 15204
rect 10848 15260 10912 15264
rect 10848 15204 10852 15260
rect 10852 15204 10908 15260
rect 10908 15204 10912 15260
rect 10848 15200 10912 15204
rect 10928 15260 10992 15264
rect 10928 15204 10932 15260
rect 10932 15204 10988 15260
rect 10988 15204 10992 15260
rect 10928 15200 10992 15204
rect 11008 15260 11072 15264
rect 11008 15204 11012 15260
rect 11012 15204 11068 15260
rect 11068 15204 11072 15260
rect 11008 15200 11072 15204
rect 11088 15260 11152 15264
rect 11088 15204 11092 15260
rect 11092 15204 11148 15260
rect 11148 15204 11152 15260
rect 11088 15200 11152 15204
rect 17445 15260 17509 15264
rect 17445 15204 17449 15260
rect 17449 15204 17505 15260
rect 17505 15204 17509 15260
rect 17445 15200 17509 15204
rect 17525 15260 17589 15264
rect 17525 15204 17529 15260
rect 17529 15204 17585 15260
rect 17585 15204 17589 15260
rect 17525 15200 17589 15204
rect 17605 15260 17669 15264
rect 17605 15204 17609 15260
rect 17609 15204 17665 15260
rect 17665 15204 17669 15260
rect 17605 15200 17669 15204
rect 17685 15260 17749 15264
rect 17685 15204 17689 15260
rect 17689 15204 17745 15260
rect 17745 15204 17749 15260
rect 17685 15200 17749 15204
rect 7549 14716 7613 14720
rect 7549 14660 7553 14716
rect 7553 14660 7609 14716
rect 7609 14660 7613 14716
rect 7549 14656 7613 14660
rect 7629 14716 7693 14720
rect 7629 14660 7633 14716
rect 7633 14660 7689 14716
rect 7689 14660 7693 14716
rect 7629 14656 7693 14660
rect 7709 14716 7773 14720
rect 7709 14660 7713 14716
rect 7713 14660 7769 14716
rect 7769 14660 7773 14716
rect 7709 14656 7773 14660
rect 7789 14716 7853 14720
rect 7789 14660 7793 14716
rect 7793 14660 7849 14716
rect 7849 14660 7853 14716
rect 7789 14656 7853 14660
rect 14146 14716 14210 14720
rect 14146 14660 14150 14716
rect 14150 14660 14206 14716
rect 14206 14660 14210 14716
rect 14146 14656 14210 14660
rect 14226 14716 14290 14720
rect 14226 14660 14230 14716
rect 14230 14660 14286 14716
rect 14286 14660 14290 14716
rect 14226 14656 14290 14660
rect 14306 14716 14370 14720
rect 14306 14660 14310 14716
rect 14310 14660 14366 14716
rect 14366 14660 14370 14716
rect 14306 14656 14370 14660
rect 14386 14716 14450 14720
rect 14386 14660 14390 14716
rect 14390 14660 14446 14716
rect 14446 14660 14450 14716
rect 14386 14656 14450 14660
rect 4250 14172 4314 14176
rect 4250 14116 4254 14172
rect 4254 14116 4310 14172
rect 4310 14116 4314 14172
rect 4250 14112 4314 14116
rect 4330 14172 4394 14176
rect 4330 14116 4334 14172
rect 4334 14116 4390 14172
rect 4390 14116 4394 14172
rect 4330 14112 4394 14116
rect 4410 14172 4474 14176
rect 4410 14116 4414 14172
rect 4414 14116 4470 14172
rect 4470 14116 4474 14172
rect 4410 14112 4474 14116
rect 4490 14172 4554 14176
rect 4490 14116 4494 14172
rect 4494 14116 4550 14172
rect 4550 14116 4554 14172
rect 4490 14112 4554 14116
rect 10848 14172 10912 14176
rect 10848 14116 10852 14172
rect 10852 14116 10908 14172
rect 10908 14116 10912 14172
rect 10848 14112 10912 14116
rect 10928 14172 10992 14176
rect 10928 14116 10932 14172
rect 10932 14116 10988 14172
rect 10988 14116 10992 14172
rect 10928 14112 10992 14116
rect 11008 14172 11072 14176
rect 11008 14116 11012 14172
rect 11012 14116 11068 14172
rect 11068 14116 11072 14172
rect 11008 14112 11072 14116
rect 11088 14172 11152 14176
rect 11088 14116 11092 14172
rect 11092 14116 11148 14172
rect 11148 14116 11152 14172
rect 11088 14112 11152 14116
rect 17445 14172 17509 14176
rect 17445 14116 17449 14172
rect 17449 14116 17505 14172
rect 17505 14116 17509 14172
rect 17445 14112 17509 14116
rect 17525 14172 17589 14176
rect 17525 14116 17529 14172
rect 17529 14116 17585 14172
rect 17585 14116 17589 14172
rect 17525 14112 17589 14116
rect 17605 14172 17669 14176
rect 17605 14116 17609 14172
rect 17609 14116 17665 14172
rect 17665 14116 17669 14172
rect 17605 14112 17669 14116
rect 17685 14172 17749 14176
rect 17685 14116 17689 14172
rect 17689 14116 17745 14172
rect 17745 14116 17749 14172
rect 17685 14112 17749 14116
rect 7549 13628 7613 13632
rect 7549 13572 7553 13628
rect 7553 13572 7609 13628
rect 7609 13572 7613 13628
rect 7549 13568 7613 13572
rect 7629 13628 7693 13632
rect 7629 13572 7633 13628
rect 7633 13572 7689 13628
rect 7689 13572 7693 13628
rect 7629 13568 7693 13572
rect 7709 13628 7773 13632
rect 7709 13572 7713 13628
rect 7713 13572 7769 13628
rect 7769 13572 7773 13628
rect 7709 13568 7773 13572
rect 7789 13628 7853 13632
rect 7789 13572 7793 13628
rect 7793 13572 7849 13628
rect 7849 13572 7853 13628
rect 7789 13568 7853 13572
rect 14146 13628 14210 13632
rect 14146 13572 14150 13628
rect 14150 13572 14206 13628
rect 14206 13572 14210 13628
rect 14146 13568 14210 13572
rect 14226 13628 14290 13632
rect 14226 13572 14230 13628
rect 14230 13572 14286 13628
rect 14286 13572 14290 13628
rect 14226 13568 14290 13572
rect 14306 13628 14370 13632
rect 14306 13572 14310 13628
rect 14310 13572 14366 13628
rect 14366 13572 14370 13628
rect 14306 13568 14370 13572
rect 14386 13628 14450 13632
rect 14386 13572 14390 13628
rect 14390 13572 14446 13628
rect 14446 13572 14450 13628
rect 14386 13568 14450 13572
rect 4250 13084 4314 13088
rect 4250 13028 4254 13084
rect 4254 13028 4310 13084
rect 4310 13028 4314 13084
rect 4250 13024 4314 13028
rect 4330 13084 4394 13088
rect 4330 13028 4334 13084
rect 4334 13028 4390 13084
rect 4390 13028 4394 13084
rect 4330 13024 4394 13028
rect 4410 13084 4474 13088
rect 4410 13028 4414 13084
rect 4414 13028 4470 13084
rect 4470 13028 4474 13084
rect 4410 13024 4474 13028
rect 4490 13084 4554 13088
rect 4490 13028 4494 13084
rect 4494 13028 4550 13084
rect 4550 13028 4554 13084
rect 4490 13024 4554 13028
rect 10848 13084 10912 13088
rect 10848 13028 10852 13084
rect 10852 13028 10908 13084
rect 10908 13028 10912 13084
rect 10848 13024 10912 13028
rect 10928 13084 10992 13088
rect 10928 13028 10932 13084
rect 10932 13028 10988 13084
rect 10988 13028 10992 13084
rect 10928 13024 10992 13028
rect 11008 13084 11072 13088
rect 11008 13028 11012 13084
rect 11012 13028 11068 13084
rect 11068 13028 11072 13084
rect 11008 13024 11072 13028
rect 11088 13084 11152 13088
rect 11088 13028 11092 13084
rect 11092 13028 11148 13084
rect 11148 13028 11152 13084
rect 11088 13024 11152 13028
rect 17445 13084 17509 13088
rect 17445 13028 17449 13084
rect 17449 13028 17505 13084
rect 17505 13028 17509 13084
rect 17445 13024 17509 13028
rect 17525 13084 17589 13088
rect 17525 13028 17529 13084
rect 17529 13028 17585 13084
rect 17585 13028 17589 13084
rect 17525 13024 17589 13028
rect 17605 13084 17669 13088
rect 17605 13028 17609 13084
rect 17609 13028 17665 13084
rect 17665 13028 17669 13084
rect 17605 13024 17669 13028
rect 17685 13084 17749 13088
rect 17685 13028 17689 13084
rect 17689 13028 17745 13084
rect 17745 13028 17749 13084
rect 17685 13024 17749 13028
rect 7549 12540 7613 12544
rect 7549 12484 7553 12540
rect 7553 12484 7609 12540
rect 7609 12484 7613 12540
rect 7549 12480 7613 12484
rect 7629 12540 7693 12544
rect 7629 12484 7633 12540
rect 7633 12484 7689 12540
rect 7689 12484 7693 12540
rect 7629 12480 7693 12484
rect 7709 12540 7773 12544
rect 7709 12484 7713 12540
rect 7713 12484 7769 12540
rect 7769 12484 7773 12540
rect 7709 12480 7773 12484
rect 7789 12540 7853 12544
rect 7789 12484 7793 12540
rect 7793 12484 7849 12540
rect 7849 12484 7853 12540
rect 7789 12480 7853 12484
rect 14146 12540 14210 12544
rect 14146 12484 14150 12540
rect 14150 12484 14206 12540
rect 14206 12484 14210 12540
rect 14146 12480 14210 12484
rect 14226 12540 14290 12544
rect 14226 12484 14230 12540
rect 14230 12484 14286 12540
rect 14286 12484 14290 12540
rect 14226 12480 14290 12484
rect 14306 12540 14370 12544
rect 14306 12484 14310 12540
rect 14310 12484 14366 12540
rect 14366 12484 14370 12540
rect 14306 12480 14370 12484
rect 14386 12540 14450 12544
rect 14386 12484 14390 12540
rect 14390 12484 14446 12540
rect 14446 12484 14450 12540
rect 14386 12480 14450 12484
rect 4250 11996 4314 12000
rect 4250 11940 4254 11996
rect 4254 11940 4310 11996
rect 4310 11940 4314 11996
rect 4250 11936 4314 11940
rect 4330 11996 4394 12000
rect 4330 11940 4334 11996
rect 4334 11940 4390 11996
rect 4390 11940 4394 11996
rect 4330 11936 4394 11940
rect 4410 11996 4474 12000
rect 4410 11940 4414 11996
rect 4414 11940 4470 11996
rect 4470 11940 4474 11996
rect 4410 11936 4474 11940
rect 4490 11996 4554 12000
rect 4490 11940 4494 11996
rect 4494 11940 4550 11996
rect 4550 11940 4554 11996
rect 4490 11936 4554 11940
rect 10848 11996 10912 12000
rect 10848 11940 10852 11996
rect 10852 11940 10908 11996
rect 10908 11940 10912 11996
rect 10848 11936 10912 11940
rect 10928 11996 10992 12000
rect 10928 11940 10932 11996
rect 10932 11940 10988 11996
rect 10988 11940 10992 11996
rect 10928 11936 10992 11940
rect 11008 11996 11072 12000
rect 11008 11940 11012 11996
rect 11012 11940 11068 11996
rect 11068 11940 11072 11996
rect 11008 11936 11072 11940
rect 11088 11996 11152 12000
rect 11088 11940 11092 11996
rect 11092 11940 11148 11996
rect 11148 11940 11152 11996
rect 11088 11936 11152 11940
rect 17445 11996 17509 12000
rect 17445 11940 17449 11996
rect 17449 11940 17505 11996
rect 17505 11940 17509 11996
rect 17445 11936 17509 11940
rect 17525 11996 17589 12000
rect 17525 11940 17529 11996
rect 17529 11940 17585 11996
rect 17585 11940 17589 11996
rect 17525 11936 17589 11940
rect 17605 11996 17669 12000
rect 17605 11940 17609 11996
rect 17609 11940 17665 11996
rect 17665 11940 17669 11996
rect 17605 11936 17669 11940
rect 17685 11996 17749 12000
rect 17685 11940 17689 11996
rect 17689 11940 17745 11996
rect 17745 11940 17749 11996
rect 17685 11936 17749 11940
rect 7549 11452 7613 11456
rect 7549 11396 7553 11452
rect 7553 11396 7609 11452
rect 7609 11396 7613 11452
rect 7549 11392 7613 11396
rect 7629 11452 7693 11456
rect 7629 11396 7633 11452
rect 7633 11396 7689 11452
rect 7689 11396 7693 11452
rect 7629 11392 7693 11396
rect 7709 11452 7773 11456
rect 7709 11396 7713 11452
rect 7713 11396 7769 11452
rect 7769 11396 7773 11452
rect 7709 11392 7773 11396
rect 7789 11452 7853 11456
rect 7789 11396 7793 11452
rect 7793 11396 7849 11452
rect 7849 11396 7853 11452
rect 7789 11392 7853 11396
rect 14146 11452 14210 11456
rect 14146 11396 14150 11452
rect 14150 11396 14206 11452
rect 14206 11396 14210 11452
rect 14146 11392 14210 11396
rect 14226 11452 14290 11456
rect 14226 11396 14230 11452
rect 14230 11396 14286 11452
rect 14286 11396 14290 11452
rect 14226 11392 14290 11396
rect 14306 11452 14370 11456
rect 14306 11396 14310 11452
rect 14310 11396 14366 11452
rect 14366 11396 14370 11452
rect 14306 11392 14370 11396
rect 14386 11452 14450 11456
rect 14386 11396 14390 11452
rect 14390 11396 14446 11452
rect 14446 11396 14450 11452
rect 14386 11392 14450 11396
rect 4250 10908 4314 10912
rect 4250 10852 4254 10908
rect 4254 10852 4310 10908
rect 4310 10852 4314 10908
rect 4250 10848 4314 10852
rect 4330 10908 4394 10912
rect 4330 10852 4334 10908
rect 4334 10852 4390 10908
rect 4390 10852 4394 10908
rect 4330 10848 4394 10852
rect 4410 10908 4474 10912
rect 4410 10852 4414 10908
rect 4414 10852 4470 10908
rect 4470 10852 4474 10908
rect 4410 10848 4474 10852
rect 4490 10908 4554 10912
rect 4490 10852 4494 10908
rect 4494 10852 4550 10908
rect 4550 10852 4554 10908
rect 4490 10848 4554 10852
rect 10848 10908 10912 10912
rect 10848 10852 10852 10908
rect 10852 10852 10908 10908
rect 10908 10852 10912 10908
rect 10848 10848 10912 10852
rect 10928 10908 10992 10912
rect 10928 10852 10932 10908
rect 10932 10852 10988 10908
rect 10988 10852 10992 10908
rect 10928 10848 10992 10852
rect 11008 10908 11072 10912
rect 11008 10852 11012 10908
rect 11012 10852 11068 10908
rect 11068 10852 11072 10908
rect 11008 10848 11072 10852
rect 11088 10908 11152 10912
rect 11088 10852 11092 10908
rect 11092 10852 11148 10908
rect 11148 10852 11152 10908
rect 11088 10848 11152 10852
rect 17445 10908 17509 10912
rect 17445 10852 17449 10908
rect 17449 10852 17505 10908
rect 17505 10852 17509 10908
rect 17445 10848 17509 10852
rect 17525 10908 17589 10912
rect 17525 10852 17529 10908
rect 17529 10852 17585 10908
rect 17585 10852 17589 10908
rect 17525 10848 17589 10852
rect 17605 10908 17669 10912
rect 17605 10852 17609 10908
rect 17609 10852 17665 10908
rect 17665 10852 17669 10908
rect 17605 10848 17669 10852
rect 17685 10908 17749 10912
rect 17685 10852 17689 10908
rect 17689 10852 17745 10908
rect 17745 10852 17749 10908
rect 17685 10848 17749 10852
rect 7549 10364 7613 10368
rect 7549 10308 7553 10364
rect 7553 10308 7609 10364
rect 7609 10308 7613 10364
rect 7549 10304 7613 10308
rect 7629 10364 7693 10368
rect 7629 10308 7633 10364
rect 7633 10308 7689 10364
rect 7689 10308 7693 10364
rect 7629 10304 7693 10308
rect 7709 10364 7773 10368
rect 7709 10308 7713 10364
rect 7713 10308 7769 10364
rect 7769 10308 7773 10364
rect 7709 10304 7773 10308
rect 7789 10364 7853 10368
rect 7789 10308 7793 10364
rect 7793 10308 7849 10364
rect 7849 10308 7853 10364
rect 7789 10304 7853 10308
rect 14146 10364 14210 10368
rect 14146 10308 14150 10364
rect 14150 10308 14206 10364
rect 14206 10308 14210 10364
rect 14146 10304 14210 10308
rect 14226 10364 14290 10368
rect 14226 10308 14230 10364
rect 14230 10308 14286 10364
rect 14286 10308 14290 10364
rect 14226 10304 14290 10308
rect 14306 10364 14370 10368
rect 14306 10308 14310 10364
rect 14310 10308 14366 10364
rect 14366 10308 14370 10364
rect 14306 10304 14370 10308
rect 14386 10364 14450 10368
rect 14386 10308 14390 10364
rect 14390 10308 14446 10364
rect 14446 10308 14450 10364
rect 14386 10304 14450 10308
rect 4250 9820 4314 9824
rect 4250 9764 4254 9820
rect 4254 9764 4310 9820
rect 4310 9764 4314 9820
rect 4250 9760 4314 9764
rect 4330 9820 4394 9824
rect 4330 9764 4334 9820
rect 4334 9764 4390 9820
rect 4390 9764 4394 9820
rect 4330 9760 4394 9764
rect 4410 9820 4474 9824
rect 4410 9764 4414 9820
rect 4414 9764 4470 9820
rect 4470 9764 4474 9820
rect 4410 9760 4474 9764
rect 4490 9820 4554 9824
rect 4490 9764 4494 9820
rect 4494 9764 4550 9820
rect 4550 9764 4554 9820
rect 4490 9760 4554 9764
rect 10848 9820 10912 9824
rect 10848 9764 10852 9820
rect 10852 9764 10908 9820
rect 10908 9764 10912 9820
rect 10848 9760 10912 9764
rect 10928 9820 10992 9824
rect 10928 9764 10932 9820
rect 10932 9764 10988 9820
rect 10988 9764 10992 9820
rect 10928 9760 10992 9764
rect 11008 9820 11072 9824
rect 11008 9764 11012 9820
rect 11012 9764 11068 9820
rect 11068 9764 11072 9820
rect 11008 9760 11072 9764
rect 11088 9820 11152 9824
rect 11088 9764 11092 9820
rect 11092 9764 11148 9820
rect 11148 9764 11152 9820
rect 11088 9760 11152 9764
rect 17445 9820 17509 9824
rect 17445 9764 17449 9820
rect 17449 9764 17505 9820
rect 17505 9764 17509 9820
rect 17445 9760 17509 9764
rect 17525 9820 17589 9824
rect 17525 9764 17529 9820
rect 17529 9764 17585 9820
rect 17585 9764 17589 9820
rect 17525 9760 17589 9764
rect 17605 9820 17669 9824
rect 17605 9764 17609 9820
rect 17609 9764 17665 9820
rect 17665 9764 17669 9820
rect 17605 9760 17669 9764
rect 17685 9820 17749 9824
rect 17685 9764 17689 9820
rect 17689 9764 17745 9820
rect 17745 9764 17749 9820
rect 17685 9760 17749 9764
rect 11836 9556 11900 9620
rect 7549 9276 7613 9280
rect 7549 9220 7553 9276
rect 7553 9220 7609 9276
rect 7609 9220 7613 9276
rect 7549 9216 7613 9220
rect 7629 9276 7693 9280
rect 7629 9220 7633 9276
rect 7633 9220 7689 9276
rect 7689 9220 7693 9276
rect 7629 9216 7693 9220
rect 7709 9276 7773 9280
rect 7709 9220 7713 9276
rect 7713 9220 7769 9276
rect 7769 9220 7773 9276
rect 7709 9216 7773 9220
rect 7789 9276 7853 9280
rect 7789 9220 7793 9276
rect 7793 9220 7849 9276
rect 7849 9220 7853 9276
rect 7789 9216 7853 9220
rect 14146 9276 14210 9280
rect 14146 9220 14150 9276
rect 14150 9220 14206 9276
rect 14206 9220 14210 9276
rect 14146 9216 14210 9220
rect 14226 9276 14290 9280
rect 14226 9220 14230 9276
rect 14230 9220 14286 9276
rect 14286 9220 14290 9276
rect 14226 9216 14290 9220
rect 14306 9276 14370 9280
rect 14306 9220 14310 9276
rect 14310 9220 14366 9276
rect 14366 9220 14370 9276
rect 14306 9216 14370 9220
rect 14386 9276 14450 9280
rect 14386 9220 14390 9276
rect 14390 9220 14446 9276
rect 14446 9220 14450 9276
rect 14386 9216 14450 9220
rect 12388 9012 12452 9076
rect 4250 8732 4314 8736
rect 4250 8676 4254 8732
rect 4254 8676 4310 8732
rect 4310 8676 4314 8732
rect 4250 8672 4314 8676
rect 4330 8732 4394 8736
rect 4330 8676 4334 8732
rect 4334 8676 4390 8732
rect 4390 8676 4394 8732
rect 4330 8672 4394 8676
rect 4410 8732 4474 8736
rect 4410 8676 4414 8732
rect 4414 8676 4470 8732
rect 4470 8676 4474 8732
rect 4410 8672 4474 8676
rect 4490 8732 4554 8736
rect 4490 8676 4494 8732
rect 4494 8676 4550 8732
rect 4550 8676 4554 8732
rect 4490 8672 4554 8676
rect 7972 8604 8036 8668
rect 11836 8876 11900 8940
rect 10848 8732 10912 8736
rect 10848 8676 10852 8732
rect 10852 8676 10908 8732
rect 10908 8676 10912 8732
rect 10848 8672 10912 8676
rect 10928 8732 10992 8736
rect 10928 8676 10932 8732
rect 10932 8676 10988 8732
rect 10988 8676 10992 8732
rect 10928 8672 10992 8676
rect 11008 8732 11072 8736
rect 11008 8676 11012 8732
rect 11012 8676 11068 8732
rect 11068 8676 11072 8732
rect 11008 8672 11072 8676
rect 11088 8732 11152 8736
rect 11088 8676 11092 8732
rect 11092 8676 11148 8732
rect 11148 8676 11152 8732
rect 11088 8672 11152 8676
rect 17445 8732 17509 8736
rect 17445 8676 17449 8732
rect 17449 8676 17505 8732
rect 17505 8676 17509 8732
rect 17445 8672 17509 8676
rect 17525 8732 17589 8736
rect 17525 8676 17529 8732
rect 17529 8676 17585 8732
rect 17585 8676 17589 8732
rect 17525 8672 17589 8676
rect 17605 8732 17669 8736
rect 17605 8676 17609 8732
rect 17609 8676 17665 8732
rect 17665 8676 17669 8732
rect 17605 8672 17669 8676
rect 17685 8732 17749 8736
rect 17685 8676 17689 8732
rect 17689 8676 17745 8732
rect 17745 8676 17749 8732
rect 17685 8672 17749 8676
rect 8156 8332 8220 8396
rect 12388 8332 12452 8396
rect 7549 8188 7613 8192
rect 7549 8132 7553 8188
rect 7553 8132 7609 8188
rect 7609 8132 7613 8188
rect 7549 8128 7613 8132
rect 7629 8188 7693 8192
rect 7629 8132 7633 8188
rect 7633 8132 7689 8188
rect 7689 8132 7693 8188
rect 7629 8128 7693 8132
rect 7709 8188 7773 8192
rect 7709 8132 7713 8188
rect 7713 8132 7769 8188
rect 7769 8132 7773 8188
rect 7709 8128 7773 8132
rect 7789 8188 7853 8192
rect 7789 8132 7793 8188
rect 7793 8132 7849 8188
rect 7849 8132 7853 8188
rect 7789 8128 7853 8132
rect 14146 8188 14210 8192
rect 14146 8132 14150 8188
rect 14150 8132 14206 8188
rect 14206 8132 14210 8188
rect 14146 8128 14210 8132
rect 14226 8188 14290 8192
rect 14226 8132 14230 8188
rect 14230 8132 14286 8188
rect 14286 8132 14290 8188
rect 14226 8128 14290 8132
rect 14306 8188 14370 8192
rect 14306 8132 14310 8188
rect 14310 8132 14366 8188
rect 14366 8132 14370 8188
rect 14306 8128 14370 8132
rect 14386 8188 14450 8192
rect 14386 8132 14390 8188
rect 14390 8132 14446 8188
rect 14446 8132 14450 8188
rect 14386 8128 14450 8132
rect 4250 7644 4314 7648
rect 4250 7588 4254 7644
rect 4254 7588 4310 7644
rect 4310 7588 4314 7644
rect 4250 7584 4314 7588
rect 4330 7644 4394 7648
rect 4330 7588 4334 7644
rect 4334 7588 4390 7644
rect 4390 7588 4394 7644
rect 4330 7584 4394 7588
rect 4410 7644 4474 7648
rect 4410 7588 4414 7644
rect 4414 7588 4470 7644
rect 4470 7588 4474 7644
rect 4410 7584 4474 7588
rect 4490 7644 4554 7648
rect 4490 7588 4494 7644
rect 4494 7588 4550 7644
rect 4550 7588 4554 7644
rect 4490 7584 4554 7588
rect 10848 7644 10912 7648
rect 10848 7588 10852 7644
rect 10852 7588 10908 7644
rect 10908 7588 10912 7644
rect 10848 7584 10912 7588
rect 10928 7644 10992 7648
rect 10928 7588 10932 7644
rect 10932 7588 10988 7644
rect 10988 7588 10992 7644
rect 10928 7584 10992 7588
rect 11008 7644 11072 7648
rect 11008 7588 11012 7644
rect 11012 7588 11068 7644
rect 11068 7588 11072 7644
rect 11008 7584 11072 7588
rect 11088 7644 11152 7648
rect 11088 7588 11092 7644
rect 11092 7588 11148 7644
rect 11148 7588 11152 7644
rect 11088 7584 11152 7588
rect 17445 7644 17509 7648
rect 17445 7588 17449 7644
rect 17449 7588 17505 7644
rect 17505 7588 17509 7644
rect 17445 7584 17509 7588
rect 17525 7644 17589 7648
rect 17525 7588 17529 7644
rect 17529 7588 17585 7644
rect 17585 7588 17589 7644
rect 17525 7584 17589 7588
rect 17605 7644 17669 7648
rect 17605 7588 17609 7644
rect 17609 7588 17665 7644
rect 17665 7588 17669 7644
rect 17605 7584 17669 7588
rect 17685 7644 17749 7648
rect 17685 7588 17689 7644
rect 17689 7588 17745 7644
rect 17745 7588 17749 7644
rect 17685 7584 17749 7588
rect 7549 7100 7613 7104
rect 7549 7044 7553 7100
rect 7553 7044 7609 7100
rect 7609 7044 7613 7100
rect 7549 7040 7613 7044
rect 7629 7100 7693 7104
rect 7629 7044 7633 7100
rect 7633 7044 7689 7100
rect 7689 7044 7693 7100
rect 7629 7040 7693 7044
rect 7709 7100 7773 7104
rect 7709 7044 7713 7100
rect 7713 7044 7769 7100
rect 7769 7044 7773 7100
rect 7709 7040 7773 7044
rect 7789 7100 7853 7104
rect 7789 7044 7793 7100
rect 7793 7044 7849 7100
rect 7849 7044 7853 7100
rect 7789 7040 7853 7044
rect 14146 7100 14210 7104
rect 14146 7044 14150 7100
rect 14150 7044 14206 7100
rect 14206 7044 14210 7100
rect 14146 7040 14210 7044
rect 14226 7100 14290 7104
rect 14226 7044 14230 7100
rect 14230 7044 14286 7100
rect 14286 7044 14290 7100
rect 14226 7040 14290 7044
rect 14306 7100 14370 7104
rect 14306 7044 14310 7100
rect 14310 7044 14366 7100
rect 14366 7044 14370 7100
rect 14306 7040 14370 7044
rect 14386 7100 14450 7104
rect 14386 7044 14390 7100
rect 14390 7044 14446 7100
rect 14446 7044 14450 7100
rect 14386 7040 14450 7044
rect 4250 6556 4314 6560
rect 4250 6500 4254 6556
rect 4254 6500 4310 6556
rect 4310 6500 4314 6556
rect 4250 6496 4314 6500
rect 4330 6556 4394 6560
rect 4330 6500 4334 6556
rect 4334 6500 4390 6556
rect 4390 6500 4394 6556
rect 4330 6496 4394 6500
rect 4410 6556 4474 6560
rect 4410 6500 4414 6556
rect 4414 6500 4470 6556
rect 4470 6500 4474 6556
rect 4410 6496 4474 6500
rect 4490 6556 4554 6560
rect 4490 6500 4494 6556
rect 4494 6500 4550 6556
rect 4550 6500 4554 6556
rect 4490 6496 4554 6500
rect 10848 6556 10912 6560
rect 10848 6500 10852 6556
rect 10852 6500 10908 6556
rect 10908 6500 10912 6556
rect 10848 6496 10912 6500
rect 10928 6556 10992 6560
rect 10928 6500 10932 6556
rect 10932 6500 10988 6556
rect 10988 6500 10992 6556
rect 10928 6496 10992 6500
rect 11008 6556 11072 6560
rect 11008 6500 11012 6556
rect 11012 6500 11068 6556
rect 11068 6500 11072 6556
rect 11008 6496 11072 6500
rect 11088 6556 11152 6560
rect 11088 6500 11092 6556
rect 11092 6500 11148 6556
rect 11148 6500 11152 6556
rect 11088 6496 11152 6500
rect 17445 6556 17509 6560
rect 17445 6500 17449 6556
rect 17449 6500 17505 6556
rect 17505 6500 17509 6556
rect 17445 6496 17509 6500
rect 17525 6556 17589 6560
rect 17525 6500 17529 6556
rect 17529 6500 17585 6556
rect 17585 6500 17589 6556
rect 17525 6496 17589 6500
rect 17605 6556 17669 6560
rect 17605 6500 17609 6556
rect 17609 6500 17665 6556
rect 17665 6500 17669 6556
rect 17605 6496 17669 6500
rect 17685 6556 17749 6560
rect 17685 6500 17689 6556
rect 17689 6500 17745 6556
rect 17745 6500 17749 6556
rect 17685 6496 17749 6500
rect 7549 6012 7613 6016
rect 7549 5956 7553 6012
rect 7553 5956 7609 6012
rect 7609 5956 7613 6012
rect 7549 5952 7613 5956
rect 7629 6012 7693 6016
rect 7629 5956 7633 6012
rect 7633 5956 7689 6012
rect 7689 5956 7693 6012
rect 7629 5952 7693 5956
rect 7709 6012 7773 6016
rect 7709 5956 7713 6012
rect 7713 5956 7769 6012
rect 7769 5956 7773 6012
rect 7709 5952 7773 5956
rect 7789 6012 7853 6016
rect 7789 5956 7793 6012
rect 7793 5956 7849 6012
rect 7849 5956 7853 6012
rect 7789 5952 7853 5956
rect 14146 6012 14210 6016
rect 14146 5956 14150 6012
rect 14150 5956 14206 6012
rect 14206 5956 14210 6012
rect 14146 5952 14210 5956
rect 14226 6012 14290 6016
rect 14226 5956 14230 6012
rect 14230 5956 14286 6012
rect 14286 5956 14290 6012
rect 14226 5952 14290 5956
rect 14306 6012 14370 6016
rect 14306 5956 14310 6012
rect 14310 5956 14366 6012
rect 14366 5956 14370 6012
rect 14306 5952 14370 5956
rect 14386 6012 14450 6016
rect 14386 5956 14390 6012
rect 14390 5956 14446 6012
rect 14446 5956 14450 6012
rect 14386 5952 14450 5956
rect 11468 5536 11532 5540
rect 11468 5480 11482 5536
rect 11482 5480 11532 5536
rect 11468 5476 11532 5480
rect 4250 5468 4314 5472
rect 4250 5412 4254 5468
rect 4254 5412 4310 5468
rect 4310 5412 4314 5468
rect 4250 5408 4314 5412
rect 4330 5468 4394 5472
rect 4330 5412 4334 5468
rect 4334 5412 4390 5468
rect 4390 5412 4394 5468
rect 4330 5408 4394 5412
rect 4410 5468 4474 5472
rect 4410 5412 4414 5468
rect 4414 5412 4470 5468
rect 4470 5412 4474 5468
rect 4410 5408 4474 5412
rect 4490 5468 4554 5472
rect 4490 5412 4494 5468
rect 4494 5412 4550 5468
rect 4550 5412 4554 5468
rect 4490 5408 4554 5412
rect 10848 5468 10912 5472
rect 10848 5412 10852 5468
rect 10852 5412 10908 5468
rect 10908 5412 10912 5468
rect 10848 5408 10912 5412
rect 10928 5468 10992 5472
rect 10928 5412 10932 5468
rect 10932 5412 10988 5468
rect 10988 5412 10992 5468
rect 10928 5408 10992 5412
rect 11008 5468 11072 5472
rect 11008 5412 11012 5468
rect 11012 5412 11068 5468
rect 11068 5412 11072 5468
rect 11008 5408 11072 5412
rect 11088 5468 11152 5472
rect 11088 5412 11092 5468
rect 11092 5412 11148 5468
rect 11148 5412 11152 5468
rect 11088 5408 11152 5412
rect 17445 5468 17509 5472
rect 17445 5412 17449 5468
rect 17449 5412 17505 5468
rect 17505 5412 17509 5468
rect 17445 5408 17509 5412
rect 17525 5468 17589 5472
rect 17525 5412 17529 5468
rect 17529 5412 17585 5468
rect 17585 5412 17589 5468
rect 17525 5408 17589 5412
rect 17605 5468 17669 5472
rect 17605 5412 17609 5468
rect 17609 5412 17665 5468
rect 17665 5412 17669 5468
rect 17605 5408 17669 5412
rect 17685 5468 17749 5472
rect 17685 5412 17689 5468
rect 17689 5412 17745 5468
rect 17745 5412 17749 5468
rect 17685 5408 17749 5412
rect 7549 4924 7613 4928
rect 7549 4868 7553 4924
rect 7553 4868 7609 4924
rect 7609 4868 7613 4924
rect 7549 4864 7613 4868
rect 7629 4924 7693 4928
rect 7629 4868 7633 4924
rect 7633 4868 7689 4924
rect 7689 4868 7693 4924
rect 7629 4864 7693 4868
rect 7709 4924 7773 4928
rect 7709 4868 7713 4924
rect 7713 4868 7769 4924
rect 7769 4868 7773 4924
rect 7709 4864 7773 4868
rect 7789 4924 7853 4928
rect 7789 4868 7793 4924
rect 7793 4868 7849 4924
rect 7849 4868 7853 4924
rect 7789 4864 7853 4868
rect 14146 4924 14210 4928
rect 14146 4868 14150 4924
rect 14150 4868 14206 4924
rect 14206 4868 14210 4924
rect 14146 4864 14210 4868
rect 14226 4924 14290 4928
rect 14226 4868 14230 4924
rect 14230 4868 14286 4924
rect 14286 4868 14290 4924
rect 14226 4864 14290 4868
rect 14306 4924 14370 4928
rect 14306 4868 14310 4924
rect 14310 4868 14366 4924
rect 14366 4868 14370 4924
rect 14306 4864 14370 4868
rect 14386 4924 14450 4928
rect 14386 4868 14390 4924
rect 14390 4868 14446 4924
rect 14446 4868 14450 4924
rect 14386 4864 14450 4868
rect 4250 4380 4314 4384
rect 4250 4324 4254 4380
rect 4254 4324 4310 4380
rect 4310 4324 4314 4380
rect 4250 4320 4314 4324
rect 4330 4380 4394 4384
rect 4330 4324 4334 4380
rect 4334 4324 4390 4380
rect 4390 4324 4394 4380
rect 4330 4320 4394 4324
rect 4410 4380 4474 4384
rect 4410 4324 4414 4380
rect 4414 4324 4470 4380
rect 4470 4324 4474 4380
rect 4410 4320 4474 4324
rect 4490 4380 4554 4384
rect 4490 4324 4494 4380
rect 4494 4324 4550 4380
rect 4550 4324 4554 4380
rect 4490 4320 4554 4324
rect 10848 4380 10912 4384
rect 10848 4324 10852 4380
rect 10852 4324 10908 4380
rect 10908 4324 10912 4380
rect 10848 4320 10912 4324
rect 10928 4380 10992 4384
rect 10928 4324 10932 4380
rect 10932 4324 10988 4380
rect 10988 4324 10992 4380
rect 10928 4320 10992 4324
rect 11008 4380 11072 4384
rect 11008 4324 11012 4380
rect 11012 4324 11068 4380
rect 11068 4324 11072 4380
rect 11008 4320 11072 4324
rect 11088 4380 11152 4384
rect 11088 4324 11092 4380
rect 11092 4324 11148 4380
rect 11148 4324 11152 4380
rect 11088 4320 11152 4324
rect 17445 4380 17509 4384
rect 17445 4324 17449 4380
rect 17449 4324 17505 4380
rect 17505 4324 17509 4380
rect 17445 4320 17509 4324
rect 17525 4380 17589 4384
rect 17525 4324 17529 4380
rect 17529 4324 17585 4380
rect 17585 4324 17589 4380
rect 17525 4320 17589 4324
rect 17605 4380 17669 4384
rect 17605 4324 17609 4380
rect 17609 4324 17665 4380
rect 17665 4324 17669 4380
rect 17605 4320 17669 4324
rect 17685 4380 17749 4384
rect 17685 4324 17689 4380
rect 17689 4324 17745 4380
rect 17745 4324 17749 4380
rect 17685 4320 17749 4324
rect 7549 3836 7613 3840
rect 7549 3780 7553 3836
rect 7553 3780 7609 3836
rect 7609 3780 7613 3836
rect 7549 3776 7613 3780
rect 7629 3836 7693 3840
rect 7629 3780 7633 3836
rect 7633 3780 7689 3836
rect 7689 3780 7693 3836
rect 7629 3776 7693 3780
rect 7709 3836 7773 3840
rect 7709 3780 7713 3836
rect 7713 3780 7769 3836
rect 7769 3780 7773 3836
rect 7709 3776 7773 3780
rect 7789 3836 7853 3840
rect 7789 3780 7793 3836
rect 7793 3780 7849 3836
rect 7849 3780 7853 3836
rect 7789 3776 7853 3780
rect 14146 3836 14210 3840
rect 14146 3780 14150 3836
rect 14150 3780 14206 3836
rect 14206 3780 14210 3836
rect 14146 3776 14210 3780
rect 14226 3836 14290 3840
rect 14226 3780 14230 3836
rect 14230 3780 14286 3836
rect 14286 3780 14290 3836
rect 14226 3776 14290 3780
rect 14306 3836 14370 3840
rect 14306 3780 14310 3836
rect 14310 3780 14366 3836
rect 14366 3780 14370 3836
rect 14306 3776 14370 3780
rect 14386 3836 14450 3840
rect 14386 3780 14390 3836
rect 14390 3780 14446 3836
rect 14446 3780 14450 3836
rect 14386 3776 14450 3780
rect 11468 3436 11532 3500
rect 4250 3292 4314 3296
rect 4250 3236 4254 3292
rect 4254 3236 4310 3292
rect 4310 3236 4314 3292
rect 4250 3232 4314 3236
rect 4330 3292 4394 3296
rect 4330 3236 4334 3292
rect 4334 3236 4390 3292
rect 4390 3236 4394 3292
rect 4330 3232 4394 3236
rect 4410 3292 4474 3296
rect 4410 3236 4414 3292
rect 4414 3236 4470 3292
rect 4470 3236 4474 3292
rect 4410 3232 4474 3236
rect 4490 3292 4554 3296
rect 4490 3236 4494 3292
rect 4494 3236 4550 3292
rect 4550 3236 4554 3292
rect 4490 3232 4554 3236
rect 10848 3292 10912 3296
rect 10848 3236 10852 3292
rect 10852 3236 10908 3292
rect 10908 3236 10912 3292
rect 10848 3232 10912 3236
rect 10928 3292 10992 3296
rect 10928 3236 10932 3292
rect 10932 3236 10988 3292
rect 10988 3236 10992 3292
rect 10928 3232 10992 3236
rect 11008 3292 11072 3296
rect 11008 3236 11012 3292
rect 11012 3236 11068 3292
rect 11068 3236 11072 3292
rect 11008 3232 11072 3236
rect 11088 3292 11152 3296
rect 11088 3236 11092 3292
rect 11092 3236 11148 3292
rect 11148 3236 11152 3292
rect 11088 3232 11152 3236
rect 17445 3292 17509 3296
rect 17445 3236 17449 3292
rect 17449 3236 17505 3292
rect 17505 3236 17509 3292
rect 17445 3232 17509 3236
rect 17525 3292 17589 3296
rect 17525 3236 17529 3292
rect 17529 3236 17585 3292
rect 17585 3236 17589 3292
rect 17525 3232 17589 3236
rect 17605 3292 17669 3296
rect 17605 3236 17609 3292
rect 17609 3236 17665 3292
rect 17665 3236 17669 3292
rect 17605 3232 17669 3236
rect 17685 3292 17749 3296
rect 17685 3236 17689 3292
rect 17689 3236 17745 3292
rect 17745 3236 17749 3292
rect 17685 3232 17749 3236
rect 7549 2748 7613 2752
rect 7549 2692 7553 2748
rect 7553 2692 7609 2748
rect 7609 2692 7613 2748
rect 7549 2688 7613 2692
rect 7629 2748 7693 2752
rect 7629 2692 7633 2748
rect 7633 2692 7689 2748
rect 7689 2692 7693 2748
rect 7629 2688 7693 2692
rect 7709 2748 7773 2752
rect 7709 2692 7713 2748
rect 7713 2692 7769 2748
rect 7769 2692 7773 2748
rect 7709 2688 7773 2692
rect 7789 2748 7853 2752
rect 7789 2692 7793 2748
rect 7793 2692 7849 2748
rect 7849 2692 7853 2748
rect 7789 2688 7853 2692
rect 14146 2748 14210 2752
rect 14146 2692 14150 2748
rect 14150 2692 14206 2748
rect 14206 2692 14210 2748
rect 14146 2688 14210 2692
rect 14226 2748 14290 2752
rect 14226 2692 14230 2748
rect 14230 2692 14286 2748
rect 14286 2692 14290 2748
rect 14226 2688 14290 2692
rect 14306 2748 14370 2752
rect 14306 2692 14310 2748
rect 14310 2692 14366 2748
rect 14366 2692 14370 2748
rect 14306 2688 14370 2692
rect 14386 2748 14450 2752
rect 14386 2692 14390 2748
rect 14390 2692 14446 2748
rect 14446 2692 14450 2748
rect 14386 2688 14450 2692
rect 4250 2204 4314 2208
rect 4250 2148 4254 2204
rect 4254 2148 4310 2204
rect 4310 2148 4314 2204
rect 4250 2144 4314 2148
rect 4330 2204 4394 2208
rect 4330 2148 4334 2204
rect 4334 2148 4390 2204
rect 4390 2148 4394 2204
rect 4330 2144 4394 2148
rect 4410 2204 4474 2208
rect 4410 2148 4414 2204
rect 4414 2148 4470 2204
rect 4470 2148 4474 2204
rect 4410 2144 4474 2148
rect 4490 2204 4554 2208
rect 4490 2148 4494 2204
rect 4494 2148 4550 2204
rect 4550 2148 4554 2204
rect 4490 2144 4554 2148
rect 10848 2204 10912 2208
rect 10848 2148 10852 2204
rect 10852 2148 10908 2204
rect 10908 2148 10912 2204
rect 10848 2144 10912 2148
rect 10928 2204 10992 2208
rect 10928 2148 10932 2204
rect 10932 2148 10988 2204
rect 10988 2148 10992 2204
rect 10928 2144 10992 2148
rect 11008 2204 11072 2208
rect 11008 2148 11012 2204
rect 11012 2148 11068 2204
rect 11068 2148 11072 2204
rect 11008 2144 11072 2148
rect 11088 2204 11152 2208
rect 11088 2148 11092 2204
rect 11092 2148 11148 2204
rect 11148 2148 11152 2204
rect 11088 2144 11152 2148
rect 17445 2204 17509 2208
rect 17445 2148 17449 2204
rect 17449 2148 17505 2204
rect 17505 2148 17509 2204
rect 17445 2144 17509 2148
rect 17525 2204 17589 2208
rect 17525 2148 17529 2204
rect 17529 2148 17585 2204
rect 17585 2148 17589 2204
rect 17525 2144 17589 2148
rect 17605 2204 17669 2208
rect 17605 2148 17609 2204
rect 17609 2148 17665 2204
rect 17665 2148 17669 2204
rect 17605 2144 17669 2148
rect 17685 2204 17749 2208
rect 17685 2148 17689 2204
rect 17689 2148 17745 2204
rect 17745 2148 17749 2204
rect 17685 2144 17749 2148
<< metal4 >>
rect 4242 19616 4563 19632
rect 4242 19552 4250 19616
rect 4314 19552 4330 19616
rect 4394 19552 4410 19616
rect 4474 19552 4490 19616
rect 4554 19552 4563 19616
rect 4242 18528 4563 19552
rect 4242 18464 4250 18528
rect 4314 18464 4330 18528
rect 4394 18464 4410 18528
rect 4474 18464 4490 18528
rect 4554 18464 4563 18528
rect 4242 17440 4563 18464
rect 4242 17376 4250 17440
rect 4314 17376 4330 17440
rect 4394 17376 4410 17440
rect 4474 17376 4490 17440
rect 4554 17376 4563 17440
rect 4242 16352 4563 17376
rect 4242 16288 4250 16352
rect 4314 16288 4330 16352
rect 4394 16288 4410 16352
rect 4474 16288 4490 16352
rect 4554 16288 4563 16352
rect 4242 15264 4563 16288
rect 4242 15200 4250 15264
rect 4314 15200 4330 15264
rect 4394 15200 4410 15264
rect 4474 15200 4490 15264
rect 4554 15200 4563 15264
rect 4242 14176 4563 15200
rect 4242 14112 4250 14176
rect 4314 14112 4330 14176
rect 4394 14112 4410 14176
rect 4474 14112 4490 14176
rect 4554 14112 4563 14176
rect 4242 13088 4563 14112
rect 4242 13024 4250 13088
rect 4314 13024 4330 13088
rect 4394 13024 4410 13088
rect 4474 13024 4490 13088
rect 4554 13024 4563 13088
rect 4242 12000 4563 13024
rect 4242 11936 4250 12000
rect 4314 11936 4330 12000
rect 4394 11936 4410 12000
rect 4474 11936 4490 12000
rect 4554 11936 4563 12000
rect 4242 10912 4563 11936
rect 4242 10848 4250 10912
rect 4314 10848 4330 10912
rect 4394 10848 4410 10912
rect 4474 10848 4490 10912
rect 4554 10848 4563 10912
rect 4242 9824 4563 10848
rect 4242 9760 4250 9824
rect 4314 9760 4330 9824
rect 4394 9760 4410 9824
rect 4474 9760 4490 9824
rect 4554 9760 4563 9824
rect 4242 8736 4563 9760
rect 4242 8672 4250 8736
rect 4314 8672 4330 8736
rect 4394 8672 4410 8736
rect 4474 8672 4490 8736
rect 4554 8672 4563 8736
rect 4242 7648 4563 8672
rect 4242 7584 4250 7648
rect 4314 7584 4330 7648
rect 4394 7584 4410 7648
rect 4474 7584 4490 7648
rect 4554 7584 4563 7648
rect 4242 6560 4563 7584
rect 4242 6496 4250 6560
rect 4314 6496 4330 6560
rect 4394 6496 4410 6560
rect 4474 6496 4490 6560
rect 4554 6496 4563 6560
rect 4242 5472 4563 6496
rect 4242 5408 4250 5472
rect 4314 5408 4330 5472
rect 4394 5408 4410 5472
rect 4474 5408 4490 5472
rect 4554 5408 4563 5472
rect 4242 4384 4563 5408
rect 4242 4320 4250 4384
rect 4314 4320 4330 4384
rect 4394 4320 4410 4384
rect 4474 4320 4490 4384
rect 4554 4320 4563 4384
rect 4242 3296 4563 4320
rect 4242 3232 4250 3296
rect 4314 3232 4330 3296
rect 4394 3232 4410 3296
rect 4474 3232 4490 3296
rect 4554 3232 4563 3296
rect 4242 2208 4563 3232
rect 4242 2144 4250 2208
rect 4314 2144 4330 2208
rect 4394 2144 4410 2208
rect 4474 2144 4490 2208
rect 4554 2144 4563 2208
rect 4242 2128 4563 2144
rect 7541 19072 7861 19632
rect 7541 19008 7549 19072
rect 7613 19008 7629 19072
rect 7693 19008 7709 19072
rect 7773 19008 7789 19072
rect 7853 19008 7861 19072
rect 7541 17984 7861 19008
rect 7541 17920 7549 17984
rect 7613 17920 7629 17984
rect 7693 17920 7709 17984
rect 7773 17920 7789 17984
rect 7853 17920 7861 17984
rect 7541 16896 7861 17920
rect 7541 16832 7549 16896
rect 7613 16832 7629 16896
rect 7693 16832 7709 16896
rect 7773 16832 7789 16896
rect 7853 16832 7861 16896
rect 7541 15808 7861 16832
rect 7541 15744 7549 15808
rect 7613 15744 7629 15808
rect 7693 15744 7709 15808
rect 7773 15744 7789 15808
rect 7853 15744 7861 15808
rect 7541 14720 7861 15744
rect 7541 14656 7549 14720
rect 7613 14656 7629 14720
rect 7693 14656 7709 14720
rect 7773 14656 7789 14720
rect 7853 14656 7861 14720
rect 7541 13632 7861 14656
rect 7541 13568 7549 13632
rect 7613 13568 7629 13632
rect 7693 13568 7709 13632
rect 7773 13568 7789 13632
rect 7853 13568 7861 13632
rect 7541 12544 7861 13568
rect 7541 12480 7549 12544
rect 7613 12480 7629 12544
rect 7693 12480 7709 12544
rect 7773 12480 7789 12544
rect 7853 12480 7861 12544
rect 7541 11456 7861 12480
rect 7541 11392 7549 11456
rect 7613 11392 7629 11456
rect 7693 11392 7709 11456
rect 7773 11392 7789 11456
rect 7853 11392 7861 11456
rect 7541 10368 7861 11392
rect 7541 10304 7549 10368
rect 7613 10304 7629 10368
rect 7693 10304 7709 10368
rect 7773 10304 7789 10368
rect 7853 10304 7861 10368
rect 7541 9280 7861 10304
rect 7541 9216 7549 9280
rect 7613 9216 7629 9280
rect 7693 9216 7709 9280
rect 7773 9216 7789 9280
rect 7853 9216 7861 9280
rect 7541 8192 7861 9216
rect 10840 19616 11160 19632
rect 10840 19552 10848 19616
rect 10912 19552 10928 19616
rect 10992 19552 11008 19616
rect 11072 19552 11088 19616
rect 11152 19552 11160 19616
rect 10840 18528 11160 19552
rect 10840 18464 10848 18528
rect 10912 18464 10928 18528
rect 10992 18464 11008 18528
rect 11072 18464 11088 18528
rect 11152 18464 11160 18528
rect 10840 17440 11160 18464
rect 10840 17376 10848 17440
rect 10912 17376 10928 17440
rect 10992 17376 11008 17440
rect 11072 17376 11088 17440
rect 11152 17376 11160 17440
rect 10840 16352 11160 17376
rect 10840 16288 10848 16352
rect 10912 16288 10928 16352
rect 10992 16288 11008 16352
rect 11072 16288 11088 16352
rect 11152 16288 11160 16352
rect 10840 15264 11160 16288
rect 10840 15200 10848 15264
rect 10912 15200 10928 15264
rect 10992 15200 11008 15264
rect 11072 15200 11088 15264
rect 11152 15200 11160 15264
rect 10840 14176 11160 15200
rect 10840 14112 10848 14176
rect 10912 14112 10928 14176
rect 10992 14112 11008 14176
rect 11072 14112 11088 14176
rect 11152 14112 11160 14176
rect 10840 13088 11160 14112
rect 10840 13024 10848 13088
rect 10912 13024 10928 13088
rect 10992 13024 11008 13088
rect 11072 13024 11088 13088
rect 11152 13024 11160 13088
rect 10840 12000 11160 13024
rect 10840 11936 10848 12000
rect 10912 11936 10928 12000
rect 10992 11936 11008 12000
rect 11072 11936 11088 12000
rect 11152 11936 11160 12000
rect 10840 10912 11160 11936
rect 10840 10848 10848 10912
rect 10912 10848 10928 10912
rect 10992 10848 11008 10912
rect 11072 10848 11088 10912
rect 11152 10848 11160 10912
rect 10840 9824 11160 10848
rect 10840 9760 10848 9824
rect 10912 9760 10928 9824
rect 10992 9760 11008 9824
rect 11072 9760 11088 9824
rect 11152 9760 11160 9824
rect 10840 8736 11160 9760
rect 14138 19072 14458 19632
rect 14138 19008 14146 19072
rect 14210 19008 14226 19072
rect 14290 19008 14306 19072
rect 14370 19008 14386 19072
rect 14450 19008 14458 19072
rect 14138 17984 14458 19008
rect 17437 19616 17757 19632
rect 17437 19552 17445 19616
rect 17509 19552 17525 19616
rect 17589 19552 17605 19616
rect 17669 19552 17685 19616
rect 17749 19552 17757 19616
rect 17437 18528 17757 19552
rect 17437 18464 17445 18528
rect 17509 18464 17525 18528
rect 17589 18464 17605 18528
rect 17669 18464 17685 18528
rect 17749 18464 17757 18528
rect 14963 18052 15029 18053
rect 14963 17988 14964 18052
rect 15028 17988 15029 18052
rect 14963 17987 15029 17988
rect 14138 17920 14146 17984
rect 14210 17920 14226 17984
rect 14290 17920 14306 17984
rect 14370 17920 14386 17984
rect 14450 17920 14458 17984
rect 14138 16896 14458 17920
rect 14138 16832 14146 16896
rect 14210 16832 14226 16896
rect 14290 16832 14306 16896
rect 14370 16832 14386 16896
rect 14450 16832 14458 16896
rect 14138 15808 14458 16832
rect 14966 16557 15026 17987
rect 17437 17440 17757 18464
rect 17437 17376 17445 17440
rect 17509 17376 17525 17440
rect 17589 17376 17605 17440
rect 17669 17376 17685 17440
rect 17749 17376 17757 17440
rect 14963 16556 15029 16557
rect 14963 16492 14964 16556
rect 15028 16492 15029 16556
rect 14963 16491 15029 16492
rect 14138 15744 14146 15808
rect 14210 15744 14226 15808
rect 14290 15744 14306 15808
rect 14370 15744 14386 15808
rect 14450 15744 14458 15808
rect 14138 14720 14458 15744
rect 14138 14656 14146 14720
rect 14210 14656 14226 14720
rect 14290 14656 14306 14720
rect 14370 14656 14386 14720
rect 14450 14656 14458 14720
rect 14138 13632 14458 14656
rect 14138 13568 14146 13632
rect 14210 13568 14226 13632
rect 14290 13568 14306 13632
rect 14370 13568 14386 13632
rect 14450 13568 14458 13632
rect 14138 12544 14458 13568
rect 14138 12480 14146 12544
rect 14210 12480 14226 12544
rect 14290 12480 14306 12544
rect 14370 12480 14386 12544
rect 14450 12480 14458 12544
rect 14138 11456 14458 12480
rect 14138 11392 14146 11456
rect 14210 11392 14226 11456
rect 14290 11392 14306 11456
rect 14370 11392 14386 11456
rect 14450 11392 14458 11456
rect 14138 10368 14458 11392
rect 14138 10304 14146 10368
rect 14210 10304 14226 10368
rect 14290 10304 14306 10368
rect 14370 10304 14386 10368
rect 14450 10304 14458 10368
rect 11835 9620 11901 9621
rect 11835 9556 11836 9620
rect 11900 9556 11901 9620
rect 11835 9555 11901 9556
rect 11838 8941 11898 9555
rect 14138 9280 14458 10304
rect 14138 9216 14146 9280
rect 14210 9216 14226 9280
rect 14290 9216 14306 9280
rect 14370 9216 14386 9280
rect 14450 9216 14458 9280
rect 12387 9076 12453 9077
rect 12387 9012 12388 9076
rect 12452 9012 12453 9076
rect 12387 9011 12453 9012
rect 11835 8940 11901 8941
rect 11835 8876 11836 8940
rect 11900 8876 11901 8940
rect 11835 8875 11901 8876
rect 10840 8672 10848 8736
rect 10912 8672 10928 8736
rect 10992 8672 11008 8736
rect 11072 8672 11088 8736
rect 11152 8672 11160 8736
rect 7971 8668 8037 8669
rect 7971 8604 7972 8668
rect 8036 8604 8037 8668
rect 7971 8603 8037 8604
rect 7974 8394 8034 8603
rect 8155 8396 8221 8397
rect 8155 8394 8156 8396
rect 7974 8334 8156 8394
rect 8155 8332 8156 8334
rect 8220 8332 8221 8396
rect 8155 8331 8221 8332
rect 7541 8128 7549 8192
rect 7613 8128 7629 8192
rect 7693 8128 7709 8192
rect 7773 8128 7789 8192
rect 7853 8128 7861 8192
rect 7541 7104 7861 8128
rect 7541 7040 7549 7104
rect 7613 7040 7629 7104
rect 7693 7040 7709 7104
rect 7773 7040 7789 7104
rect 7853 7040 7861 7104
rect 7541 6016 7861 7040
rect 7541 5952 7549 6016
rect 7613 5952 7629 6016
rect 7693 5952 7709 6016
rect 7773 5952 7789 6016
rect 7853 5952 7861 6016
rect 7541 4928 7861 5952
rect 7541 4864 7549 4928
rect 7613 4864 7629 4928
rect 7693 4864 7709 4928
rect 7773 4864 7789 4928
rect 7853 4864 7861 4928
rect 7541 3840 7861 4864
rect 7541 3776 7549 3840
rect 7613 3776 7629 3840
rect 7693 3776 7709 3840
rect 7773 3776 7789 3840
rect 7853 3776 7861 3840
rect 7541 2752 7861 3776
rect 7541 2688 7549 2752
rect 7613 2688 7629 2752
rect 7693 2688 7709 2752
rect 7773 2688 7789 2752
rect 7853 2688 7861 2752
rect 7541 2128 7861 2688
rect 10840 7648 11160 8672
rect 12390 8397 12450 9011
rect 12387 8396 12453 8397
rect 12387 8332 12388 8396
rect 12452 8332 12453 8396
rect 12387 8331 12453 8332
rect 10840 7584 10848 7648
rect 10912 7584 10928 7648
rect 10992 7584 11008 7648
rect 11072 7584 11088 7648
rect 11152 7584 11160 7648
rect 10840 6560 11160 7584
rect 10840 6496 10848 6560
rect 10912 6496 10928 6560
rect 10992 6496 11008 6560
rect 11072 6496 11088 6560
rect 11152 6496 11160 6560
rect 10840 5472 11160 6496
rect 14138 8192 14458 9216
rect 14138 8128 14146 8192
rect 14210 8128 14226 8192
rect 14290 8128 14306 8192
rect 14370 8128 14386 8192
rect 14450 8128 14458 8192
rect 14138 7104 14458 8128
rect 14138 7040 14146 7104
rect 14210 7040 14226 7104
rect 14290 7040 14306 7104
rect 14370 7040 14386 7104
rect 14450 7040 14458 7104
rect 14138 6016 14458 7040
rect 14138 5952 14146 6016
rect 14210 5952 14226 6016
rect 14290 5952 14306 6016
rect 14370 5952 14386 6016
rect 14450 5952 14458 6016
rect 11467 5540 11533 5541
rect 11467 5476 11468 5540
rect 11532 5476 11533 5540
rect 11467 5475 11533 5476
rect 10840 5408 10848 5472
rect 10912 5408 10928 5472
rect 10992 5408 11008 5472
rect 11072 5408 11088 5472
rect 11152 5408 11160 5472
rect 10840 4384 11160 5408
rect 10840 4320 10848 4384
rect 10912 4320 10928 4384
rect 10992 4320 11008 4384
rect 11072 4320 11088 4384
rect 11152 4320 11160 4384
rect 10840 3296 11160 4320
rect 11470 3501 11530 5475
rect 14138 4928 14458 5952
rect 14138 4864 14146 4928
rect 14210 4864 14226 4928
rect 14290 4864 14306 4928
rect 14370 4864 14386 4928
rect 14450 4864 14458 4928
rect 14138 3840 14458 4864
rect 14138 3776 14146 3840
rect 14210 3776 14226 3840
rect 14290 3776 14306 3840
rect 14370 3776 14386 3840
rect 14450 3776 14458 3840
rect 11467 3500 11533 3501
rect 11467 3436 11468 3500
rect 11532 3436 11533 3500
rect 11467 3435 11533 3436
rect 10840 3232 10848 3296
rect 10912 3232 10928 3296
rect 10992 3232 11008 3296
rect 11072 3232 11088 3296
rect 11152 3232 11160 3296
rect 10840 2208 11160 3232
rect 10840 2144 10848 2208
rect 10912 2144 10928 2208
rect 10992 2144 11008 2208
rect 11072 2144 11088 2208
rect 11152 2144 11160 2208
rect 10840 2128 11160 2144
rect 14138 2752 14458 3776
rect 14138 2688 14146 2752
rect 14210 2688 14226 2752
rect 14290 2688 14306 2752
rect 14370 2688 14386 2752
rect 14450 2688 14458 2752
rect 14138 2128 14458 2688
rect 17437 16352 17757 17376
rect 17437 16288 17445 16352
rect 17509 16288 17525 16352
rect 17589 16288 17605 16352
rect 17669 16288 17685 16352
rect 17749 16288 17757 16352
rect 17437 15264 17757 16288
rect 17437 15200 17445 15264
rect 17509 15200 17525 15264
rect 17589 15200 17605 15264
rect 17669 15200 17685 15264
rect 17749 15200 17757 15264
rect 17437 14176 17757 15200
rect 17437 14112 17445 14176
rect 17509 14112 17525 14176
rect 17589 14112 17605 14176
rect 17669 14112 17685 14176
rect 17749 14112 17757 14176
rect 17437 13088 17757 14112
rect 17437 13024 17445 13088
rect 17509 13024 17525 13088
rect 17589 13024 17605 13088
rect 17669 13024 17685 13088
rect 17749 13024 17757 13088
rect 17437 12000 17757 13024
rect 17437 11936 17445 12000
rect 17509 11936 17525 12000
rect 17589 11936 17605 12000
rect 17669 11936 17685 12000
rect 17749 11936 17757 12000
rect 17437 10912 17757 11936
rect 17437 10848 17445 10912
rect 17509 10848 17525 10912
rect 17589 10848 17605 10912
rect 17669 10848 17685 10912
rect 17749 10848 17757 10912
rect 17437 9824 17757 10848
rect 17437 9760 17445 9824
rect 17509 9760 17525 9824
rect 17589 9760 17605 9824
rect 17669 9760 17685 9824
rect 17749 9760 17757 9824
rect 17437 8736 17757 9760
rect 17437 8672 17445 8736
rect 17509 8672 17525 8736
rect 17589 8672 17605 8736
rect 17669 8672 17685 8736
rect 17749 8672 17757 8736
rect 17437 7648 17757 8672
rect 17437 7584 17445 7648
rect 17509 7584 17525 7648
rect 17589 7584 17605 7648
rect 17669 7584 17685 7648
rect 17749 7584 17757 7648
rect 17437 6560 17757 7584
rect 17437 6496 17445 6560
rect 17509 6496 17525 6560
rect 17589 6496 17605 6560
rect 17669 6496 17685 6560
rect 17749 6496 17757 6560
rect 17437 5472 17757 6496
rect 17437 5408 17445 5472
rect 17509 5408 17525 5472
rect 17589 5408 17605 5472
rect 17669 5408 17685 5472
rect 17749 5408 17757 5472
rect 17437 4384 17757 5408
rect 17437 4320 17445 4384
rect 17509 4320 17525 4384
rect 17589 4320 17605 4384
rect 17669 4320 17685 4384
rect 17749 4320 17757 4384
rect 17437 3296 17757 4320
rect 17437 3232 17445 3296
rect 17509 3232 17525 3296
rect 17589 3232 17605 3296
rect 17669 3232 17685 3296
rect 17749 3232 17757 3296
rect 17437 2208 17757 3232
rect 17437 2144 17445 2208
rect 17509 2144 17525 2208
rect 17589 2144 17605 2208
rect 17669 2144 17685 2208
rect 17749 2144 17757 2208
rect 17437 2128 17757 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _64_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5060 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4416 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40
timestamp 1604681595
transform 1 0 4784 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_35 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 5980 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5244 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5336 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52
timestamp 1604681595
transform 1 0 5888 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8372 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 8280 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10304 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10212 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1604681595
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1604681595
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98
timestamp 1604681595
transform 1 0 10120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_94
timestamp 1604681595
transform 1 0 9752 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11684 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp 1604681595
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13892 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13892 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16928 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 15456 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 15916 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_160
timestamp 1604681595
transform 1 0 15824 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_155
timestamp 1604681595
transform 1 0 15364 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _67_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18308 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 18676 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 19780 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 20884 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 20884 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1604681595
transform 1 0 20148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1604681595
transform 1 0 20516 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_52
timestamp 1604681595
transform 1 0 5888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 8096 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_71
timestamp 1604681595
transform 1 0 7636 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_75
timestamp 1604681595
transform 1 0 8004 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_102
timestamp 1604681595
transform 1 0 10488 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 12696 0 -1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_147
timestamp 1604681595
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 15548 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 17020 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 18492 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 19136 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1604681595
transform 1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 4416 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_35
timestamp 1604681595
transform 1 0 4324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 5888 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8372 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_75
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 13892 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14996 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14168 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 17112 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 15916 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_160
timestamp 1604681595
transform 1 0 15824 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_193
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 20884 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 4508 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1604681595
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5980 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 7636 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11592 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_123
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13432 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_prog_clk
timestamp 1604681595
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 16100 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 19136 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 17572 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1604681595
transform 1 0 19044 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 4600 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_35
timestamp 1604681595
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 6900 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 6256 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1604681595
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1604681595
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7268 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 8924 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8096 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9292 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1604681595
transform 1 0 11040 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11408 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1604681595
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13616 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17112 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 19504 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 20884 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_209
timestamp 1604681595
transform 1 0 20332 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_21
timestamp 1604681595
transform 1 0 3036 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3128 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 4508 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_prog_clk
timestamp 1604681595
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6348 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 5980 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8096 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9108 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_6_75
timestamp 1604681595
transform 1 0 8004 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 11040 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10580 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_prog_clk
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_103
timestamp 1604681595
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1604681595
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13616 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_148
timestamp 1604681595
transform 1 0 14720 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_152
timestamp 1604681595
transform 1 0 15088 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16744 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15180 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 17572 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 18124 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 18676 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_prog_clk
timestamp 1604681595
transform 1 0 18400 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_183
timestamp 1604681595
transform 1 0 17940 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 19596 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 20148 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 20884 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_210
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 4876 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_40
timestamp 1604681595
transform 1 0 4784 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 6624 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7084 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 6348 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8740 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_81
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10028 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11500 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1604681595
transform 1 0 13340 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1604681595
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17020 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16192 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_163
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 19136 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 18768 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 18492 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 1604681595
transform 1 0 20332 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1604681595
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 5244 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8556 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10856 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 9384 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_9_139
timestamp 1604681595
transform 1 0 13892 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16100 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1604681595
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 20332 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19504 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 20884 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_21
timestamp 1604681595
transform 1 0 3036 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4600 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3128 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 5428 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1604681595
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 8096 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 9752 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12236 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1604681595
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13708 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 16100 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18308 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19136 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 4876 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3220 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 6900 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 8464 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_79
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_96
timestamp 1604681595
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 14076 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 14904 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16928 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1604681595
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1604681595
transform 1 0 20332 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 20884 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1604681595
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_205
timestamp 1604681595
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2300 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1604681595
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 4324 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3128 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_prog_clk
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 5796 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 7268 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 8740 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10212 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 11040 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1604681595
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 12512 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 14352 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16744 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 18768 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 18400 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17572 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19136 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1604681595
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1604681595
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 3772 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_prog_clk
timestamp 1604681595
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5520 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 6532 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 5244 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_57
timestamp 1604681595
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_63
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 7820 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 7820 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 8740 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1604681595
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_82
timestamp 1604681595
transform 1 0 8648 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 9752 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 9292 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 10120 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11592 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12880 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1604681595
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_127
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 13708 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_136
timestamp 1604681595
transform 1 0 13616 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604681595
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 15548 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15364 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16008 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1604681595
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 17848 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 18216 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18584 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 20056 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19780 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 20884 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_210
timestamp 1604681595
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 4324 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1604681595
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 8648 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_80
timestamp 1604681595
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk
timestamp 1604681595
transform 1 0 10304 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 13892 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15364 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_prog_clk
timestamp 1604681595
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1604681595
transform 1 0 20332 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19504 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 20884 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2852 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_prog_clk
timestamp 1604681595
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 5704 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6072 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1604681595
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 8740 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 7544 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 9936 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 11408 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 12236 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 13064 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 14536 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 17020 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_prog_clk
timestamp 1604681595
transform 1 0 16744 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1604681595
transform 1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19136 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17388 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2668 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 3496 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5888 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 5520 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_47
timestamp 1604681595
transform 1 0 5428 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8280 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1604681595
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 10304 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10672 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_98
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 12512 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 14904 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_149
timestamp 1604681595
transform 1 0 14812 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 16468 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_166
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19780 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 20884 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_200
timestamp 1604681595
transform 1 0 19504 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_prog_clk
timestamp 1604681595
transform 1 0 2852 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 3128 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 4140 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 5612 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 5980 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 7728 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 10580 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1604681595
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 12512 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16744 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17572 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18860 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_192
timestamp 1604681595
transform 1 0 18768 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1604681595
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 2852 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 2944 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 1472 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4232 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 4416 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 5060 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5888 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8188 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8280 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 11040 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_109
timestamp 1604681595
transform 1 0 11132 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 12696 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11500 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12880 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 13064 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1604681595
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14444 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_144
timestamp 1604681595
transform 1 0 14352 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16744 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16744 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15640 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 15272 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 16468 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 17572 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18400 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18124 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19044 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_194
timestamp 1604681595
transform 1 0 18952 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 20884 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_211
timestamp 1604681595
transform 1 0 20516 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1604681595
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 1656 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 3128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 3496 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 6900 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604681595
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7452 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_21_68
timestamp 1604681595
transform 1 0 7360 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1604681595
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10672 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _61_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 13156 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 12788 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_126
timestamp 1604681595
transform 1 0 12696 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_130
timestamp 1604681595
transform 1 0 13064 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 15088 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 16928 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 15456 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18216 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 19044 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 20884 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_211
timestamp 1604681595
transform 1 0 20516 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 2852 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 5796 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_50
timestamp 1604681595
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7268 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _62_
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10304 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11776 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13524 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 15364 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 15732 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 18676 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 17204 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 20148 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 3036 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 1472 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_20
timestamp 1604681595
transform 1 0 2944 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4876 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 3404 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8280 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _60_
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10856 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9752 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 12788 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13156 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_prog_clk
timestamp 1604681595
transform 1 0 11684 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_prog_clk
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_126
timestamp 1604681595
transform 1 0 12696 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 14996 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 15364 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 16192 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18308 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_prog_clk
timestamp 1604681595
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 20884 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5520 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6992 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1604681595
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_109
timestamp 1604681595
transform 1 0 11132 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11500 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 15456 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 17112 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_172
timestamp 1604681595
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 1840 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_prog_clk
timestamp 1604681595
transform 1 0 3312 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 6900 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 6256 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1604681595
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 8096 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7268 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1604681595
transform 1 0 10028 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 10304 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1604681595
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 14536 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 16008 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1604681595
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 19504 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_209
timestamp 1604681595
transform 1 0 20332 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 1748 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4508 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4048 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 3220 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4876 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 4140 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1604681595
transform 1 0 6532 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5336 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 6164 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5704 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6900 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 7636 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 8372 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1604681595
transform 1 0 10580 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10856 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 10212 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11592 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12512 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_123
timestamp 1604681595
transform 1 0 12420 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13984 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16560 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_163
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_158
timestamp 1604681595
transform 1 0 15640 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 17572 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 17848 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 20148 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19504 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 19320 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 20884 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_211
timestamp 1604681595
transform 1 0 20516 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_209
timestamp 1604681595
transform 1 0 20332 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_19
timestamp 1604681595
transform 1 0 2852 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 3128 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4324 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5244 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 6072 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6624 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_59
timestamp 1604681595
transform 1 0 6532 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 8924 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8096 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1604681595
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9844 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11316 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _63_
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14352 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 13708 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_136
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 15640 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 17112 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 16008 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_171
timestamp 1604681595
transform 1 0 16836 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 17940 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19412 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 2944 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_19
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 4416 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5244 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7820 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_71
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9292 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1604681595
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15088 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 14720 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13892 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 15916 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_177
timestamp 1604681595
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 19504 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 20884 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_209
timestamp 1604681595
transform 1 0 20332 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 2116 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5520 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_64
timestamp 1604681595
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7176 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8740 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_82
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 12144 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_124
timestamp 1604681595
transform 1 0 12512 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1604681595
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 15732 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 17204 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 17572 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 18400 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 19872 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 1656 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 3312 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 4876 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 4048 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 3956 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_28
timestamp 1604681595
transform 1 0 3680 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 6900 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_50
timestamp 1604681595
transform 1 0 5704 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 7268 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 8464 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8832 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10304 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 9752 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9660 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12696 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12512 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_125
timestamp 1604681595
transform 1 0 12604 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 14996 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14168 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 17112 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 15640 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_156
timestamp 1604681595
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18308 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 18216 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_183
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 20884 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_209
timestamp 1604681595
transform 1 0 20332 0 1 19040
box -38 -48 314 592
<< labels >>
rlabel metal2 s 16394 0 16450 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 20994 21520 21050 22000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 20074 0 20130 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 21638 21520 21694 22000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 9034 0 9090 480 6 Test_en
port 4 nsew default input
rlabel metal2 s 1766 0 1822 480 6 bottom_width_0_height_0__pin_50_
port 5 nsew default tristate
rlabel metal2 s 5354 0 5410 480 6 bottom_width_0_height_0__pin_51_
port 6 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 ccff_head
port 7 nsew default input
rlabel metal3 s 21520 5584 22000 5704 6 ccff_tail
port 8 nsew default tristate
rlabel metal2 s 12714 0 12770 480 6 clk
port 9 nsew default input
rlabel metal3 s 0 18368 480 18488 6 left_width_0_height_0__pin_52_
port 10 nsew default input
rlabel metal3 s 0 3680 480 3800 6 prog_clk
port 11 nsew default input
rlabel metal3 s 21520 6264 22000 6384 6 right_width_0_height_0__pin_16_
port 12 nsew default input
rlabel metal3 s 21520 6944 22000 7064 6 right_width_0_height_0__pin_17_
port 13 nsew default input
rlabel metal3 s 21520 7624 22000 7744 6 right_width_0_height_0__pin_18_
port 14 nsew default input
rlabel metal3 s 21520 8168 22000 8288 6 right_width_0_height_0__pin_19_
port 15 nsew default input
rlabel metal3 s 21520 8848 22000 8968 6 right_width_0_height_0__pin_20_
port 16 nsew default input
rlabel metal3 s 21520 9528 22000 9648 6 right_width_0_height_0__pin_21_
port 17 nsew default input
rlabel metal3 s 21520 10208 22000 10328 6 right_width_0_height_0__pin_22_
port 18 nsew default input
rlabel metal3 s 21520 10888 22000 11008 6 right_width_0_height_0__pin_23_
port 19 nsew default input
rlabel metal3 s 21520 11568 22000 11688 6 right_width_0_height_0__pin_24_
port 20 nsew default input
rlabel metal3 s 21520 12248 22000 12368 6 right_width_0_height_0__pin_25_
port 21 nsew default input
rlabel metal3 s 21520 12928 22000 13048 6 right_width_0_height_0__pin_26_
port 22 nsew default input
rlabel metal3 s 21520 13608 22000 13728 6 right_width_0_height_0__pin_27_
port 23 nsew default input
rlabel metal3 s 21520 14288 22000 14408 6 right_width_0_height_0__pin_28_
port 24 nsew default input
rlabel metal3 s 21520 14968 22000 15088 6 right_width_0_height_0__pin_29_
port 25 nsew default input
rlabel metal3 s 21520 15512 22000 15632 6 right_width_0_height_0__pin_30_
port 26 nsew default input
rlabel metal3 s 21520 16192 22000 16312 6 right_width_0_height_0__pin_31_
port 27 nsew default input
rlabel metal3 s 21520 280 22000 400 6 right_width_0_height_0__pin_42_lower
port 28 nsew default tristate
rlabel metal3 s 21520 16872 22000 16992 6 right_width_0_height_0__pin_42_upper
port 29 nsew default tristate
rlabel metal3 s 21520 824 22000 944 6 right_width_0_height_0__pin_43_lower
port 30 nsew default tristate
rlabel metal3 s 21520 17552 22000 17672 6 right_width_0_height_0__pin_43_upper
port 31 nsew default tristate
rlabel metal3 s 21520 1504 22000 1624 6 right_width_0_height_0__pin_44_lower
port 32 nsew default tristate
rlabel metal3 s 21520 18232 22000 18352 6 right_width_0_height_0__pin_44_upper
port 33 nsew default tristate
rlabel metal3 s 21520 2184 22000 2304 6 right_width_0_height_0__pin_45_lower
port 34 nsew default tristate
rlabel metal3 s 21520 18912 22000 19032 6 right_width_0_height_0__pin_45_upper
port 35 nsew default tristate
rlabel metal3 s 21520 2864 22000 2984 6 right_width_0_height_0__pin_46_lower
port 36 nsew default tristate
rlabel metal3 s 21520 19592 22000 19712 6 right_width_0_height_0__pin_46_upper
port 37 nsew default tristate
rlabel metal3 s 21520 3544 22000 3664 6 right_width_0_height_0__pin_47_lower
port 38 nsew default tristate
rlabel metal3 s 21520 20272 22000 20392 6 right_width_0_height_0__pin_47_upper
port 39 nsew default tristate
rlabel metal3 s 21520 4224 22000 4344 6 right_width_0_height_0__pin_48_lower
port 40 nsew default tristate
rlabel metal3 s 21520 20952 22000 21072 6 right_width_0_height_0__pin_48_upper
port 41 nsew default tristate
rlabel metal3 s 21520 4904 22000 5024 6 right_width_0_height_0__pin_49_lower
port 42 nsew default tristate
rlabel metal3 s 21520 21632 22000 21752 6 right_width_0_height_0__pin_49_upper
port 43 nsew default tristate
rlabel metal2 s 5170 21520 5226 22000 6 top_width_0_height_0__pin_0_
port 44 nsew default input
rlabel metal2 s 11242 21520 11298 22000 6 top_width_0_height_0__pin_10_
port 45 nsew default input
rlabel metal2 s 11886 21520 11942 22000 6 top_width_0_height_0__pin_11_
port 46 nsew default input
rlabel metal2 s 12438 21520 12494 22000 6 top_width_0_height_0__pin_12_
port 47 nsew default input
rlabel metal2 s 13082 21520 13138 22000 6 top_width_0_height_0__pin_13_
port 48 nsew default input
rlabel metal2 s 13726 21520 13782 22000 6 top_width_0_height_0__pin_14_
port 49 nsew default input
rlabel metal2 s 14278 21520 14334 22000 6 top_width_0_height_0__pin_15_
port 50 nsew default input
rlabel metal2 s 5722 21520 5778 22000 6 top_width_0_height_0__pin_1_
port 51 nsew default input
rlabel metal2 s 6366 21520 6422 22000 6 top_width_0_height_0__pin_2_
port 52 nsew default input
rlabel metal2 s 14922 21520 14978 22000 6 top_width_0_height_0__pin_32_
port 53 nsew default input
rlabel metal2 s 15474 21520 15530 22000 6 top_width_0_height_0__pin_33_
port 54 nsew default input
rlabel metal2 s 16118 21520 16174 22000 6 top_width_0_height_0__pin_34_lower
port 55 nsew default tristate
rlabel metal2 s 294 21520 350 22000 6 top_width_0_height_0__pin_34_upper
port 56 nsew default tristate
rlabel metal2 s 16762 21520 16818 22000 6 top_width_0_height_0__pin_35_lower
port 57 nsew default tristate
rlabel metal2 s 846 21520 902 22000 6 top_width_0_height_0__pin_35_upper
port 58 nsew default tristate
rlabel metal2 s 17314 21520 17370 22000 6 top_width_0_height_0__pin_36_lower
port 59 nsew default tristate
rlabel metal2 s 1490 21520 1546 22000 6 top_width_0_height_0__pin_36_upper
port 60 nsew default tristate
rlabel metal2 s 17958 21520 18014 22000 6 top_width_0_height_0__pin_37_lower
port 61 nsew default tristate
rlabel metal2 s 2042 21520 2098 22000 6 top_width_0_height_0__pin_37_upper
port 62 nsew default tristate
rlabel metal2 s 18602 21520 18658 22000 6 top_width_0_height_0__pin_38_lower
port 63 nsew default tristate
rlabel metal2 s 2686 21520 2742 22000 6 top_width_0_height_0__pin_38_upper
port 64 nsew default tristate
rlabel metal2 s 19154 21520 19210 22000 6 top_width_0_height_0__pin_39_lower
port 65 nsew default tristate
rlabel metal2 s 3330 21520 3386 22000 6 top_width_0_height_0__pin_39_upper
port 66 nsew default tristate
rlabel metal2 s 7010 21520 7066 22000 6 top_width_0_height_0__pin_3_
port 67 nsew default input
rlabel metal2 s 19798 21520 19854 22000 6 top_width_0_height_0__pin_40_lower
port 68 nsew default tristate
rlabel metal2 s 3882 21520 3938 22000 6 top_width_0_height_0__pin_40_upper
port 69 nsew default tristate
rlabel metal2 s 20442 21520 20498 22000 6 top_width_0_height_0__pin_41_lower
port 70 nsew default tristate
rlabel metal2 s 4526 21520 4582 22000 6 top_width_0_height_0__pin_41_upper
port 71 nsew default tristate
rlabel metal2 s 7562 21520 7618 22000 6 top_width_0_height_0__pin_4_
port 72 nsew default input
rlabel metal2 s 8206 21520 8262 22000 6 top_width_0_height_0__pin_5_
port 73 nsew default input
rlabel metal2 s 8758 21520 8814 22000 6 top_width_0_height_0__pin_6_
port 74 nsew default input
rlabel metal2 s 9402 21520 9458 22000 6 top_width_0_height_0__pin_7_
port 75 nsew default input
rlabel metal2 s 10046 21520 10102 22000 6 top_width_0_height_0__pin_8_
port 76 nsew default input
rlabel metal2 s 10598 21520 10654 22000 6 top_width_0_height_0__pin_9_
port 77 nsew default input
rlabel metal4 s 4243 2128 4563 19632 6 VPWR
port 78 nsew default input
rlabel metal4 s 7541 2128 7861 19632 6 VGND
port 79 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22000 22000
<< end >>
