VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decoder6to61
  CLASS BLOCK ;
  FOREIGN decoder6to61 ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.270 BY 120.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 117.600 10.030 120.000 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 117.600 29.810 120.000 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 117.600 50.050 120.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 117.600 69.830 120.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 117.600 90.070 120.000 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.570 117.600 109.850 120.000 ;
    END
  END address[5]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 2.400 1.320 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 2.400 20.360 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 2.400 24.440 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.400 26.480 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 2.400 30.560 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 2.400 32.600 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 2.400 34.640 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 2.400 36.000 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 2.400 38.040 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 2.400 40.080 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 2.400 42.120 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 2.400 46.200 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 2.400 48.240 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 2.400 50.280 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.400 52.320 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.400 53.680 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 2.400 57.760 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.400 61.840 ;
    END
  END data_out[31]
  PIN data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.400 63.880 ;
    END
  END data_out[32]
  PIN data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END data_out[33]
  PIN data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 2.400 67.960 ;
    END
  END data_out[34]
  PIN data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 2.400 69.320 ;
    END
  END data_out[35]
  PIN data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.400 71.360 ;
    END
  END data_out[36]
  PIN data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END data_out[37]
  PIN data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 2.400 75.440 ;
    END
  END data_out[38]
  PIN data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END data_out[39]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 2.400 6.760 ;
    END
  END data_out[3]
  PIN data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END data_out[40]
  PIN data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 2.400 81.560 ;
    END
  END data_out[41]
  PIN data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.400 83.600 ;
    END
  END data_out[42]
  PIN data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END data_out[43]
  PIN data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END data_out[44]
  PIN data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 2.400 89.040 ;
    END
  END data_out[45]
  PIN data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 2.400 91.080 ;
    END
  END data_out[46]
  PIN data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.400 93.120 ;
    END
  END data_out[47]
  PIN data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 2.400 95.160 ;
    END
  END data_out[48]
  PIN data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 2.400 97.200 ;
    END
  END data_out[49]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END data_out[4]
  PIN data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 2.400 99.240 ;
    END
  END data_out[50]
  PIN data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.400 101.280 ;
    END
  END data_out[51]
  PIN data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 2.400 103.320 ;
    END
  END data_out[52]
  PIN data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 2.400 104.680 ;
    END
  END data_out[53]
  PIN data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.400 106.720 ;
    END
  END data_out[54]
  PIN data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.400 108.760 ;
    END
  END data_out[55]
  PIN data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.400 110.800 ;
    END
  END data_out[56]
  PIN data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.400 112.840 ;
    END
  END data_out[57]
  PIN data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 2.400 114.880 ;
    END
  END data_out[58]
  PIN data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 2.400 116.920 ;
    END
  END data_out[59]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END data_out[5]
  PIN data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 2.400 118.960 ;
    END
  END data_out[60]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 2.400 14.920 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 2.400 16.960 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 2.400 18.320 ;
    END
  END data_out[9]
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END enable
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 24.720 10.640 26.320 109.040 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 44.720 10.640 46.320 109.040 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 0.145 10.795 114.080 108.885 ;
      LAYER met1 ;
        RECT 0.070 6.500 114.080 117.940 ;
      LAYER met2 ;
        RECT 0.090 117.320 9.470 118.845 ;
        RECT 10.310 117.320 29.250 118.845 ;
        RECT 30.090 117.320 49.490 118.845 ;
        RECT 50.330 117.320 69.270 118.845 ;
        RECT 70.110 117.320 89.510 118.845 ;
        RECT 90.350 117.320 109.290 118.845 ;
        RECT 110.130 117.320 110.310 118.845 ;
        RECT 0.090 2.680 110.310 117.320 ;
        RECT 0.090 0.270 59.610 2.680 ;
        RECT 60.450 0.270 110.310 2.680 ;
      LAYER met3 ;
        RECT 2.800 107.760 110.335 108.965 ;
        RECT 0.270 107.120 110.335 107.760 ;
        RECT 2.800 105.720 110.335 107.120 ;
        RECT 0.270 105.080 110.335 105.720 ;
        RECT 2.800 102.320 110.335 105.080 ;
        RECT 0.270 101.680 110.335 102.320 ;
        RECT 2.800 100.280 110.335 101.680 ;
        RECT 0.270 99.640 110.335 100.280 ;
        RECT 2.800 98.240 110.335 99.640 ;
        RECT 0.270 97.600 110.335 98.240 ;
        RECT 2.800 96.200 110.335 97.600 ;
        RECT 0.270 95.560 110.335 96.200 ;
        RECT 2.800 94.160 110.335 95.560 ;
        RECT 0.270 93.520 110.335 94.160 ;
        RECT 2.800 92.120 110.335 93.520 ;
        RECT 0.270 91.480 110.335 92.120 ;
        RECT 2.800 90.080 110.335 91.480 ;
        RECT 0.270 89.440 110.335 90.080 ;
        RECT 2.800 88.040 110.335 89.440 ;
        RECT 0.270 87.400 110.335 88.040 ;
        RECT 2.800 84.640 110.335 87.400 ;
        RECT 0.270 84.000 110.335 84.640 ;
        RECT 2.800 82.600 110.335 84.000 ;
        RECT 0.270 81.960 110.335 82.600 ;
        RECT 2.800 80.560 110.335 81.960 ;
        RECT 0.270 79.920 110.335 80.560 ;
        RECT 2.800 78.520 110.335 79.920 ;
        RECT 0.270 77.880 110.335 78.520 ;
        RECT 2.800 76.480 110.335 77.880 ;
        RECT 0.270 75.840 110.335 76.480 ;
        RECT 2.800 74.440 110.335 75.840 ;
        RECT 0.270 73.800 110.335 74.440 ;
        RECT 2.800 72.400 110.335 73.800 ;
        RECT 0.270 71.760 110.335 72.400 ;
        RECT 2.800 70.360 110.335 71.760 ;
        RECT 0.270 69.720 110.335 70.360 ;
        RECT 2.800 66.960 110.335 69.720 ;
        RECT 0.270 66.320 110.335 66.960 ;
        RECT 2.800 64.920 110.335 66.320 ;
        RECT 0.270 64.280 110.335 64.920 ;
        RECT 2.800 62.880 110.335 64.280 ;
        RECT 0.270 62.240 110.335 62.880 ;
        RECT 2.800 60.840 110.335 62.240 ;
        RECT 0.270 60.200 110.335 60.840 ;
        RECT 2.800 58.800 110.335 60.200 ;
        RECT 0.270 58.160 110.335 58.800 ;
        RECT 2.800 56.760 110.335 58.160 ;
        RECT 0.270 56.120 110.335 56.760 ;
        RECT 2.800 54.720 110.335 56.120 ;
        RECT 0.270 54.080 110.335 54.720 ;
        RECT 2.800 51.320 110.335 54.080 ;
        RECT 0.270 50.680 110.335 51.320 ;
        RECT 2.800 49.280 110.335 50.680 ;
        RECT 0.270 48.640 110.335 49.280 ;
        RECT 2.800 47.240 110.335 48.640 ;
        RECT 0.270 46.600 110.335 47.240 ;
        RECT 2.800 45.200 110.335 46.600 ;
        RECT 0.270 44.560 110.335 45.200 ;
        RECT 2.800 43.160 110.335 44.560 ;
        RECT 0.270 42.520 110.335 43.160 ;
        RECT 2.800 41.120 110.335 42.520 ;
        RECT 0.270 40.480 110.335 41.120 ;
        RECT 2.800 39.080 110.335 40.480 ;
        RECT 0.270 38.440 110.335 39.080 ;
        RECT 2.800 37.040 110.335 38.440 ;
        RECT 0.270 36.400 110.335 37.040 ;
        RECT 2.800 33.640 110.335 36.400 ;
        RECT 0.270 33.000 110.335 33.640 ;
        RECT 2.800 31.600 110.335 33.000 ;
        RECT 0.270 30.960 110.335 31.600 ;
        RECT 2.800 29.560 110.335 30.960 ;
        RECT 0.270 28.920 110.335 29.560 ;
        RECT 2.800 27.520 110.335 28.920 ;
        RECT 0.270 26.880 110.335 27.520 ;
        RECT 2.800 25.480 110.335 26.880 ;
        RECT 0.270 24.840 110.335 25.480 ;
        RECT 2.800 23.440 110.335 24.840 ;
        RECT 0.270 22.800 110.335 23.440 ;
        RECT 2.800 21.400 110.335 22.800 ;
        RECT 0.270 20.760 110.335 21.400 ;
        RECT 2.800 19.360 110.335 20.760 ;
        RECT 0.270 18.720 110.335 19.360 ;
        RECT 2.800 15.960 110.335 18.720 ;
        RECT 0.270 15.320 110.335 15.960 ;
        RECT 2.800 13.920 110.335 15.320 ;
        RECT 0.270 13.280 110.335 13.920 ;
        RECT 2.800 11.880 110.335 13.280 ;
        RECT 0.270 11.240 110.335 11.880 ;
        RECT 2.800 9.840 110.335 11.240 ;
        RECT 0.270 9.200 110.335 9.840 ;
        RECT 2.800 7.800 110.335 9.200 ;
        RECT 0.270 7.160 110.335 7.800 ;
        RECT 2.800 5.760 110.335 7.160 ;
        RECT 0.270 5.120 110.335 5.760 ;
        RECT 2.800 3.720 110.335 5.120 ;
        RECT 0.270 3.080 110.335 3.720 ;
        RECT 2.800 2.680 110.335 3.080 ;
      LAYER met4 ;
        RECT 0.295 109.440 106.320 110.665 ;
        RECT 0.295 10.640 24.320 109.440 ;
        RECT 26.720 10.640 44.320 109.440 ;
        RECT 46.720 10.640 106.320 109.440 ;
  END
END decoder6to61
END LIBRARY

