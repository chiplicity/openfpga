magic
tech sky130A
magscale 1 2
timestamp 1608135360
<< obsli1 >>
rect 1104 2159 15824 17425
<< obsm1 >>
rect 198 1300 16822 19168
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 938 19200 994 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2226 19200 2282 20000
rect 2594 19200 2650 20000
rect 2962 19200 3018 20000
rect 3422 19200 3478 20000
rect 3790 19200 3846 20000
rect 4250 19200 4306 20000
rect 4618 19200 4674 20000
rect 4986 19200 5042 20000
rect 5446 19200 5502 20000
rect 5814 19200 5870 20000
rect 6274 19200 6330 20000
rect 6642 19200 6698 20000
rect 7010 19200 7066 20000
rect 7470 19200 7526 20000
rect 7838 19200 7894 20000
rect 8298 19200 8354 20000
rect 8666 19200 8722 20000
rect 9034 19200 9090 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 10322 19200 10378 20000
rect 10690 19200 10746 20000
rect 11058 19200 11114 20000
rect 11518 19200 11574 20000
rect 11886 19200 11942 20000
rect 12346 19200 12402 20000
rect 12714 19200 12770 20000
rect 13082 19200 13138 20000
rect 13542 19200 13598 20000
rect 13910 19200 13966 20000
rect 14370 19200 14426 20000
rect 14738 19200 14794 20000
rect 15106 19200 15162 20000
rect 15566 19200 15622 20000
rect 15934 19200 15990 20000
rect 16394 19200 16450 20000
rect 16762 19200 16818 20000
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16762 0 16818 800
<< obsm2 >>
rect 314 19144 514 19553
rect 682 19144 882 19553
rect 1050 19144 1342 19553
rect 1510 19144 1710 19553
rect 1878 19144 2170 19553
rect 2338 19144 2538 19553
rect 2706 19144 2906 19553
rect 3074 19144 3366 19553
rect 3534 19144 3734 19553
rect 3902 19144 4194 19553
rect 4362 19144 4562 19553
rect 4730 19144 4930 19553
rect 5098 19144 5390 19553
rect 5558 19144 5758 19553
rect 5926 19144 6218 19553
rect 6386 19144 6586 19553
rect 6754 19144 6954 19553
rect 7122 19144 7414 19553
rect 7582 19144 7782 19553
rect 7950 19144 8242 19553
rect 8410 19144 8610 19553
rect 8778 19144 8978 19553
rect 9146 19144 9438 19553
rect 9606 19144 9806 19553
rect 9974 19144 10266 19553
rect 10434 19144 10634 19553
rect 10802 19144 11002 19553
rect 11170 19144 11462 19553
rect 11630 19144 11830 19553
rect 11998 19144 12290 19553
rect 12458 19144 12658 19553
rect 12826 19144 13026 19553
rect 13194 19144 13486 19553
rect 13654 19144 13854 19553
rect 14022 19144 14314 19553
rect 14482 19144 14682 19553
rect 14850 19144 15050 19553
rect 15218 19144 15510 19553
rect 15678 19144 15878 19553
rect 16046 19144 16338 19553
rect 16506 19144 16706 19553
rect 202 856 16816 19144
rect 314 800 514 856
rect 682 800 974 856
rect 1142 800 1342 856
rect 1510 800 1802 856
rect 1970 800 2170 856
rect 2338 800 2630 856
rect 2798 800 2998 856
rect 3166 800 3458 856
rect 3626 800 3826 856
rect 3994 800 4286 856
rect 4454 800 4654 856
rect 4822 800 5114 856
rect 5282 800 5482 856
rect 5650 800 5942 856
rect 6110 800 6310 856
rect 6478 800 6770 856
rect 6938 800 7138 856
rect 7306 800 7598 856
rect 7766 800 7966 856
rect 8134 800 8426 856
rect 8594 800 8794 856
rect 8962 800 9254 856
rect 9422 800 9622 856
rect 9790 800 10082 856
rect 10250 800 10450 856
rect 10618 800 10910 856
rect 11078 800 11278 856
rect 11446 800 11738 856
rect 11906 800 12106 856
rect 12274 800 12566 856
rect 12734 800 12934 856
rect 13102 800 13394 856
rect 13562 800 13762 856
rect 13930 800 14222 856
rect 14390 800 14590 856
rect 14758 800 15050 856
rect 15218 800 15418 856
rect 15586 800 15878 856
rect 16046 800 16246 856
rect 16414 800 16706 856
<< metal3 >>
rect 0 19456 800 19576
rect 0 18504 800 18624
rect 16200 17824 17000 17944
rect 0 17552 800 17672
rect 0 16600 800 16720
rect 0 15648 800 15768
rect 0 14696 800 14816
rect 0 13744 800 13864
rect 16200 13880 17000 14000
rect 0 12792 800 12912
rect 0 11840 800 11960
rect 0 10888 800 11008
rect 0 9936 800 10056
rect 16200 9800 17000 9920
rect 0 8984 800 9104
rect 0 8032 800 8152
rect 0 7080 800 7200
rect 0 6128 800 6248
rect 16200 5856 17000 5976
rect 0 5176 800 5296
rect 0 4224 800 4344
rect 0 3272 800 3392
rect 0 2320 800 2440
rect 16200 1912 17000 2032
rect 0 1368 800 1488
rect 0 416 800 536
<< obsm3 >>
rect 880 19376 16200 19549
rect 197 18704 16200 19376
rect 880 18424 16200 18704
rect 197 18024 16200 18424
rect 197 17752 16120 18024
rect 880 17744 16120 17752
rect 880 17472 16200 17744
rect 197 16800 16200 17472
rect 880 16520 16200 16800
rect 197 15848 16200 16520
rect 880 15568 16200 15848
rect 197 14896 16200 15568
rect 880 14616 16200 14896
rect 197 14080 16200 14616
rect 197 13944 16120 14080
rect 880 13800 16120 13944
rect 880 13664 16200 13800
rect 197 12992 16200 13664
rect 880 12712 16200 12992
rect 197 12040 16200 12712
rect 880 11760 16200 12040
rect 197 11088 16200 11760
rect 880 10808 16200 11088
rect 197 10136 16200 10808
rect 880 10000 16200 10136
rect 880 9856 16120 10000
rect 197 9720 16120 9856
rect 197 9184 16200 9720
rect 880 8904 16200 9184
rect 197 8232 16200 8904
rect 880 7952 16200 8232
rect 197 7280 16200 7952
rect 880 7000 16200 7280
rect 197 6328 16200 7000
rect 880 6056 16200 6328
rect 880 6048 16120 6056
rect 197 5776 16120 6048
rect 197 5376 16200 5776
rect 880 5096 16200 5376
rect 197 4424 16200 5096
rect 880 4144 16200 4424
rect 197 3472 16200 4144
rect 880 3192 16200 3472
rect 197 2520 16200 3192
rect 880 2240 16200 2520
rect 197 2112 16200 2240
rect 197 1832 16120 2112
rect 197 1568 16200 1832
rect 880 1288 16200 1568
rect 197 616 16200 1288
rect 880 444 16200 616
<< metal4 >>
rect 3409 2128 3729 17456
rect 5875 2128 6195 17456
<< obsm4 >>
rect 2819 2048 3329 17456
rect 3809 2048 5795 17456
rect 6275 2048 14661 17456
rect 2819 443 14661 2048
<< labels >>
rlabel metal2 s 202 19200 258 20000 6 IO_ISOL_N
port 1 nsew default input
rlabel metal3 s 0 1368 800 1488 6 ccff_head
port 2 nsew default input
rlabel metal3 s 16200 1912 17000 2032 6 ccff_tail
port 3 nsew default output
rlabel metal2 s 8482 0 8538 800 6 chany_bottom_in[0]
port 4 nsew default input
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_in[10]
port 5 nsew default input
rlabel metal2 s 12990 0 13046 800 6 chany_bottom_in[11]
port 6 nsew default input
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_in[12]
port 7 nsew default input
rlabel metal2 s 13818 0 13874 800 6 chany_bottom_in[13]
port 8 nsew default input
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_in[14]
port 9 nsew default input
rlabel metal2 s 14646 0 14702 800 6 chany_bottom_in[15]
port 10 nsew default input
rlabel metal2 s 15106 0 15162 800 6 chany_bottom_in[16]
port 11 nsew default input
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_in[17]
port 12 nsew default input
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_in[18]
port 13 nsew default input
rlabel metal2 s 16302 0 16358 800 6 chany_bottom_in[19]
port 14 nsew default input
rlabel metal2 s 8850 0 8906 800 6 chany_bottom_in[1]
port 15 nsew default input
rlabel metal2 s 9310 0 9366 800 6 chany_bottom_in[2]
port 16 nsew default input
rlabel metal2 s 9678 0 9734 800 6 chany_bottom_in[3]
port 17 nsew default input
rlabel metal2 s 10138 0 10194 800 6 chany_bottom_in[4]
port 18 nsew default input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[5]
port 19 nsew default input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[6]
port 20 nsew default input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_in[7]
port 21 nsew default input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[8]
port 22 nsew default input
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_in[9]
port 23 nsew default input
rlabel metal2 s 202 0 258 800 6 chany_bottom_out[0]
port 24 nsew default output
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_out[10]
port 25 nsew default output
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_out[11]
port 26 nsew default output
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_out[12]
port 27 nsew default output
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_out[13]
port 28 nsew default output
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_out[14]
port 29 nsew default output
rlabel metal2 s 6366 0 6422 800 6 chany_bottom_out[15]
port 30 nsew default output
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_out[16]
port 31 nsew default output
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_out[17]
port 32 nsew default output
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_out[18]
port 33 nsew default output
rlabel metal2 s 8022 0 8078 800 6 chany_bottom_out[19]
port 34 nsew default output
rlabel metal2 s 570 0 626 800 6 chany_bottom_out[1]
port 35 nsew default output
rlabel metal2 s 1030 0 1086 800 6 chany_bottom_out[2]
port 36 nsew default output
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_out[3]
port 37 nsew default output
rlabel metal2 s 1858 0 1914 800 6 chany_bottom_out[4]
port 38 nsew default output
rlabel metal2 s 2226 0 2282 800 6 chany_bottom_out[5]
port 39 nsew default output
rlabel metal2 s 2686 0 2742 800 6 chany_bottom_out[6]
port 40 nsew default output
rlabel metal2 s 3054 0 3110 800 6 chany_bottom_out[7]
port 41 nsew default output
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_out[8]
port 42 nsew default output
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_out[9]
port 43 nsew default output
rlabel metal2 s 8666 19200 8722 20000 6 chany_top_in[0]
port 44 nsew default input
rlabel metal2 s 12714 19200 12770 20000 6 chany_top_in[10]
port 45 nsew default input
rlabel metal2 s 13082 19200 13138 20000 6 chany_top_in[11]
port 46 nsew default input
rlabel metal2 s 13542 19200 13598 20000 6 chany_top_in[12]
port 47 nsew default input
rlabel metal2 s 13910 19200 13966 20000 6 chany_top_in[13]
port 48 nsew default input
rlabel metal2 s 14370 19200 14426 20000 6 chany_top_in[14]
port 49 nsew default input
rlabel metal2 s 14738 19200 14794 20000 6 chany_top_in[15]
port 50 nsew default input
rlabel metal2 s 15106 19200 15162 20000 6 chany_top_in[16]
port 51 nsew default input
rlabel metal2 s 15566 19200 15622 20000 6 chany_top_in[17]
port 52 nsew default input
rlabel metal2 s 15934 19200 15990 20000 6 chany_top_in[18]
port 53 nsew default input
rlabel metal2 s 16394 19200 16450 20000 6 chany_top_in[19]
port 54 nsew default input
rlabel metal2 s 9034 19200 9090 20000 6 chany_top_in[1]
port 55 nsew default input
rlabel metal2 s 9494 19200 9550 20000 6 chany_top_in[2]
port 56 nsew default input
rlabel metal2 s 9862 19200 9918 20000 6 chany_top_in[3]
port 57 nsew default input
rlabel metal2 s 10322 19200 10378 20000 6 chany_top_in[4]
port 58 nsew default input
rlabel metal2 s 10690 19200 10746 20000 6 chany_top_in[5]
port 59 nsew default input
rlabel metal2 s 11058 19200 11114 20000 6 chany_top_in[6]
port 60 nsew default input
rlabel metal2 s 11518 19200 11574 20000 6 chany_top_in[7]
port 61 nsew default input
rlabel metal2 s 11886 19200 11942 20000 6 chany_top_in[8]
port 62 nsew default input
rlabel metal2 s 12346 19200 12402 20000 6 chany_top_in[9]
port 63 nsew default input
rlabel metal2 s 570 19200 626 20000 6 chany_top_out[0]
port 64 nsew default output
rlabel metal2 s 4618 19200 4674 20000 6 chany_top_out[10]
port 65 nsew default output
rlabel metal2 s 4986 19200 5042 20000 6 chany_top_out[11]
port 66 nsew default output
rlabel metal2 s 5446 19200 5502 20000 6 chany_top_out[12]
port 67 nsew default output
rlabel metal2 s 5814 19200 5870 20000 6 chany_top_out[13]
port 68 nsew default output
rlabel metal2 s 6274 19200 6330 20000 6 chany_top_out[14]
port 69 nsew default output
rlabel metal2 s 6642 19200 6698 20000 6 chany_top_out[15]
port 70 nsew default output
rlabel metal2 s 7010 19200 7066 20000 6 chany_top_out[16]
port 71 nsew default output
rlabel metal2 s 7470 19200 7526 20000 6 chany_top_out[17]
port 72 nsew default output
rlabel metal2 s 7838 19200 7894 20000 6 chany_top_out[18]
port 73 nsew default output
rlabel metal2 s 8298 19200 8354 20000 6 chany_top_out[19]
port 74 nsew default output
rlabel metal2 s 938 19200 994 20000 6 chany_top_out[1]
port 75 nsew default output
rlabel metal2 s 1398 19200 1454 20000 6 chany_top_out[2]
port 76 nsew default output
rlabel metal2 s 1766 19200 1822 20000 6 chany_top_out[3]
port 77 nsew default output
rlabel metal2 s 2226 19200 2282 20000 6 chany_top_out[4]
port 78 nsew default output
rlabel metal2 s 2594 19200 2650 20000 6 chany_top_out[5]
port 79 nsew default output
rlabel metal2 s 2962 19200 3018 20000 6 chany_top_out[6]
port 80 nsew default output
rlabel metal2 s 3422 19200 3478 20000 6 chany_top_out[7]
port 81 nsew default output
rlabel metal2 s 3790 19200 3846 20000 6 chany_top_out[8]
port 82 nsew default output
rlabel metal2 s 4250 19200 4306 20000 6 chany_top_out[9]
port 83 nsew default output
rlabel metal3 s 16200 9800 17000 9920 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 84 nsew default output
rlabel metal3 s 16200 13880 17000 14000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 85 nsew default input
rlabel metal3 s 16200 17824 17000 17944 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 86 nsew default output
rlabel metal3 s 0 3272 800 3392 6 left_grid_pin_16_
port 87 nsew default output
rlabel metal3 s 0 4224 800 4344 6 left_grid_pin_17_
port 88 nsew default output
rlabel metal3 s 0 5176 800 5296 6 left_grid_pin_18_
port 89 nsew default output
rlabel metal3 s 0 6128 800 6248 6 left_grid_pin_19_
port 90 nsew default output
rlabel metal3 s 0 7080 800 7200 6 left_grid_pin_20_
port 91 nsew default output
rlabel metal3 s 0 8032 800 8152 6 left_grid_pin_21_
port 92 nsew default output
rlabel metal3 s 0 8984 800 9104 6 left_grid_pin_22_
port 93 nsew default output
rlabel metal3 s 0 9936 800 10056 6 left_grid_pin_23_
port 94 nsew default output
rlabel metal3 s 0 10888 800 11008 6 left_grid_pin_24_
port 95 nsew default output
rlabel metal3 s 0 11840 800 11960 6 left_grid_pin_25_
port 96 nsew default output
rlabel metal3 s 0 12792 800 12912 6 left_grid_pin_26_
port 97 nsew default output
rlabel metal3 s 0 13744 800 13864 6 left_grid_pin_27_
port 98 nsew default output
rlabel metal3 s 0 14696 800 14816 6 left_grid_pin_28_
port 99 nsew default output
rlabel metal3 s 0 15648 800 15768 6 left_grid_pin_29_
port 100 nsew default output
rlabel metal3 s 0 16600 800 16720 6 left_grid_pin_30_
port 101 nsew default output
rlabel metal3 s 0 17552 800 17672 6 left_grid_pin_31_
port 102 nsew default output
rlabel metal3 s 0 18504 800 18624 6 left_width_0_height_0__pin_0_
port 103 nsew default input
rlabel metal3 s 0 416 800 536 6 left_width_0_height_0__pin_1_lower
port 104 nsew default output
rlabel metal3 s 0 19456 800 19576 6 left_width_0_height_0__pin_1_upper
port 105 nsew default output
rlabel metal2 s 16762 19200 16818 20000 6 prog_clk_0_N_out
port 106 nsew default output
rlabel metal2 s 16762 0 16818 800 6 prog_clk_0_S_out
port 107 nsew default output
rlabel metal3 s 0 2320 800 2440 6 prog_clk_0_W_in
port 108 nsew default input
rlabel metal3 s 16200 5856 17000 5976 6 right_grid_pin_0_
port 109 nsew default output
rlabel metal4 s 3409 2128 3729 17456 6 VPWR
port 110 nsew power input
rlabel metal4 s 5875 2128 6195 17456 6 VGND
port 111 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 17000 20000
string LEFview TRUE
<< end >>
