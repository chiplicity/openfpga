VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_2__0_
  CLASS BLOCK ;
  FOREIGN sb_2__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.000 BY 114.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 57.160 114.000 57.760 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 2.400 45.520 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 2.400 47.560 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 2.400 50.280 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.400 52.320 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.400 61.840 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.400 63.880 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.400 66.600 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 2.400 24.440 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.400 26.480 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.400 29.200 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 2.400 31.240 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 2.400 36.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 2.400 38.040 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 2.400 40.760 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 2.400 42.800 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 2.400 91.760 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 2.400 94.480 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 2.400 96.520 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 2.400 99.240 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.400 101.280 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 2.400 103.320 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.400 106.040 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 2.400 108.080 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.400 110.800 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.400 112.840 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 2.400 75.440 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 2.400 78.160 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 2.400 82.920 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 2.400 84.960 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 2.400 89.720 ;
    END
  END chanx_left_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 111.600 19.230 114.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 111.600 42.230 114.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 111.600 44.530 114.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 111.600 46.830 114.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 111.600 49.130 114.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 111.600 51.430 114.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 111.600 53.730 114.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 111.600 56.030 114.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 111.600 58.330 114.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 111.600 60.170 114.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 111.600 62.470 114.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 111.600 21.530 114.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 111.600 23.830 114.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 111.600 26.130 114.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 111.600 28.430 114.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 111.600 30.730 114.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 111.600 33.030 114.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 111.600 35.330 114.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 111.600 37.630 114.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 111.600 39.930 114.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 111.600 64.770 114.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 111.600 87.770 114.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 111.600 90.070 114.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 111.600 92.370 114.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.390 111.600 94.670 114.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 111.600 96.970 114.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 111.600 99.270 114.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 111.600 101.570 114.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 111.600 103.870 114.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 111.600 106.170 114.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 111.600 108.470 114.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.790 111.600 67.070 114.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 111.600 69.370 114.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 111.600 71.670 114.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 111.600 73.970 114.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.990 111.600 76.270 114.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 111.600 78.570 114.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.590 111.600 80.870 114.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 111.600 83.170 114.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 111.600 85.470 114.000 ;
    END
  END chany_top_out[9]
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 2.400 14.920 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 2.400 19.680 ;
    END
  END left_bottom_grid_pin_17_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 2.400 1.320 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 2.400 5.400 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 2.400 8.120 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 2.400 10.160 ;
    END
  END left_bottom_grid_pin_9_
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 111.600 110.770 114.000 ;
    END
  END prog_clk_0_N_in
  PIN top_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 111.600 1.290 114.000 ;
    END
  END top_left_grid_pin_42_
  PIN top_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 111.600 3.130 114.000 ;
    END
  END top_left_grid_pin_43_
  PIN top_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 111.600 5.430 114.000 ;
    END
  END top_left_grid_pin_44_
  PIN top_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 111.600 7.730 114.000 ;
    END
  END top_left_grid_pin_45_
  PIN top_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 111.600 10.030 114.000 ;
    END
  END top_left_grid_pin_46_
  PIN top_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 111.600 12.330 114.000 ;
    END
  END top_left_grid_pin_47_
  PIN top_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 111.600 14.630 114.000 ;
    END
  END top_left_grid_pin_48_
  PIN top_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 111.600 16.930 114.000 ;
    END
  END top_left_grid_pin_49_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.790 111.600 113.070 114.000 ;
    END
  END top_right_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.880 10.640 23.480 100.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.040 10.640 40.640 100.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.100 100.725 ;
      LAYER met1 ;
        RECT 0.990 2.080 113.090 100.880 ;
      LAYER met2 ;
        RECT 1.570 111.320 2.570 112.725 ;
        RECT 3.410 111.320 4.870 112.725 ;
        RECT 5.710 111.320 7.170 112.725 ;
        RECT 8.010 111.320 9.470 112.725 ;
        RECT 10.310 111.320 11.770 112.725 ;
        RECT 12.610 111.320 14.070 112.725 ;
        RECT 14.910 111.320 16.370 112.725 ;
        RECT 17.210 111.320 18.670 112.725 ;
        RECT 19.510 111.320 20.970 112.725 ;
        RECT 21.810 111.320 23.270 112.725 ;
        RECT 24.110 111.320 25.570 112.725 ;
        RECT 26.410 111.320 27.870 112.725 ;
        RECT 28.710 111.320 30.170 112.725 ;
        RECT 31.010 111.320 32.470 112.725 ;
        RECT 33.310 111.320 34.770 112.725 ;
        RECT 35.610 111.320 37.070 112.725 ;
        RECT 37.910 111.320 39.370 112.725 ;
        RECT 40.210 111.320 41.670 112.725 ;
        RECT 42.510 111.320 43.970 112.725 ;
        RECT 44.810 111.320 46.270 112.725 ;
        RECT 47.110 111.320 48.570 112.725 ;
        RECT 49.410 111.320 50.870 112.725 ;
        RECT 51.710 111.320 53.170 112.725 ;
        RECT 54.010 111.320 55.470 112.725 ;
        RECT 56.310 111.320 57.770 112.725 ;
        RECT 58.610 111.320 59.610 112.725 ;
        RECT 60.450 111.320 61.910 112.725 ;
        RECT 62.750 111.320 64.210 112.725 ;
        RECT 65.050 111.320 66.510 112.725 ;
        RECT 67.350 111.320 68.810 112.725 ;
        RECT 69.650 111.320 71.110 112.725 ;
        RECT 71.950 111.320 73.410 112.725 ;
        RECT 74.250 111.320 75.710 112.725 ;
        RECT 76.550 111.320 78.010 112.725 ;
        RECT 78.850 111.320 80.310 112.725 ;
        RECT 81.150 111.320 82.610 112.725 ;
        RECT 83.450 111.320 84.910 112.725 ;
        RECT 85.750 111.320 87.210 112.725 ;
        RECT 88.050 111.320 89.510 112.725 ;
        RECT 90.350 111.320 91.810 112.725 ;
        RECT 92.650 111.320 94.110 112.725 ;
        RECT 94.950 111.320 96.410 112.725 ;
        RECT 97.250 111.320 98.710 112.725 ;
        RECT 99.550 111.320 101.010 112.725 ;
        RECT 101.850 111.320 103.310 112.725 ;
        RECT 104.150 111.320 105.610 112.725 ;
        RECT 106.450 111.320 107.910 112.725 ;
        RECT 108.750 111.320 110.210 112.725 ;
        RECT 111.050 111.320 112.510 112.725 ;
        RECT 1.020 2.680 113.060 111.320 ;
        RECT 1.020 0.835 56.850 2.680 ;
        RECT 57.690 0.835 113.060 2.680 ;
      LAYER met3 ;
        RECT 2.800 111.840 111.600 112.705 ;
        RECT 2.400 111.200 111.600 111.840 ;
        RECT 2.800 109.800 111.600 111.200 ;
        RECT 2.400 108.480 111.600 109.800 ;
        RECT 2.800 107.080 111.600 108.480 ;
        RECT 2.400 106.440 111.600 107.080 ;
        RECT 2.800 105.040 111.600 106.440 ;
        RECT 2.400 103.720 111.600 105.040 ;
        RECT 2.800 102.320 111.600 103.720 ;
        RECT 2.400 101.680 111.600 102.320 ;
        RECT 2.800 100.280 111.600 101.680 ;
        RECT 2.400 99.640 111.600 100.280 ;
        RECT 2.800 98.240 111.600 99.640 ;
        RECT 2.400 96.920 111.600 98.240 ;
        RECT 2.800 95.520 111.600 96.920 ;
        RECT 2.400 94.880 111.600 95.520 ;
        RECT 2.800 93.480 111.600 94.880 ;
        RECT 2.400 92.160 111.600 93.480 ;
        RECT 2.800 90.760 111.600 92.160 ;
        RECT 2.400 90.120 111.600 90.760 ;
        RECT 2.800 88.720 111.600 90.120 ;
        RECT 2.400 87.400 111.600 88.720 ;
        RECT 2.800 86.000 111.600 87.400 ;
        RECT 2.400 85.360 111.600 86.000 ;
        RECT 2.800 83.960 111.600 85.360 ;
        RECT 2.400 83.320 111.600 83.960 ;
        RECT 2.800 81.920 111.600 83.320 ;
        RECT 2.400 80.600 111.600 81.920 ;
        RECT 2.800 79.200 111.600 80.600 ;
        RECT 2.400 78.560 111.600 79.200 ;
        RECT 2.800 77.160 111.600 78.560 ;
        RECT 2.400 75.840 111.600 77.160 ;
        RECT 2.800 74.440 111.600 75.840 ;
        RECT 2.400 73.800 111.600 74.440 ;
        RECT 2.800 72.400 111.600 73.800 ;
        RECT 2.400 71.080 111.600 72.400 ;
        RECT 2.800 69.680 111.600 71.080 ;
        RECT 2.400 69.040 111.600 69.680 ;
        RECT 2.800 67.640 111.600 69.040 ;
        RECT 2.400 67.000 111.600 67.640 ;
        RECT 2.800 65.600 111.600 67.000 ;
        RECT 2.400 64.280 111.600 65.600 ;
        RECT 2.800 62.880 111.600 64.280 ;
        RECT 2.400 62.240 111.600 62.880 ;
        RECT 2.800 60.840 111.600 62.240 ;
        RECT 2.400 59.520 111.600 60.840 ;
        RECT 2.800 58.160 111.600 59.520 ;
        RECT 2.800 58.120 111.200 58.160 ;
        RECT 2.400 57.480 111.200 58.120 ;
        RECT 2.800 56.760 111.200 57.480 ;
        RECT 2.800 56.080 111.600 56.760 ;
        RECT 2.400 54.760 111.600 56.080 ;
        RECT 2.800 53.360 111.600 54.760 ;
        RECT 2.400 52.720 111.600 53.360 ;
        RECT 2.800 51.320 111.600 52.720 ;
        RECT 2.400 50.680 111.600 51.320 ;
        RECT 2.800 49.280 111.600 50.680 ;
        RECT 2.400 47.960 111.600 49.280 ;
        RECT 2.800 46.560 111.600 47.960 ;
        RECT 2.400 45.920 111.600 46.560 ;
        RECT 2.800 44.520 111.600 45.920 ;
        RECT 2.400 43.200 111.600 44.520 ;
        RECT 2.800 41.800 111.600 43.200 ;
        RECT 2.400 41.160 111.600 41.800 ;
        RECT 2.800 39.760 111.600 41.160 ;
        RECT 2.400 38.440 111.600 39.760 ;
        RECT 2.800 37.040 111.600 38.440 ;
        RECT 2.400 36.400 111.600 37.040 ;
        RECT 2.800 35.000 111.600 36.400 ;
        RECT 2.400 34.360 111.600 35.000 ;
        RECT 2.800 32.960 111.600 34.360 ;
        RECT 2.400 31.640 111.600 32.960 ;
        RECT 2.800 30.240 111.600 31.640 ;
        RECT 2.400 29.600 111.600 30.240 ;
        RECT 2.800 28.200 111.600 29.600 ;
        RECT 2.400 26.880 111.600 28.200 ;
        RECT 2.800 25.480 111.600 26.880 ;
        RECT 2.400 24.840 111.600 25.480 ;
        RECT 2.800 23.440 111.600 24.840 ;
        RECT 2.400 22.120 111.600 23.440 ;
        RECT 2.800 20.720 111.600 22.120 ;
        RECT 2.400 20.080 111.600 20.720 ;
        RECT 2.800 18.680 111.600 20.080 ;
        RECT 2.400 18.040 111.600 18.680 ;
        RECT 2.800 16.640 111.600 18.040 ;
        RECT 2.400 15.320 111.600 16.640 ;
        RECT 2.800 13.920 111.600 15.320 ;
        RECT 2.400 13.280 111.600 13.920 ;
        RECT 2.800 11.880 111.600 13.280 ;
        RECT 2.400 10.560 111.600 11.880 ;
        RECT 2.800 9.160 111.600 10.560 ;
        RECT 2.400 8.520 111.600 9.160 ;
        RECT 2.800 7.120 111.600 8.520 ;
        RECT 2.400 5.800 111.600 7.120 ;
        RECT 2.800 4.400 111.600 5.800 ;
        RECT 2.400 3.760 111.600 4.400 ;
        RECT 2.800 2.360 111.600 3.760 ;
        RECT 2.400 1.720 111.600 2.360 ;
        RECT 2.800 0.855 111.600 1.720 ;
      LAYER met4 ;
        RECT 56.200 10.640 92.120 100.880 ;
  END
END sb_2__0_
END LIBRARY

