magic
tech EFS8A
magscale 1 2
timestamp 1602527098
<< locali >>
rect 23155 43809 23190 43843
rect 24995 43809 25122 43843
rect 25271 42721 25306 42755
rect 32447 42721 32482 42755
rect 38151 42721 38186 42755
rect 39899 42721 39934 42755
rect 34069 42143 34103 42245
rect 22195 39593 22201 39627
rect 32499 39593 32505 39627
rect 22195 39525 22229 39593
rect 32499 39525 32533 39593
rect 25179 39457 25214 39491
rect 37099 38743 37133 38811
rect 42901 38743 42935 38981
rect 37099 38709 37105 38743
rect 43499 38505 43545 38539
rect 19015 38369 19142 38403
rect 25329 37723 25363 37825
rect 26887 37655 26921 37723
rect 26887 37621 26893 37655
rect 43303 37281 43430 37315
rect 5043 36125 5181 36159
rect 20545 35547 20579 35785
rect 4715 35241 4721 35275
rect 13087 35241 13093 35275
rect 21275 35241 21281 35275
rect 4715 35173 4749 35241
rect 11667 35173 11713 35207
rect 13087 35173 13121 35241
rect 21275 35173 21309 35241
rect 40635 35105 40670 35139
rect 43303 35105 43430 35139
rect 7239 34493 7274 34527
rect 4807 34391 4841 34459
rect 4807 34357 4813 34391
rect 32275 34153 32413 34187
rect 32079 34017 32206 34051
rect 33459 34017 33494 34051
rect 34471 34017 34506 34051
rect 16543 33609 16589 33643
rect 9367 33541 9505 33575
rect 31953 33303 31987 33609
rect 7843 33065 7849 33099
rect 23575 33065 23581 33099
rect 7843 32997 7877 33065
rect 23575 32997 23609 33065
rect 32447 32997 32492 33031
rect 43303 32929 43430 32963
rect 26663 32725 26801 32759
rect 23023 31977 23029 32011
rect 29923 31977 29929 32011
rect 23023 31909 23057 31977
rect 29923 31909 29957 31977
rect 21499 31841 21626 31875
rect 40647 31433 40785 31467
rect 38243 31229 38278 31263
rect 24041 31127 24075 31229
rect 4623 30889 4629 30923
rect 19251 30889 19257 30923
rect 4623 30821 4657 30889
rect 11287 30821 11332 30855
rect 19251 30821 19285 30889
rect 41187 30753 41222 30787
rect 32781 30039 32815 30209
rect 4623 28951 4657 29019
rect 38479 28997 38513 29019
rect 4623 28917 4629 28951
rect 38479 28936 38513 28963
rect 18279 28577 18314 28611
rect 21275 27625 21281 27659
rect 29739 27625 29745 27659
rect 21275 27557 21309 27625
rect 29739 27557 29773 27625
rect 19843 27489 19878 27523
rect 40601 26911 40635 26945
rect 40601 26877 40762 26911
rect 7015 26537 7021 26571
rect 36271 26537 36277 26571
rect 7015 26469 7049 26537
rect 36271 26469 36305 26537
rect 34839 26401 34874 26435
rect 21275 25449 21281 25483
rect 21275 25381 21309 25449
rect 23523 25313 23650 25347
rect 30699 25313 30826 25347
rect 36369 25313 36530 25347
rect 43303 25313 43430 25347
rect 36369 25211 36403 25313
rect 2145 24735 2179 24837
rect 33333 24599 33367 24905
rect 32689 24259 32723 24293
rect 32689 24225 32850 24259
rect 37565 24225 37818 24259
rect 37565 24123 37599 24225
rect 4353 23511 4387 23749
rect 30941 23579 30975 23817
rect 32499 23273 32505 23307
rect 32499 23205 32533 23273
rect 44959 23137 44994 23171
rect 33149 22967 33183 23137
rect 22845 22559 22879 22661
rect 13731 22423 13765 22491
rect 13731 22389 13737 22423
rect 5543 22185 5549 22219
rect 23299 22185 23305 22219
rect 4445 21879 4479 22185
rect 5543 22117 5577 22185
rect 23299 22117 23333 22185
rect 14231 22049 14266 22083
rect 31861 21471 31895 21641
rect 14283 21335 14317 21403
rect 14283 21301 14289 21335
rect 33327 21097 33333 21131
rect 33327 21029 33361 21097
rect 38485 20961 38646 20995
rect 38485 20859 38519 20961
rect 30481 20383 30515 20553
rect 37657 20383 37691 20485
rect 14191 20247 14225 20315
rect 31677 20247 31711 20349
rect 14191 20213 14197 20247
rect 4715 20009 4721 20043
rect 13823 20009 13829 20043
rect 32591 20009 32597 20043
rect 4715 19941 4749 20009
rect 13823 19941 13857 20009
rect 32591 19941 32625 20009
rect 45051 19873 45086 19907
rect 4715 19159 4749 19227
rect 13277 19159 13311 19397
rect 4715 19125 4721 19159
rect 7199 18921 7205 18955
rect 10879 18921 10885 18955
rect 21051 18921 21189 18955
rect 7199 18853 7233 18921
rect 10879 18853 10913 18921
rect 31067 18785 31102 18819
rect 15663 17833 15669 17867
rect 15663 17765 15697 17833
rect 33057 17119 33091 17221
rect 35357 17085 35518 17119
rect 35357 17051 35391 17085
rect 12167 16745 12173 16779
rect 34339 16745 34345 16779
rect 12167 16677 12201 16745
rect 34339 16677 34373 16745
rect 24535 16609 24662 16643
rect 44959 16609 44994 16643
rect 23305 16099 23339 16201
rect 38393 15963 38427 16201
rect 5083 15895 5117 15963
rect 42619 15895 42653 15963
rect 5083 15861 5089 15895
rect 42619 15861 42625 15895
rect 21683 15521 21718 15555
rect 34195 15521 34230 15555
rect 35115 15521 35242 15555
rect 36219 15521 36254 15555
rect 23811 15113 23949 15147
rect 9689 14807 9723 15045
rect 23397 14807 23431 14977
rect 6975 14773 7113 14807
rect 26467 14433 26594 14467
rect 38485 14433 38646 14467
rect 38485 14263 38519 14433
rect 12587 14025 12725 14059
rect 24811 13345 24846 13379
rect 28675 13345 28802 13379
rect 37691 13345 37818 13379
rect 43303 13345 43430 13379
rect 17693 12631 17727 12801
rect 18423 12631 18457 12699
rect 18423 12597 18429 12631
rect 29003 12393 29009 12427
rect 29003 12325 29037 12393
rect 8527 12257 8654 12291
rect 11621 12257 11782 12291
rect 36679 12257 36714 12291
rect 11621 12087 11655 12257
rect 20079 11543 20113 11611
rect 20079 11509 20085 11543
rect 28675 11169 28802 11203
rect 18003 10557 18130 10591
rect 25415 10455 25449 10523
rect 25415 10421 25421 10455
rect 36087 10217 36093 10251
rect 36087 10149 36121 10217
rect 25053 9435 25087 9673
rect 20079 9367 20113 9435
rect 20079 9333 20085 9367
rect 11247 9129 11253 9163
rect 11247 9061 11281 9129
rect 33643 8993 33678 9027
rect 36587 8993 36622 9027
rect 21051 8041 21189 8075
rect 14105 7939 14139 7973
rect 13127 7905 13162 7939
rect 14105 7905 14266 7939
<< viali >>
rect 30732 44285 30766 44319
rect 31125 44285 31159 44319
rect 33216 44285 33250 44319
rect 33609 44285 33643 44319
rect 30803 44149 30837 44183
rect 33287 44149 33321 44183
rect 32505 43945 32539 43979
rect 33425 43877 33459 43911
rect 23121 43809 23155 43843
rect 24961 43809 24995 43843
rect 30456 43809 30490 43843
rect 33333 43741 33367 43775
rect 33609 43741 33643 43775
rect 23259 43605 23293 43639
rect 23765 43605 23799 43639
rect 24041 43605 24075 43639
rect 25191 43605 25225 43639
rect 25605 43605 25639 43639
rect 30527 43605 30561 43639
rect 31033 43605 31067 43639
rect 31309 43605 31343 43639
rect 23121 43401 23155 43435
rect 25053 43401 25087 43435
rect 30389 43401 30423 43435
rect 30849 43401 30883 43435
rect 33885 43401 33919 43435
rect 24317 43333 24351 43367
rect 23765 43265 23799 43299
rect 25789 43265 25823 43299
rect 30067 43265 30101 43299
rect 31033 43265 31067 43299
rect 32597 43265 32631 43299
rect 32873 43265 32907 43299
rect 22604 43197 22638 43231
rect 27445 43197 27479 43231
rect 27537 43197 27571 43231
rect 27997 43197 28031 43231
rect 29980 43197 30014 43231
rect 34964 43197 34998 43231
rect 23857 43129 23891 43163
rect 24777 43129 24811 43163
rect 25513 43129 25547 43163
rect 25605 43129 25639 43163
rect 31125 43129 31159 43163
rect 31677 43129 31711 43163
rect 32689 43129 32723 43163
rect 22385 43061 22419 43095
rect 22707 43061 22741 43095
rect 27629 43061 27663 43095
rect 32321 43061 32355 43095
rect 33609 43061 33643 43095
rect 35035 43061 35069 43095
rect 35449 43061 35483 43095
rect 27629 42857 27663 42891
rect 23581 42789 23615 42823
rect 23673 42789 23707 42823
rect 24225 42789 24259 42823
rect 26617 42789 26651 42823
rect 26709 42789 26743 42823
rect 30573 42789 30607 42823
rect 30665 42789 30699 42823
rect 31217 42789 31251 42823
rect 33609 42789 33643 42823
rect 35081 42789 35115 42823
rect 35173 42789 35207 42823
rect 22452 42721 22486 42755
rect 25237 42721 25271 42755
rect 29193 42721 29227 42755
rect 29469 42721 29503 42755
rect 32413 42721 32447 42755
rect 38117 42721 38151 42755
rect 39865 42721 39899 42755
rect 26893 42653 26927 42687
rect 29653 42653 29687 42687
rect 33517 42653 33551 42687
rect 35541 42653 35575 42687
rect 34069 42585 34103 42619
rect 22523 42517 22557 42551
rect 24501 42517 24535 42551
rect 25375 42517 25409 42551
rect 25697 42517 25731 42551
rect 32551 42517 32585 42551
rect 38255 42517 38289 42551
rect 38577 42517 38611 42551
rect 40003 42517 40037 42551
rect 25329 42313 25363 42347
rect 30665 42313 30699 42347
rect 31033 42313 31067 42347
rect 33103 42313 33137 42347
rect 34253 42313 34287 42347
rect 34713 42313 34747 42347
rect 35725 42313 35759 42347
rect 39865 42313 39899 42347
rect 21925 42245 21959 42279
rect 26617 42245 26651 42279
rect 28365 42245 28399 42279
rect 31309 42245 31343 42279
rect 32091 42245 32125 42279
rect 33793 42245 33827 42279
rect 34069 42245 34103 42279
rect 22109 42177 22143 42211
rect 23765 42177 23799 42211
rect 24409 42177 24443 42211
rect 25605 42177 25639 42211
rect 26985 42177 27019 42211
rect 27445 42177 27479 42211
rect 29745 42177 29779 42211
rect 33425 42177 33459 42211
rect 36369 42177 36403 42211
rect 38485 42177 38519 42211
rect 39405 42177 39439 42211
rect 21072 42109 21106 42143
rect 21465 42109 21499 42143
rect 32020 42109 32054 42143
rect 33032 42109 33066 42143
rect 34069 42109 34103 42143
rect 34964 42109 34998 42143
rect 35944 42109 35978 42143
rect 37448 42109 37482 42143
rect 40544 42109 40578 42143
rect 40969 42109 41003 42143
rect 22201 42041 22235 42075
rect 22753 42041 22787 42075
rect 23857 42041 23891 42075
rect 25697 42041 25731 42075
rect 26249 42041 26283 42075
rect 27766 42041 27800 42075
rect 29009 42041 29043 42075
rect 30066 42041 30100 42075
rect 36047 42041 36081 42075
rect 37933 42041 37967 42075
rect 38577 42041 38611 42075
rect 39129 42041 39163 42075
rect 21143 41973 21177 42007
rect 23121 41973 23155 42007
rect 23489 41973 23523 42007
rect 24685 41973 24719 42007
rect 27261 41973 27295 42007
rect 29561 41973 29595 42007
rect 32505 41973 32539 42007
rect 32873 41973 32907 42007
rect 35035 41973 35069 42007
rect 35449 41973 35483 42007
rect 37519 41973 37553 42007
rect 38209 41973 38243 42007
rect 40647 41973 40681 42007
rect 22109 41769 22143 41803
rect 22339 41769 22373 41803
rect 24225 41769 24259 41803
rect 25283 41769 25317 41803
rect 25697 41769 25731 41803
rect 26249 41769 26283 41803
rect 29929 41769 29963 41803
rect 34897 41769 34931 41803
rect 23305 41701 23339 41735
rect 23397 41701 23431 41735
rect 23949 41701 23983 41735
rect 26709 41701 26743 41735
rect 30665 41701 30699 41735
rect 33701 41701 33735 41735
rect 33793 41701 33827 41735
rect 35265 41701 35299 41735
rect 35357 41701 35391 41735
rect 38669 41701 38703 41735
rect 40325 41701 40359 41735
rect 40417 41701 40451 41735
rect 42257 41701 42291 41735
rect 22236 41633 22270 41667
rect 25212 41633 25246 41667
rect 29193 41633 29227 41667
rect 29469 41633 29503 41667
rect 32632 41633 32666 41667
rect 41864 41633 41898 41667
rect 26617 41565 26651 41599
rect 26893 41565 26927 41599
rect 28825 41565 28859 41599
rect 29653 41565 29687 41599
rect 30297 41565 30331 41599
rect 30573 41565 30607 41599
rect 31217 41565 31251 41599
rect 34069 41565 34103 41599
rect 35541 41565 35575 41599
rect 38577 41565 38611 41599
rect 40601 41565 40635 41599
rect 39129 41497 39163 41531
rect 32735 41429 32769 41463
rect 36645 41429 36679 41463
rect 41935 41429 41969 41463
rect 23305 41225 23339 41259
rect 24777 41225 24811 41259
rect 28181 41225 28215 41259
rect 29929 41225 29963 41259
rect 31033 41225 31067 41259
rect 31309 41225 31343 41259
rect 33333 41225 33367 41259
rect 37841 41225 37875 41259
rect 26525 41157 26559 41191
rect 27905 41157 27939 41191
rect 25053 41089 25087 41123
rect 26985 41089 27019 41123
rect 30113 41089 30147 41123
rect 31953 41089 31987 41123
rect 32229 41089 32263 41123
rect 34989 41089 35023 41123
rect 35265 41089 35299 41123
rect 38485 41089 38519 41123
rect 39405 41089 39439 41123
rect 40601 41089 40635 41123
rect 40877 41089 40911 41123
rect 42441 41089 42475 41123
rect 21868 41021 21902 41055
rect 22293 41021 22327 41055
rect 23740 41021 23774 41055
rect 24133 41021 24167 41055
rect 25237 41021 25271 41055
rect 33492 41021 33526 41055
rect 33885 41021 33919 41055
rect 36645 41021 36679 41055
rect 37565 41021 37599 41055
rect 21971 40953 22005 40987
rect 25558 40953 25592 40987
rect 26801 40953 26835 40987
rect 27306 40953 27340 40987
rect 30435 40953 30469 40987
rect 32045 40953 32079 40987
rect 34713 40953 34747 40987
rect 35081 40953 35115 40987
rect 37007 40953 37041 40987
rect 38301 40953 38335 40987
rect 38577 40953 38611 40987
rect 39129 40953 39163 40987
rect 40693 40953 40727 40987
rect 42165 40953 42199 40987
rect 42257 40953 42291 40987
rect 22661 40885 22695 40919
rect 23811 40885 23845 40919
rect 26157 40885 26191 40919
rect 29009 40885 29043 40919
rect 29561 40885 29595 40919
rect 31677 40885 31711 40919
rect 32873 40885 32907 40919
rect 33563 40885 33597 40919
rect 34345 40885 34379 40919
rect 35909 40885 35943 40919
rect 36553 40885 36587 40919
rect 39957 40885 39991 40919
rect 40233 40885 40267 40919
rect 41889 40885 41923 40919
rect 43085 40885 43119 40919
rect 23397 40681 23431 40715
rect 25329 40681 25363 40715
rect 27445 40681 27479 40715
rect 29929 40681 29963 40715
rect 30941 40681 30975 40715
rect 31953 40681 31987 40715
rect 35725 40681 35759 40715
rect 38255 40681 38289 40715
rect 40417 40681 40451 40715
rect 40785 40681 40819 40715
rect 43545 40681 43579 40715
rect 22569 40613 22603 40647
rect 24133 40613 24167 40647
rect 30383 40613 30417 40647
rect 33425 40613 33459 40647
rect 33517 40613 33551 40647
rect 34069 40613 34103 40647
rect 36645 40613 36679 40647
rect 40095 40613 40129 40647
rect 41797 40613 41831 40647
rect 42349 40613 42383 40647
rect 21408 40545 21442 40579
rect 27629 40545 27663 40579
rect 27905 40545 27939 40579
rect 29009 40545 29043 40579
rect 32137 40545 32171 40579
rect 34932 40545 34966 40579
rect 35909 40545 35943 40579
rect 36369 40545 36403 40579
rect 38152 40545 38186 40579
rect 38577 40545 38611 40579
rect 39992 40545 40026 40579
rect 22477 40477 22511 40511
rect 22753 40477 22787 40511
rect 24041 40477 24075 40511
rect 24409 40477 24443 40511
rect 30021 40477 30055 40511
rect 35449 40477 35483 40511
rect 41705 40477 41739 40511
rect 21511 40409 21545 40443
rect 29193 40409 29227 40443
rect 27077 40341 27111 40375
rect 29561 40341 29595 40375
rect 31217 40341 31251 40375
rect 32321 40341 32355 40375
rect 35035 40341 35069 40375
rect 38945 40341 38979 40375
rect 41521 40341 41555 40375
rect 23397 40137 23431 40171
rect 24869 40137 24903 40171
rect 32137 40137 32171 40171
rect 35081 40137 35115 40171
rect 36277 40137 36311 40171
rect 38117 40137 38151 40171
rect 39681 40137 39715 40171
rect 21419 40069 21453 40103
rect 30665 40069 30699 40103
rect 39957 40069 39991 40103
rect 25513 40001 25547 40035
rect 25789 40001 25823 40035
rect 30021 40001 30055 40035
rect 33333 40001 33367 40035
rect 33609 40001 33643 40035
rect 38669 40001 38703 40035
rect 41981 40001 42015 40035
rect 43269 40001 43303 40035
rect 43545 40001 43579 40035
rect 12516 39933 12550 39967
rect 21348 39933 21382 39967
rect 23740 39933 23774 39967
rect 24133 39933 24167 39967
rect 26801 39933 26835 39967
rect 27537 39933 27571 39967
rect 27813 39933 27847 39967
rect 28273 39933 28307 39967
rect 29469 39933 29503 39967
rect 29745 39933 29779 39967
rect 30849 39933 30883 39967
rect 31309 39933 31343 39967
rect 35265 39933 35299 39967
rect 35725 39933 35759 39967
rect 36001 39933 36035 39967
rect 36829 39933 36863 39967
rect 40636 39933 40670 39967
rect 41061 39933 41095 39967
rect 22201 39865 22235 39899
rect 25605 39865 25639 39899
rect 27169 39865 27203 39899
rect 29101 39865 29135 39899
rect 31585 39865 31619 39899
rect 32781 39865 32815 39899
rect 33149 39865 33183 39899
rect 33425 39865 33459 39899
rect 37150 39865 37184 39899
rect 38761 39865 38795 39899
rect 39313 39865 39347 39899
rect 41705 39865 41739 39899
rect 41797 39865 41831 39899
rect 43085 39865 43119 39899
rect 43361 39865 43395 39899
rect 12587 39797 12621 39831
rect 13001 39797 13035 39831
rect 21741 39797 21775 39831
rect 22293 39797 22327 39831
rect 22845 39797 22879 39831
rect 23811 39797 23845 39831
rect 24501 39797 24535 39831
rect 25329 39797 25363 39831
rect 27353 39797 27387 39831
rect 28733 39797 28767 39831
rect 30297 39797 30331 39831
rect 36737 39797 36771 39831
rect 37749 39797 37783 39831
rect 40739 39797 40773 39831
rect 41521 39797 41555 39831
rect 42625 39797 42659 39831
rect 22201 39593 22235 39627
rect 23029 39593 23063 39627
rect 27629 39593 27663 39627
rect 28181 39593 28215 39627
rect 30021 39593 30055 39627
rect 32505 39593 32539 39627
rect 33057 39593 33091 39627
rect 33701 39593 33735 39627
rect 36921 39593 36955 39627
rect 41613 39593 41647 39627
rect 43499 39593 43533 39627
rect 23765 39525 23799 39559
rect 26709 39525 26743 39559
rect 30665 39525 30699 39559
rect 33425 39525 33459 39559
rect 33977 39525 34011 39559
rect 34069 39525 34103 39559
rect 38669 39525 38703 39559
rect 40233 39525 40267 39559
rect 41797 39525 41831 39559
rect 41889 39525 41923 39559
rect 11989 39457 12023 39491
rect 14013 39457 14047 39491
rect 15368 39457 15402 39491
rect 25145 39457 25179 39491
rect 28365 39457 28399 39491
rect 28549 39457 28583 39491
rect 32137 39457 32171 39491
rect 36185 39457 36219 39491
rect 36369 39457 36403 39491
rect 42441 39457 42475 39491
rect 43396 39457 43430 39491
rect 12357 39389 12391 39423
rect 21833 39389 21867 39423
rect 23673 39389 23707 39423
rect 25605 39389 25639 39423
rect 26617 39389 26651 39423
rect 26893 39389 26927 39423
rect 30573 39389 30607 39423
rect 35265 39389 35299 39423
rect 36645 39389 36679 39423
rect 38577 39389 38611 39423
rect 40141 39389 40175 39423
rect 40417 39389 40451 39423
rect 24225 39321 24259 39355
rect 31125 39321 31159 39355
rect 31585 39321 31619 39355
rect 34529 39321 34563 39355
rect 39129 39321 39163 39355
rect 14197 39253 14231 39287
rect 15439 39253 15473 39287
rect 22753 39253 22787 39287
rect 25283 39253 25317 39287
rect 29561 39253 29595 39287
rect 35725 39253 35759 39287
rect 22201 39049 22235 39083
rect 23489 39049 23523 39083
rect 24685 39049 24719 39083
rect 30481 39049 30515 39083
rect 30757 39049 30791 39083
rect 32689 39049 32723 39083
rect 38577 39049 38611 39083
rect 39773 39049 39807 39083
rect 40831 39049 40865 39083
rect 43177 39049 43211 39083
rect 26617 38981 26651 39015
rect 28365 38981 28399 39015
rect 31953 38981 31987 39015
rect 37657 38981 37691 39015
rect 39313 38981 39347 39015
rect 42809 38981 42843 39015
rect 42901 38981 42935 39015
rect 11161 38913 11195 38947
rect 21189 38913 21223 38947
rect 24225 38913 24259 38947
rect 25789 38913 25823 38947
rect 26985 38913 27019 38947
rect 27445 38913 27479 38947
rect 31401 38913 31435 38947
rect 34345 38913 34379 38947
rect 36737 38913 36771 38947
rect 42073 38913 42107 38947
rect 11897 38845 11931 38879
rect 12516 38845 12550 38879
rect 12909 38845 12943 38879
rect 13645 38845 13679 38879
rect 14381 38845 14415 38879
rect 14841 38845 14875 38879
rect 15352 38845 15386 38879
rect 16380 38845 16414 38879
rect 20704 38845 20738 38879
rect 21716 38845 21750 38879
rect 29101 38845 29135 38879
rect 29561 38845 29595 38879
rect 35265 38845 35299 38879
rect 35725 38845 35759 38879
rect 40760 38845 40794 38879
rect 10885 38777 10919 38811
rect 10977 38777 11011 38811
rect 13737 38777 13771 38811
rect 15439 38777 15473 38811
rect 23765 38777 23799 38811
rect 23857 38777 23891 38811
rect 25513 38777 25547 38811
rect 25605 38777 25639 38811
rect 27766 38777 27800 38811
rect 29882 38777 29916 38811
rect 31493 38777 31527 38811
rect 33333 38777 33367 38811
rect 33425 38777 33459 38811
rect 33977 38777 34011 38811
rect 34713 38777 34747 38811
rect 35909 38777 35943 38811
rect 38761 38777 38795 38811
rect 38853 38777 38887 38811
rect 41797 38777 41831 38811
rect 41889 38777 41923 38811
rect 43637 38913 43671 38947
rect 43361 38777 43395 38811
rect 43453 38777 43487 38811
rect 10701 38709 10735 38743
rect 12587 38709 12621 38743
rect 15853 38709 15887 38743
rect 16129 38709 16163 38743
rect 16451 38709 16485 38743
rect 16865 38709 16899 38743
rect 20775 38709 20809 38743
rect 21465 38709 21499 38743
rect 21787 38709 21821 38743
rect 22477 38709 22511 38743
rect 23029 38709 23063 38743
rect 25237 38709 25271 38743
rect 27261 38709 27295 38743
rect 28733 38709 28767 38743
rect 31125 38709 31159 38743
rect 32321 38709 32355 38743
rect 33057 38709 33091 38743
rect 36277 38709 36311 38743
rect 36645 38709 36679 38743
rect 37105 38709 37139 38743
rect 38117 38709 38151 38743
rect 40049 38709 40083 38743
rect 41153 38709 41187 38743
rect 41613 38709 41647 38743
rect 42901 38709 42935 38743
rect 44281 38709 44315 38743
rect 23765 38505 23799 38539
rect 26249 38505 26283 38539
rect 28089 38505 28123 38539
rect 29285 38505 29319 38539
rect 30757 38505 30791 38539
rect 32597 38505 32631 38539
rect 33333 38505 33367 38539
rect 34621 38505 34655 38539
rect 37105 38505 37139 38539
rect 38669 38505 38703 38539
rect 41521 38505 41555 38539
rect 42165 38505 42199 38539
rect 43545 38505 43579 38539
rect 9873 38437 9907 38471
rect 13829 38437 13863 38471
rect 15485 38437 15519 38471
rect 21005 38437 21039 38471
rect 21097 38437 21131 38471
rect 22845 38437 22879 38471
rect 22937 38437 22971 38471
rect 24225 38437 24259 38471
rect 24409 38437 24443 38471
rect 24501 38437 24535 38471
rect 26617 38437 26651 38471
rect 26709 38437 26743 38471
rect 33701 38437 33735 38471
rect 33793 38437 33827 38471
rect 36001 38437 36035 38471
rect 38070 38437 38104 38471
rect 38945 38437 38979 38471
rect 39818 38437 39852 38471
rect 11897 38369 11931 38403
rect 16932 38369 16966 38403
rect 18981 38369 19015 38403
rect 29285 38369 29319 38403
rect 29561 38369 29595 38403
rect 30573 38369 30607 38403
rect 36093 38369 36127 38403
rect 36553 38369 36587 38403
rect 36829 38369 36863 38403
rect 39497 38369 39531 38403
rect 40417 38369 40451 38403
rect 43428 38369 43462 38403
rect 9781 38301 9815 38335
rect 10057 38301 10091 38335
rect 10793 38301 10827 38335
rect 11253 38301 11287 38335
rect 13737 38301 13771 38335
rect 15393 38301 15427 38335
rect 15669 38301 15703 38335
rect 21649 38301 21683 38335
rect 24685 38301 24719 38335
rect 26893 38301 26927 38335
rect 34345 38301 34379 38335
rect 37749 38301 37783 38335
rect 39313 38301 39347 38335
rect 41705 38301 41739 38335
rect 9413 38233 9447 38267
rect 14289 38233 14323 38267
rect 17003 38233 17037 38267
rect 23397 38233 23431 38267
rect 31401 38233 31435 38267
rect 42533 38233 42567 38267
rect 7665 38165 7699 38199
rect 19211 38165 19245 38199
rect 19625 38165 19659 38199
rect 21925 38165 21959 38199
rect 25513 38165 25547 38199
rect 30205 38165 30239 38199
rect 35265 38165 35299 38199
rect 11897 37961 11931 37995
rect 12633 37961 12667 37995
rect 12909 37961 12943 37995
rect 13645 37961 13679 37995
rect 14197 37961 14231 37995
rect 15209 37961 15243 37995
rect 17785 37961 17819 37995
rect 19073 37961 19107 37995
rect 20637 37961 20671 37995
rect 22845 37961 22879 37995
rect 23489 37961 23523 37995
rect 25145 37961 25179 37995
rect 27445 37961 27479 37995
rect 29101 37961 29135 37995
rect 29929 37961 29963 37995
rect 31033 37961 31067 37995
rect 34069 37961 34103 37995
rect 37013 37961 37047 37995
rect 38117 37961 38151 37995
rect 38853 37961 38887 37995
rect 39865 37961 39899 37995
rect 40923 37961 40957 37995
rect 41705 37961 41739 37995
rect 10241 37893 10275 37927
rect 28089 37893 28123 37927
rect 33425 37893 33459 37927
rect 33793 37893 33827 37927
rect 8309 37825 8343 37859
rect 9873 37825 9907 37859
rect 15301 37825 15335 37859
rect 19533 37825 19567 37859
rect 21005 37825 21039 37859
rect 21649 37825 21683 37859
rect 21925 37825 21959 37859
rect 25329 37825 25363 37859
rect 26341 37825 26375 37859
rect 31309 37825 31343 37859
rect 35265 37825 35299 37859
rect 37197 37825 37231 37859
rect 39083 37825 39117 37859
rect 41889 37825 41923 37859
rect 42165 37825 42199 37859
rect 12449 37757 12483 37791
rect 13829 37757 13863 37791
rect 15945 37757 15979 37791
rect 16865 37757 16899 37791
rect 17325 37757 17359 37791
rect 18096 37757 18130 37791
rect 18521 37757 18555 37791
rect 24225 37757 24259 37791
rect 26525 37757 26559 37791
rect 27721 37757 27755 37791
rect 29561 37757 29595 37791
rect 30113 37757 30147 37791
rect 32505 37757 32539 37791
rect 38393 37757 38427 37791
rect 38996 37757 39030 37791
rect 40820 37757 40854 37791
rect 41245 37757 41279 37791
rect 43428 37757 43462 37791
rect 44189 37757 44223 37791
rect 7665 37689 7699 37723
rect 7757 37689 7791 37723
rect 9045 37689 9079 37723
rect 9229 37689 9263 37723
rect 9330 37689 9364 37723
rect 10885 37689 10919 37723
rect 10977 37689 11011 37723
rect 11529 37689 11563 37723
rect 14841 37689 14875 37723
rect 19625 37689 19659 37723
rect 20177 37689 20211 37723
rect 21741 37689 21775 37723
rect 24546 37689 24580 37723
rect 25329 37689 25363 37723
rect 30434 37689 30468 37723
rect 32321 37689 32355 37723
rect 32826 37689 32860 37723
rect 34989 37689 35023 37723
rect 35081 37689 35115 37723
rect 36553 37689 36587 37723
rect 37519 37689 37553 37723
rect 39497 37689 39531 37723
rect 41981 37689 42015 37723
rect 7481 37621 7515 37655
rect 10701 37621 10735 37655
rect 17049 37621 17083 37655
rect 18199 37621 18233 37655
rect 21465 37621 21499 37655
rect 24041 37621 24075 37655
rect 25513 37621 25547 37655
rect 25973 37621 26007 37655
rect 26893 37621 26927 37655
rect 34621 37621 34655 37655
rect 36093 37621 36127 37655
rect 43499 37621 43533 37655
rect 43821 37621 43855 37655
rect 9229 37417 9263 37451
rect 10885 37417 10919 37451
rect 13829 37417 13863 37451
rect 15485 37417 15519 37451
rect 19901 37417 19935 37451
rect 23167 37417 23201 37451
rect 25053 37417 25087 37451
rect 26893 37417 26927 37451
rect 33793 37417 33827 37451
rect 37933 37417 37967 37451
rect 39589 37417 39623 37451
rect 40509 37417 40543 37451
rect 41705 37417 41739 37451
rect 41981 37417 42015 37451
rect 42441 37417 42475 37451
rect 7021 37349 7055 37383
rect 9873 37349 9907 37383
rect 11437 37349 11471 37383
rect 13001 37349 13035 37383
rect 19073 37349 19107 37383
rect 21373 37349 21407 37383
rect 21557 37349 21591 37383
rect 21649 37349 21683 37383
rect 22845 37349 22879 37383
rect 24454 37349 24488 37383
rect 30205 37349 30239 37383
rect 33235 37349 33269 37383
rect 39031 37349 39065 37383
rect 41106 37349 41140 37383
rect 16313 37281 16347 37315
rect 17928 37281 17962 37315
rect 23064 37281 23098 37315
rect 27077 37281 27111 37315
rect 27353 37281 27387 37315
rect 28365 37281 28399 37315
rect 29469 37281 29503 37315
rect 29929 37281 29963 37315
rect 31100 37281 31134 37315
rect 35725 37281 35759 37315
rect 36001 37281 36035 37315
rect 43269 37281 43303 37315
rect 6929 37213 6963 37247
rect 7205 37213 7239 37247
rect 9781 37213 9815 37247
rect 11345 37213 11379 37247
rect 11621 37213 11655 37247
rect 12909 37213 12943 37247
rect 13185 37213 13219 37247
rect 14197 37213 14231 37247
rect 15761 37213 15795 37247
rect 18015 37213 18049 37247
rect 18981 37213 19015 37247
rect 19349 37213 19383 37247
rect 21833 37213 21867 37247
rect 24133 37213 24167 37247
rect 32873 37213 32907 37247
rect 36185 37213 36219 37247
rect 38669 37213 38703 37247
rect 40785 37213 40819 37247
rect 10333 37145 10367 37179
rect 43499 37145 43533 37179
rect 18429 37077 18463 37111
rect 28549 37077 28583 37111
rect 29285 37077 29319 37111
rect 31171 37077 31205 37111
rect 32505 37077 32539 37111
rect 34897 37077 34931 37111
rect 37105 37077 37139 37111
rect 37473 37077 37507 37111
rect 5779 36873 5813 36907
rect 8125 36873 8159 36907
rect 8953 36873 8987 36907
rect 9321 36873 9355 36907
rect 9689 36873 9723 36907
rect 11621 36873 11655 36907
rect 12909 36873 12943 36907
rect 13829 36873 13863 36907
rect 16497 36873 16531 36907
rect 17877 36873 17911 36907
rect 27813 36873 27847 36907
rect 31125 36873 31159 36907
rect 32873 36873 32907 36907
rect 33793 36873 33827 36907
rect 34713 36873 34747 36907
rect 40233 36873 40267 36907
rect 41521 36873 41555 36907
rect 41889 36873 41923 36907
rect 26617 36805 26651 36839
rect 38485 36805 38519 36839
rect 7849 36737 7883 36771
rect 10517 36737 10551 36771
rect 13461 36737 13495 36771
rect 14013 36737 14047 36771
rect 14657 36737 14691 36771
rect 15853 36737 15887 36771
rect 17509 36737 17543 36771
rect 18337 36737 18371 36771
rect 22201 36737 22235 36771
rect 23029 36737 23063 36771
rect 24133 36737 24167 36771
rect 25697 36737 25731 36771
rect 27261 36737 27295 36771
rect 31493 36737 31527 36771
rect 32413 36737 32447 36771
rect 36185 36737 36219 36771
rect 37565 36737 37599 36771
rect 39129 36737 39163 36771
rect 39957 36737 39991 36771
rect 40601 36737 40635 36771
rect 40877 36737 40911 36771
rect 42165 36737 42199 36771
rect 42441 36737 42475 36771
rect 5676 36669 5710 36703
rect 23740 36669 23774 36703
rect 25053 36669 25087 36703
rect 25145 36669 25179 36703
rect 25605 36669 25639 36703
rect 26249 36669 26283 36703
rect 26801 36669 26835 36703
rect 27169 36669 27203 36703
rect 29561 36669 29595 36703
rect 29745 36669 29779 36703
rect 31677 36669 31711 36703
rect 32137 36669 32171 36703
rect 33292 36669 33326 36703
rect 35449 36669 35483 36703
rect 36001 36669 36035 36703
rect 37013 36669 37047 36703
rect 37473 36669 37507 36703
rect 38736 36669 38770 36703
rect 7205 36601 7239 36635
rect 7297 36601 7331 36635
rect 9873 36601 9907 36635
rect 9965 36601 9999 36635
rect 14105 36601 14139 36635
rect 15577 36601 15611 36635
rect 15669 36601 15703 36635
rect 18429 36601 18463 36635
rect 18981 36601 19015 36635
rect 19901 36601 19935 36635
rect 19993 36601 20027 36635
rect 20545 36601 20579 36635
rect 21925 36601 21959 36635
rect 22017 36601 22051 36635
rect 23397 36601 23431 36635
rect 29101 36601 29135 36635
rect 33379 36601 33413 36635
rect 40693 36601 40727 36635
rect 42257 36601 42291 36635
rect 5549 36533 5583 36567
rect 6193 36533 6227 36567
rect 6653 36533 6687 36567
rect 11345 36533 11379 36567
rect 15393 36533 15427 36567
rect 19257 36533 19291 36567
rect 19625 36533 19659 36567
rect 21189 36533 21223 36567
rect 21465 36533 21499 36567
rect 23811 36533 23845 36567
rect 24593 36533 24627 36567
rect 28365 36533 28399 36567
rect 29377 36533 29411 36567
rect 30297 36533 30331 36567
rect 35357 36533 35391 36567
rect 36553 36533 36587 36567
rect 36829 36533 36863 36567
rect 38807 36533 38841 36567
rect 39589 36533 39623 36567
rect 43361 36533 43395 36567
rect 12909 36329 12943 36363
rect 18521 36329 18555 36363
rect 18981 36329 19015 36363
rect 22201 36329 22235 36363
rect 25237 36329 25271 36363
rect 27629 36329 27663 36363
rect 29745 36329 29779 36363
rect 31769 36329 31803 36363
rect 34897 36329 34931 36363
rect 35817 36329 35851 36363
rect 37933 36329 37967 36363
rect 6101 36261 6135 36295
rect 6653 36261 6687 36295
rect 7665 36261 7699 36295
rect 8217 36261 8251 36295
rect 10241 36261 10275 36295
rect 10793 36261 10827 36295
rect 11805 36261 11839 36295
rect 17922 36261 17956 36295
rect 19487 36261 19521 36295
rect 19901 36261 19935 36295
rect 21373 36261 21407 36295
rect 24317 36261 24351 36295
rect 26709 36261 26743 36295
rect 30573 36261 30607 36295
rect 32873 36261 32907 36295
rect 33149 36261 33183 36295
rect 35449 36261 35483 36295
rect 39129 36261 39163 36295
rect 39221 36261 39255 36295
rect 40785 36261 40819 36295
rect 4972 36193 5006 36227
rect 5365 36193 5399 36227
rect 13896 36193 13930 36227
rect 16221 36193 16255 36227
rect 19400 36193 19434 36227
rect 22804 36193 22838 36227
rect 28917 36193 28951 36227
rect 29101 36193 29135 36227
rect 32413 36193 32447 36227
rect 32597 36193 32631 36227
rect 33736 36193 33770 36227
rect 34713 36193 34747 36227
rect 36093 36193 36127 36227
rect 36553 36193 36587 36227
rect 37749 36193 37783 36227
rect 42200 36193 42234 36227
rect 43428 36193 43462 36227
rect 5181 36125 5215 36159
rect 6009 36125 6043 36159
rect 7573 36125 7607 36159
rect 10149 36125 10183 36159
rect 11713 36125 11747 36159
rect 11989 36125 12023 36159
rect 16037 36125 16071 36159
rect 17601 36125 17635 36159
rect 21281 36125 21315 36159
rect 22891 36125 22925 36159
rect 24225 36125 24259 36159
rect 24501 36125 24535 36159
rect 26617 36125 26651 36159
rect 29377 36125 29411 36159
rect 30481 36125 30515 36159
rect 36829 36125 36863 36159
rect 39405 36125 39439 36159
rect 40693 36125 40727 36159
rect 41337 36125 41371 36159
rect 21833 36057 21867 36091
rect 27169 36057 27203 36091
rect 30021 36057 30055 36091
rect 31033 36057 31067 36091
rect 43499 36057 43533 36091
rect 4629 35989 4663 36023
rect 7113 35989 7147 36023
rect 9873 35989 9907 36023
rect 13645 35989 13679 36023
rect 13967 35989 14001 36023
rect 15577 35989 15611 36023
rect 24041 35989 24075 36023
rect 33839 35989 33873 36023
rect 42303 35989 42337 36023
rect 42993 35989 43027 36023
rect 5549 35785 5583 35819
rect 6009 35785 6043 35819
rect 10149 35785 10183 35819
rect 12173 35785 12207 35819
rect 16221 35785 16255 35819
rect 16865 35785 16899 35819
rect 19257 35785 19291 35819
rect 20545 35785 20579 35819
rect 20729 35785 20763 35819
rect 22845 35785 22879 35819
rect 28319 35785 28353 35819
rect 30573 35785 30607 35819
rect 31217 35785 31251 35819
rect 31585 35785 31619 35819
rect 32781 35785 32815 35819
rect 37105 35785 37139 35819
rect 38485 35785 38519 35819
rect 38945 35785 38979 35819
rect 39175 35785 39209 35819
rect 40325 35785 40359 35819
rect 40785 35785 40819 35819
rect 42441 35785 42475 35819
rect 3755 35717 3789 35751
rect 11897 35717 11931 35751
rect 14933 35717 14967 35751
rect 19993 35717 20027 35751
rect 6929 35649 6963 35683
rect 7573 35649 7607 35683
rect 11529 35649 11563 35683
rect 13645 35649 13679 35683
rect 14289 35649 14323 35683
rect 15485 35649 15519 35683
rect 3684 35581 3718 35615
rect 4629 35581 4663 35615
rect 12608 35581 12642 35615
rect 16681 35581 16715 35615
rect 21833 35717 21867 35751
rect 28089 35717 28123 35751
rect 34253 35717 34287 35751
rect 39957 35717 39991 35751
rect 21281 35649 21315 35683
rect 22201 35649 22235 35683
rect 23489 35649 23523 35683
rect 24133 35649 24167 35683
rect 24961 35649 24995 35683
rect 26985 35649 27019 35683
rect 31769 35649 31803 35683
rect 32413 35649 32447 35683
rect 41245 35649 41279 35683
rect 43085 35649 43119 35683
rect 43361 35649 43395 35683
rect 28248 35581 28282 35615
rect 29285 35581 29319 35615
rect 35909 35581 35943 35615
rect 36277 35581 36311 35615
rect 36461 35581 36495 35615
rect 37289 35581 37323 35615
rect 39072 35581 39106 35615
rect 39497 35581 39531 35615
rect 4950 35513 4984 35547
rect 6653 35513 6687 35547
rect 7021 35513 7055 35547
rect 9781 35513 9815 35547
rect 10885 35513 10919 35547
rect 10977 35513 11011 35547
rect 13093 35513 13127 35547
rect 13737 35513 13771 35547
rect 15209 35513 15243 35547
rect 15301 35513 15335 35547
rect 18337 35513 18371 35547
rect 18889 35513 18923 35547
rect 19441 35513 19475 35547
rect 19533 35513 19567 35547
rect 20545 35513 20579 35547
rect 21097 35513 21131 35547
rect 21373 35513 21407 35547
rect 24317 35513 24351 35547
rect 24409 35513 24443 35547
rect 26525 35513 26559 35547
rect 26617 35513 26651 35547
rect 29101 35513 29135 35547
rect 29606 35513 29640 35547
rect 31861 35513 31895 35547
rect 33333 35513 33367 35547
rect 33425 35513 33459 35547
rect 33977 35513 34011 35547
rect 35633 35513 35667 35547
rect 37610 35513 37644 35547
rect 41566 35513 41600 35547
rect 42809 35513 42843 35547
rect 43177 35513 43211 35547
rect 4169 35445 4203 35479
rect 4537 35445 4571 35479
rect 7849 35445 7883 35479
rect 8217 35445 8251 35479
rect 10701 35445 10735 35479
rect 12679 35445 12713 35479
rect 13369 35445 13403 35479
rect 14565 35445 14599 35479
rect 17233 35445 17267 35479
rect 17693 35445 17727 35479
rect 25237 35445 25271 35479
rect 25973 35445 26007 35479
rect 26249 35445 26283 35479
rect 27537 35445 27571 35479
rect 28641 35445 28675 35479
rect 30205 35445 30239 35479
rect 33057 35445 33091 35479
rect 35081 35445 35115 35479
rect 36737 35445 36771 35479
rect 38209 35445 38243 35479
rect 41061 35445 41095 35479
rect 42165 35445 42199 35479
rect 44005 35445 44039 35479
rect 4721 35241 4755 35275
rect 5273 35241 5307 35275
rect 6009 35241 6043 35275
rect 13093 35241 13127 35275
rect 13645 35241 13679 35275
rect 14013 35241 14047 35275
rect 19349 35241 19383 35275
rect 20729 35241 20763 35275
rect 21281 35241 21315 35275
rect 21833 35241 21867 35275
rect 22799 35241 22833 35275
rect 28917 35241 28951 35275
rect 30941 35241 30975 35275
rect 37289 35241 37323 35275
rect 41245 35241 41279 35275
rect 6422 35173 6456 35207
rect 8033 35173 8067 35207
rect 8585 35173 8619 35207
rect 9873 35173 9907 35207
rect 11713 35173 11747 35207
rect 15577 35173 15611 35207
rect 18791 35173 18825 35207
rect 19717 35173 19751 35207
rect 24317 35173 24351 35207
rect 24869 35173 24903 35207
rect 26709 35173 26743 35207
rect 29698 35173 29732 35207
rect 30665 35173 30699 35207
rect 32321 35173 32355 35207
rect 33885 35173 33919 35207
rect 35357 35173 35391 35207
rect 35449 35173 35483 35207
rect 39221 35173 39255 35207
rect 41889 35173 41923 35207
rect 7021 35105 7055 35139
rect 11596 35105 11630 35139
rect 17024 35105 17058 35139
rect 22728 35105 22762 35139
rect 28400 35105 28434 35139
rect 29377 35105 29411 35139
rect 30297 35105 30331 35139
rect 31677 35105 31711 35139
rect 38071 35105 38105 35139
rect 40601 35105 40635 35139
rect 43269 35105 43303 35139
rect 4353 35037 4387 35071
rect 6101 35037 6135 35071
rect 7941 35037 7975 35071
rect 9781 35037 9815 35071
rect 10425 35037 10459 35071
rect 12725 35037 12759 35071
rect 15485 35037 15519 35071
rect 18429 35037 18463 35071
rect 20913 35037 20947 35071
rect 22109 35037 22143 35071
rect 24225 35037 24259 35071
rect 26617 35037 26651 35071
rect 26893 35037 26927 35071
rect 32229 35037 32263 35071
rect 33793 35037 33827 35071
rect 34069 35037 34103 35071
rect 35633 35037 35667 35071
rect 38163 35037 38197 35071
rect 39129 35037 39163 35071
rect 40739 35037 40773 35071
rect 41797 35037 41831 35071
rect 42441 35037 42475 35071
rect 16037 34969 16071 35003
rect 32781 34969 32815 35003
rect 38853 34969 38887 35003
rect 39681 34969 39715 35003
rect 7297 34901 7331 34935
rect 8861 34901 8895 34935
rect 10885 34901 10919 34935
rect 17095 34901 17129 34935
rect 17601 34901 17635 34935
rect 18153 34901 18187 34935
rect 23765 34901 23799 34935
rect 26341 34901 26375 34935
rect 28503 34901 28537 34935
rect 33333 34901 33367 34935
rect 36277 34901 36311 34935
rect 42809 34901 42843 34935
rect 43499 34901 43533 34935
rect 7343 34697 7377 34731
rect 9321 34697 9355 34731
rect 11483 34697 11517 34731
rect 14657 34697 14691 34731
rect 15393 34697 15427 34731
rect 16589 34697 16623 34731
rect 17049 34697 17083 34731
rect 20269 34697 20303 34731
rect 21281 34697 21315 34731
rect 22845 34697 22879 34731
rect 24593 34697 24627 34731
rect 24869 34697 24903 34731
rect 28319 34697 28353 34731
rect 30113 34697 30147 34731
rect 31677 34697 31711 34731
rect 31953 34697 31987 34731
rect 33609 34697 33643 34731
rect 33839 34697 33873 34731
rect 35035 34697 35069 34731
rect 36093 34697 36127 34731
rect 36921 34697 36955 34731
rect 39773 34697 39807 34731
rect 41429 34697 41463 34731
rect 41797 34697 41831 34731
rect 42257 34697 42291 34731
rect 43453 34697 43487 34731
rect 10425 34629 10459 34663
rect 11161 34629 11195 34663
rect 15117 34629 15151 34663
rect 19165 34629 19199 34663
rect 22385 34629 22419 34663
rect 23489 34629 23523 34663
rect 25743 34629 25777 34663
rect 27261 34629 27295 34663
rect 29101 34629 29135 34663
rect 29745 34629 29779 34663
rect 32781 34629 32815 34663
rect 35725 34629 35759 34663
rect 40969 34629 41003 34663
rect 3571 34561 3605 34595
rect 7021 34561 7055 34595
rect 8309 34561 8343 34595
rect 9873 34561 9907 34595
rect 10793 34561 10827 34595
rect 13277 34561 13311 34595
rect 15669 34561 15703 34595
rect 16037 34561 16071 34595
rect 18613 34561 18647 34595
rect 19855 34561 19889 34595
rect 26709 34561 26743 34595
rect 27997 34561 28031 34595
rect 30389 34561 30423 34595
rect 31033 34561 31067 34595
rect 33149 34561 33183 34595
rect 34621 34561 34655 34595
rect 38853 34561 38887 34595
rect 42533 34561 42567 34595
rect 42809 34561 42843 34595
rect 3341 34493 3375 34527
rect 3468 34493 3502 34527
rect 4445 34493 4479 34527
rect 5641 34493 5675 34527
rect 7205 34493 7239 34527
rect 11412 34493 11446 34527
rect 12173 34493 12207 34527
rect 17877 34493 17911 34527
rect 18245 34493 18279 34527
rect 18521 34493 18555 34527
rect 19768 34493 19802 34527
rect 20796 34493 20830 34527
rect 23673 34493 23707 34527
rect 25672 34493 25706 34527
rect 26157 34493 26191 34527
rect 28248 34493 28282 34527
rect 29352 34493 29386 34527
rect 33768 34493 33802 34527
rect 34964 34493 34998 34527
rect 35449 34493 35483 34527
rect 36553 34493 36587 34527
rect 37013 34493 37047 34527
rect 40576 34493 40610 34527
rect 8401 34425 8435 34459
rect 8953 34425 8987 34459
rect 9965 34425 9999 34459
rect 12817 34425 12851 34459
rect 13185 34425 13219 34459
rect 13639 34425 13673 34459
rect 15761 34425 15795 34459
rect 20545 34425 20579 34459
rect 21833 34425 21867 34459
rect 21925 34425 21959 34459
rect 23994 34425 24028 34459
rect 26801 34425 26835 34459
rect 30481 34425 30515 34459
rect 32229 34425 32263 34459
rect 32321 34425 32355 34459
rect 34253 34425 34287 34459
rect 37375 34425 37409 34459
rect 38945 34425 38979 34459
rect 39497 34425 39531 34459
rect 42625 34425 42659 34459
rect 3985 34357 4019 34391
rect 4353 34357 4387 34391
rect 4813 34357 4847 34391
rect 5365 34357 5399 34391
rect 6101 34357 6135 34391
rect 6469 34357 6503 34391
rect 7941 34357 7975 34391
rect 9689 34357 9723 34391
rect 11897 34357 11931 34391
rect 14197 34357 14231 34391
rect 20867 34357 20901 34391
rect 21649 34357 21683 34391
rect 26433 34357 26467 34391
rect 27629 34357 27663 34391
rect 28733 34357 28767 34391
rect 29423 34357 29457 34391
rect 37933 34357 37967 34391
rect 38209 34357 38243 34391
rect 38669 34357 38703 34391
rect 40647 34357 40681 34391
rect 6147 34153 6181 34187
rect 7711 34153 7745 34187
rect 8723 34153 8757 34187
rect 12265 34153 12299 34187
rect 13507 34153 13541 34187
rect 17417 34153 17451 34187
rect 18429 34153 18463 34187
rect 22615 34153 22649 34187
rect 23995 34153 24029 34187
rect 24317 34153 24351 34187
rect 25559 34153 25593 34187
rect 26341 34153 26375 34187
rect 30849 34153 30883 34187
rect 32413 34153 32447 34187
rect 32689 34153 32723 34187
rect 32965 34153 32999 34187
rect 34575 34153 34609 34187
rect 38669 34153 38703 34187
rect 39129 34153 39163 34187
rect 39405 34153 39439 34187
rect 41797 34153 41831 34187
rect 8309 34085 8343 34119
rect 9873 34085 9907 34119
rect 11707 34085 11741 34119
rect 15577 34085 15611 34119
rect 19441 34085 19475 34119
rect 21097 34085 21131 34119
rect 21925 34085 21959 34119
rect 26893 34085 26927 34119
rect 29285 34085 29319 34119
rect 36829 34085 36863 34119
rect 38070 34085 38104 34119
rect 40601 34085 40635 34119
rect 41153 34085 41187 34119
rect 43545 34085 43579 34119
rect 4721 34017 4755 34051
rect 4905 34017 4939 34051
rect 6044 34017 6078 34051
rect 7640 34017 7674 34051
rect 8620 34017 8654 34051
rect 13436 34017 13470 34051
rect 16221 34017 16255 34051
rect 17141 34017 17175 34051
rect 17693 34017 17727 34051
rect 21649 34017 21683 34051
rect 22512 34017 22546 34051
rect 23892 34017 23926 34051
rect 25456 34017 25490 34051
rect 28549 34017 28583 34051
rect 29101 34017 29135 34051
rect 32045 34017 32079 34051
rect 33425 34017 33459 34051
rect 34437 34017 34471 34051
rect 36369 34017 36403 34051
rect 36553 34017 36587 34051
rect 42292 34017 42326 34051
rect 4997 33949 5031 33983
rect 9781 33949 9815 33983
rect 10057 33949 10091 33983
rect 11345 33949 11379 33983
rect 19165 33949 19199 33983
rect 19349 33949 19383 33983
rect 21005 33949 21039 33983
rect 26801 33949 26835 33983
rect 27077 33949 27111 33983
rect 30389 33949 30423 33983
rect 37749 33949 37783 33983
rect 40509 33949 40543 33983
rect 42395 33949 42429 33983
rect 43453 33949 43487 33983
rect 43729 33949 43763 33983
rect 19901 33881 19935 33915
rect 4261 33813 4295 33847
rect 7297 33813 7331 33847
rect 12817 33813 12851 33847
rect 13829 33813 13863 33847
rect 23765 33813 23799 33847
rect 29561 33813 29595 33847
rect 33563 33813 33597 33847
rect 42717 33813 42751 33847
rect 5917 33609 5951 33643
rect 6193 33609 6227 33643
rect 7757 33609 7791 33643
rect 8033 33609 8067 33643
rect 9137 33609 9171 33643
rect 10379 33609 10413 33643
rect 11253 33609 11287 33643
rect 14013 33609 14047 33643
rect 15945 33609 15979 33643
rect 16589 33609 16623 33643
rect 17141 33609 17175 33643
rect 19533 33609 19567 33643
rect 19809 33609 19843 33643
rect 20269 33609 20303 33643
rect 20499 33609 20533 33643
rect 21281 33609 21315 33643
rect 22477 33609 22511 33643
rect 24685 33609 24719 33643
rect 25421 33609 25455 33643
rect 28319 33609 28353 33643
rect 29009 33609 29043 33643
rect 30481 33609 30515 33643
rect 31953 33609 31987 33643
rect 33517 33609 33551 33643
rect 34437 33609 34471 33643
rect 37197 33609 37231 33643
rect 37841 33609 37875 33643
rect 38577 33609 38611 33643
rect 39957 33609 39991 33643
rect 40325 33609 40359 33643
rect 41521 33609 41555 33643
rect 42257 33609 42291 33643
rect 9505 33541 9539 33575
rect 9689 33541 9723 33575
rect 22017 33541 22051 33575
rect 27261 33541 27295 33575
rect 28733 33541 28767 33575
rect 4997 33473 5031 33507
rect 13645 33473 13679 33507
rect 21465 33473 21499 33507
rect 22845 33473 22879 33507
rect 25743 33473 25777 33507
rect 26709 33473 26743 33507
rect 27997 33473 28031 33507
rect 30757 33473 30791 33507
rect 31033 33473 31067 33507
rect 3341 33405 3375 33439
rect 3709 33405 3743 33439
rect 3985 33405 4019 33439
rect 4169 33405 4203 33439
rect 6837 33405 6871 33439
rect 9296 33405 9330 33439
rect 10057 33405 10091 33439
rect 10308 33405 10342 33439
rect 11412 33405 11446 33439
rect 12173 33405 12207 33439
rect 12817 33405 12851 33439
rect 13185 33405 13219 33439
rect 13461 33405 13495 33439
rect 14657 33405 14691 33439
rect 15577 33405 15611 33439
rect 16221 33405 16255 33439
rect 16440 33405 16474 33439
rect 18613 33405 18647 33439
rect 20428 33405 20462 33439
rect 23397 33405 23431 33439
rect 23673 33405 23707 33439
rect 24133 33405 24167 33439
rect 25640 33405 25674 33439
rect 26065 33405 26099 33439
rect 28248 33405 28282 33439
rect 29336 33405 29370 33439
rect 4905 33337 4939 33371
rect 5359 33337 5393 33371
rect 6653 33337 6687 33371
rect 7199 33337 7233 33371
rect 10701 33337 10735 33371
rect 11897 33337 11931 33371
rect 14565 33337 14599 33371
rect 15019 33337 15053 33371
rect 17601 33337 17635 33371
rect 18975 33337 19009 33371
rect 21557 33337 21591 33371
rect 26433 33337 26467 33371
rect 26801 33337 26835 33371
rect 29423 33337 29457 33371
rect 30205 33337 30239 33371
rect 30849 33337 30883 33371
rect 31861 33337 31895 33371
rect 41153 33541 41187 33575
rect 32505 33473 32539 33507
rect 32781 33473 32815 33507
rect 35357 33473 35391 33507
rect 36093 33473 36127 33507
rect 36921 33473 36955 33507
rect 38117 33473 38151 33507
rect 38853 33473 38887 33507
rect 39497 33473 39531 33507
rect 40601 33473 40635 33507
rect 41889 33473 41923 33507
rect 42717 33473 42751 33507
rect 42993 33473 43027 33507
rect 44557 33473 44591 33507
rect 34932 33405 34966 33439
rect 36461 33405 36495 33439
rect 36645 33405 36679 33439
rect 32597 33337 32631 33371
rect 38945 33337 38979 33371
rect 40693 33337 40727 33371
rect 42809 33337 42843 33371
rect 43729 33337 43763 33371
rect 44281 33337 44315 33371
rect 44373 33337 44407 33371
rect 4537 33269 4571 33303
rect 8585 33269 8619 33303
rect 11483 33269 11517 33303
rect 18429 33269 18463 33303
rect 20913 33269 20947 33303
rect 23765 33269 23799 33303
rect 27629 33269 27663 33303
rect 29837 33269 29871 33303
rect 31953 33269 31987 33303
rect 32137 33269 32171 33303
rect 35035 33269 35069 33303
rect 44005 33269 44039 33303
rect 4169 33065 4203 33099
rect 5457 33065 5491 33099
rect 7849 33065 7883 33099
rect 8401 33065 8435 33099
rect 10609 33065 10643 33099
rect 12357 33065 12391 33099
rect 13277 33065 13311 33099
rect 14657 33065 14691 33099
rect 18613 33065 18647 33099
rect 19073 33065 19107 33099
rect 20269 33065 20303 33099
rect 23581 33065 23615 33099
rect 27445 33065 27479 33099
rect 33057 33065 33091 33099
rect 43085 33065 43119 33099
rect 44281 33065 44315 33099
rect 10051 32997 10085 33031
rect 11758 32997 11792 33031
rect 15622 32997 15656 33031
rect 17738 32997 17772 33031
rect 19257 32997 19291 33031
rect 19349 32997 19383 33031
rect 30665 32997 30699 33031
rect 31217 32997 31251 33031
rect 32413 32997 32447 33031
rect 34069 32997 34103 33031
rect 35633 32997 35667 33031
rect 36921 32997 36955 33031
rect 39037 32997 39071 33031
rect 40601 32997 40635 33031
rect 42809 32997 42843 33031
rect 43499 32997 43533 33031
rect 4077 32929 4111 32963
rect 4629 32929 4663 32963
rect 6101 32929 6135 32963
rect 6377 32929 6411 32963
rect 6561 32929 6595 32963
rect 6837 32929 6871 32963
rect 13461 32929 13495 32963
rect 13645 32929 13679 32963
rect 16221 32929 16255 32963
rect 21925 32929 21959 32963
rect 22201 32929 22235 32963
rect 25488 32929 25522 32963
rect 26560 32929 26594 32963
rect 27588 32929 27622 32963
rect 29193 32929 29227 32963
rect 29377 32929 29411 32963
rect 37749 32929 37783 32963
rect 43269 32929 43303 32963
rect 7481 32861 7515 32895
rect 9689 32861 9723 32895
rect 11437 32861 11471 32895
rect 15301 32861 15335 32895
rect 17417 32861 17451 32895
rect 19901 32861 19935 32895
rect 22385 32861 22419 32895
rect 23213 32861 23247 32895
rect 27675 32861 27709 32895
rect 29561 32861 29595 32895
rect 30573 32861 30607 32895
rect 32137 32861 32171 32895
rect 33977 32861 34011 32895
rect 34253 32861 34287 32895
rect 35541 32861 35575 32895
rect 35817 32861 35851 32895
rect 38945 32861 38979 32895
rect 40509 32861 40543 32895
rect 42257 32861 42291 32895
rect 18337 32793 18371 32827
rect 26985 32793 27019 32827
rect 36553 32793 36587 32827
rect 37933 32793 37967 32827
rect 39497 32793 39531 32827
rect 41061 32793 41095 32827
rect 3433 32725 3467 32759
rect 5181 32725 5215 32759
rect 13001 32725 13035 32759
rect 17325 32725 17359 32759
rect 21373 32725 21407 32759
rect 24133 32725 24167 32759
rect 25237 32725 25271 32759
rect 25559 32725 25593 32759
rect 26801 32725 26835 32759
rect 28641 32725 28675 32759
rect 29929 32725 29963 32759
rect 42073 32725 42107 32759
rect 43913 32725 43947 32759
rect 3249 32521 3283 32555
rect 5181 32521 5215 32555
rect 5641 32521 5675 32555
rect 7021 32521 7055 32555
rect 8861 32521 8895 32555
rect 15393 32521 15427 32555
rect 17417 32521 17451 32555
rect 19257 32521 19291 32555
rect 22845 32521 22879 32555
rect 26157 32521 26191 32555
rect 26525 32521 26559 32555
rect 29009 32521 29043 32555
rect 29653 32521 29687 32555
rect 30757 32521 30791 32555
rect 33057 32521 33091 32555
rect 34253 32521 34287 32555
rect 34621 32521 34655 32555
rect 36829 32521 36863 32555
rect 38301 32521 38335 32555
rect 39037 32521 39071 32555
rect 39865 32521 39899 32555
rect 40325 32521 40359 32555
rect 10609 32453 10643 32487
rect 21189 32453 21223 32487
rect 24685 32453 24719 32487
rect 27629 32453 27663 32487
rect 28089 32453 28123 32487
rect 35633 32453 35667 32487
rect 39543 32453 39577 32487
rect 44281 32453 44315 32487
rect 4629 32385 4663 32419
rect 7941 32385 7975 32419
rect 14657 32385 14691 32419
rect 16405 32385 16439 32419
rect 17049 32385 17083 32419
rect 17877 32385 17911 32419
rect 18613 32385 18647 32419
rect 19809 32385 19843 32419
rect 21741 32385 21775 32419
rect 23765 32385 23799 32419
rect 24225 32385 24259 32419
rect 27077 32385 27111 32419
rect 29837 32385 29871 32419
rect 32597 32385 32631 32419
rect 33333 32385 33367 32419
rect 33793 32385 33827 32419
rect 40601 32385 40635 32419
rect 41521 32385 41555 32419
rect 42165 32385 42199 32419
rect 42441 32385 42475 32419
rect 43729 32385 43763 32419
rect 44649 32385 44683 32419
rect 3985 32317 4019 32351
rect 4077 32317 4111 32351
rect 4537 32317 4571 32351
rect 5800 32317 5834 32351
rect 6653 32317 6687 32351
rect 6837 32317 6871 32351
rect 9689 32317 9723 32351
rect 12173 32317 12207 32351
rect 12449 32317 12483 32351
rect 13001 32317 13035 32351
rect 14013 32317 14047 32351
rect 14105 32317 14139 32351
rect 14565 32317 14599 32351
rect 15669 32317 15703 32351
rect 16221 32317 16255 32351
rect 16681 32317 16715 32351
rect 18337 32317 18371 32351
rect 18521 32317 18555 32351
rect 25237 32317 25271 32351
rect 31493 32317 31527 32351
rect 31861 32317 31895 32351
rect 32045 32317 32079 32351
rect 35817 32317 35851 32351
rect 36369 32317 36403 32351
rect 36553 32317 36587 32351
rect 37381 32317 37415 32351
rect 39472 32317 39506 32351
rect 7481 32249 7515 32283
rect 7849 32249 7883 32283
rect 8303 32249 8337 32283
rect 9229 32249 9263 32283
rect 9597 32249 9631 32283
rect 10010 32249 10044 32283
rect 11437 32249 11471 32283
rect 11897 32249 11931 32283
rect 19901 32249 19935 32283
rect 20453 32249 20487 32283
rect 20821 32249 20855 32283
rect 21373 32249 21407 32283
rect 21465 32249 21499 32283
rect 23857 32249 23891 32283
rect 25053 32249 25087 32283
rect 25558 32249 25592 32283
rect 27169 32249 27203 32283
rect 30158 32249 30192 32283
rect 31033 32249 31067 32283
rect 32321 32249 32355 32283
rect 33425 32249 33459 32283
rect 35357 32249 35391 32283
rect 37743 32249 37777 32283
rect 40693 32249 40727 32283
rect 41245 32249 41279 32283
rect 42257 32249 42291 32283
rect 43821 32249 43855 32283
rect 3525 32181 3559 32215
rect 5871 32181 5905 32215
rect 6285 32181 6319 32215
rect 10885 32181 10919 32215
rect 12541 32181 12575 32215
rect 13461 32181 13495 32215
rect 19625 32181 19659 32215
rect 22385 32181 22419 32215
rect 23213 32181 23247 32215
rect 28641 32181 28675 32215
rect 37289 32181 37323 32215
rect 38669 32181 38703 32215
rect 41889 32181 41923 32215
rect 43361 32181 43395 32215
rect 9505 31977 9539 32011
rect 9781 31977 9815 32011
rect 11437 31977 11471 32011
rect 14197 31977 14231 32011
rect 15669 31977 15703 32011
rect 17325 31977 17359 32011
rect 22109 31977 22143 32011
rect 23029 31977 23063 32011
rect 23949 31977 23983 32011
rect 27537 31977 27571 32011
rect 29929 31977 29963 32011
rect 30481 31977 30515 32011
rect 30757 31977 30791 32011
rect 32321 31977 32355 32011
rect 33011 31977 33045 32011
rect 33793 31977 33827 32011
rect 37381 31977 37415 32011
rect 38669 31977 38703 32011
rect 40693 31977 40727 32011
rect 42441 31977 42475 32011
rect 4813 31909 4847 31943
rect 8723 31909 8757 31943
rect 19441 31909 19475 31943
rect 21695 31909 21729 31943
rect 24593 31909 24627 31943
rect 26709 31909 26743 31943
rect 27261 31909 27295 31943
rect 33425 31909 33459 31943
rect 34069 31909 34103 31943
rect 38111 31909 38145 31943
rect 38945 31909 38979 31943
rect 39818 31909 39852 31943
rect 41842 31909 41876 31943
rect 43545 31909 43579 31943
rect 4077 31841 4111 31875
rect 4537 31841 4571 31875
rect 5708 31841 5742 31875
rect 6929 31841 6963 31875
rect 7389 31841 7423 31875
rect 8620 31841 8654 31875
rect 9689 31841 9723 31875
rect 10149 31841 10183 31875
rect 11437 31841 11471 31875
rect 11897 31841 11931 31875
rect 13461 31841 13495 31875
rect 16104 31841 16138 31875
rect 17325 31841 17359 31875
rect 17601 31841 17635 31875
rect 21465 31841 21499 31875
rect 23581 31841 23615 31875
rect 29561 31841 29595 31875
rect 32908 31841 32942 31875
rect 35541 31841 35575 31875
rect 36093 31841 36127 31875
rect 36277 31841 36311 31875
rect 40417 31841 40451 31875
rect 7481 31773 7515 31807
rect 7941 31773 7975 31807
rect 19349 31773 19383 31807
rect 19625 31773 19659 31807
rect 22661 31773 22695 31807
rect 24501 31773 24535 31807
rect 24777 31773 24811 31807
rect 26617 31773 26651 31807
rect 28089 31773 28123 31807
rect 33977 31773 34011 31807
rect 34253 31773 34287 31807
rect 37749 31773 37783 31807
rect 39497 31773 39531 31807
rect 41521 31773 41555 31807
rect 43453 31773 43487 31807
rect 43729 31773 43763 31807
rect 5779 31705 5813 31739
rect 16175 31705 16209 31739
rect 41153 31705 41187 31739
rect 5457 31637 5491 31671
rect 6193 31637 6227 31671
rect 8309 31637 8343 31671
rect 12449 31637 12483 31671
rect 13185 31637 13219 31671
rect 13645 31637 13679 31671
rect 18061 31637 18095 31671
rect 18981 31637 19015 31671
rect 21373 31637 21407 31671
rect 25513 31637 25547 31671
rect 29377 31637 29411 31671
rect 31585 31637 31619 31671
rect 35357 31637 35391 31671
rect 4905 31433 4939 31467
rect 16497 31433 16531 31467
rect 18521 31433 18555 31467
rect 19901 31433 19935 31467
rect 21557 31433 21591 31467
rect 25329 31433 25363 31467
rect 25973 31433 26007 31467
rect 27813 31433 27847 31467
rect 30297 31433 30331 31467
rect 32873 31433 32907 31467
rect 33747 31433 33781 31467
rect 34161 31433 34195 31467
rect 36001 31433 36035 31467
rect 36369 31433 36403 31467
rect 38669 31433 38703 31467
rect 39405 31433 39439 31467
rect 40785 31433 40819 31467
rect 41889 31433 41923 31467
rect 42395 31433 42429 31467
rect 43177 31433 43211 31467
rect 43729 31433 43763 31467
rect 44097 31433 44131 31467
rect 14657 31365 14691 31399
rect 18797 31365 18831 31399
rect 20269 31365 20303 31399
rect 32505 31365 32539 31399
rect 39681 31365 39715 31399
rect 41521 31365 41555 31399
rect 6653 31297 6687 31331
rect 13461 31297 13495 31331
rect 22661 31297 22695 31331
rect 23305 31297 23339 31331
rect 25053 31297 25087 31331
rect 26709 31297 26743 31331
rect 26893 31297 26927 31331
rect 27169 31297 27203 31331
rect 29929 31297 29963 31331
rect 31953 31297 31987 31331
rect 37197 31297 37231 31331
rect 37841 31297 37875 31331
rect 43407 31297 43441 31331
rect 4512 31229 4546 31263
rect 5492 31229 5526 31263
rect 10701 31229 10735 31263
rect 10793 31229 10827 31263
rect 11253 31229 11287 31263
rect 14473 31229 14507 31263
rect 14933 31229 14967 31263
rect 15393 31229 15427 31263
rect 15577 31229 15611 31263
rect 18981 31229 19015 31263
rect 20729 31229 20763 31263
rect 21925 31229 21959 31263
rect 22385 31229 22419 31263
rect 24041 31229 24075 31263
rect 24317 31229 24351 31263
rect 24777 31229 24811 31263
rect 29101 31229 29135 31263
rect 29469 31229 29503 31263
rect 29837 31229 29871 31263
rect 30849 31229 30883 31263
rect 31309 31229 31343 31263
rect 33676 31229 33710 31263
rect 35173 31229 35207 31263
rect 35357 31229 35391 31263
rect 36461 31229 36495 31263
rect 36921 31229 36955 31263
rect 38209 31229 38243 31263
rect 39221 31229 39255 31263
rect 40049 31229 40083 31263
rect 40576 31229 40610 31263
rect 42324 31229 42358 31263
rect 43320 31229 43354 31263
rect 5595 31161 5629 31195
rect 6929 31161 6963 31195
rect 7021 31161 7055 31195
rect 7573 31161 7607 31195
rect 8861 31161 8895 31195
rect 8953 31161 8987 31195
rect 9505 31161 9539 31195
rect 12541 31161 12575 31195
rect 12633 31161 12667 31195
rect 13185 31161 13219 31195
rect 15485 31161 15519 31195
rect 17141 31161 17175 31195
rect 19302 31161 19336 31195
rect 26985 31161 27019 31195
rect 32045 31161 32079 31195
rect 34713 31161 34747 31195
rect 35633 31161 35667 31195
rect 39037 31161 39071 31195
rect 4077 31093 4111 31127
rect 4583 31093 4617 31127
rect 5365 31093 5399 31127
rect 6285 31093 6319 31127
rect 7849 31093 7883 31127
rect 8309 31093 8343 31127
rect 8677 31093 8711 31127
rect 9781 31093 9815 31127
rect 10149 31093 10183 31127
rect 10885 31093 10919 31127
rect 11805 31093 11839 31127
rect 12265 31093 12299 31127
rect 17509 31093 17543 31127
rect 20913 31093 20947 31127
rect 21281 31093 21315 31127
rect 22937 31093 22971 31127
rect 24041 31093 24075 31127
rect 24133 31093 24167 31127
rect 26341 31093 26375 31127
rect 31033 31093 31067 31127
rect 31677 31093 31711 31127
rect 33517 31093 33551 31127
rect 38347 31093 38381 31127
rect 41061 31093 41095 31127
rect 42717 31093 42751 31127
rect 4629 30889 4663 30923
rect 5181 30889 5215 30923
rect 5733 30889 5767 30923
rect 6929 30889 6963 30923
rect 8861 30889 8895 30923
rect 10103 30889 10137 30923
rect 12541 30889 12575 30923
rect 19257 30889 19291 30923
rect 25053 30889 25087 30923
rect 29561 30889 29595 30923
rect 31953 30889 31987 30923
rect 33425 30889 33459 30923
rect 34989 30889 35023 30923
rect 36461 30889 36495 30923
rect 38301 30889 38335 30923
rect 6330 30821 6364 30855
rect 7849 30821 7883 30855
rect 7941 30821 7975 30855
rect 11253 30821 11287 30855
rect 12265 30821 12299 30855
rect 23857 30821 23891 30855
rect 26709 30821 26743 30855
rect 27261 30821 27295 30855
rect 32413 30821 32447 30855
rect 32965 30821 32999 30855
rect 34069 30821 34103 30855
rect 35265 30821 35299 30855
rect 35633 30821 35667 30855
rect 7573 30753 7607 30787
rect 10032 30753 10066 30787
rect 11897 30753 11931 30787
rect 13277 30753 13311 30787
rect 13737 30753 13771 30787
rect 15485 30753 15519 30787
rect 17141 30753 17175 30787
rect 19809 30753 19843 30787
rect 20913 30753 20947 30787
rect 22636 30753 22670 30787
rect 25456 30753 25490 30787
rect 28917 30753 28951 30787
rect 30205 30753 30239 30787
rect 30481 30753 30515 30787
rect 37749 30753 37783 30787
rect 38761 30753 38795 30787
rect 39773 30753 39807 30787
rect 41153 30753 41187 30787
rect 4261 30685 4295 30719
rect 6009 30685 6043 30719
rect 8125 30685 8159 30719
rect 10977 30685 11011 30719
rect 13829 30685 13863 30719
rect 15393 30685 15427 30719
rect 16957 30685 16991 30719
rect 18889 30685 18923 30719
rect 23765 30685 23799 30719
rect 24133 30685 24167 30719
rect 26617 30685 26651 30719
rect 30665 30685 30699 30719
rect 30941 30685 30975 30719
rect 32321 30685 32355 30719
rect 33793 30685 33827 30719
rect 33977 30685 34011 30719
rect 34253 30685 34287 30719
rect 35541 30685 35575 30719
rect 35817 30685 35851 30719
rect 21925 30617 21959 30651
rect 25559 30617 25593 30651
rect 26249 30617 26283 30651
rect 29101 30617 29135 30651
rect 39957 30617 39991 30651
rect 7205 30549 7239 30583
rect 10793 30549 10827 30583
rect 18337 30549 18371 30583
rect 21097 30549 21131 30583
rect 22707 30549 22741 30583
rect 24685 30549 24719 30583
rect 37933 30549 37967 30583
rect 38945 30549 38979 30583
rect 39221 30549 39255 30583
rect 40969 30549 41003 30583
rect 41291 30549 41325 30583
rect 6377 30345 6411 30379
rect 10057 30345 10091 30379
rect 11529 30345 11563 30379
rect 15485 30345 15519 30379
rect 19349 30345 19383 30379
rect 20269 30345 20303 30379
rect 21373 30345 21407 30379
rect 23029 30345 23063 30379
rect 23489 30345 23523 30379
rect 24869 30345 24903 30379
rect 28457 30345 28491 30379
rect 30481 30345 30515 30379
rect 31585 30345 31619 30379
rect 32229 30345 32263 30379
rect 33977 30345 34011 30379
rect 36461 30345 36495 30379
rect 40785 30345 40819 30379
rect 13093 30277 13127 30311
rect 26249 30277 26283 30311
rect 27077 30277 27111 30311
rect 29469 30277 29503 30311
rect 30205 30277 30239 30311
rect 7481 30209 7515 30243
rect 8125 30209 8159 30243
rect 9045 30209 9079 30243
rect 10609 30209 10643 30243
rect 13645 30209 13679 30243
rect 17877 30209 17911 30243
rect 19073 30209 19107 30243
rect 19717 30209 19751 30243
rect 22477 30209 22511 30243
rect 24133 30209 24167 30243
rect 26525 30209 26559 30243
rect 28135 30209 28169 30243
rect 30665 30209 30699 30243
rect 32781 30209 32815 30243
rect 35725 30209 35759 30243
rect 40969 30209 41003 30243
rect 3249 30141 3283 30175
rect 3709 30141 3743 30175
rect 4721 30141 4755 30175
rect 5089 30141 5123 30175
rect 5273 30141 5307 30175
rect 12265 30141 12299 30175
rect 12700 30141 12734 30175
rect 14565 30141 14599 30175
rect 15117 30141 15151 30175
rect 15761 30141 15795 30175
rect 18337 30141 18371 30175
rect 18797 30141 18831 30175
rect 20453 30141 20487 30175
rect 22636 30141 22670 30175
rect 25488 30141 25522 30175
rect 28048 30141 28082 30175
rect 29285 30141 29319 30175
rect 32597 30141 32631 30175
rect 3985 30073 4019 30107
rect 6009 30073 6043 30107
rect 7297 30073 7331 30107
rect 7573 30073 7607 30107
rect 8861 30073 8895 30107
rect 9137 30073 9171 30107
rect 9689 30073 9723 30107
rect 10517 30073 10551 30107
rect 10971 30073 11005 30107
rect 11897 30073 11931 30107
rect 13553 30073 13587 30107
rect 13966 30073 14000 30107
rect 15669 30073 15703 30107
rect 20775 30073 20809 30107
rect 23857 30073 23891 30107
rect 23949 30073 23983 30107
rect 26617 30073 26651 30107
rect 29745 30073 29779 30107
rect 30986 30073 31020 30107
rect 33057 30141 33091 30175
rect 34713 30141 34747 30175
rect 35265 30141 35299 30175
rect 35541 30141 35575 30175
rect 36553 30141 36587 30175
rect 37105 30141 37139 30175
rect 38184 30141 38218 30175
rect 38577 30141 38611 30175
rect 39129 30141 39163 30175
rect 42752 30141 42786 30175
rect 43177 30141 43211 30175
rect 33419 30073 33453 30107
rect 34345 30073 34379 30107
rect 37289 30073 37323 30107
rect 41290 30073 41324 30107
rect 3065 30005 3099 30039
rect 4353 30005 4387 30039
rect 4905 30005 4939 30039
rect 8493 30005 8527 30039
rect 12771 30005 12805 30039
rect 17049 30005 17083 30039
rect 21741 30005 21775 30039
rect 22707 30005 22741 30039
rect 25559 30005 25593 30039
rect 25973 30005 26007 30039
rect 27445 30005 27479 30039
rect 27905 30005 27939 30039
rect 29009 30005 29043 30039
rect 32781 30005 32815 30039
rect 32873 30005 32907 30039
rect 36001 30005 36035 30039
rect 37749 30005 37783 30039
rect 38255 30005 38289 30039
rect 38945 30005 38979 30039
rect 39313 30005 39347 30039
rect 39773 30005 39807 30039
rect 41889 30005 41923 30039
rect 42855 30005 42889 30039
rect 3893 29801 3927 29835
rect 5273 29801 5307 29835
rect 6101 29801 6135 29835
rect 8401 29801 8435 29835
rect 9045 29801 9079 29835
rect 10701 29801 10735 29835
rect 11069 29801 11103 29835
rect 11805 29801 11839 29835
rect 13829 29801 13863 29835
rect 18337 29801 18371 29835
rect 23489 29801 23523 29835
rect 26341 29801 26375 29835
rect 31953 29801 31987 29835
rect 34161 29801 34195 29835
rect 34621 29801 34655 29835
rect 34897 29801 34931 29835
rect 41429 29801 41463 29835
rect 42533 29801 42567 29835
rect 4439 29733 4473 29767
rect 7573 29733 7607 29767
rect 8125 29733 8159 29767
rect 12550 29733 12584 29767
rect 13093 29733 13127 29767
rect 15485 29733 15519 29767
rect 17049 29733 17083 29767
rect 22890 29733 22924 29767
rect 24638 29733 24672 29767
rect 26617 29733 26651 29767
rect 26709 29733 26743 29767
rect 30021 29733 30055 29767
rect 32873 29733 32907 29767
rect 33839 29733 33873 29767
rect 35633 29733 35667 29767
rect 36001 29733 36035 29767
rect 38990 29733 39024 29767
rect 40601 29733 40635 29767
rect 43545 29733 43579 29767
rect 5825 29665 5859 29699
rect 6285 29665 6319 29699
rect 9848 29665 9882 29699
rect 10793 29665 10827 29699
rect 11345 29665 11379 29699
rect 13988 29665 14022 29699
rect 14381 29665 14415 29699
rect 18705 29665 18739 29699
rect 18889 29665 18923 29699
rect 21097 29665 21131 29699
rect 21557 29665 21591 29699
rect 23857 29665 23891 29699
rect 25237 29665 25271 29699
rect 28181 29665 28215 29699
rect 28641 29665 28675 29699
rect 30573 29665 30607 29699
rect 30941 29665 30975 29699
rect 32137 29665 32171 29699
rect 32689 29665 32723 29699
rect 33736 29665 33770 29699
rect 34713 29665 34747 29699
rect 35173 29665 35207 29699
rect 36093 29665 36127 29699
rect 36645 29665 36679 29699
rect 42016 29665 42050 29699
rect 4077 29597 4111 29631
rect 7481 29597 7515 29631
rect 12449 29597 12483 29631
rect 15393 29597 15427 29631
rect 16037 29597 16071 29631
rect 16957 29597 16991 29631
rect 17601 29597 17635 29631
rect 18981 29597 19015 29631
rect 21741 29597 21775 29631
rect 22569 29597 22603 29631
rect 24317 29597 24351 29631
rect 28917 29597 28951 29631
rect 31217 29597 31251 29631
rect 36829 29597 36863 29631
rect 38669 29597 38703 29631
rect 40509 29597 40543 29631
rect 41153 29597 41187 29631
rect 42119 29597 42153 29631
rect 43453 29597 43487 29631
rect 43729 29597 43763 29631
rect 14059 29529 14093 29563
rect 24225 29529 24259 29563
rect 27169 29529 27203 29563
rect 3249 29461 3283 29495
rect 4997 29461 5031 29495
rect 6929 29461 6963 29495
rect 9919 29461 9953 29495
rect 13369 29461 13403 29495
rect 19993 29461 20027 29495
rect 20453 29461 20487 29495
rect 25513 29461 25547 29495
rect 39589 29461 39623 29495
rect 40325 29461 40359 29495
rect 5181 29257 5215 29291
rect 8217 29257 8251 29291
rect 10793 29257 10827 29291
rect 13737 29257 13771 29291
rect 15393 29257 15427 29291
rect 17877 29257 17911 29291
rect 21465 29257 21499 29291
rect 23121 29257 23155 29291
rect 23397 29257 23431 29291
rect 23949 29257 23983 29291
rect 24593 29257 24627 29291
rect 24869 29257 24903 29291
rect 25237 29257 25271 29291
rect 26341 29257 26375 29291
rect 26709 29257 26743 29291
rect 28089 29257 28123 29291
rect 30205 29257 30239 29291
rect 32137 29257 32171 29291
rect 32505 29257 32539 29291
rect 32781 29257 32815 29291
rect 33747 29257 33781 29291
rect 37565 29257 37599 29291
rect 40233 29257 40267 29291
rect 41613 29257 41647 29291
rect 43453 29257 43487 29291
rect 12265 29189 12299 29223
rect 39681 29189 39715 29223
rect 3433 29121 3467 29155
rect 7205 29121 7239 29155
rect 9781 29121 9815 29155
rect 12817 29121 12851 29155
rect 14381 29121 14415 29155
rect 14657 29121 14691 29155
rect 15669 29121 15703 29155
rect 20453 29121 20487 29155
rect 22753 29121 22787 29155
rect 25421 29121 25455 29155
rect 31217 29121 31251 29155
rect 37197 29121 37231 29155
rect 38117 29121 38151 29155
rect 40601 29121 40635 29155
rect 42165 29121 42199 29155
rect 42441 29121 42475 29155
rect 43729 29121 43763 29155
rect 2605 29053 2639 29087
rect 2973 29053 3007 29087
rect 3249 29053 3283 29087
rect 4261 29053 4295 29087
rect 5457 29053 5491 29087
rect 11012 29053 11046 29087
rect 11805 29053 11839 29087
rect 18889 29053 18923 29087
rect 19809 29053 19843 29087
rect 20177 29053 20211 29087
rect 20361 29053 20395 29087
rect 22017 29053 22051 29087
rect 22477 29053 22511 29087
rect 24409 29053 24443 29087
rect 27169 29053 27203 29087
rect 29285 29053 29319 29087
rect 29745 29053 29779 29087
rect 33676 29053 33710 29087
rect 35265 29053 35299 29087
rect 35541 29053 35575 29087
rect 36829 29053 36863 29087
rect 37105 29053 37139 29087
rect 39037 29053 39071 29087
rect 6929 28985 6963 29019
rect 7021 28985 7055 29019
rect 9137 28985 9171 29019
rect 9229 28985 9263 29019
rect 12541 28985 12575 29019
rect 12633 28985 12667 29019
rect 14197 28985 14231 29019
rect 14473 28985 14507 29019
rect 16497 28985 16531 29019
rect 16589 28985 16623 29019
rect 17141 28985 17175 29019
rect 17509 28985 17543 29019
rect 18245 28985 18279 29019
rect 25742 28985 25776 29019
rect 26985 28985 27019 29019
rect 27490 28985 27524 29019
rect 28733 28985 28767 29019
rect 30573 28985 30607 29019
rect 31538 28985 31572 29019
rect 34437 28985 34471 29019
rect 35725 28985 35759 29019
rect 36093 28985 36127 29019
rect 38479 28963 38513 28997
rect 40693 28985 40727 29019
rect 41245 28985 41279 29019
rect 42257 28985 42291 29019
rect 3801 28917 3835 28951
rect 4077 28917 4111 28951
rect 4629 28917 4663 28951
rect 5825 28917 5859 28951
rect 6193 28917 6227 28951
rect 6653 28917 6687 28951
rect 7941 28917 7975 28951
rect 8953 28917 8987 28951
rect 10149 28917 10183 28951
rect 11115 28917 11149 28951
rect 11437 28917 11471 28951
rect 16313 28917 16347 28951
rect 19349 28917 19383 28951
rect 21097 28917 21131 28951
rect 21833 28917 21867 28951
rect 24317 28917 24351 28951
rect 28365 28917 28399 28951
rect 29469 28917 29503 28951
rect 31125 28917 31159 28951
rect 34161 28917 34195 28951
rect 38025 28917 38059 28951
rect 39313 28917 39347 28951
rect 41889 28917 41923 28951
rect 4491 28713 4525 28747
rect 12449 28713 12483 28747
rect 17693 28713 17727 28747
rect 22109 28713 22143 28747
rect 26249 28713 26283 28747
rect 31493 28713 31527 28747
rect 34989 28713 35023 28747
rect 36921 28713 36955 28747
rect 38117 28713 38151 28747
rect 39313 28713 39347 28747
rect 41153 28713 41187 28747
rect 5503 28645 5537 28679
rect 6561 28645 6595 28679
rect 7113 28645 7147 28679
rect 9045 28645 9079 28679
rect 9873 28645 9907 28679
rect 11529 28645 11563 28679
rect 11621 28645 11655 28679
rect 13185 28645 13219 28679
rect 13829 28645 13863 28679
rect 14381 28645 14415 28679
rect 16405 28645 16439 28679
rect 16865 28645 16899 28679
rect 19993 28645 20027 28679
rect 25605 28645 25639 28679
rect 27169 28645 27203 28679
rect 29647 28645 29681 28679
rect 33425 28645 33459 28679
rect 35265 28645 35299 28679
rect 38714 28645 38748 28679
rect 40049 28645 40083 28679
rect 40325 28645 40359 28679
rect 41797 28645 41831 28679
rect 41889 28645 41923 28679
rect 4420 28577 4454 28611
rect 5400 28577 5434 28611
rect 7976 28577 8010 28611
rect 12817 28577 12851 28611
rect 15336 28577 15370 28611
rect 18245 28577 18279 28611
rect 19257 28577 19291 28611
rect 19809 28577 19843 28611
rect 20913 28577 20947 28611
rect 21465 28577 21499 28611
rect 22477 28577 22511 28611
rect 23029 28577 23063 28611
rect 25145 28577 25179 28611
rect 25421 28577 25455 28611
rect 26592 28577 26626 28611
rect 27997 28577 28031 28611
rect 28273 28577 28307 28611
rect 31033 28577 31067 28611
rect 32296 28577 32330 28611
rect 34805 28577 34839 28611
rect 35909 28577 35943 28611
rect 36369 28577 36403 28611
rect 38393 28577 38427 28611
rect 4813 28509 4847 28543
rect 6469 28509 6503 28543
rect 9781 28509 9815 28543
rect 10425 28509 10459 28543
rect 12173 28509 12207 28543
rect 13737 28509 13771 28543
rect 16773 28509 16807 28543
rect 17233 28509 17267 28543
rect 21557 28509 21591 28543
rect 23213 28509 23247 28543
rect 28457 28509 28491 28543
rect 29285 28509 29319 28543
rect 33333 28509 33367 28543
rect 33701 28509 33735 28543
rect 36461 28509 36495 28543
rect 40233 28509 40267 28543
rect 42441 28509 42475 28543
rect 32367 28441 32401 28475
rect 40785 28441 40819 28475
rect 2789 28373 2823 28407
rect 8079 28373 8113 28407
rect 8401 28373 8435 28407
rect 15439 28373 15473 28407
rect 15853 28373 15887 28407
rect 18383 28373 18417 28407
rect 26663 28373 26697 28407
rect 27629 28373 27663 28407
rect 30205 28373 30239 28407
rect 30481 28373 30515 28407
rect 31217 28373 31251 28407
rect 32689 28373 32723 28407
rect 5181 28169 5215 28203
rect 6377 28169 6411 28203
rect 7665 28169 7699 28203
rect 9321 28169 9355 28203
rect 10241 28169 10275 28203
rect 12173 28169 12207 28203
rect 13737 28169 13771 28203
rect 14013 28169 14047 28203
rect 14381 28169 14415 28203
rect 15301 28169 15335 28203
rect 16773 28169 16807 28203
rect 17141 28169 17175 28203
rect 17877 28169 17911 28203
rect 26755 28169 26789 28203
rect 27169 28169 27203 28203
rect 27537 28169 27571 28203
rect 31861 28169 31895 28203
rect 33885 28169 33919 28203
rect 35035 28169 35069 28203
rect 35725 28169 35759 28203
rect 38853 28169 38887 28203
rect 40141 28169 40175 28203
rect 42809 28169 42843 28203
rect 5503 28101 5537 28135
rect 8769 28101 8803 28135
rect 11805 28101 11839 28135
rect 17509 28101 17543 28135
rect 21189 28101 21223 28135
rect 21557 28101 21591 28135
rect 23121 28101 23155 28135
rect 24685 28101 24719 28135
rect 25881 28101 25915 28135
rect 34621 28101 34655 28135
rect 35449 28101 35483 28135
rect 4077 28033 4111 28067
rect 8217 28033 8251 28067
rect 10885 28033 10919 28067
rect 16129 28033 16163 28067
rect 18153 28033 18187 28067
rect 22109 28033 22143 28067
rect 22753 28033 22787 28067
rect 25513 28033 25547 28067
rect 29653 28033 29687 28067
rect 36277 28033 36311 28067
rect 41889 28033 41923 28067
rect 3433 27965 3467 27999
rect 3801 27965 3835 27999
rect 3985 27965 4019 27999
rect 5432 27965 5466 27999
rect 5825 27965 5859 27999
rect 7180 27965 7214 27999
rect 9781 27965 9815 27999
rect 12817 27965 12851 27999
rect 16957 27965 16991 27999
rect 18245 27965 18279 27999
rect 20085 27965 20119 27999
rect 20637 27965 20671 27999
rect 20821 27965 20855 27999
rect 23832 27965 23866 27999
rect 25053 27965 25087 27999
rect 25329 27965 25363 27999
rect 26525 27965 26559 27999
rect 26652 27965 26686 27999
rect 27813 27965 27847 27999
rect 28181 27965 28215 27999
rect 28365 27965 28399 27999
rect 32321 27965 32355 27999
rect 34964 27965 34998 27999
rect 37197 27965 37231 27999
rect 39288 27965 39322 27999
rect 40544 27965 40578 27999
rect 40969 27965 41003 27999
rect 43412 27965 43446 27999
rect 8033 27897 8067 27931
rect 8309 27897 8343 27931
rect 10701 27897 10735 27931
rect 10977 27897 11011 27931
rect 11529 27897 11563 27931
rect 12725 27897 12759 27931
rect 13138 27897 13172 27931
rect 15485 27897 15519 27931
rect 15577 27897 15611 27931
rect 19901 27897 19935 27931
rect 21833 27897 21867 27931
rect 21925 27897 21959 27931
rect 28641 27897 28675 27931
rect 29101 27897 29135 27931
rect 29561 27897 29595 27931
rect 30015 27897 30049 27931
rect 32229 27897 32263 27931
rect 32683 27897 32717 27931
rect 36598 27897 36632 27931
rect 38485 27897 38519 27931
rect 40647 27897 40681 27931
rect 41981 27897 42015 27931
rect 42533 27897 42567 27931
rect 43269 27897 43303 27931
rect 43499 27897 43533 27931
rect 4629 27829 4663 27863
rect 7251 27829 7285 27863
rect 9689 27829 9723 27863
rect 9965 27829 9999 27863
rect 14933 27829 14967 27863
rect 19257 27829 19291 27863
rect 23903 27829 23937 27863
rect 24317 27829 24351 27863
rect 30573 27829 30607 27863
rect 31033 27829 31067 27863
rect 33241 27829 33275 27863
rect 33609 27829 33643 27863
rect 36185 27829 36219 27863
rect 38025 27829 38059 27863
rect 39359 27829 39393 27863
rect 39681 27829 39715 27863
rect 41613 27829 41647 27863
rect 43913 27829 43947 27863
rect 4997 27625 5031 27659
rect 6929 27625 6963 27659
rect 9781 27625 9815 27659
rect 10885 27625 10919 27659
rect 16681 27625 16715 27659
rect 18245 27625 18279 27659
rect 19349 27625 19383 27659
rect 20361 27625 20395 27659
rect 21281 27625 21315 27659
rect 21833 27625 21867 27659
rect 22109 27625 22143 27659
rect 23673 27625 23707 27659
rect 25053 27625 25087 27659
rect 25421 27625 25455 27659
rect 27721 27625 27755 27659
rect 29193 27625 29227 27659
rect 29745 27625 29779 27659
rect 36277 27625 36311 27659
rect 36645 27625 36679 27659
rect 41613 27625 41647 27659
rect 4439 27557 4473 27591
rect 8125 27557 8159 27591
rect 8217 27557 8251 27591
rect 8769 27557 8803 27591
rect 12909 27557 12943 27591
rect 13185 27557 13219 27591
rect 15393 27557 15427 27591
rect 15485 27557 15519 27591
rect 17049 27557 17083 27591
rect 17601 27557 17635 27591
rect 24133 27557 24167 27591
rect 32321 27557 32355 27591
rect 33885 27557 33919 27591
rect 38209 27557 38243 27591
rect 38301 27557 38335 27591
rect 39773 27557 39807 27591
rect 39865 27557 39899 27591
rect 41889 27557 41923 27591
rect 42441 27557 42475 27591
rect 4077 27489 4111 27523
rect 5917 27489 5951 27523
rect 6469 27489 6503 27523
rect 9873 27489 9907 27523
rect 10149 27489 10183 27523
rect 12265 27489 12299 27523
rect 12725 27489 12759 27523
rect 13737 27489 13771 27523
rect 18588 27489 18622 27523
rect 19809 27489 19843 27523
rect 26560 27489 26594 27523
rect 27997 27489 28031 27523
rect 28273 27489 28307 27523
rect 35357 27489 35391 27523
rect 35817 27489 35851 27523
rect 43428 27489 43462 27523
rect 6653 27421 6687 27455
rect 7665 27421 7699 27455
rect 16037 27421 16071 27455
rect 16957 27421 16991 27455
rect 20913 27421 20947 27455
rect 22937 27421 22971 27455
rect 24041 27421 24075 27455
rect 24317 27421 24351 27455
rect 28549 27421 28583 27455
rect 29377 27421 29411 27455
rect 32229 27421 32263 27455
rect 32505 27421 32539 27455
rect 33793 27421 33827 27455
rect 34437 27421 34471 27455
rect 35909 27421 35943 27455
rect 38577 27421 38611 27455
rect 40049 27421 40083 27455
rect 41797 27421 41831 27455
rect 19947 27353 19981 27387
rect 40785 27353 40819 27387
rect 3617 27285 3651 27319
rect 7389 27285 7423 27319
rect 13921 27285 13955 27319
rect 14197 27285 14231 27319
rect 18659 27285 18693 27319
rect 22477 27285 22511 27319
rect 26663 27285 26697 27319
rect 30297 27285 30331 27319
rect 30849 27285 30883 27319
rect 39129 27285 39163 27319
rect 43499 27285 43533 27319
rect 5181 27081 5215 27115
rect 5641 27081 5675 27115
rect 7757 27081 7791 27115
rect 8401 27081 8435 27115
rect 10793 27081 10827 27115
rect 12173 27081 12207 27115
rect 14105 27081 14139 27115
rect 15761 27081 15795 27115
rect 17417 27081 17451 27115
rect 19073 27081 19107 27115
rect 24593 27081 24627 27115
rect 27813 27081 27847 27115
rect 29009 27081 29043 27115
rect 29745 27081 29779 27115
rect 30573 27081 30607 27115
rect 32137 27081 32171 27115
rect 33425 27081 33459 27115
rect 36277 27081 36311 27115
rect 38117 27081 38151 27115
rect 40049 27081 40083 27115
rect 43177 27081 43211 27115
rect 43821 27081 43855 27115
rect 8125 27013 8159 27047
rect 16773 27013 16807 27047
rect 20453 27013 20487 27047
rect 29423 27013 29457 27047
rect 31769 27013 31803 27047
rect 41521 27013 41555 27047
rect 42349 27013 42383 27047
rect 3801 26945 3835 26979
rect 6837 26945 6871 26979
rect 9873 26945 9907 26979
rect 11437 26945 11471 26979
rect 12817 26945 12851 26979
rect 14197 26945 14231 26979
rect 15485 26945 15519 26979
rect 18153 26945 18187 26979
rect 18429 26945 18463 26979
rect 21557 26945 21591 26979
rect 23673 26945 23707 26979
rect 26893 26945 26927 26979
rect 27353 26945 27387 26979
rect 30849 26945 30883 26979
rect 31125 26945 31159 26979
rect 32413 26945 32447 26979
rect 32781 26945 32815 26979
rect 34345 26945 34379 26979
rect 36737 26945 36771 26979
rect 38577 26945 38611 26979
rect 40601 26945 40635 26979
rect 41797 26945 41831 26979
rect 43407 26945 43441 26979
rect 3433 26877 3467 26911
rect 4261 26877 4295 26911
rect 8585 26877 8619 26911
rect 9045 26877 9079 26911
rect 11069 26877 11103 26911
rect 11897 26877 11931 26911
rect 15117 26877 15151 26911
rect 15980 26877 16014 26911
rect 16405 26877 16439 26911
rect 16992 26877 17026 26911
rect 20612 26877 20646 26911
rect 26249 26877 26283 26911
rect 26617 26877 26651 26911
rect 26801 26877 26835 26911
rect 27940 26877 27974 26911
rect 28365 26877 28399 26911
rect 29352 26877 29386 26911
rect 34713 26877 34747 26911
rect 35449 26877 35483 26911
rect 35725 26877 35759 26911
rect 41153 26877 41187 26911
rect 43320 26877 43354 26911
rect 44097 26877 44131 26911
rect 4169 26809 4203 26843
rect 4623 26809 4657 26843
rect 6653 26809 6687 26843
rect 7199 26809 7233 26843
rect 9781 26809 9815 26843
rect 10235 26809 10269 26843
rect 12541 26809 12575 26843
rect 12633 26809 12667 26843
rect 14518 26809 14552 26843
rect 18245 26809 18279 26843
rect 19901 26809 19935 26843
rect 21465 26809 21499 26843
rect 21919 26809 21953 26843
rect 23489 26809 23523 26843
rect 23994 26809 24028 26843
rect 25881 26809 25915 26843
rect 30941 26809 30975 26843
rect 32505 26809 32539 26843
rect 35909 26809 35943 26843
rect 37058 26809 37092 26843
rect 38669 26809 38703 26843
rect 39221 26809 39255 26843
rect 41889 26809 41923 26843
rect 5917 26741 5951 26775
rect 8769 26741 8803 26775
rect 13645 26741 13679 26775
rect 16083 26741 16117 26775
rect 17095 26741 17129 26775
rect 17877 26741 17911 26775
rect 20683 26741 20717 26775
rect 21097 26741 21131 26775
rect 22477 26741 22511 26775
rect 28043 26741 28077 26775
rect 30205 26741 30239 26775
rect 33793 26741 33827 26775
rect 36553 26741 36587 26775
rect 37657 26741 37691 26775
rect 39773 26741 39807 26775
rect 40831 26741 40865 26775
rect 42717 26741 42751 26775
rect 3893 26537 3927 26571
rect 4353 26537 4387 26571
rect 5825 26537 5859 26571
rect 7021 26537 7055 26571
rect 7573 26537 7607 26571
rect 8769 26537 8803 26571
rect 11161 26537 11195 26571
rect 13001 26537 13035 26571
rect 16865 26537 16899 26571
rect 18429 26537 18463 26571
rect 21097 26537 21131 26571
rect 22201 26537 22235 26571
rect 24041 26537 24075 26571
rect 24409 26537 24443 26571
rect 27813 26537 27847 26571
rect 32367 26537 32401 26571
rect 35357 26537 35391 26571
rect 35725 26537 35759 26571
rect 36277 26537 36311 26571
rect 10603 26469 10637 26503
rect 14289 26469 14323 26503
rect 15485 26469 15519 26503
rect 16037 26469 16071 26503
rect 17601 26469 17635 26503
rect 18981 26469 19015 26503
rect 22569 26469 22603 26503
rect 24685 26469 24719 26503
rect 27214 26469 27248 26503
rect 28825 26469 28859 26503
rect 33425 26469 33459 26503
rect 38117 26469 38151 26503
rect 38945 26469 38979 26503
rect 39589 26469 39623 26503
rect 39681 26469 39715 26503
rect 40233 26469 40267 26503
rect 41613 26469 41647 26503
rect 41889 26469 41923 26503
rect 42441 26469 42475 26503
rect 43453 26469 43487 26503
rect 43545 26469 43579 26503
rect 4353 26401 4387 26435
rect 4629 26401 4663 26435
rect 5641 26401 5675 26435
rect 8585 26401 8619 26435
rect 12541 26401 12575 26435
rect 13553 26401 13587 26435
rect 14013 26401 14047 26435
rect 19073 26401 19107 26435
rect 21408 26401 21442 26435
rect 30884 26401 30918 26435
rect 32264 26401 32298 26435
rect 34805 26401 34839 26435
rect 35909 26401 35943 26435
rect 6653 26333 6687 26367
rect 10241 26333 10275 26367
rect 13461 26333 13495 26367
rect 15393 26333 15427 26367
rect 17509 26333 17543 26367
rect 18153 26333 18187 26367
rect 22477 26333 22511 26367
rect 24593 26333 24627 26367
rect 26893 26333 26927 26367
rect 28733 26333 28767 26367
rect 33333 26333 33367 26367
rect 38025 26333 38059 26367
rect 41797 26333 41831 26367
rect 43729 26333 43763 26367
rect 21511 26265 21545 26299
rect 23029 26265 23063 26299
rect 25145 26265 25179 26299
rect 29285 26265 29319 26299
rect 31953 26265 31987 26299
rect 33885 26265 33919 26299
rect 38577 26265 38611 26299
rect 39313 26265 39347 26299
rect 9873 26197 9907 26231
rect 12265 26197 12299 26231
rect 12725 26197 12759 26231
rect 14565 26197 14599 26231
rect 19993 26197 20027 26231
rect 21833 26197 21867 26231
rect 28181 26197 28215 26231
rect 30987 26197 31021 26231
rect 31309 26197 31343 26231
rect 32689 26197 32723 26231
rect 34943 26197 34977 26231
rect 36829 26197 36863 26231
rect 4721 25993 4755 26027
rect 5365 25993 5399 26027
rect 6653 25993 6687 26027
rect 8585 25993 8619 26027
rect 11529 25993 11563 26027
rect 13553 25993 13587 26027
rect 14105 25993 14139 26027
rect 15209 25993 15243 26027
rect 15485 25993 15519 26027
rect 15945 25993 15979 26027
rect 16865 25993 16899 26027
rect 17509 25993 17543 26027
rect 18337 25993 18371 26027
rect 19073 25993 19107 26027
rect 21373 25993 21407 26027
rect 22661 25993 22695 26027
rect 23029 25993 23063 26027
rect 24041 25993 24075 26027
rect 25145 25993 25179 26027
rect 25605 25993 25639 26027
rect 27813 25993 27847 26027
rect 28641 25993 28675 26027
rect 33793 25993 33827 26027
rect 35357 25993 35391 26027
rect 37749 25993 37783 26027
rect 39865 25993 39899 26027
rect 42625 25993 42659 26027
rect 43085 25993 43119 26027
rect 4353 25925 4387 25959
rect 10609 25925 10643 25959
rect 20821 25925 20855 25959
rect 22293 25925 22327 25959
rect 26341 25925 26375 25959
rect 32229 25925 32263 25959
rect 34161 25925 34195 25959
rect 38577 25925 38611 25959
rect 42257 25925 42291 25959
rect 5733 25857 5767 25891
rect 8953 25857 8987 25891
rect 14289 25857 14323 25891
rect 19901 25857 19935 25891
rect 24501 25857 24535 25891
rect 25973 25857 26007 25891
rect 27445 25857 27479 25891
rect 31309 25857 31343 25891
rect 31585 25857 31619 25891
rect 35817 25857 35851 25891
rect 38025 25857 38059 25891
rect 39037 25857 39071 25891
rect 44327 25857 44361 25891
rect 3157 25789 3191 25823
rect 4169 25789 4203 25823
rect 4997 25789 5031 25823
rect 5181 25789 5215 25823
rect 7021 25789 7055 25823
rect 7389 25789 7423 25823
rect 7849 25789 7883 25823
rect 8401 25789 8435 25823
rect 9413 25789 9447 25823
rect 9689 25789 9723 25823
rect 10057 25789 10091 25823
rect 10885 25789 10919 25823
rect 11345 25789 11379 25823
rect 12633 25789 12667 25823
rect 13093 25789 13127 25823
rect 16957 25789 16991 25823
rect 18153 25789 18187 25823
rect 26617 25789 26651 25823
rect 26985 25789 27019 25823
rect 30272 25789 30306 25823
rect 30757 25789 30791 25823
rect 34964 25789 34998 25823
rect 36093 25789 36127 25823
rect 40576 25789 40610 25823
rect 40969 25789 41003 25823
rect 43244 25789 43278 25823
rect 43637 25789 43671 25823
rect 44240 25789 44274 25823
rect 44649 25789 44683 25823
rect 10241 25721 10275 25755
rect 14610 25721 14644 25755
rect 19809 25721 19843 25755
rect 20263 25721 20297 25755
rect 21741 25721 21775 25755
rect 21833 25721 21867 25755
rect 24225 25721 24259 25755
rect 24317 25721 24351 25755
rect 27169 25721 27203 25755
rect 31401 25721 31435 25755
rect 32597 25721 32631 25755
rect 32873 25721 32907 25755
rect 32965 25721 32999 25755
rect 33517 25721 33551 25755
rect 36455 25721 36489 25755
rect 38117 25721 38151 25755
rect 41429 25721 41463 25755
rect 41705 25721 41739 25755
rect 41797 25721 41831 25755
rect 44005 25721 44039 25755
rect 3341 25653 3375 25687
rect 3709 25653 3743 25687
rect 4077 25653 4111 25687
rect 6009 25653 6043 25687
rect 6929 25653 6963 25687
rect 8217 25653 8251 25687
rect 11897 25653 11931 25687
rect 12265 25653 12299 25687
rect 12817 25653 12851 25687
rect 17141 25653 17175 25687
rect 17877 25653 17911 25687
rect 27997 25653 28031 25687
rect 29101 25653 29135 25687
rect 30343 25653 30377 25687
rect 31033 25653 31067 25687
rect 35035 25653 35069 25687
rect 37013 25653 37047 25687
rect 37381 25653 37415 25687
rect 39589 25653 39623 25687
rect 40647 25653 40681 25687
rect 43315 25653 43349 25687
rect 4353 25449 4387 25483
rect 6561 25449 6595 25483
rect 7389 25449 7423 25483
rect 10701 25449 10735 25483
rect 16681 25449 16715 25483
rect 17693 25449 17727 25483
rect 18061 25449 18095 25483
rect 21281 25449 21315 25483
rect 24225 25449 24259 25483
rect 27169 25449 27203 25483
rect 28181 25449 28215 25483
rect 33149 25449 33183 25483
rect 36921 25449 36955 25483
rect 38393 25449 38427 25483
rect 41613 25449 41647 25483
rect 41981 25449 42015 25483
rect 44557 25449 44591 25483
rect 5457 25381 5491 25415
rect 6009 25381 6043 25415
rect 6837 25381 6871 25415
rect 8217 25381 8251 25415
rect 10425 25381 10459 25415
rect 12357 25381 12391 25415
rect 14197 25381 14231 25415
rect 19993 25381 20027 25415
rect 24777 25381 24811 25415
rect 27582 25381 27616 25415
rect 29101 25381 29135 25415
rect 29193 25381 29227 25415
rect 33425 25381 33459 25415
rect 33517 25381 33551 25415
rect 35081 25381 35115 25415
rect 36185 25381 36219 25415
rect 38025 25381 38059 25415
rect 39773 25381 39807 25415
rect 40325 25381 40359 25415
rect 43499 25381 43533 25415
rect 1961 25313 1995 25347
rect 2973 25313 3007 25347
rect 4077 25313 4111 25347
rect 4261 25313 4295 25347
rect 5641 25313 5675 25347
rect 7665 25313 7699 25347
rect 8033 25313 8067 25347
rect 9965 25313 9999 25347
rect 10241 25313 10275 25347
rect 11805 25313 11839 25347
rect 11989 25313 12023 25347
rect 13553 25313 13587 25347
rect 14013 25313 14047 25347
rect 14473 25313 14507 25347
rect 15301 25313 15335 25347
rect 16497 25313 16531 25347
rect 17509 25313 17543 25347
rect 19441 25313 19475 25347
rect 19809 25313 19843 25347
rect 23489 25313 23523 25347
rect 27261 25313 27295 25347
rect 30665 25313 30699 25347
rect 32172 25313 32206 25347
rect 38577 25313 38611 25347
rect 41188 25313 41222 25347
rect 42200 25313 42234 25347
rect 43269 25313 43303 25347
rect 44373 25313 44407 25347
rect 9505 25245 9539 25279
rect 20913 25245 20947 25279
rect 23719 25245 23753 25279
rect 24685 25245 24719 25279
rect 30895 25245 30929 25279
rect 32781 25245 32815 25279
rect 33701 25245 33735 25279
rect 34989 25245 35023 25279
rect 35265 25245 35299 25279
rect 39681 25245 39715 25279
rect 22201 25177 22235 25211
rect 25237 25177 25271 25211
rect 29653 25177 29687 25211
rect 36369 25177 36403 25211
rect 2145 25109 2179 25143
rect 3157 25109 3191 25143
rect 4997 25109 5031 25143
rect 8769 25109 8803 25143
rect 15485 25109 15519 25143
rect 21833 25109 21867 25143
rect 28457 25109 28491 25143
rect 31217 25109 31251 25143
rect 31677 25109 31711 25143
rect 32275 25109 32309 25143
rect 34713 25109 34747 25143
rect 36599 25109 36633 25143
rect 38761 25109 38795 25143
rect 41061 25109 41095 25143
rect 41291 25109 41325 25143
rect 42303 25109 42337 25143
rect 3893 24905 3927 24939
rect 9781 24905 9815 24939
rect 13093 24905 13127 24939
rect 14013 24905 14047 24939
rect 15945 24905 15979 24939
rect 18245 24905 18279 24939
rect 19349 24905 19383 24939
rect 21005 24905 21039 24939
rect 22109 24905 22143 24939
rect 23029 24905 23063 24939
rect 23489 24905 23523 24939
rect 24685 24905 24719 24939
rect 25053 24905 25087 24939
rect 26157 24905 26191 24939
rect 29101 24905 29135 24939
rect 33333 24905 33367 24939
rect 33793 24905 33827 24939
rect 35909 24905 35943 24939
rect 39313 24905 39347 24939
rect 40233 24905 40267 24939
rect 41981 24905 42015 24939
rect 43361 24905 43395 24939
rect 2145 24837 2179 24871
rect 2329 24837 2363 24871
rect 6285 24837 6319 24871
rect 11897 24837 11931 24871
rect 17509 24837 17543 24871
rect 24317 24837 24351 24871
rect 27353 24837 27387 24871
rect 28733 24837 28767 24871
rect 1961 24769 1995 24803
rect 3525 24769 3559 24803
rect 4077 24769 4111 24803
rect 4721 24769 4755 24803
rect 7849 24769 7883 24803
rect 8769 24769 8803 24803
rect 9413 24769 9447 24803
rect 18981 24769 19015 24803
rect 20269 24769 20303 24803
rect 20637 24769 20671 24803
rect 21833 24769 21867 24803
rect 23765 24769 23799 24803
rect 25743 24769 25777 24803
rect 27721 24769 27755 24803
rect 29653 24769 29687 24803
rect 30941 24769 30975 24803
rect 32137 24769 32171 24803
rect 32505 24769 32539 24803
rect 33149 24769 33183 24803
rect 2145 24701 2179 24735
rect 2513 24701 2547 24735
rect 3985 24701 4019 24735
rect 4261 24701 4295 24735
rect 5733 24701 5767 24735
rect 7481 24701 7515 24735
rect 8125 24701 8159 24735
rect 8677 24701 8711 24735
rect 8953 24701 8987 24735
rect 10609 24701 10643 24735
rect 12173 24701 12207 24735
rect 12633 24701 12667 24735
rect 13001 24701 13035 24735
rect 14473 24701 14507 24735
rect 14657 24701 14691 24735
rect 14933 24701 14967 24735
rect 15761 24701 15795 24735
rect 17024 24701 17058 24735
rect 18061 24701 18095 24735
rect 18521 24701 18555 24735
rect 19809 24701 19843 24735
rect 20085 24701 20119 24735
rect 25640 24701 25674 24735
rect 26652 24701 26686 24735
rect 28365 24701 28399 24735
rect 31585 24701 31619 24735
rect 2421 24633 2455 24667
rect 4997 24633 5031 24667
rect 7205 24633 7239 24667
rect 7297 24633 7331 24667
rect 10241 24633 10275 24667
rect 10425 24633 10459 24667
rect 12817 24633 12851 24667
rect 13645 24633 13679 24667
rect 15577 24633 15611 24667
rect 16589 24633 16623 24667
rect 21189 24633 21223 24667
rect 21281 24633 21315 24667
rect 23857 24633 23891 24667
rect 26755 24633 26789 24667
rect 27813 24633 27847 24667
rect 29377 24633 29411 24667
rect 29469 24633 29503 24667
rect 31033 24633 31067 24667
rect 32597 24633 32631 24667
rect 36277 24837 36311 24871
rect 35265 24769 35299 24803
rect 36829 24769 36863 24803
rect 38025 24701 38059 24735
rect 38485 24701 38519 24735
rect 39440 24701 39474 24735
rect 39865 24701 39899 24735
rect 42844 24701 42878 24735
rect 43888 24701 43922 24735
rect 44868 24701 44902 24735
rect 45293 24701 45327 24735
rect 34989 24633 35023 24667
rect 35081 24633 35115 24667
rect 36553 24633 36587 24667
rect 36645 24633 36679 24667
rect 41061 24633 41095 24667
rect 41153 24633 41187 24667
rect 41705 24633 41739 24667
rect 44281 24633 44315 24667
rect 5549 24565 5583 24599
rect 5917 24565 5951 24599
rect 6653 24565 6687 24599
rect 8493 24565 8527 24599
rect 10701 24565 10735 24599
rect 11253 24565 11287 24599
rect 15209 24565 15243 24599
rect 17095 24565 17129 24599
rect 22477 24565 22511 24599
rect 26525 24565 26559 24599
rect 30297 24565 30331 24599
rect 30757 24565 30791 24599
rect 33333 24565 33367 24599
rect 33517 24565 33551 24599
rect 34345 24565 34379 24599
rect 34713 24565 34747 24599
rect 37565 24565 37599 24599
rect 38209 24565 38243 24599
rect 38853 24565 38887 24599
rect 39543 24565 39577 24599
rect 40877 24565 40911 24599
rect 42625 24565 42659 24599
rect 42947 24565 42981 24599
rect 43959 24565 43993 24599
rect 44649 24565 44683 24599
rect 44971 24565 45005 24599
rect 2237 24361 2271 24395
rect 3341 24361 3375 24395
rect 4721 24361 4755 24395
rect 7481 24361 7515 24395
rect 10057 24361 10091 24395
rect 10425 24361 10459 24395
rect 11161 24361 11195 24395
rect 12541 24361 12575 24395
rect 14565 24361 14599 24395
rect 19073 24361 19107 24395
rect 19993 24361 20027 24395
rect 24409 24361 24443 24395
rect 27721 24361 27755 24395
rect 28917 24361 28951 24395
rect 29653 24361 29687 24395
rect 32919 24361 32953 24395
rect 34713 24361 34747 24395
rect 42165 24361 42199 24395
rect 45109 24361 45143 24395
rect 4077 24293 4111 24327
rect 6377 24293 6411 24327
rect 6745 24293 6779 24327
rect 10885 24293 10919 24327
rect 13645 24293 13679 24327
rect 14197 24293 14231 24327
rect 15663 24293 15697 24327
rect 17049 24293 17083 24327
rect 19625 24293 19659 24327
rect 21189 24293 21223 24327
rect 22845 24293 22879 24327
rect 22937 24293 22971 24327
rect 24777 24293 24811 24327
rect 28318 24293 28352 24327
rect 30665 24293 30699 24327
rect 32689 24293 32723 24327
rect 33333 24293 33367 24327
rect 34989 24293 35023 24327
rect 39542 24293 39576 24327
rect 41153 24293 41187 24327
rect 43545 24293 43579 24327
rect 1869 24225 1903 24259
rect 2973 24225 3007 24259
rect 5641 24225 5675 24259
rect 5917 24225 5951 24259
rect 7205 24225 7239 24259
rect 7389 24225 7423 24259
rect 8585 24225 8619 24259
rect 9873 24225 9907 24259
rect 11069 24225 11103 24259
rect 12265 24225 12299 24259
rect 12449 24225 12483 24259
rect 13829 24225 13863 24259
rect 17969 24225 18003 24259
rect 18889 24225 18923 24259
rect 26525 24225 26559 24259
rect 33860 24225 33894 24259
rect 36404 24225 36438 24259
rect 40141 24225 40175 24259
rect 44925 24225 44959 24259
rect 3893 24157 3927 24191
rect 4445 24157 4479 24191
rect 15301 24157 15335 24191
rect 17325 24157 17359 24191
rect 21097 24157 21131 24191
rect 21741 24157 21775 24191
rect 23121 24157 23155 24191
rect 24685 24157 24719 24191
rect 24961 24157 24995 24191
rect 27997 24157 28031 24191
rect 30573 24157 30607 24191
rect 32413 24157 32447 24191
rect 34897 24157 34931 24191
rect 39221 24157 39255 24191
rect 41061 24157 41095 24191
rect 41705 24157 41739 24191
rect 43453 24157 43487 24191
rect 43729 24157 43763 24191
rect 4353 24089 4387 24123
rect 5457 24089 5491 24123
rect 5733 24089 5767 24123
rect 8125 24089 8159 24123
rect 13185 24089 13219 24123
rect 14841 24089 14875 24123
rect 31125 24089 31159 24123
rect 33931 24089 33965 24123
rect 35449 24089 35483 24123
rect 37565 24089 37599 24123
rect 37887 24089 37921 24123
rect 38577 24089 38611 24123
rect 4242 24021 4276 24055
rect 5089 24021 5123 24055
rect 7113 24021 7147 24055
rect 8769 24021 8803 24055
rect 9137 24021 9171 24055
rect 13553 24021 13587 24055
rect 16221 24021 16255 24055
rect 23857 24021 23891 24055
rect 26709 24021 26743 24055
rect 27077 24021 27111 24055
rect 29285 24021 29319 24055
rect 31493 24021 31527 24055
rect 36507 24021 36541 24055
rect 36921 24021 36955 24055
rect 38209 24021 38243 24055
rect 2421 23817 2455 23851
rect 2789 23817 2823 23851
rect 3433 23817 3467 23851
rect 4169 23817 4203 23851
rect 7389 23817 7423 23851
rect 7849 23817 7883 23851
rect 8585 23817 8619 23851
rect 11529 23817 11563 23851
rect 12265 23817 12299 23851
rect 13461 23817 13495 23851
rect 14749 23817 14783 23851
rect 15025 23817 15059 23851
rect 16405 23817 16439 23851
rect 17785 23817 17819 23851
rect 19809 23817 19843 23851
rect 22477 23817 22511 23851
rect 25605 23817 25639 23851
rect 28365 23817 28399 23851
rect 30941 23817 30975 23851
rect 31033 23817 31067 23851
rect 34253 23817 34287 23851
rect 34621 23817 34655 23851
rect 36369 23817 36403 23851
rect 37749 23817 37783 23851
rect 41981 23817 42015 23851
rect 45477 23817 45511 23851
rect 3249 23749 3283 23783
rect 4353 23749 4387 23783
rect 5089 23749 5123 23783
rect 19073 23749 19107 23783
rect 25145 23749 25179 23783
rect 26249 23749 26283 23783
rect 26525 23749 26559 23783
rect 30343 23749 30377 23783
rect 3341 23681 3375 23715
rect 1961 23613 1995 23647
rect 2973 23613 3007 23647
rect 3120 23613 3154 23647
rect 4445 23681 4479 23715
rect 7021 23681 7055 23715
rect 7720 23681 7754 23715
rect 7941 23681 7975 23715
rect 8953 23681 8987 23715
rect 9873 23681 9907 23715
rect 10241 23681 10275 23715
rect 14381 23681 14415 23715
rect 15209 23681 15243 23715
rect 21189 23681 21223 23715
rect 24593 23681 24627 23715
rect 27997 23681 28031 23715
rect 4997 23613 5031 23647
rect 5273 23613 5307 23647
rect 7573 23613 7607 23647
rect 9137 23613 9171 23647
rect 9229 23613 9263 23647
rect 9413 23613 9447 23647
rect 10885 23613 10919 23647
rect 11253 23613 11287 23647
rect 12449 23613 12483 23647
rect 12909 23613 12943 23647
rect 13645 23613 13679 23647
rect 14105 23613 14139 23647
rect 16129 23613 16163 23647
rect 16773 23613 16807 23647
rect 16992 23613 17026 23647
rect 18153 23613 18187 23647
rect 19625 23613 19659 23647
rect 20085 23613 20119 23647
rect 22636 23613 22670 23647
rect 23029 23613 23063 23647
rect 26709 23613 26743 23647
rect 27169 23613 27203 23647
rect 30240 23613 30274 23647
rect 30665 23613 30699 23647
rect 32229 23749 32263 23783
rect 32781 23749 32815 23783
rect 42625 23749 42659 23783
rect 31309 23681 31343 23715
rect 31585 23681 31619 23715
rect 35449 23681 35483 23715
rect 36553 23681 36587 23715
rect 38117 23681 38151 23715
rect 38393 23681 38427 23715
rect 39589 23681 39623 23715
rect 40325 23681 40359 23715
rect 41061 23681 41095 23715
rect 43177 23681 43211 23715
rect 43545 23681 43579 23715
rect 44684 23613 44718 23647
rect 45109 23613 45143 23647
rect 5733 23545 5767 23579
rect 8309 23545 8343 23579
rect 10701 23545 10735 23579
rect 15530 23545 15564 23579
rect 17095 23545 17129 23579
rect 20729 23545 20763 23579
rect 20821 23545 20855 23579
rect 24685 23545 24719 23579
rect 27445 23545 27479 23579
rect 30941 23545 30975 23579
rect 31401 23545 31435 23579
rect 33333 23545 33367 23579
rect 33425 23545 33459 23579
rect 33977 23545 34011 23579
rect 34989 23545 35023 23579
rect 35081 23545 35115 23579
rect 36645 23545 36679 23579
rect 37197 23545 37231 23579
rect 38209 23545 38243 23579
rect 40877 23545 40911 23579
rect 41153 23545 41187 23579
rect 41705 23545 41739 23579
rect 43269 23545 43303 23579
rect 44097 23545 44131 23579
rect 1777 23477 1811 23511
rect 2145 23477 2179 23511
rect 4353 23477 4387 23511
rect 4813 23477 4847 23511
rect 6009 23477 6043 23511
rect 6653 23477 6687 23511
rect 10517 23477 10551 23511
rect 12633 23477 12667 23511
rect 17509 23477 17543 23511
rect 18521 23477 18555 23511
rect 20545 23477 20579 23511
rect 21649 23477 21683 23511
rect 22707 23477 22741 23511
rect 23489 23477 23523 23511
rect 24041 23477 24075 23511
rect 24409 23477 24443 23511
rect 29745 23477 29779 23511
rect 35909 23477 35943 23511
rect 39313 23477 39347 23511
rect 42901 23477 42935 23511
rect 44787 23477 44821 23511
rect 2513 23273 2547 23307
rect 7665 23273 7699 23307
rect 9229 23273 9263 23307
rect 10701 23273 10735 23307
rect 12357 23273 12391 23307
rect 14197 23273 14231 23307
rect 15485 23273 15519 23307
rect 20729 23273 20763 23307
rect 21051 23273 21085 23307
rect 28917 23273 28951 23307
rect 31309 23273 31343 23307
rect 32505 23273 32539 23307
rect 33057 23273 33091 23307
rect 35265 23273 35299 23307
rect 37105 23273 37139 23307
rect 43177 23273 43211 23307
rect 45063 23273 45097 23307
rect 4261 23205 4295 23239
rect 11621 23205 11655 23239
rect 17049 23205 17083 23239
rect 18613 23205 18647 23239
rect 21373 23205 21407 23239
rect 23121 23205 23155 23239
rect 24685 23205 24719 23239
rect 28359 23205 28393 23239
rect 30987 23205 31021 23239
rect 34069 23205 34103 23239
rect 34897 23205 34931 23239
rect 36277 23205 36311 23239
rect 38577 23205 38611 23239
rect 39726 23205 39760 23239
rect 41061 23205 41095 23239
rect 41337 23205 41371 23239
rect 41889 23205 41923 23239
rect 43545 23205 43579 23239
rect 2329 23137 2363 23171
rect 4445 23137 4479 23171
rect 5641 23137 5675 23171
rect 6745 23137 6779 23171
rect 7205 23137 7239 23171
rect 8217 23137 8251 23171
rect 8401 23137 8435 23171
rect 8769 23137 8803 23171
rect 9689 23137 9723 23171
rect 9873 23137 9907 23171
rect 11069 23137 11103 23171
rect 11253 23137 11287 23171
rect 13461 23137 13495 23171
rect 13645 23137 13679 23171
rect 15920 23137 15954 23171
rect 20980 23137 21014 23171
rect 21925 23137 21959 23171
rect 26709 23137 26743 23171
rect 27997 23137 28031 23171
rect 29745 23137 29779 23171
rect 30884 23137 30918 23171
rect 33149 23137 33183 23171
rect 37841 23137 37875 23171
rect 38301 23137 38335 23171
rect 38853 23137 38887 23171
rect 44925 23137 44959 23171
rect 6009 23069 6043 23103
rect 8125 23069 8159 23103
rect 10241 23069 10275 23103
rect 13921 23069 13955 23103
rect 16957 23069 16991 23103
rect 18521 23069 18555 23103
rect 23029 23069 23063 23103
rect 23305 23069 23339 23103
rect 24593 23069 24627 23103
rect 24869 23069 24903 23103
rect 32137 23069 32171 23103
rect 5181 23001 5215 23035
rect 5549 23001 5583 23035
rect 6285 23001 6319 23035
rect 7389 23001 7423 23035
rect 15991 23001 16025 23035
rect 17509 23001 17543 23035
rect 19073 23001 19107 23035
rect 26893 23001 26927 23035
rect 29929 23001 29963 23035
rect 33333 23069 33367 23103
rect 33977 23069 34011 23103
rect 34253 23069 34287 23103
rect 36185 23069 36219 23103
rect 39405 23069 39439 23103
rect 41245 23069 41279 23103
rect 43453 23069 43487 23103
rect 43729 23069 43763 23103
rect 35633 23001 35667 23035
rect 36737 23001 36771 23035
rect 40325 23001 40359 23035
rect 2973 22933 3007 22967
rect 3341 22933 3375 22967
rect 3801 22933 3835 22967
rect 4537 22933 4571 22967
rect 5779 22933 5813 22967
rect 5917 22933 5951 22967
rect 7021 22933 7055 22967
rect 18153 22933 18187 22967
rect 22109 22933 22143 22967
rect 27169 22933 27203 22967
rect 29285 22933 29319 22967
rect 30481 22933 30515 22967
rect 33149 22933 33183 22967
rect 3985 22729 4019 22763
rect 4353 22729 4387 22763
rect 6377 22729 6411 22763
rect 7021 22729 7055 22763
rect 7297 22729 7331 22763
rect 7849 22729 7883 22763
rect 8217 22729 8251 22763
rect 9781 22729 9815 22763
rect 11437 22729 11471 22763
rect 16037 22729 16071 22763
rect 16773 22729 16807 22763
rect 17417 22729 17451 22763
rect 21005 22729 21039 22763
rect 21281 22729 21315 22763
rect 23397 22729 23431 22763
rect 25513 22729 25547 22763
rect 26249 22729 26283 22763
rect 26617 22729 26651 22763
rect 28365 22729 28399 22763
rect 29469 22729 29503 22763
rect 32965 22729 32999 22763
rect 33701 22729 33735 22763
rect 33931 22729 33965 22763
rect 34713 22729 34747 22763
rect 35035 22729 35069 22763
rect 35817 22729 35851 22763
rect 37427 22729 37461 22763
rect 38117 22729 38151 22763
rect 40325 22729 40359 22763
rect 40647 22729 40681 22763
rect 41337 22729 41371 22763
rect 42625 22729 42659 22763
rect 5641 22661 5675 22695
rect 6101 22661 6135 22695
rect 15301 22661 15335 22695
rect 17141 22661 17175 22695
rect 22845 22661 22879 22695
rect 23121 22661 23155 22695
rect 36093 22661 36127 22695
rect 37197 22661 37231 22695
rect 41981 22661 42015 22695
rect 2881 22593 2915 22627
rect 9413 22593 9447 22627
rect 13277 22593 13311 22627
rect 17877 22593 17911 22627
rect 24593 22593 24627 22627
rect 27445 22593 27479 22627
rect 39129 22593 39163 22627
rect 39773 22593 39807 22627
rect 43177 22593 43211 22627
rect 2237 22525 2271 22559
rect 3157 22525 3191 22559
rect 4445 22525 4479 22559
rect 4905 22525 4939 22559
rect 6837 22525 6871 22559
rect 8585 22525 8619 22559
rect 8769 22525 8803 22559
rect 10793 22525 10827 22559
rect 13369 22525 13403 22559
rect 14565 22525 14599 22559
rect 15117 22525 15151 22559
rect 15577 22525 15611 22559
rect 16957 22525 16991 22559
rect 18705 22525 18739 22559
rect 20085 22525 20119 22559
rect 22017 22525 22051 22559
rect 22477 22525 22511 22559
rect 22845 22525 22879 22559
rect 23673 22525 23707 22559
rect 24685 22525 24719 22559
rect 25145 22525 25179 22559
rect 25697 22525 25731 22559
rect 26801 22525 26835 22559
rect 27169 22525 27203 22559
rect 28089 22525 28123 22559
rect 29285 22525 29319 22559
rect 30481 22525 30515 22559
rect 31033 22525 31067 22559
rect 31217 22525 31251 22559
rect 32045 22525 32079 22559
rect 33241 22525 33275 22559
rect 33828 22525 33862 22559
rect 34253 22525 34287 22559
rect 34932 22525 34966 22559
rect 36344 22525 36378 22559
rect 36737 22525 36771 22559
rect 37356 22525 37390 22559
rect 38393 22525 38427 22559
rect 38853 22525 38887 22559
rect 40576 22525 40610 22559
rect 41556 22525 41590 22559
rect 3617 22457 3651 22491
rect 5181 22457 5215 22491
rect 9137 22457 9171 22491
rect 10609 22457 10643 22491
rect 11161 22457 11195 22491
rect 12909 22457 12943 22491
rect 18061 22457 18095 22491
rect 19993 22457 20027 22491
rect 20406 22457 20440 22491
rect 22753 22457 22787 22491
rect 24225 22457 24259 22491
rect 30021 22457 30055 22491
rect 32407 22457 32441 22491
rect 37841 22457 37875 22491
rect 43269 22457 43303 22491
rect 43821 22457 43855 22491
rect 1961 22389 1995 22423
rect 10149 22389 10183 22423
rect 11805 22389 11839 22423
rect 13737 22389 13771 22423
rect 14289 22389 14323 22423
rect 19073 22389 19107 22423
rect 21833 22389 21867 22423
rect 23857 22389 23891 22423
rect 24869 22389 24903 22423
rect 25881 22389 25915 22423
rect 29009 22389 29043 22423
rect 30297 22389 30331 22423
rect 31585 22389 31619 22423
rect 31861 22389 31895 22423
rect 35357 22389 35391 22423
rect 36415 22389 36449 22423
rect 39497 22389 39531 22423
rect 41061 22389 41095 22423
rect 41659 22389 41693 22423
rect 42993 22389 43027 22423
rect 44097 22389 44131 22423
rect 44925 22389 44959 22423
rect 4353 22185 4387 22219
rect 4445 22185 4479 22219
rect 4629 22185 4663 22219
rect 5549 22185 5583 22219
rect 6469 22185 6503 22219
rect 8309 22185 8343 22219
rect 8677 22185 8711 22219
rect 10701 22185 10735 22219
rect 14013 22185 14047 22219
rect 19487 22185 19521 22219
rect 23305 22185 23339 22219
rect 23857 22185 23891 22219
rect 24593 22185 24627 22219
rect 26801 22185 26835 22219
rect 32919 22185 32953 22219
rect 38393 22185 38427 22219
rect 42257 22185 42291 22219
rect 43177 22185 43211 22219
rect 2789 22117 2823 22151
rect 2145 22049 2179 22083
rect 4169 22049 4203 22083
rect 7113 22117 7147 22151
rect 13369 22117 13403 22151
rect 15485 22117 15519 22151
rect 17877 22117 17911 22151
rect 17969 22117 18003 22151
rect 18797 22117 18831 22151
rect 21097 22117 21131 22151
rect 21649 22117 21683 22151
rect 24869 22117 24903 22151
rect 28825 22117 28859 22151
rect 31217 22117 31251 22151
rect 32321 22117 32355 22151
rect 33977 22117 34011 22151
rect 36001 22117 36035 22151
rect 36185 22117 36219 22151
rect 36277 22117 36311 22151
rect 41429 22117 41463 22151
rect 8493 22049 8527 22083
rect 9689 22049 9723 22083
rect 11529 22049 11563 22083
rect 12633 22049 12667 22083
rect 13093 22049 13127 22083
rect 14197 22049 14231 22083
rect 19384 22049 19418 22083
rect 27077 22049 27111 22083
rect 28089 22049 28123 22083
rect 30481 22049 30515 22083
rect 31033 22049 31067 22083
rect 32848 22049 32882 22083
rect 37816 22049 37850 22083
rect 38761 22049 38795 22083
rect 39221 22049 39255 22083
rect 43396 22049 43430 22083
rect 44373 22049 44407 22083
rect 5181 21981 5215 22015
rect 7021 21981 7055 22015
rect 15393 21981 15427 22015
rect 18521 21981 18555 22015
rect 21005 21981 21039 22015
rect 22937 21981 22971 22015
rect 24777 21981 24811 22015
rect 25053 21981 25087 22015
rect 28457 21981 28491 22015
rect 30389 21981 30423 22015
rect 33885 21981 33919 22015
rect 34161 21981 34195 22015
rect 36829 21981 36863 22015
rect 39497 21981 39531 22015
rect 41337 21981 41371 22015
rect 41613 21981 41647 22015
rect 43913 21981 43947 22015
rect 6101 21913 6135 21947
rect 7573 21913 7607 21947
rect 9873 21913 9907 21947
rect 13645 21913 13679 21947
rect 14335 21913 14369 21947
rect 15945 21913 15979 21947
rect 27629 21913 27663 21947
rect 29377 21913 29411 21947
rect 43499 21913 43533 21947
rect 4445 21845 4479 21879
rect 4997 21845 5031 21879
rect 10977 21845 11011 21879
rect 11713 21845 11747 21879
rect 20177 21845 20211 21879
rect 22109 21845 22143 21879
rect 22385 21845 22419 21879
rect 25789 21845 25823 21879
rect 27261 21845 27295 21879
rect 27905 21845 27939 21879
rect 28227 21845 28261 21879
rect 28365 21845 28399 21879
rect 29653 21845 29687 21879
rect 35357 21845 35391 21879
rect 37887 21845 37921 21879
rect 40509 21845 40543 21879
rect 44189 21845 44223 21879
rect 44557 21845 44591 21879
rect 2513 21641 2547 21675
rect 3525 21641 3559 21675
rect 4077 21641 4111 21675
rect 4537 21641 4571 21675
rect 5825 21641 5859 21675
rect 8033 21641 8067 21675
rect 8401 21641 8435 21675
rect 11805 21641 11839 21675
rect 12909 21641 12943 21675
rect 15209 21641 15243 21675
rect 17509 21641 17543 21675
rect 19257 21641 19291 21675
rect 19533 21641 19567 21675
rect 21005 21641 21039 21675
rect 21649 21641 21683 21675
rect 22753 21641 22787 21675
rect 23397 21641 23431 21675
rect 25513 21641 25547 21675
rect 25881 21641 25915 21675
rect 26985 21641 27019 21675
rect 27997 21641 28031 21675
rect 31861 21641 31895 21675
rect 31953 21641 31987 21675
rect 34161 21641 34195 21675
rect 43361 21641 43395 21675
rect 9321 21573 9355 21607
rect 10701 21573 10735 21607
rect 17785 21573 17819 21607
rect 27813 21573 27847 21607
rect 29423 21573 29457 21607
rect 29561 21573 29595 21607
rect 31033 21573 31067 21607
rect 4629 21505 4663 21539
rect 9045 21505 9079 21539
rect 9689 21505 9723 21539
rect 13921 21505 13955 21539
rect 16037 21505 16071 21539
rect 18153 21505 18187 21539
rect 18613 21505 18647 21539
rect 20269 21505 20303 21539
rect 24409 21505 24443 21539
rect 25605 21505 25639 21539
rect 26249 21505 26283 21539
rect 26617 21505 26651 21539
rect 27905 21505 27939 21539
rect 29653 21505 29687 21539
rect 30021 21505 30055 21539
rect 37473 21573 37507 21607
rect 33701 21505 33735 21539
rect 35357 21505 35391 21539
rect 35633 21505 35667 21539
rect 36921 21505 36955 21539
rect 39589 21505 39623 21539
rect 40509 21505 40543 21539
rect 42349 21505 42383 21539
rect 42993 21505 43027 21539
rect 43913 21505 43947 21539
rect 44189 21505 44223 21539
rect 2329 21437 2363 21471
rect 2789 21437 2823 21471
rect 3652 21437 3686 21471
rect 3755 21437 3789 21471
rect 6193 21437 6227 21471
rect 8493 21437 8527 21471
rect 8677 21437 8711 21471
rect 12484 21437 12518 21471
rect 13737 21437 13771 21471
rect 19717 21437 19751 21471
rect 20177 21437 20211 21471
rect 21373 21437 21407 21471
rect 21833 21437 21867 21471
rect 25384 21437 25418 21471
rect 27684 21437 27718 21471
rect 30849 21437 30883 21471
rect 31309 21437 31343 21471
rect 31861 21437 31895 21471
rect 32137 21437 32171 21471
rect 32597 21437 32631 21471
rect 37933 21437 37967 21471
rect 38853 21437 38887 21471
rect 39313 21437 39347 21471
rect 39865 21437 39899 21471
rect 4991 21369 5025 21403
rect 6929 21369 6963 21403
rect 7021 21369 7055 21403
rect 7573 21369 7607 21403
rect 10333 21369 10367 21403
rect 10885 21369 10919 21403
rect 10977 21369 11011 21403
rect 11529 21369 11563 21403
rect 15761 21369 15795 21403
rect 15853 21369 15887 21403
rect 18245 21369 18279 21403
rect 22154 21369 22188 21403
rect 23029 21369 23063 21403
rect 23765 21369 23799 21403
rect 23857 21369 23891 21403
rect 24777 21369 24811 21403
rect 25237 21369 25271 21403
rect 27537 21369 27571 21403
rect 29101 21369 29135 21403
rect 29284 21369 29318 21403
rect 30481 21369 30515 21403
rect 32873 21369 32907 21403
rect 33241 21369 33275 21403
rect 35449 21369 35483 21403
rect 37013 21369 37047 21403
rect 38669 21369 38703 21403
rect 40830 21369 40864 21403
rect 42441 21369 42475 21403
rect 44005 21369 44039 21403
rect 2053 21301 2087 21335
rect 5549 21301 5583 21335
rect 6653 21301 6687 21335
rect 12173 21301 12207 21335
rect 12587 21301 12621 21335
rect 13277 21301 13311 21335
rect 14289 21301 14323 21335
rect 14841 21301 14875 21335
rect 15577 21301 15611 21335
rect 25145 21301 25179 21335
rect 27445 21301 27479 21335
rect 28549 21301 28583 21335
rect 34529 21301 34563 21335
rect 35081 21301 35115 21335
rect 36277 21301 36311 21335
rect 36645 21301 36679 21335
rect 38301 21301 38335 21335
rect 40325 21301 40359 21335
rect 41429 21301 41463 21335
rect 41705 21301 41739 21335
rect 42073 21301 42107 21335
rect 44833 21301 44867 21335
rect 5181 21097 5215 21131
rect 5963 21097 5997 21131
rect 7297 21097 7331 21131
rect 10609 21097 10643 21131
rect 14289 21097 14323 21131
rect 15439 21097 15473 21131
rect 15761 21097 15795 21131
rect 16129 21097 16163 21131
rect 18521 21097 18555 21131
rect 19809 21097 19843 21131
rect 21741 21097 21775 21131
rect 22937 21097 22971 21131
rect 23765 21097 23799 21131
rect 24409 21097 24443 21131
rect 28227 21097 28261 21131
rect 29745 21097 29779 21131
rect 32413 21097 32447 21131
rect 33333 21097 33367 21131
rect 33885 21097 33919 21131
rect 35127 21097 35161 21131
rect 37013 21097 37047 21131
rect 38715 21097 38749 21131
rect 41153 21097 41187 21131
rect 4813 21029 4847 21063
rect 10051 21029 10085 21063
rect 11621 21029 11655 21063
rect 17325 21029 17359 21063
rect 25605 21029 25639 21063
rect 30113 21029 30147 21063
rect 36185 21029 36219 21063
rect 39129 21029 39163 21063
rect 39951 21029 39985 21063
rect 41521 21029 41555 21063
rect 42073 21029 42107 21063
rect 43545 21029 43579 21063
rect 44097 21029 44131 21063
rect 4077 20961 4111 20995
rect 4629 20961 4663 20995
rect 5860 20961 5894 20995
rect 7757 20961 7791 20995
rect 8217 20961 8251 20995
rect 13001 20961 13035 20995
rect 13461 20961 13495 20995
rect 15336 20961 15370 20995
rect 18797 20961 18831 20995
rect 21925 20961 21959 20995
rect 22109 20961 22143 20995
rect 23213 20961 23247 20995
rect 24869 20961 24903 20995
rect 26525 20961 26559 20995
rect 28124 20961 28158 20995
rect 29101 20961 29135 20995
rect 30665 20961 30699 20995
rect 32965 20961 32999 20995
rect 35056 20961 35090 20995
rect 39589 20961 39623 20995
rect 44976 20961 45010 20995
rect 8493 20893 8527 20927
rect 9689 20893 9723 20927
rect 11529 20893 11563 20927
rect 13553 20893 13587 20927
rect 17233 20893 17267 20927
rect 17877 20893 17911 20927
rect 25016 20893 25050 20927
rect 25237 20893 25271 20927
rect 26893 20893 26927 20927
rect 28917 20893 28951 20927
rect 29469 20893 29503 20927
rect 30481 20893 30515 20927
rect 36093 20893 36127 20927
rect 36369 20893 36403 20927
rect 41429 20893 41463 20927
rect 43453 20893 43487 20927
rect 45063 20893 45097 20927
rect 12081 20825 12115 20859
rect 14565 20825 14599 20859
rect 20637 20825 20671 20859
rect 23397 20825 23431 20859
rect 26341 20825 26375 20859
rect 26985 20825 27019 20859
rect 29248 20825 29282 20859
rect 30849 20825 30883 20859
rect 31125 20825 31159 20859
rect 38485 20825 38519 20859
rect 7021 20757 7055 20791
rect 18245 20757 18279 20791
rect 18981 20757 19015 20791
rect 21281 20757 21315 20791
rect 24777 20757 24811 20791
rect 25145 20757 25179 20791
rect 25881 20757 25915 20791
rect 26663 20757 26697 20791
rect 26801 20757 26835 20791
rect 27629 20757 27663 20791
rect 27997 20757 28031 20791
rect 28641 20757 28675 20791
rect 29377 20757 29411 20791
rect 31585 20757 31619 20791
rect 40509 20757 40543 20791
rect 3801 20553 3835 20587
rect 4169 20553 4203 20587
rect 5825 20553 5859 20587
rect 7665 20553 7699 20587
rect 11207 20553 11241 20587
rect 11989 20553 12023 20587
rect 13277 20553 13311 20587
rect 13645 20553 13679 20587
rect 15301 20553 15335 20587
rect 19073 20553 19107 20587
rect 21097 20553 21131 20587
rect 23121 20553 23155 20587
rect 25973 20553 26007 20587
rect 26893 20553 26927 20587
rect 27261 20553 27295 20587
rect 30297 20553 30331 20587
rect 30481 20553 30515 20587
rect 30665 20553 30699 20587
rect 30987 20553 31021 20587
rect 31493 20553 31527 20587
rect 31953 20553 31987 20587
rect 35633 20553 35667 20587
rect 35863 20553 35897 20587
rect 36553 20553 36587 20587
rect 38117 20553 38151 20587
rect 39313 20553 39347 20587
rect 40785 20553 40819 20587
rect 41061 20553 41095 20587
rect 42625 20553 42659 20587
rect 42993 20553 43027 20587
rect 43361 20553 43395 20587
rect 2605 20485 2639 20519
rect 22201 20485 22235 20519
rect 25789 20485 25823 20519
rect 29423 20485 29457 20519
rect 29561 20485 29595 20519
rect 11529 20417 11563 20451
rect 18153 20417 18187 20451
rect 19717 20417 19751 20451
rect 24225 20417 24259 20451
rect 25881 20417 25915 20451
rect 27537 20417 27571 20451
rect 29653 20417 29687 20451
rect 31125 20485 31159 20519
rect 37657 20485 37691 20519
rect 44097 20485 44131 20519
rect 33149 20417 33183 20451
rect 38577 20417 38611 20451
rect 39543 20417 39577 20451
rect 43545 20417 43579 20451
rect 44465 20417 44499 20451
rect 45477 20417 45511 20451
rect 2697 20349 2731 20383
rect 3249 20349 3283 20383
rect 3433 20349 3467 20383
rect 4261 20349 4295 20383
rect 7757 20349 7791 20383
rect 8217 20349 8251 20383
rect 8493 20349 8527 20383
rect 9321 20349 9355 20383
rect 10241 20349 10275 20383
rect 10885 20349 10919 20383
rect 11104 20349 11138 20383
rect 12817 20349 12851 20383
rect 13829 20349 13863 20383
rect 14749 20349 14783 20383
rect 15612 20349 15646 20383
rect 16037 20349 16071 20383
rect 16624 20349 16658 20383
rect 21281 20349 21315 20383
rect 23397 20349 23431 20383
rect 23857 20349 23891 20383
rect 25660 20349 25694 20383
rect 26525 20349 26559 20383
rect 27077 20349 27111 20383
rect 28181 20349 28215 20383
rect 30481 20349 30515 20383
rect 30849 20349 30883 20383
rect 31188 20349 31222 20383
rect 31677 20349 31711 20383
rect 32229 20349 32263 20383
rect 35792 20349 35826 20383
rect 36185 20349 36219 20383
rect 36988 20349 37022 20383
rect 37381 20349 37415 20383
rect 37657 20349 37691 20383
rect 37933 20349 37967 20383
rect 39456 20349 39490 20383
rect 4623 20281 4657 20315
rect 5549 20281 5583 20315
rect 9229 20281 9263 20315
rect 9683 20281 9717 20315
rect 18245 20281 18279 20315
rect 18797 20281 18831 20315
rect 19809 20281 19843 20315
rect 20361 20281 20395 20315
rect 21189 20281 21223 20315
rect 23673 20281 23707 20315
rect 24501 20281 24535 20315
rect 25513 20281 25547 20315
rect 29009 20281 29043 20315
rect 29285 20281 29319 20315
rect 30021 20281 30055 20315
rect 33241 20281 33275 20315
rect 33793 20281 33827 20315
rect 40233 20281 40267 20315
rect 41337 20281 41371 20315
rect 41429 20281 41463 20315
rect 41981 20281 42015 20315
rect 43637 20281 43671 20315
rect 5181 20213 5215 20247
rect 7297 20213 7331 20247
rect 8861 20213 8895 20247
rect 10609 20213 10643 20247
rect 12725 20213 12759 20247
rect 13001 20213 13035 20247
rect 14197 20213 14231 20247
rect 15715 20213 15749 20247
rect 16405 20213 16439 20247
rect 16727 20213 16761 20247
rect 17233 20213 17267 20247
rect 17785 20213 17819 20247
rect 19533 20213 19567 20247
rect 24961 20213 24995 20247
rect 25329 20213 25363 20247
rect 27997 20213 28031 20247
rect 28365 20213 28399 20247
rect 28733 20213 28767 20247
rect 31677 20213 31711 20247
rect 32873 20213 32907 20247
rect 34069 20213 34103 20247
rect 35173 20213 35207 20247
rect 37059 20213 37093 20247
rect 37749 20213 37783 20247
rect 39957 20213 39991 20247
rect 45017 20213 45051 20247
rect 2789 20009 2823 20043
rect 3801 20009 3835 20043
rect 4721 20009 4755 20043
rect 7757 20009 7791 20043
rect 8309 20009 8343 20043
rect 9321 20009 9355 20043
rect 10517 20009 10551 20043
rect 13829 20009 13863 20043
rect 14381 20009 14415 20043
rect 16957 20009 16991 20043
rect 18153 20009 18187 20043
rect 20085 20009 20119 20043
rect 26341 20009 26375 20043
rect 27169 20009 27203 20043
rect 27629 20009 27663 20043
rect 28825 20009 28859 20043
rect 30757 20009 30791 20043
rect 31769 20009 31803 20043
rect 32597 20009 32631 20043
rect 33425 20009 33459 20043
rect 33885 20009 33919 20043
rect 40969 20009 41003 20043
rect 41337 20009 41371 20043
rect 6745 19941 6779 19975
rect 12633 19941 12667 19975
rect 15485 19941 15519 19975
rect 15577 19941 15611 19975
rect 17325 19941 17359 19975
rect 18889 19941 18923 19975
rect 25605 19941 25639 19975
rect 29285 19941 29319 19975
rect 31401 19941 31435 19975
rect 34161 19941 34195 19975
rect 36277 19941 36311 19975
rect 37841 19941 37875 19975
rect 37933 19941 37967 19975
rect 41797 19941 41831 19975
rect 43545 19941 43579 19975
rect 43637 19941 43671 19975
rect 45155 19941 45189 19975
rect 3040 19873 3074 19907
rect 8125 19873 8159 19907
rect 9689 19873 9723 19907
rect 10952 19873 10986 19907
rect 11897 19873 11931 19907
rect 12357 19873 12391 19907
rect 13001 19873 13035 19907
rect 13461 19873 13495 19907
rect 21005 19873 21039 19907
rect 22753 19873 22787 19907
rect 23305 19873 23339 19907
rect 25329 19873 25363 19907
rect 26709 19873 26743 19907
rect 27997 19873 28031 19907
rect 28089 19873 28123 19907
rect 28365 19873 28399 19907
rect 29432 19873 29466 19907
rect 30916 19873 30950 19907
rect 33149 19873 33183 19907
rect 39313 19873 39347 19907
rect 39773 19873 39807 19907
rect 45017 19873 45051 19907
rect 4353 19805 4387 19839
rect 6653 19805 6687 19839
rect 7297 19805 7331 19839
rect 16129 19805 16163 19839
rect 17233 19805 17267 19839
rect 18797 19805 18831 19839
rect 19073 19805 19107 19839
rect 23121 19805 23155 19839
rect 29653 19805 29687 19839
rect 30297 19805 30331 19839
rect 32229 19805 32263 19839
rect 34069 19805 34103 19839
rect 36185 19805 36219 19839
rect 36829 19805 36863 19839
rect 38117 19805 38151 19839
rect 40049 19805 40083 19839
rect 41705 19805 41739 19839
rect 41981 19805 42015 19839
rect 43821 19805 43855 19839
rect 3111 19737 3145 19771
rect 9873 19737 9907 19771
rect 17785 19737 17819 19771
rect 24777 19737 24811 19771
rect 29929 19737 29963 19771
rect 34621 19737 34655 19771
rect 5273 19669 5307 19703
rect 6377 19669 6411 19703
rect 10149 19669 10183 19703
rect 11023 19669 11057 19703
rect 19717 19669 19751 19703
rect 21189 19669 21223 19703
rect 24317 19669 24351 19703
rect 25881 19669 25915 19703
rect 26893 19669 26927 19703
rect 29101 19669 29135 19703
rect 29561 19669 29595 19703
rect 30987 19669 31021 19703
rect 35081 19669 35115 19703
rect 40509 19669 40543 19703
rect 3801 19465 3835 19499
rect 5549 19465 5583 19499
rect 6285 19465 6319 19499
rect 7941 19465 7975 19499
rect 9689 19465 9723 19499
rect 11529 19465 11563 19499
rect 13461 19465 13495 19499
rect 13921 19465 13955 19499
rect 15117 19465 15151 19499
rect 16589 19465 16623 19499
rect 17233 19465 17267 19499
rect 17877 19465 17911 19499
rect 19073 19465 19107 19499
rect 20729 19465 20763 19499
rect 21097 19465 21131 19499
rect 22753 19465 22787 19499
rect 27353 19465 27387 19499
rect 29009 19465 29043 19499
rect 29515 19465 29549 19499
rect 29653 19465 29687 19499
rect 30849 19465 30883 19499
rect 32873 19465 32907 19499
rect 33609 19465 33643 19499
rect 36001 19465 36035 19499
rect 36277 19465 36311 19499
rect 38209 19465 38243 19499
rect 39865 19465 39899 19499
rect 41429 19465 41463 19499
rect 41797 19465 41831 19499
rect 43361 19465 43395 19499
rect 43729 19465 43763 19499
rect 4261 19397 4295 19431
rect 6653 19397 6687 19431
rect 11897 19397 11931 19431
rect 13277 19397 13311 19431
rect 15393 19397 15427 19431
rect 16221 19397 16255 19431
rect 37473 19397 37507 19431
rect 37933 19397 37967 19431
rect 44005 19397 44039 19431
rect 2697 19329 2731 19363
rect 8861 19329 8895 19363
rect 2789 19261 2823 19295
rect 3249 19261 3283 19295
rect 3525 19261 3559 19295
rect 4353 19261 4387 19295
rect 9965 19261 9999 19295
rect 10517 19261 10551 19295
rect 12173 19261 12207 19295
rect 6929 19193 6963 19227
rect 7021 19193 7055 19227
rect 7573 19193 7607 19227
rect 8493 19193 8527 19227
rect 8585 19193 8619 19227
rect 10701 19193 10735 19227
rect 12541 19193 12575 19227
rect 12633 19193 12667 19227
rect 13185 19193 13219 19227
rect 14381 19329 14415 19363
rect 15669 19329 15703 19363
rect 18797 19329 18831 19363
rect 19717 19329 19751 19363
rect 20361 19329 20395 19363
rect 21281 19329 21315 19363
rect 21557 19329 21591 19363
rect 23949 19329 23983 19363
rect 25329 19329 25363 19363
rect 29745 19329 29779 19363
rect 39589 19329 39623 19363
rect 40509 19329 40543 19363
rect 42441 19329 42475 19363
rect 24685 19261 24719 19295
rect 26341 19261 26375 19295
rect 26985 19261 27019 19295
rect 27537 19261 27571 19295
rect 29377 19261 29411 19295
rect 30389 19261 30423 19295
rect 30849 19261 30883 19295
rect 30976 19261 31010 19295
rect 31953 19261 31987 19295
rect 33768 19261 33802 19295
rect 34161 19261 34195 19295
rect 35081 19261 35115 19295
rect 38761 19261 38795 19295
rect 38853 19261 38887 19295
rect 39313 19261 39347 19295
rect 14105 19193 14139 19227
rect 14197 19193 14231 19227
rect 15761 19193 15795 19227
rect 18153 19193 18187 19227
rect 18245 19193 18279 19227
rect 19533 19193 19567 19227
rect 19809 19193 19843 19227
rect 21373 19193 21407 19227
rect 26065 19193 26099 19227
rect 26157 19193 26191 19227
rect 30113 19193 30147 19227
rect 32274 19193 32308 19227
rect 34621 19193 34655 19227
rect 35402 19193 35436 19227
rect 36921 19193 36955 19227
rect 37013 19193 37047 19227
rect 40830 19193 40864 19227
rect 42762 19193 42796 19227
rect 4721 19125 4755 19159
rect 5273 19125 5307 19159
rect 8217 19125 8251 19159
rect 11069 19125 11103 19159
rect 13277 19125 13311 19159
rect 23121 19125 23155 19159
rect 24409 19125 24443 19159
rect 25605 19125 25639 19159
rect 26433 19125 26467 19159
rect 27721 19125 27755 19159
rect 27997 19125 28031 19159
rect 28457 19125 28491 19159
rect 31079 19125 31113 19159
rect 31401 19125 31435 19159
rect 31769 19125 31803 19159
rect 33149 19125 33183 19159
rect 33839 19125 33873 19159
rect 36645 19125 36679 19159
rect 40325 19125 40359 19159
rect 42257 19125 42291 19159
rect 45017 19125 45051 19159
rect 2881 18921 2915 18955
rect 4721 18921 4755 18955
rect 6561 18921 6595 18955
rect 7205 18921 7239 18955
rect 9965 18921 9999 18955
rect 10885 18921 10919 18955
rect 12173 18921 12207 18955
rect 13553 18921 13587 18955
rect 14105 18921 14139 18955
rect 14381 18921 14415 18955
rect 16267 18921 16301 18955
rect 18153 18921 18187 18955
rect 18705 18921 18739 18955
rect 21189 18921 21223 18955
rect 21373 18921 21407 18955
rect 25605 18921 25639 18955
rect 29285 18921 29319 18955
rect 30573 18921 30607 18955
rect 31585 18921 31619 18955
rect 32229 18921 32263 18955
rect 34805 18921 34839 18955
rect 36185 18921 36219 18955
rect 38945 18921 38979 18955
rect 39313 18921 39347 18955
rect 41705 18921 41739 18955
rect 12586 18853 12620 18887
rect 15577 18853 15611 18887
rect 17233 18853 17267 18887
rect 17325 18853 17359 18887
rect 17877 18853 17911 18887
rect 19349 18853 19383 18887
rect 19441 18853 19475 18887
rect 19993 18853 20027 18887
rect 23029 18853 23063 18887
rect 28181 18853 28215 18887
rect 34437 18853 34471 18887
rect 35586 18853 35620 18887
rect 37933 18853 37967 18887
rect 40554 18853 40588 18887
rect 42441 18853 42475 18887
rect 43545 18853 43579 18887
rect 4445 18785 4479 18819
rect 5273 18785 5307 18819
rect 5733 18785 5767 18819
rect 7757 18785 7791 18819
rect 8620 18785 8654 18819
rect 13185 18785 13219 18819
rect 14197 18785 14231 18819
rect 16196 18785 16230 18819
rect 20980 18785 21014 18819
rect 22937 18785 22971 18819
rect 23397 18785 23431 18819
rect 23857 18785 23891 18819
rect 24961 18785 24995 18819
rect 25421 18785 25455 18819
rect 26617 18785 26651 18819
rect 28328 18785 28362 18819
rect 29812 18785 29846 18819
rect 31033 18785 31067 18819
rect 32413 18785 32447 18819
rect 32597 18785 32631 18819
rect 33701 18785 33735 18819
rect 34253 18785 34287 18819
rect 36461 18785 36495 18819
rect 41981 18785 42015 18819
rect 6009 18717 6043 18751
rect 6837 18717 6871 18751
rect 10517 18717 10551 18751
rect 12265 18717 12299 18751
rect 24225 18717 24259 18751
rect 26985 18717 27019 18751
rect 27721 18717 27755 18751
rect 28549 18717 28583 18751
rect 28917 18717 28951 18751
rect 33333 18717 33367 18751
rect 35265 18717 35299 18751
rect 37841 18717 37875 18751
rect 40233 18717 40267 18751
rect 43453 18717 43487 18751
rect 43729 18717 43763 18751
rect 24022 18649 24056 18683
rect 26341 18649 26375 18683
rect 26782 18649 26816 18683
rect 31171 18649 31205 18683
rect 36921 18649 36955 18683
rect 38393 18649 38427 18683
rect 41153 18649 41187 18683
rect 8401 18581 8435 18615
rect 8723 18581 8757 18615
rect 11437 18581 11471 18615
rect 16037 18581 16071 18615
rect 16957 18581 16991 18615
rect 23765 18581 23799 18615
rect 24133 18581 24167 18615
rect 24317 18581 24351 18615
rect 25237 18581 25271 18615
rect 26893 18581 26927 18615
rect 27077 18581 27111 18615
rect 28089 18581 28123 18615
rect 28457 18581 28491 18615
rect 29883 18581 29917 18615
rect 30205 18581 30239 18615
rect 31953 18581 31987 18615
rect 35173 18581 35207 18615
rect 40049 18581 40083 18615
rect 42165 18581 42199 18615
rect 5273 18377 5307 18411
rect 5871 18377 5905 18411
rect 7389 18377 7423 18411
rect 9597 18377 9631 18411
rect 11253 18377 11287 18411
rect 13461 18377 13495 18411
rect 13829 18377 13863 18411
rect 15761 18377 15795 18411
rect 17325 18377 17359 18411
rect 19441 18377 19475 18411
rect 19809 18377 19843 18411
rect 24133 18377 24167 18411
rect 26341 18377 26375 18411
rect 27077 18377 27111 18411
rect 27905 18377 27939 18411
rect 29450 18377 29484 18411
rect 34253 18377 34287 18411
rect 35357 18377 35391 18411
rect 36461 18377 36495 18411
rect 37105 18377 37139 18411
rect 41981 18377 42015 18411
rect 43453 18377 43487 18411
rect 4997 18309 5031 18343
rect 7941 18309 7975 18343
rect 23949 18309 23983 18343
rect 25513 18309 25547 18343
rect 28641 18309 28675 18343
rect 29009 18309 29043 18343
rect 29561 18309 29595 18343
rect 31125 18309 31159 18343
rect 41429 18309 41463 18343
rect 43821 18309 43855 18343
rect 4537 18241 4571 18275
rect 8217 18241 8251 18275
rect 8861 18241 8895 18275
rect 9229 18241 9263 18275
rect 11483 18241 11517 18275
rect 20177 18241 20211 18275
rect 21741 18241 21775 18275
rect 23489 18241 23523 18275
rect 24041 18241 24075 18275
rect 25605 18241 25639 18275
rect 27997 18241 28031 18275
rect 29653 18241 29687 18275
rect 31953 18241 31987 18275
rect 38393 18241 38427 18275
rect 39589 18241 39623 18275
rect 42993 18241 43027 18275
rect 3709 18173 3743 18207
rect 4077 18173 4111 18207
rect 4353 18173 4387 18207
rect 5768 18173 5802 18207
rect 6193 18173 6227 18207
rect 9781 18173 9815 18207
rect 10241 18173 10275 18207
rect 11380 18173 11414 18207
rect 11897 18173 11931 18207
rect 12633 18173 12667 18207
rect 12909 18173 12943 18207
rect 14381 18173 14415 18207
rect 14933 18173 14967 18207
rect 15945 18173 15979 18207
rect 16405 18173 16439 18207
rect 18337 18173 18371 18207
rect 19625 18173 19659 18207
rect 20729 18173 20763 18207
rect 22236 18173 22270 18207
rect 23820 18173 23854 18207
rect 25237 18173 25271 18207
rect 25384 18173 25418 18207
rect 27776 18173 27810 18207
rect 29285 18173 29319 18207
rect 30665 18173 30699 18207
rect 31401 18173 31435 18207
rect 31861 18173 31895 18207
rect 33241 18173 33275 18207
rect 33793 18173 33827 18207
rect 33977 18173 34011 18207
rect 35541 18173 35575 18207
rect 36737 18173 36771 18207
rect 37340 18173 37374 18207
rect 38853 18173 38887 18207
rect 39313 18173 39347 18207
rect 40509 18173 40543 18207
rect 8309 18105 8343 18139
rect 10425 18105 10459 18139
rect 13185 18105 13219 18139
rect 15117 18105 15151 18139
rect 17785 18105 17819 18139
rect 18153 18105 18187 18139
rect 20637 18105 20671 18139
rect 23673 18105 23707 18139
rect 27629 18105 27663 18139
rect 28365 18105 28399 18139
rect 33057 18105 33091 18139
rect 35862 18105 35896 18139
rect 37427 18105 37461 18139
rect 40830 18105 40864 18139
rect 42349 18105 42383 18139
rect 42441 18105 42475 18139
rect 7113 18037 7147 18071
rect 10701 18037 10735 18071
rect 12173 18037 12207 18071
rect 14289 18037 14323 18071
rect 16221 18037 16255 18071
rect 16957 18037 16991 18071
rect 18429 18037 18463 18071
rect 18981 18037 19015 18071
rect 20453 18037 20487 18071
rect 22017 18037 22051 18071
rect 22339 18037 22373 18071
rect 22753 18037 22787 18071
rect 23121 18037 23155 18071
rect 24777 18037 24811 18071
rect 25053 18037 25087 18071
rect 25881 18037 25915 18071
rect 26617 18037 26651 18071
rect 27445 18037 27479 18071
rect 29929 18037 29963 18071
rect 30297 18037 30331 18071
rect 32505 18037 32539 18071
rect 34713 18037 34747 18071
rect 37749 18037 37783 18071
rect 38669 18037 38703 18071
rect 39865 18037 39899 18071
rect 40233 18037 40267 18071
rect 3801 17833 3835 17867
rect 4169 17833 4203 17867
rect 5779 17833 5813 17867
rect 8217 17833 8251 17867
rect 8585 17833 8619 17867
rect 9781 17833 9815 17867
rect 10701 17833 10735 17867
rect 11805 17833 11839 17867
rect 14657 17833 14691 17867
rect 15669 17833 15703 17867
rect 17509 17833 17543 17867
rect 18337 17833 18371 17867
rect 19349 17833 19383 17867
rect 19717 17833 19751 17867
rect 22845 17833 22879 17867
rect 24685 17833 24719 17867
rect 25329 17833 25363 17867
rect 25881 17833 25915 17867
rect 27721 17833 27755 17867
rect 29377 17833 29411 17867
rect 31033 17833 31067 17867
rect 31493 17833 31527 17867
rect 31861 17833 31895 17867
rect 32781 17833 32815 17867
rect 35173 17833 35207 17867
rect 35909 17833 35943 17867
rect 37933 17833 37967 17867
rect 40417 17833 40451 17867
rect 41153 17833 41187 17867
rect 42625 17833 42659 17867
rect 21097 17765 21131 17799
rect 27077 17765 27111 17799
rect 28733 17765 28767 17799
rect 4077 17697 4111 17731
rect 4629 17697 4663 17731
rect 5676 17697 5710 17731
rect 7389 17697 7423 17731
rect 7573 17697 7607 17731
rect 9965 17697 9999 17731
rect 10149 17697 10183 17731
rect 11989 17697 12023 17731
rect 12173 17697 12207 17731
rect 12725 17697 12759 17731
rect 13553 17697 13587 17731
rect 14105 17697 14139 17731
rect 17049 17697 17083 17731
rect 18061 17697 18095 17731
rect 18245 17697 18279 17731
rect 19441 17697 19475 17731
rect 19625 17697 19659 17731
rect 22661 17697 22695 17731
rect 23581 17697 23615 17731
rect 23673 17697 23707 17731
rect 25421 17697 25455 17731
rect 26525 17697 26559 17731
rect 26709 17697 26743 17731
rect 28089 17697 28123 17731
rect 29653 17697 29687 17731
rect 30021 17697 30055 17731
rect 32321 17697 32355 17731
rect 33609 17697 33643 17731
rect 33793 17697 33827 17731
rect 35173 17697 35207 17731
rect 35449 17697 35483 17731
rect 36496 17697 36530 17731
rect 38577 17697 38611 17731
rect 39129 17697 39163 17731
rect 40141 17697 40175 17731
rect 40601 17697 40635 17731
rect 41772 17697 41806 17731
rect 42349 17697 42383 17731
rect 7021 17629 7055 17663
rect 7757 17629 7791 17663
rect 14289 17629 14323 17663
rect 15301 17629 15335 17663
rect 21005 17629 21039 17663
rect 21281 17629 21315 17663
rect 23213 17629 23247 17663
rect 24041 17629 24075 17663
rect 30297 17629 30331 17663
rect 30573 17629 30607 17663
rect 34069 17629 34103 17663
rect 39313 17629 39347 17663
rect 17233 17561 17267 17595
rect 24133 17561 24167 17595
rect 25605 17561 25639 17595
rect 26249 17561 26283 17595
rect 16221 17493 16255 17527
rect 23820 17493 23854 17527
rect 23949 17493 23983 17527
rect 32505 17493 32539 17527
rect 36599 17493 36633 17527
rect 36921 17493 36955 17527
rect 41843 17493 41877 17527
rect 3617 17289 3651 17323
rect 3985 17289 4019 17323
rect 5549 17289 5583 17323
rect 7941 17289 7975 17323
rect 10333 17289 10367 17323
rect 11437 17289 11471 17323
rect 13553 17289 13587 17323
rect 14197 17289 14231 17323
rect 16405 17289 16439 17323
rect 16865 17289 16899 17323
rect 19349 17289 19383 17323
rect 21465 17289 21499 17323
rect 23489 17289 23523 17323
rect 24593 17289 24627 17323
rect 25513 17289 25547 17323
rect 26249 17289 26283 17323
rect 28641 17289 28675 17323
rect 29101 17289 29135 17323
rect 33333 17289 33367 17323
rect 34713 17289 34747 17323
rect 35173 17289 35207 17323
rect 42349 17289 42383 17323
rect 11805 17221 11839 17255
rect 19579 17221 19613 17255
rect 21833 17221 21867 17255
rect 23949 17221 23983 17255
rect 32873 17221 32907 17255
rect 33057 17221 33091 17255
rect 36277 17221 36311 17255
rect 37841 17221 37875 17255
rect 39037 17221 39071 17255
rect 39773 17221 39807 17255
rect 40141 17221 40175 17255
rect 6653 17153 6687 17187
rect 15209 17153 15243 17187
rect 20545 17153 20579 17187
rect 21189 17153 21223 17187
rect 30113 17153 30147 17187
rect 31953 17153 31987 17187
rect 35587 17153 35621 17187
rect 36553 17153 36587 17187
rect 38485 17153 38519 17187
rect 4169 17085 4203 17119
rect 4629 17085 4663 17119
rect 5181 17085 5215 17119
rect 5733 17085 5767 17119
rect 7205 17085 7239 17119
rect 7481 17085 7515 17119
rect 9229 17085 9263 17119
rect 9597 17085 9631 17119
rect 9873 17085 9907 17119
rect 10793 17085 10827 17119
rect 10920 17085 10954 17119
rect 12173 17085 12207 17119
rect 12449 17085 12483 17119
rect 12909 17085 12943 17119
rect 14013 17085 14047 17119
rect 16957 17085 16991 17119
rect 18061 17085 18095 17119
rect 18245 17085 18279 17119
rect 19508 17085 19542 17119
rect 22344 17085 22378 17119
rect 22845 17085 22879 17119
rect 24501 17085 24535 17119
rect 25145 17085 25179 17119
rect 26617 17085 26651 17119
rect 26893 17085 26927 17119
rect 28181 17085 28215 17119
rect 33057 17085 33091 17119
rect 33476 17085 33510 17119
rect 40576 17085 40610 17119
rect 41556 17085 41590 17119
rect 41981 17085 42015 17119
rect 43152 17085 43186 17119
rect 43545 17085 43579 17119
rect 4905 17017 4939 17051
rect 6285 17017 6319 17051
rect 7665 17017 7699 17051
rect 8861 17017 8895 17051
rect 15530 17017 15564 17051
rect 20637 17017 20671 17051
rect 22431 17017 22465 17051
rect 24317 17017 24351 17051
rect 27445 17017 27479 17051
rect 30434 17017 30468 17051
rect 32045 17017 32079 17051
rect 32597 17017 32631 17051
rect 33563 17017 33597 17051
rect 35357 17017 35391 17051
rect 36001 17017 36035 17051
rect 36645 17017 36679 17051
rect 37197 17017 37231 17051
rect 38117 17017 38151 17051
rect 38209 17017 38243 17051
rect 41659 17017 41693 17051
rect 3249 16949 3283 16983
rect 5917 16949 5951 16983
rect 9597 16949 9631 16983
rect 11023 16949 11057 16983
rect 12541 16949 12575 16983
rect 14657 16949 14691 16983
rect 15025 16949 15059 16983
rect 16129 16949 16163 16983
rect 17141 16949 17175 16983
rect 17509 16949 17543 16983
rect 17877 16949 17911 16983
rect 18337 16949 18371 16983
rect 18889 16949 18923 16983
rect 19901 16949 19935 16983
rect 20361 16949 20395 16983
rect 26433 16949 26467 16983
rect 27997 16949 28031 16983
rect 28365 16949 28399 16983
rect 29653 16949 29687 16983
rect 30021 16949 30055 16983
rect 31033 16949 31067 16983
rect 31677 16949 31711 16983
rect 33977 16949 34011 16983
rect 37473 16949 37507 16983
rect 39497 16949 39531 16983
rect 40647 16949 40681 16983
rect 40969 16949 41003 16983
rect 43223 16949 43257 16983
rect 7573 16745 7607 16779
rect 9413 16745 9447 16779
rect 10793 16745 10827 16779
rect 12173 16745 12207 16779
rect 13001 16745 13035 16779
rect 13553 16745 13587 16779
rect 15945 16745 15979 16779
rect 18153 16745 18187 16779
rect 19441 16745 19475 16779
rect 20545 16745 20579 16779
rect 21189 16745 21223 16779
rect 22753 16745 22787 16779
rect 26617 16745 26651 16779
rect 27629 16745 27663 16779
rect 28273 16745 28307 16779
rect 29377 16745 29411 16779
rect 29745 16745 29779 16779
rect 31401 16745 31435 16779
rect 31953 16745 31987 16779
rect 33425 16745 33459 16779
rect 34345 16745 34379 16779
rect 40325 16745 40359 16779
rect 45063 16745 45097 16779
rect 8027 16677 8061 16711
rect 10235 16677 10269 16711
rect 17509 16677 17543 16711
rect 18337 16677 18371 16711
rect 23213 16677 23247 16711
rect 26249 16677 26283 16711
rect 30526 16677 30560 16711
rect 32229 16677 32263 16711
rect 32321 16677 32355 16711
rect 36087 16677 36121 16711
rect 37841 16677 37875 16711
rect 37933 16677 37967 16711
rect 38485 16677 38519 16711
rect 40693 16677 40727 16711
rect 40877 16677 40911 16711
rect 40969 16677 41003 16711
rect 43453 16677 43487 16711
rect 43545 16677 43579 16711
rect 2697 16609 2731 16643
rect 2973 16609 3007 16643
rect 4077 16609 4111 16643
rect 4629 16609 4663 16643
rect 5641 16609 5675 16643
rect 6101 16609 6135 16643
rect 7205 16609 7239 16643
rect 7665 16609 7699 16643
rect 9873 16609 9907 16643
rect 11805 16609 11839 16643
rect 14264 16609 14298 16643
rect 15552 16609 15586 16643
rect 16957 16609 16991 16643
rect 17141 16609 17175 16643
rect 18521 16609 18555 16643
rect 21557 16609 21591 16643
rect 24501 16609 24535 16643
rect 26801 16609 26835 16643
rect 27077 16609 27111 16643
rect 28825 16609 28859 16643
rect 35725 16609 35759 16643
rect 39313 16609 39347 16643
rect 44925 16609 44959 16643
rect 3157 16541 3191 16575
rect 4813 16541 4847 16575
rect 6377 16541 6411 16575
rect 14105 16541 14139 16575
rect 19901 16541 19935 16575
rect 23121 16541 23155 16575
rect 24731 16541 24765 16575
rect 25973 16541 26007 16575
rect 30205 16541 30239 16575
rect 32505 16541 32539 16575
rect 33977 16541 34011 16575
rect 43729 16541 43763 16575
rect 23673 16473 23707 16507
rect 24409 16473 24443 16507
rect 41429 16473 41463 16507
rect 8585 16405 8619 16439
rect 12725 16405 12759 16439
rect 14335 16405 14369 16439
rect 15623 16405 15657 16439
rect 22109 16405 22143 16439
rect 29009 16405 29043 16439
rect 31125 16405 31159 16439
rect 34897 16405 34931 16439
rect 36645 16405 36679 16439
rect 36921 16405 36955 16439
rect 39497 16405 39531 16439
rect 2513 16201 2547 16235
rect 2881 16201 2915 16235
rect 3709 16201 3743 16235
rect 4077 16201 4111 16235
rect 5917 16201 5951 16235
rect 6285 16201 6319 16235
rect 7113 16201 7147 16235
rect 13829 16201 13863 16235
rect 15577 16201 15611 16235
rect 17141 16201 17175 16235
rect 21097 16201 21131 16235
rect 23121 16201 23155 16235
rect 23305 16201 23339 16235
rect 27261 16201 27295 16235
rect 29009 16201 29043 16235
rect 31217 16201 31251 16235
rect 32413 16201 32447 16235
rect 33149 16201 33183 16235
rect 35265 16201 35299 16235
rect 38393 16201 38427 16235
rect 38485 16201 38519 16235
rect 39865 16201 39899 16235
rect 17877 16133 17911 16167
rect 22661 16133 22695 16167
rect 24685 16133 24719 16167
rect 7573 16065 7607 16099
rect 9597 16065 9631 16099
rect 10793 16065 10827 16099
rect 12449 16065 12483 16099
rect 14289 16065 14323 16099
rect 17509 16065 17543 16099
rect 18429 16065 18463 16099
rect 19717 16065 19751 16099
rect 23305 16065 23339 16099
rect 25973 16065 26007 16099
rect 28641 16065 28675 16099
rect 30021 16065 30055 16099
rect 30665 16065 30699 16099
rect 31493 16065 31527 16099
rect 32137 16065 32171 16099
rect 33977 16065 34011 16099
rect 34621 16065 34655 16099
rect 36369 16065 36403 16099
rect 37197 16065 37231 16099
rect 4721 15997 4755 16031
rect 10517 15997 10551 16031
rect 11161 15997 11195 16031
rect 11380 15997 11414 16031
rect 16865 15997 16899 16031
rect 16957 15997 16991 16031
rect 18981 15997 19015 16031
rect 20177 15997 20211 16031
rect 20637 15997 20671 16031
rect 27537 15997 27571 16031
rect 28216 15997 28250 16031
rect 29285 15997 29319 16031
rect 29745 15997 29779 16031
rect 33517 15997 33551 16031
rect 33701 15997 33735 16031
rect 35500 15997 35534 16031
rect 38209 15997 38243 16031
rect 41337 16133 41371 16167
rect 40785 16065 40819 16099
rect 42257 16065 42291 16099
rect 44097 16065 44131 16099
rect 44373 16065 44407 16099
rect 38669 15997 38703 16031
rect 39589 15997 39623 16031
rect 40233 15997 40267 16031
rect 7481 15929 7515 15963
rect 7935 15929 7969 15963
rect 9137 15929 9171 15963
rect 9505 15929 9539 15963
rect 9918 15929 9952 15963
rect 11897 15929 11931 15963
rect 12173 15929 12207 15963
rect 12811 15929 12845 15963
rect 14105 15929 14139 15963
rect 14610 15929 14644 15963
rect 18797 15929 18831 15963
rect 22109 15929 22143 15963
rect 22201 15929 22235 15963
rect 23489 15929 23523 15963
rect 23765 15929 23799 15963
rect 23857 15929 23891 15963
rect 24409 15929 24443 15963
rect 25881 15929 25915 15963
rect 26294 15929 26328 15963
rect 28319 15929 28353 15963
rect 31585 15929 31619 15963
rect 34253 15929 34287 15963
rect 35587 15929 35621 15963
rect 36553 15929 36587 15963
rect 36645 15929 36679 15963
rect 38393 15929 38427 15963
rect 39031 15929 39065 15963
rect 40877 15929 40911 15963
rect 44189 15929 44223 15963
rect 4629 15861 4663 15895
rect 5089 15861 5123 15895
rect 5641 15861 5675 15895
rect 8493 15861 8527 15895
rect 11483 15861 11517 15895
rect 13369 15861 13403 15895
rect 15209 15861 15243 15895
rect 19073 15861 19107 15895
rect 20361 15861 20395 15895
rect 21925 15861 21959 15895
rect 26893 15861 26927 15895
rect 30297 15861 30331 15895
rect 35909 15861 35943 15895
rect 37473 15861 37507 15895
rect 41705 15861 41739 15895
rect 42165 15861 42199 15895
rect 42625 15861 42659 15895
rect 43177 15861 43211 15895
rect 43545 15861 43579 15895
rect 43821 15861 43855 15895
rect 45017 15861 45051 15895
rect 5089 15657 5123 15691
rect 7665 15657 7699 15691
rect 9505 15657 9539 15691
rect 10793 15657 10827 15691
rect 11805 15657 11839 15691
rect 12909 15657 12943 15691
rect 14289 15657 14323 15691
rect 22569 15657 22603 15691
rect 23765 15657 23799 15691
rect 26065 15657 26099 15691
rect 28917 15657 28951 15691
rect 31953 15657 31987 15691
rect 35311 15657 35345 15691
rect 37013 15657 37047 15691
rect 37473 15657 37507 15691
rect 37933 15657 37967 15691
rect 38577 15657 38611 15691
rect 42257 15657 42291 15691
rect 43177 15657 43211 15691
rect 44373 15657 44407 15691
rect 6739 15589 6773 15623
rect 9873 15589 9907 15623
rect 13455 15589 13489 15623
rect 15853 15589 15887 15623
rect 15945 15589 15979 15623
rect 17969 15589 18003 15623
rect 19901 15589 19935 15623
rect 22845 15589 22879 15623
rect 24317 15589 24351 15623
rect 24409 15589 24443 15623
rect 26846 15589 26880 15623
rect 29285 15589 29319 15623
rect 32321 15589 32355 15623
rect 32873 15589 32907 15623
rect 41061 15589 41095 15623
rect 43545 15589 43579 15623
rect 4077 15521 4111 15555
rect 4537 15521 4571 15555
rect 6377 15521 6411 15555
rect 8192 15521 8226 15555
rect 12148 15521 12182 15555
rect 13093 15521 13127 15555
rect 18153 15521 18187 15555
rect 18797 15521 18831 15555
rect 19349 15521 19383 15555
rect 19533 15521 19567 15555
rect 21649 15521 21683 15555
rect 26525 15521 26559 15555
rect 31068 15521 31102 15555
rect 34161 15521 34195 15555
rect 35081 15521 35115 15555
rect 36185 15521 36219 15555
rect 38301 15521 38335 15555
rect 38761 15521 38795 15555
rect 39865 15521 39899 15555
rect 44960 15521 44994 15555
rect 4629 15453 4663 15487
rect 9781 15453 9815 15487
rect 10057 15453 10091 15487
rect 16129 15453 16163 15487
rect 22753 15453 22787 15487
rect 23397 15453 23431 15487
rect 24593 15453 24627 15487
rect 29193 15453 29227 15487
rect 32229 15453 32263 15487
rect 33333 15453 33367 15487
rect 40969 15453 41003 15487
rect 43453 15453 43487 15487
rect 45063 15453 45097 15487
rect 8263 15385 8297 15419
rect 29745 15385 29779 15419
rect 41521 15385 41555 15419
rect 44005 15385 44039 15419
rect 7297 15317 7331 15351
rect 8861 15317 8895 15351
rect 12219 15317 12253 15351
rect 12541 15317 12575 15351
rect 14013 15317 14047 15351
rect 18245 15317 18279 15351
rect 21787 15317 21821 15351
rect 25237 15317 25271 15351
rect 27445 15317 27479 15351
rect 31171 15317 31205 15351
rect 34299 15317 34333 15351
rect 34989 15317 35023 15351
rect 36323 15317 36357 15351
rect 36645 15317 36679 15351
rect 40049 15317 40083 15351
rect 40601 15317 40635 15351
rect 3617 15113 3651 15147
rect 3893 15113 3927 15147
rect 6101 15113 6135 15147
rect 8217 15113 8251 15147
rect 10149 15113 10183 15147
rect 11897 15113 11931 15147
rect 13829 15113 13863 15147
rect 17877 15113 17911 15147
rect 18613 15113 18647 15147
rect 19349 15113 19383 15147
rect 22293 15113 22327 15147
rect 23949 15113 23983 15147
rect 27721 15113 27755 15147
rect 28365 15113 28399 15147
rect 31033 15113 31067 15147
rect 31861 15113 31895 15147
rect 32229 15113 32263 15147
rect 33241 15113 33275 15147
rect 37933 15113 37967 15147
rect 39865 15113 39899 15147
rect 40325 15113 40359 15147
rect 42993 15113 43027 15147
rect 43269 15113 43303 15147
rect 44465 15113 44499 15147
rect 9689 15045 9723 15079
rect 18245 15045 18279 15079
rect 22523 15045 22557 15079
rect 26249 15045 26283 15079
rect 28733 15045 28767 15079
rect 34621 15045 34655 15079
rect 36277 15045 36311 15079
rect 37473 15045 37507 15079
rect 38209 15045 38243 15079
rect 4445 14977 4479 15011
rect 5641 14977 5675 15011
rect 6469 14977 6503 15011
rect 9505 14977 9539 15011
rect 6872 14909 6906 14943
rect 7297 14909 7331 14943
rect 4353 14841 4387 14875
rect 4807 14841 4841 14875
rect 8861 14841 8895 14875
rect 8953 14841 8987 14875
rect 10793 14977 10827 15011
rect 11161 14977 11195 15011
rect 12541 14977 12575 15011
rect 12817 14977 12851 15011
rect 15117 14977 15151 15011
rect 16405 14977 16439 15011
rect 16681 14977 16715 15011
rect 19073 14977 19107 15011
rect 23305 14977 23339 15011
rect 23397 14977 23431 15011
rect 25237 14977 25271 15011
rect 25881 14977 25915 15011
rect 27077 14977 27111 15011
rect 35265 14977 35299 15011
rect 36553 14977 36587 15011
rect 36829 14977 36863 15011
rect 38577 14977 38611 15011
rect 40601 14977 40635 15011
rect 42211 14977 42245 15011
rect 18061 14909 18095 14943
rect 19901 14909 19935 14943
rect 22452 14909 22486 14943
rect 22937 14909 22971 14943
rect 10885 14841 10919 14875
rect 12265 14841 12299 14875
rect 12633 14841 12667 14875
rect 14841 14841 14875 14875
rect 14933 14841 14967 14875
rect 16221 14841 16255 14875
rect 16497 14841 16531 14875
rect 19809 14841 19843 14875
rect 20222 14841 20256 14875
rect 23740 14909 23774 14943
rect 24133 14909 24167 14943
rect 29285 14909 29319 14943
rect 30481 14909 30515 14943
rect 31452 14909 31486 14943
rect 32448 14909 32482 14943
rect 32873 14909 32907 14943
rect 33425 14909 33459 14943
rect 38761 14909 38795 14943
rect 39313 14909 39347 14943
rect 42124 14909 42158 14943
rect 42533 14909 42567 14943
rect 45084 14909 45118 14943
rect 45477 14909 45511 14943
rect 24593 14841 24627 14875
rect 25053 14841 25087 14875
rect 25329 14841 25363 14875
rect 26801 14841 26835 14875
rect 26893 14841 26927 14875
rect 29606 14841 29640 14875
rect 31539 14841 31573 14875
rect 34989 14841 35023 14875
rect 35081 14841 35115 14875
rect 36645 14841 36679 14875
rect 39497 14841 39531 14875
rect 40693 14841 40727 14875
rect 41245 14841 41279 14875
rect 43545 14841 43579 14875
rect 43637 14841 43671 14875
rect 44189 14841 44223 14875
rect 44833 14841 44867 14875
rect 5365 14773 5399 14807
rect 7113 14773 7147 14807
rect 8585 14773 8619 14807
rect 9689 14773 9723 14807
rect 9873 14773 9907 14807
rect 10517 14773 10551 14807
rect 13553 14773 13587 14807
rect 14657 14773 14691 14807
rect 15853 14773 15887 14807
rect 20821 14773 20855 14807
rect 21741 14773 21775 14807
rect 23397 14773 23431 14807
rect 26525 14773 26559 14807
rect 29009 14773 29043 14807
rect 30205 14773 30239 14807
rect 32551 14773 32585 14807
rect 33609 14773 33643 14807
rect 34161 14773 34195 14807
rect 41521 14773 41555 14807
rect 45155 14773 45189 14807
rect 14841 14569 14875 14603
rect 15439 14569 15473 14603
rect 15853 14569 15887 14603
rect 16405 14569 16439 14603
rect 18153 14569 18187 14603
rect 24225 14569 24259 14603
rect 25007 14569 25041 14603
rect 31171 14569 31205 14603
rect 34069 14569 34103 14603
rect 39129 14569 39163 14603
rect 43913 14569 43947 14603
rect 4807 14501 4841 14535
rect 7021 14501 7055 14535
rect 10517 14501 10551 14535
rect 10609 14501 10643 14535
rect 11161 14501 11195 14535
rect 12173 14501 12207 14535
rect 12265 14501 12299 14535
rect 13829 14501 13863 14535
rect 14381 14501 14415 14535
rect 16865 14501 16899 14535
rect 19809 14501 19843 14535
rect 20085 14501 20119 14535
rect 21097 14501 21131 14535
rect 22753 14501 22787 14535
rect 22845 14501 22879 14535
rect 23397 14501 23431 14535
rect 28273 14501 28307 14535
rect 29285 14501 29319 14535
rect 31493 14501 31527 14535
rect 32229 14501 32263 14535
rect 32321 14501 32355 14535
rect 34345 14501 34379 14535
rect 34437 14501 34471 14535
rect 34989 14501 35023 14535
rect 36277 14501 36311 14535
rect 36829 14501 36863 14535
rect 39951 14501 39985 14535
rect 41705 14501 41739 14535
rect 42257 14501 42291 14535
rect 4445 14433 4479 14467
rect 8436 14433 8470 14467
rect 8861 14433 8895 14467
rect 15336 14433 15370 14467
rect 17233 14433 17267 14467
rect 19073 14433 19107 14467
rect 19625 14433 19659 14467
rect 24936 14433 24970 14467
rect 26433 14433 26467 14467
rect 26663 14433 26697 14467
rect 27353 14433 27387 14467
rect 27537 14433 27571 14467
rect 28089 14433 28123 14467
rect 31100 14433 31134 14467
rect 31953 14433 31987 14467
rect 38715 14433 38749 14467
rect 40877 14433 40911 14467
rect 43428 14433 43462 14467
rect 6929 14365 6963 14399
rect 12449 14365 12483 14399
rect 13737 14365 13771 14399
rect 21005 14365 21039 14399
rect 29193 14365 29227 14399
rect 29837 14365 29871 14399
rect 32505 14365 32539 14399
rect 35265 14365 35299 14399
rect 36185 14365 36219 14399
rect 7481 14297 7515 14331
rect 10057 14297 10091 14331
rect 21557 14297 21591 14331
rect 39589 14365 39623 14399
rect 41613 14365 41647 14399
rect 5365 14229 5399 14263
rect 8539 14229 8573 14263
rect 25329 14229 25363 14263
rect 26985 14229 27019 14263
rect 38485 14229 38519 14263
rect 40509 14229 40543 14263
rect 41337 14229 41371 14263
rect 43499 14229 43533 14263
rect 3709 14025 3743 14059
rect 4077 14025 4111 14059
rect 7849 14025 7883 14059
rect 11161 14025 11195 14059
rect 12173 14025 12207 14059
rect 12725 14025 12759 14059
rect 13369 14025 13403 14059
rect 13599 14025 13633 14059
rect 13921 14025 13955 14059
rect 14289 14025 14323 14059
rect 15853 14025 15887 14059
rect 20085 14025 20119 14059
rect 21373 14025 21407 14059
rect 22385 14025 22419 14059
rect 23121 14025 23155 14059
rect 23489 14025 23523 14059
rect 24961 14025 24995 14059
rect 26433 14025 26467 14059
rect 27629 14025 27663 14059
rect 28089 14025 28123 14059
rect 30665 14025 30699 14059
rect 32505 14025 32539 14059
rect 32873 14025 32907 14059
rect 34345 14025 34379 14059
rect 36093 14025 36127 14059
rect 37657 14025 37691 14059
rect 38117 14025 38151 14059
rect 39221 14025 39255 14059
rect 39957 14025 39991 14059
rect 40647 14025 40681 14059
rect 42993 14025 43027 14059
rect 7481 13957 7515 13991
rect 12909 13957 12943 13991
rect 20683 13957 20717 13991
rect 21097 13957 21131 13991
rect 29101 13957 29135 13991
rect 29929 13957 29963 13991
rect 31125 13957 31159 13991
rect 34621 13957 34655 13991
rect 39681 13957 39715 13991
rect 41429 13957 41463 13991
rect 42165 13957 42199 13991
rect 4537 13889 4571 13923
rect 6285 13889 6319 13923
rect 8217 13889 8251 13923
rect 8493 13889 8527 13923
rect 9413 13889 9447 13923
rect 10149 13889 10183 13923
rect 14933 13889 14967 13923
rect 16313 13889 16347 13923
rect 18521 13889 18555 13923
rect 22109 13889 22143 13923
rect 25145 13889 25179 13923
rect 25789 13889 25823 13923
rect 26157 13889 26191 13923
rect 28319 13889 28353 13923
rect 29377 13889 29411 13923
rect 30297 13889 30331 13923
rect 31585 13889 31619 13923
rect 31861 13889 31895 13923
rect 33425 13889 33459 13923
rect 37197 13889 37231 13923
rect 38301 13889 38335 13923
rect 38577 13889 38611 13923
rect 40969 13889 41003 13923
rect 41613 13889 41647 13923
rect 43913 13889 43947 13923
rect 4445 13821 4479 13855
rect 12516 13821 12550 13855
rect 13512 13821 13546 13855
rect 16405 13821 16439 13855
rect 17049 13821 17083 13855
rect 18981 13821 19015 13855
rect 19533 13821 19567 13855
rect 20596 13821 20630 13855
rect 21624 13821 21658 13855
rect 22636 13821 22670 13855
rect 24108 13821 24142 13855
rect 26893 13821 26927 13855
rect 27077 13821 27111 13855
rect 28232 13821 28266 13855
rect 28733 13821 28767 13855
rect 34897 13821 34931 13855
rect 40544 13821 40578 13855
rect 43120 13821 43154 13855
rect 4899 13753 4933 13787
rect 6929 13753 6963 13787
rect 7021 13753 7055 13787
rect 8585 13753 8619 13787
rect 9137 13753 9171 13787
rect 10241 13753 10275 13787
rect 10793 13753 10827 13787
rect 14749 13753 14783 13787
rect 15025 13753 15059 13787
rect 15577 13753 15611 13787
rect 18797 13753 18831 13787
rect 19717 13753 19751 13787
rect 24593 13753 24627 13787
rect 25237 13753 25271 13787
rect 29469 13753 29503 13787
rect 31677 13753 31711 13787
rect 33138 13753 33172 13787
rect 33234 13753 33268 13787
rect 35218 13753 35252 13787
rect 36737 13753 36771 13787
rect 36829 13753 36863 13787
rect 38393 13753 38427 13787
rect 41705 13753 41739 13787
rect 5457 13685 5491 13719
rect 6653 13685 6687 13719
rect 9965 13685 9999 13719
rect 17417 13685 17451 13719
rect 20361 13685 20395 13719
rect 21695 13685 21729 13719
rect 22707 13685 22741 13719
rect 24179 13685 24213 13719
rect 26709 13685 26743 13719
rect 35817 13685 35851 13719
rect 36553 13685 36587 13719
rect 42533 13685 42567 13719
rect 43223 13685 43257 13719
rect 43545 13685 43579 13719
rect 4629 13481 4663 13515
rect 5641 13481 5675 13515
rect 10517 13481 10551 13515
rect 12541 13481 12575 13515
rect 14933 13481 14967 13515
rect 24915 13481 24949 13515
rect 28871 13481 28905 13515
rect 29285 13481 29319 13515
rect 31585 13481 31619 13515
rect 31861 13481 31895 13515
rect 37105 13481 37139 13515
rect 37887 13481 37921 13515
rect 5042 13413 5076 13447
rect 7113 13413 7147 13447
rect 11253 13413 11287 13447
rect 12817 13413 12851 13447
rect 15485 13413 15519 13447
rect 19073 13413 19107 13447
rect 21189 13413 21223 13447
rect 23397 13413 23431 13447
rect 26846 13413 26880 13447
rect 32321 13413 32355 13447
rect 32873 13413 32907 13447
rect 34621 13413 34655 13447
rect 35265 13413 35299 13447
rect 36277 13413 36311 13447
rect 39910 13413 39944 13447
rect 41613 13413 41647 13447
rect 4721 13345 4755 13379
rect 8528 13345 8562 13379
rect 8953 13345 8987 13379
rect 9689 13345 9723 13379
rect 14197 13345 14231 13379
rect 18128 13345 18162 13379
rect 19257 13345 19291 13379
rect 19717 13345 19751 13379
rect 24777 13345 24811 13379
rect 26525 13345 26559 13379
rect 28641 13345 28675 13379
rect 30056 13345 30090 13379
rect 31084 13345 31118 13379
rect 33885 13345 33919 13379
rect 34345 13345 34379 13379
rect 34989 13345 35023 13379
rect 37657 13345 37691 13379
rect 43269 13345 43303 13379
rect 7021 13277 7055 13311
rect 7665 13277 7699 13311
rect 11161 13277 11195 13311
rect 11621 13277 11655 13311
rect 12725 13277 12759 13311
rect 13001 13277 13035 13311
rect 15393 13277 15427 13311
rect 15669 13277 15703 13311
rect 17049 13277 17083 13311
rect 19993 13277 20027 13311
rect 20269 13277 20303 13311
rect 21097 13277 21131 13311
rect 21557 13277 21591 13311
rect 23305 13277 23339 13311
rect 23581 13277 23615 13311
rect 30159 13277 30193 13311
rect 32229 13277 32263 13311
rect 36185 13277 36219 13311
rect 36829 13277 36863 13311
rect 39589 13277 39623 13311
rect 41521 13277 41555 13311
rect 8631 13209 8665 13243
rect 42073 13209 42107 13243
rect 6745 13141 6779 13175
rect 9873 13141 9907 13175
rect 14381 13141 14415 13175
rect 18199 13141 18233 13175
rect 18613 13141 18647 13175
rect 24225 13141 24259 13175
rect 25329 13141 25363 13175
rect 27445 13141 27479 13175
rect 29653 13141 29687 13175
rect 31171 13141 31205 13175
rect 33149 13141 33183 13175
rect 38209 13141 38243 13175
rect 40509 13141 40543 13175
rect 40785 13141 40819 13175
rect 43499 13141 43533 13175
rect 4445 12937 4479 12971
rect 5365 12937 5399 12971
rect 5687 12937 5721 12971
rect 9505 12937 9539 12971
rect 11437 12937 11471 12971
rect 11897 12937 11931 12971
rect 15301 12937 15335 12971
rect 15853 12937 15887 12971
rect 19625 12937 19659 12971
rect 20085 12937 20119 12971
rect 21373 12937 21407 12971
rect 22385 12937 22419 12971
rect 23489 12937 23523 12971
rect 27537 12937 27571 12971
rect 30573 12937 30607 12971
rect 31125 12937 31159 12971
rect 32505 12937 32539 12971
rect 32873 12937 32907 12971
rect 33701 12937 33735 12971
rect 34345 12937 34379 12971
rect 34621 12937 34655 12971
rect 36185 12937 36219 12971
rect 37841 12937 37875 12971
rect 39865 12937 39899 12971
rect 41797 12937 41831 12971
rect 42257 12937 42291 12971
rect 44097 12937 44131 12971
rect 7573 12869 7607 12903
rect 11069 12869 11103 12903
rect 21097 12869 21131 12903
rect 21741 12869 21775 12903
rect 32137 12869 32171 12903
rect 38669 12869 38703 12903
rect 4721 12801 4755 12835
rect 7021 12801 7055 12835
rect 7941 12801 7975 12835
rect 10793 12801 10827 12835
rect 12909 12801 12943 12835
rect 13829 12801 13863 12835
rect 17693 12801 17727 12835
rect 20177 12801 20211 12835
rect 23765 12801 23799 12835
rect 24409 12801 24443 12835
rect 24869 12801 24903 12835
rect 28825 12801 28859 12835
rect 29653 12801 29687 12835
rect 36645 12801 36679 12835
rect 36921 12801 36955 12835
rect 37197 12801 37231 12835
rect 39589 12801 39623 12835
rect 40233 12801 40267 12835
rect 43177 12801 43211 12835
rect 43453 12801 43487 12835
rect 5584 12733 5618 12767
rect 14749 12733 14783 12767
rect 15485 12733 15519 12767
rect 16405 12733 16439 12767
rect 16957 12733 16991 12767
rect 17141 12733 17175 12767
rect 17509 12733 17543 12767
rect 6285 12665 6319 12699
rect 6653 12665 6687 12699
rect 7113 12665 7147 12699
rect 8585 12665 8619 12699
rect 8677 12665 8711 12699
rect 9229 12665 9263 12699
rect 10149 12665 10183 12699
rect 10241 12665 10275 12699
rect 12265 12665 12299 12699
rect 13001 12665 13035 12699
rect 13553 12665 13587 12699
rect 16221 12665 16255 12699
rect 18061 12733 18095 12767
rect 19257 12733 19291 12767
rect 22636 12733 22670 12767
rect 25789 12733 25823 12767
rect 27629 12733 27663 12767
rect 28089 12733 28123 12767
rect 33844 12733 33878 12767
rect 34897 12733 34931 12767
rect 35357 12733 35391 12767
rect 38853 12733 38887 12767
rect 39313 12733 39347 12767
rect 44684 12733 44718 12767
rect 45109 12733 45143 12767
rect 20498 12665 20532 12699
rect 23857 12665 23891 12699
rect 26110 12665 26144 12699
rect 26985 12665 27019 12699
rect 28365 12665 28399 12699
rect 29745 12665 29779 12699
rect 30297 12665 30331 12699
rect 31585 12665 31619 12699
rect 31677 12665 31711 12699
rect 33931 12665 33965 12699
rect 37013 12665 37047 12699
rect 40877 12665 40911 12699
rect 40969 12665 41003 12699
rect 41521 12665 41555 12699
rect 43269 12665 43303 12699
rect 8401 12597 8435 12631
rect 9965 12597 9999 12631
rect 12633 12597 12667 12631
rect 14197 12597 14231 12631
rect 17693 12597 17727 12631
rect 17785 12597 17819 12631
rect 18429 12597 18463 12631
rect 18981 12597 19015 12631
rect 22707 12597 22741 12631
rect 23121 12597 23155 12631
rect 25605 12597 25639 12631
rect 26709 12597 26743 12631
rect 35173 12597 35207 12631
rect 42993 12597 43027 12631
rect 44787 12597 44821 12631
rect 5963 12393 5997 12427
rect 8723 12393 8757 12427
rect 10701 12393 10735 12427
rect 15117 12393 15151 12427
rect 15853 12393 15887 12427
rect 16497 12393 16531 12427
rect 19947 12393 19981 12427
rect 24317 12393 24351 12427
rect 26341 12393 26375 12427
rect 27721 12393 27755 12427
rect 29009 12393 29043 12427
rect 29561 12393 29595 12427
rect 29929 12393 29963 12427
rect 31585 12393 31619 12427
rect 35265 12393 35299 12427
rect 36185 12393 36219 12427
rect 37887 12393 37921 12427
rect 38945 12393 38979 12427
rect 40601 12393 40635 12427
rect 43177 12393 43211 12427
rect 6837 12325 6871 12359
rect 7113 12325 7147 12359
rect 7665 12325 7699 12359
rect 9045 12325 9079 12359
rect 9781 12325 9815 12359
rect 9873 12325 9907 12359
rect 12817 12325 12851 12359
rect 12909 12325 12943 12359
rect 17877 12325 17911 12359
rect 17969 12325 18003 12359
rect 20269 12325 20303 12359
rect 21097 12325 21131 12359
rect 23029 12325 23063 12359
rect 23121 12325 23155 12359
rect 23673 12325 23707 12359
rect 23949 12325 23983 12359
rect 24777 12325 24811 12359
rect 24869 12325 24903 12359
rect 25421 12325 25455 12359
rect 30573 12325 30607 12359
rect 32321 12325 32355 12359
rect 34437 12325 34471 12359
rect 34989 12325 35023 12359
rect 40002 12325 40036 12359
rect 40877 12325 40911 12359
rect 41613 12325 41647 12359
rect 43545 12325 43579 12359
rect 44097 12325 44131 12359
rect 5860 12257 5894 12291
rect 8493 12257 8527 12291
rect 15485 12257 15519 12291
rect 19844 12257 19878 12291
rect 26801 12257 26835 12291
rect 26985 12257 27019 12291
rect 31125 12257 31159 12291
rect 36645 12257 36679 12291
rect 37816 12257 37850 12291
rect 7021 12189 7055 12223
rect 10057 12189 10091 12223
rect 13461 12189 13495 12223
rect 21005 12189 21039 12223
rect 25881 12189 25915 12223
rect 27077 12189 27111 12223
rect 28641 12189 28675 12223
rect 30481 12189 30515 12223
rect 32229 12189 32263 12223
rect 32597 12189 32631 12223
rect 34345 12189 34379 12223
rect 39681 12189 39715 12223
rect 41521 12189 41555 12223
rect 41889 12189 41923 12223
rect 43453 12189 43487 12223
rect 18429 12121 18463 12155
rect 21557 12121 21591 12155
rect 41337 12121 41371 12155
rect 11621 12053 11655 12087
rect 11851 12053 11885 12087
rect 31953 12053 31987 12087
rect 36783 12053 36817 12087
rect 37105 12053 37139 12087
rect 5779 11849 5813 11883
rect 7389 11849 7423 11883
rect 8585 11849 8619 11883
rect 10057 11849 10091 11883
rect 11437 11849 11471 11883
rect 13277 11849 13311 11883
rect 14933 11849 14967 11883
rect 17877 11849 17911 11883
rect 18475 11849 18509 11883
rect 19625 11849 19659 11883
rect 20637 11849 20671 11883
rect 21005 11849 21039 11883
rect 22615 11849 22649 11883
rect 26617 11849 26651 11883
rect 30205 11849 30239 11883
rect 30573 11849 30607 11883
rect 32137 11849 32171 11883
rect 34621 11849 34655 11883
rect 38025 11849 38059 11883
rect 38669 11849 38703 11883
rect 39957 11849 39991 11883
rect 40785 11849 40819 11883
rect 42257 11849 42291 11883
rect 44465 11849 44499 11883
rect 6101 11781 6135 11815
rect 7113 11781 7147 11815
rect 11805 11781 11839 11815
rect 17509 11781 17543 11815
rect 26157 11781 26191 11815
rect 30849 11781 30883 11815
rect 36737 11781 36771 11815
rect 41889 11781 41923 11815
rect 44695 11781 44729 11815
rect 9781 11713 9815 11747
rect 12587 11713 12621 11747
rect 14289 11713 14323 11747
rect 19717 11713 19751 11747
rect 21465 11713 21499 11747
rect 24041 11713 24075 11747
rect 24317 11713 24351 11747
rect 25605 11713 25639 11747
rect 31447 11713 31481 11747
rect 32505 11713 32539 11747
rect 35265 11713 35299 11747
rect 37105 11713 37139 11747
rect 37749 11713 37783 11747
rect 39589 11713 39623 11747
rect 40233 11713 40267 11747
rect 41337 11713 41371 11747
rect 43085 11713 43119 11747
rect 43361 11713 43395 11747
rect 5676 11645 5710 11679
rect 6469 11645 6503 11679
rect 10885 11645 10919 11679
rect 12484 11645 12518 11679
rect 15577 11645 15611 11679
rect 18372 11645 18406 11679
rect 18797 11645 18831 11679
rect 22512 11645 22546 11679
rect 22937 11645 22971 11679
rect 27537 11645 27571 11679
rect 27813 11645 27847 11679
rect 28089 11645 28123 11679
rect 28365 11645 28399 11679
rect 29285 11645 29319 11679
rect 31344 11645 31378 11679
rect 31769 11645 31803 11679
rect 33241 11645 33275 11679
rect 33793 11645 33827 11679
rect 38853 11645 38887 11679
rect 39313 11645 39347 11679
rect 44592 11645 44626 11679
rect 45017 11645 45051 11679
rect 14013 11577 14047 11611
rect 14105 11577 14139 11611
rect 15485 11577 15519 11611
rect 24133 11577 24167 11611
rect 25697 11577 25731 11611
rect 27169 11577 27203 11611
rect 29606 11577 29640 11611
rect 33149 11577 33183 11611
rect 35586 11577 35620 11611
rect 37197 11577 37231 11611
rect 41429 11577 41463 11611
rect 43177 11577 43211 11611
rect 11069 11509 11103 11543
rect 12265 11509 12299 11543
rect 13001 11509 13035 11543
rect 13829 11509 13863 11543
rect 15393 11509 15427 11543
rect 19165 11509 19199 11543
rect 20085 11509 20119 11543
rect 21281 11509 21315 11543
rect 23397 11509 23431 11543
rect 25053 11509 25087 11543
rect 25421 11509 25455 11543
rect 28641 11509 28675 11543
rect 29009 11509 29043 11543
rect 33517 11509 33551 11543
rect 34253 11509 34287 11543
rect 35081 11509 35115 11543
rect 36185 11509 36219 11543
rect 41153 11509 41187 11543
rect 42901 11509 42935 11543
rect 44097 11509 44131 11543
rect 14013 11305 14047 11339
rect 19073 11305 19107 11339
rect 22937 11305 22971 11339
rect 24685 11305 24719 11339
rect 25605 11305 25639 11339
rect 25881 11305 25915 11339
rect 26341 11305 26375 11339
rect 29193 11305 29227 11339
rect 29561 11305 29595 11339
rect 30849 11305 30883 11339
rect 34621 11305 34655 11339
rect 35265 11305 35299 11339
rect 37105 11305 37139 11339
rect 37473 11305 37507 11339
rect 38945 11305 38979 11339
rect 43085 11305 43119 11339
rect 11437 11237 11471 11271
rect 13001 11237 13035 11271
rect 13093 11237 13127 11271
rect 13645 11237 13679 11271
rect 17141 11237 17175 11271
rect 23397 11237 23431 11271
rect 23489 11237 23523 11271
rect 26846 11237 26880 11271
rect 29929 11237 29963 11271
rect 32321 11237 32355 11271
rect 34022 11237 34056 11271
rect 36277 11237 36311 11271
rect 37841 11237 37875 11271
rect 37933 11237 37967 11271
rect 41429 11237 41463 11271
rect 43545 11237 43579 11271
rect 9965 11169 9999 11203
rect 10241 11169 10275 11203
rect 15669 11169 15703 11203
rect 15945 11169 15979 11203
rect 18981 11169 19015 11203
rect 19441 11169 19475 11203
rect 20913 11169 20947 11203
rect 22109 11169 22143 11203
rect 25421 11169 25455 11203
rect 28641 11169 28675 11203
rect 33701 11169 33735 11203
rect 39313 11169 39347 11203
rect 39773 11169 39807 11203
rect 10425 11101 10459 11135
rect 10701 11101 10735 11135
rect 11345 11101 11379 11135
rect 16129 11101 16163 11135
rect 17049 11101 17083 11135
rect 17693 11101 17727 11135
rect 22293 11101 22327 11135
rect 23673 11101 23707 11135
rect 26525 11101 26559 11135
rect 29837 11101 29871 11135
rect 30113 11101 30147 11135
rect 32229 11101 32263 11135
rect 32505 11101 32539 11135
rect 36185 11101 36219 11135
rect 38117 11101 38151 11135
rect 40049 11101 40083 11135
rect 41337 11101 41371 11135
rect 43453 11101 43487 11135
rect 43729 11101 43763 11135
rect 11897 11033 11931 11067
rect 24409 11033 24443 11067
rect 27445 11033 27479 11067
rect 36737 11033 36771 11067
rect 41889 11033 41923 11067
rect 19993 10965 20027 10999
rect 21097 10965 21131 10999
rect 25145 10965 25179 10999
rect 28871 10965 28905 10999
rect 33241 10965 33275 10999
rect 9873 10761 9907 10795
rect 11253 10761 11287 10795
rect 12173 10761 12207 10795
rect 13001 10761 13035 10795
rect 14749 10761 14783 10795
rect 15347 10761 15381 10795
rect 17141 10761 17175 10795
rect 17417 10761 17451 10795
rect 18199 10761 18233 10795
rect 18981 10761 19015 10795
rect 21465 10761 21499 10795
rect 25973 10761 26007 10795
rect 28181 10761 28215 10795
rect 28733 10761 28767 10795
rect 29561 10761 29595 10795
rect 30481 10761 30515 10795
rect 31769 10761 31803 10795
rect 33333 10761 33367 10795
rect 33931 10761 33965 10795
rect 34345 10761 34379 10795
rect 36185 10761 36219 10795
rect 37749 10761 37783 10795
rect 38117 10761 38151 10795
rect 38669 10761 38703 10795
rect 39865 10761 39899 10795
rect 41337 10761 41371 10795
rect 42901 10761 42935 10795
rect 43453 10761 43487 10795
rect 44189 10761 44223 10795
rect 15117 10693 15151 10727
rect 17785 10693 17819 10727
rect 22661 10693 22695 10727
rect 24501 10693 24535 10727
rect 31309 10693 31343 10727
rect 41797 10693 41831 10727
rect 10333 10625 10367 10659
rect 13185 10625 13219 10659
rect 16221 10625 16255 10659
rect 18613 10625 18647 10659
rect 21925 10625 21959 10659
rect 22109 10625 22143 10659
rect 24225 10625 24259 10659
rect 29791 10625 29825 10659
rect 32781 10625 32815 10659
rect 34989 10625 35023 10659
rect 35265 10625 35299 10659
rect 36829 10625 36863 10659
rect 37105 10625 37139 10659
rect 41981 10625 42015 10659
rect 43729 10625 43763 10659
rect 9321 10557 9355 10591
rect 11529 10557 11563 10591
rect 13277 10557 13311 10591
rect 15244 10557 15278 10591
rect 15761 10557 15795 10591
rect 17969 10557 18003 10591
rect 19349 10557 19383 10591
rect 19809 10557 19843 10591
rect 20361 10557 20395 10591
rect 23397 10557 23431 10591
rect 23740 10557 23774 10591
rect 25053 10557 25087 10591
rect 26893 10557 26927 10591
rect 27261 10557 27295 10591
rect 29704 10557 29738 10591
rect 30205 10557 30239 10591
rect 33860 10557 33894 10591
rect 38853 10557 38887 10591
rect 39313 10557 39347 10591
rect 40325 10557 40359 10591
rect 40544 10557 40578 10591
rect 9229 10489 9263 10523
rect 10654 10489 10688 10523
rect 16037 10489 16071 10523
rect 16542 10489 16576 10523
rect 20085 10489 20119 10523
rect 22201 10489 22235 10523
rect 27813 10489 27847 10523
rect 30757 10489 30791 10523
rect 30849 10489 30883 10523
rect 32137 10489 32171 10523
rect 32321 10489 32355 10523
rect 32413 10489 32447 10523
rect 35081 10489 35115 10523
rect 36921 10489 36955 10523
rect 39589 10489 39623 10523
rect 42302 10489 42336 10523
rect 10149 10421 10183 10455
rect 21005 10421 21039 10455
rect 23811 10421 23845 10455
rect 24869 10421 24903 10455
rect 25421 10421 25455 10455
rect 26525 10421 26559 10455
rect 26893 10421 26927 10455
rect 33609 10421 33643 10455
rect 34621 10421 34655 10455
rect 36645 10421 36679 10455
rect 40647 10421 40681 10455
rect 11345 10217 11379 10251
rect 11805 10217 11839 10251
rect 13277 10217 13311 10251
rect 15807 10217 15841 10251
rect 16221 10217 16255 10251
rect 18061 10217 18095 10251
rect 18981 10217 19015 10251
rect 23949 10217 23983 10251
rect 25881 10217 25915 10251
rect 27169 10217 27203 10251
rect 27445 10217 27479 10251
rect 29285 10217 29319 10251
rect 30481 10217 30515 10251
rect 30849 10217 30883 10251
rect 32137 10217 32171 10251
rect 32597 10217 32631 10251
rect 34437 10217 34471 10251
rect 34897 10217 34931 10251
rect 36093 10217 36127 10251
rect 36645 10217 36679 10251
rect 38945 10217 38979 10251
rect 39313 10217 39347 10251
rect 41061 10217 41095 10251
rect 41981 10217 42015 10251
rect 12909 10149 12943 10183
rect 13737 10149 13771 10183
rect 13829 10149 13863 10183
rect 17002 10149 17036 10183
rect 19394 10149 19428 10183
rect 21234 10149 21268 10183
rect 23350 10149 23384 10183
rect 24961 10149 24995 10183
rect 25513 10149 25547 10183
rect 26801 10149 26835 10183
rect 29882 10149 29916 10183
rect 32965 10149 32999 10183
rect 33838 10149 33872 10183
rect 36921 10149 36955 10183
rect 37933 10149 37967 10183
rect 40462 10149 40496 10183
rect 41337 10149 41371 10183
rect 10149 10081 10183 10115
rect 10609 10081 10643 10115
rect 11713 10081 11747 10115
rect 12173 10081 12207 10115
rect 15736 10081 15770 10115
rect 19073 10081 19107 10115
rect 26985 10081 27019 10115
rect 27997 10081 28031 10115
rect 28457 10081 28491 10115
rect 37289 10081 37323 10115
rect 40141 10081 40175 10115
rect 10701 10013 10735 10047
rect 16681 10013 16715 10047
rect 20913 10013 20947 10047
rect 23029 10013 23063 10047
rect 24869 10013 24903 10047
rect 28733 10013 28767 10047
rect 29561 10013 29595 10047
rect 33517 10013 33551 10047
rect 35725 10013 35759 10047
rect 37841 10013 37875 10047
rect 38117 10013 38151 10047
rect 14289 9945 14323 9979
rect 17601 9877 17635 9911
rect 19993 9877 20027 9911
rect 21833 9877 21867 9911
rect 9781 9673 9815 9707
rect 10517 9673 10551 9707
rect 11805 9673 11839 9707
rect 12173 9673 12207 9707
rect 15301 9673 15335 9707
rect 16681 9673 16715 9707
rect 18521 9673 18555 9707
rect 19165 9673 19199 9707
rect 19533 9673 19567 9707
rect 21281 9673 21315 9707
rect 22477 9673 22511 9707
rect 23029 9673 23063 9707
rect 25053 9673 25087 9707
rect 25145 9673 25179 9707
rect 26617 9673 26651 9707
rect 28181 9673 28215 9707
rect 28457 9673 28491 9707
rect 29009 9673 29043 9707
rect 30205 9673 30239 9707
rect 31953 9673 31987 9707
rect 36737 9673 36771 9707
rect 37749 9673 37783 9707
rect 38117 9673 38151 9707
rect 40141 9673 40175 9707
rect 41429 9673 41463 9707
rect 10149 9605 10183 9639
rect 24869 9605 24903 9639
rect 10609 9537 10643 9571
rect 13921 9537 13955 9571
rect 14289 9537 14323 9571
rect 17095 9537 17129 9571
rect 21557 9537 21591 9571
rect 21833 9537 21867 9571
rect 23765 9537 23799 9571
rect 24041 9537 24075 9571
rect 12516 9469 12550 9503
rect 14933 9469 14967 9503
rect 15485 9469 15519 9503
rect 17008 9469 17042 9503
rect 18128 9469 18162 9503
rect 19717 9469 19751 9503
rect 23489 9469 23523 9503
rect 26249 9605 26283 9639
rect 32873 9605 32907 9639
rect 27629 9537 27663 9571
rect 29285 9537 29319 9571
rect 30481 9537 30515 9571
rect 33793 9537 33827 9571
rect 34437 9537 34471 9571
rect 38669 9537 38703 9571
rect 25329 9469 25363 9503
rect 26985 9469 27019 9503
rect 27169 9469 27203 9503
rect 27537 9469 27571 9503
rect 31033 9469 31067 9503
rect 33057 9469 33091 9503
rect 33609 9469 33643 9503
rect 35817 9469 35851 9503
rect 38853 9469 38887 9503
rect 39313 9469 39347 9503
rect 39589 9469 39623 9503
rect 40509 9469 40543 9503
rect 10930 9401 10964 9435
rect 13001 9401 13035 9435
rect 13737 9401 13771 9435
rect 14013 9401 14047 9435
rect 15393 9401 15427 9435
rect 20913 9401 20947 9435
rect 21649 9401 21683 9435
rect 23857 9401 23891 9435
rect 25053 9401 25087 9435
rect 25650 9401 25684 9435
rect 29606 9401 29640 9435
rect 30849 9401 30883 9435
rect 31354 9401 31388 9435
rect 34069 9401 34103 9435
rect 35265 9401 35299 9435
rect 35633 9401 35667 9435
rect 36138 9401 36172 9435
rect 40830 9401 40864 9435
rect 11529 9333 11563 9367
rect 12587 9333 12621 9367
rect 13369 9333 13403 9367
rect 17509 9333 17543 9367
rect 18199 9333 18233 9367
rect 20085 9333 20119 9367
rect 20637 9333 20671 9367
rect 10701 9129 10735 9163
rect 11253 9129 11287 9163
rect 12449 9129 12483 9163
rect 13921 9129 13955 9163
rect 21925 9129 21959 9163
rect 22615 9129 22649 9163
rect 23673 9129 23707 9163
rect 24869 9129 24903 9163
rect 25421 9129 25455 9163
rect 26617 9129 26651 9163
rect 29745 9129 29779 9163
rect 33149 9129 33183 9163
rect 35725 9129 35759 9163
rect 36691 9129 36725 9163
rect 38945 9129 38979 9163
rect 40141 9129 40175 9163
rect 40877 9129 40911 9163
rect 12817 9061 12851 9095
rect 15439 9061 15473 9095
rect 17325 9061 17359 9095
rect 19717 9061 19751 9095
rect 19993 9061 20027 9095
rect 21097 9061 21131 9095
rect 21649 9061 21683 9095
rect 23029 9061 23063 9095
rect 29469 9061 29503 9095
rect 35449 9061 35483 9095
rect 36093 9061 36127 9095
rect 10885 8993 10919 9027
rect 11805 8993 11839 9027
rect 14197 8993 14231 9027
rect 15336 8993 15370 9027
rect 15761 8993 15795 9027
rect 18981 8993 19015 9027
rect 19441 8993 19475 9027
rect 22544 8993 22578 9027
rect 26709 8993 26743 9027
rect 27077 8993 27111 9027
rect 28733 8993 28767 9027
rect 29193 8993 29227 9027
rect 33609 8993 33643 9027
rect 34713 8993 34747 9027
rect 35173 8993 35207 9027
rect 36553 8993 36587 9027
rect 40509 8993 40543 9027
rect 12725 8925 12759 8959
rect 13093 8925 13127 8959
rect 17233 8925 17267 8959
rect 17693 8925 17727 8959
rect 21005 8925 21039 8959
rect 14381 8789 14415 8823
rect 16681 8789 16715 8823
rect 31033 8789 31067 8823
rect 33747 8789 33781 8823
rect 10977 8585 11011 8619
rect 12173 8585 12207 8619
rect 13461 8585 13495 8619
rect 17693 8585 17727 8619
rect 18981 8585 19015 8619
rect 19441 8585 19475 8619
rect 20039 8585 20073 8619
rect 20637 8585 20671 8619
rect 21005 8585 21039 8619
rect 27169 8585 27203 8619
rect 28457 8585 28491 8619
rect 28733 8585 28767 8619
rect 33609 8585 33643 8619
rect 34253 8585 34287 8619
rect 34621 8585 34655 8619
rect 36553 8585 36587 8619
rect 11345 8517 11379 8551
rect 13093 8517 13127 8551
rect 22569 8517 22603 8551
rect 12541 8449 12575 8483
rect 14013 8449 14047 8483
rect 21281 8449 21315 8483
rect 21925 8449 21959 8483
rect 30021 8449 30055 8483
rect 33793 8449 33827 8483
rect 35633 8449 35667 8483
rect 13921 8381 13955 8415
rect 14381 8381 14415 8415
rect 17417 8381 17451 8415
rect 18096 8381 18130 8415
rect 18521 8381 18555 8415
rect 19809 8381 19843 8415
rect 19968 8381 20002 8415
rect 26341 8381 26375 8415
rect 26617 8381 26651 8415
rect 29561 8381 29595 8415
rect 29745 8381 29779 8415
rect 34897 8381 34931 8415
rect 35357 8381 35391 8415
rect 12633 8313 12667 8347
rect 15485 8313 15519 8347
rect 15669 8313 15703 8347
rect 18199 8313 18233 8347
rect 21373 8313 21407 8347
rect 25973 8313 26007 8347
rect 15117 8245 15151 8279
rect 22201 8245 22235 8279
rect 26157 8245 26191 8279
rect 12725 8041 12759 8075
rect 13231 8041 13265 8075
rect 14335 8041 14369 8075
rect 15761 8041 15795 8075
rect 16037 8041 16071 8075
rect 16497 8041 16531 8075
rect 17233 8041 17267 8075
rect 17509 8041 17543 8075
rect 19993 8041 20027 8075
rect 21189 8041 21223 8075
rect 21373 8041 21407 8075
rect 26157 8041 26191 8075
rect 26709 8041 26743 8075
rect 29377 8041 29411 8075
rect 29745 8041 29779 8075
rect 34713 8041 34747 8075
rect 35081 8041 35115 8075
rect 14105 7973 14139 8007
rect 13093 7905 13127 7939
rect 15577 7905 15611 7939
rect 16497 7905 16531 7939
rect 16681 7905 16715 7939
rect 17049 7905 17083 7939
rect 19533 7905 19567 7939
rect 20948 7905 20982 7939
rect 17693 7837 17727 7871
rect 18061 7837 18095 7871
rect 13553 7701 13587 7735
rect 12265 7497 12299 7531
rect 15485 7497 15519 7531
rect 15945 7497 15979 7531
rect 16313 7497 16347 7531
rect 20361 7497 20395 7531
rect 20913 7497 20947 7531
rect 13185 7361 13219 7395
rect 18429 7361 18463 7395
rect 12725 7293 12759 7327
rect 13553 7293 13587 7327
rect 15025 7293 15059 7327
rect 17877 7293 17911 7327
rect 18061 7293 18095 7327
rect 19901 7293 19935 7327
rect 13001 7225 13035 7259
rect 17141 7225 17175 7259
rect 17509 7225 17543 7259
rect 16865 7157 16899 7191
rect 17693 7157 17727 7191
rect 13553 6953 13587 6987
rect 14289 6953 14323 6987
rect 17877 6953 17911 6987
rect 18521 6953 18555 6987
rect 18889 6953 18923 6987
rect 18245 6885 18279 6919
rect 13737 6817 13771 6851
rect 15945 6817 15979 6851
rect 17417 6817 17451 6851
rect 15577 6749 15611 6783
rect 13185 6613 13219 6647
rect 15209 6409 15243 6443
rect 15577 6409 15611 6443
rect 16313 6409 16347 6443
rect 17141 6409 17175 6443
rect 18337 6409 18371 6443
rect 18613 6409 18647 6443
rect 13645 6341 13679 6375
rect 17693 6341 17727 6375
rect 16037 6273 16071 6307
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 48852 47354
rect 1104 47280 48852 47302
rect 1104 46810 48852 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 48852 46810
rect 1104 46736 48852 46758
rect 1104 46266 48852 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 48852 46266
rect 1104 46192 48852 46214
rect 1104 45722 48852 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 48852 45722
rect 1104 45648 48852 45670
rect 1104 45178 48852 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 48852 45178
rect 1104 45104 48852 45126
rect 1104 44634 48852 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 48852 44634
rect 1104 44560 48852 44582
rect 38010 44384 38016 44396
rect 31128 44356 38016 44384
rect 30742 44325 30748 44328
rect 30720 44319 30748 44325
rect 30720 44316 30732 44319
rect 30655 44288 30732 44316
rect 30720 44285 30732 44288
rect 30800 44316 30806 44328
rect 31128 44325 31156 44356
rect 38010 44344 38016 44356
rect 38068 44344 38074 44396
rect 31113 44319 31171 44325
rect 31113 44316 31125 44319
rect 30800 44288 31125 44316
rect 30720 44279 30748 44285
rect 30742 44276 30748 44279
rect 30800 44276 30806 44288
rect 31113 44285 31125 44288
rect 31159 44285 31171 44319
rect 31113 44279 31171 44285
rect 31846 44276 31852 44328
rect 31904 44316 31910 44328
rect 33204 44319 33262 44325
rect 33204 44316 33216 44319
rect 31904 44288 33216 44316
rect 31904 44276 31910 44288
rect 33204 44285 33216 44288
rect 33250 44316 33262 44319
rect 33597 44319 33655 44325
rect 33597 44316 33609 44319
rect 33250 44288 33609 44316
rect 33250 44285 33262 44288
rect 33204 44279 33262 44285
rect 33597 44285 33609 44288
rect 33643 44285 33655 44319
rect 33597 44279 33655 44285
rect 30791 44183 30849 44189
rect 30791 44149 30803 44183
rect 30837 44180 30849 44183
rect 31018 44180 31024 44192
rect 30837 44152 31024 44180
rect 30837 44149 30849 44152
rect 30791 44143 30849 44149
rect 31018 44140 31024 44152
rect 31076 44140 31082 44192
rect 33275 44183 33333 44189
rect 33275 44149 33287 44183
rect 33321 44180 33333 44183
rect 34790 44180 34796 44192
rect 33321 44152 34796 44180
rect 33321 44149 33333 44152
rect 33275 44143 33333 44149
rect 34790 44140 34796 44152
rect 34848 44140 34854 44192
rect 1104 44090 48852 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 48852 44090
rect 1104 44016 48852 44038
rect 31018 43936 31024 43988
rect 31076 43976 31082 43988
rect 32493 43979 32551 43985
rect 32493 43976 32505 43979
rect 31076 43948 32505 43976
rect 31076 43936 31082 43948
rect 32493 43945 32505 43948
rect 32539 43976 32551 43979
rect 32582 43976 32588 43988
rect 32539 43948 32588 43976
rect 32539 43945 32551 43948
rect 32493 43939 32551 43945
rect 32582 43936 32588 43948
rect 32640 43936 32646 43988
rect 33413 43911 33471 43917
rect 33413 43877 33425 43911
rect 33459 43908 33471 43911
rect 33686 43908 33692 43920
rect 33459 43880 33692 43908
rect 33459 43877 33471 43880
rect 33413 43871 33471 43877
rect 33686 43868 33692 43880
rect 33744 43868 33750 43920
rect 23106 43840 23112 43852
rect 23067 43812 23112 43840
rect 23106 43800 23112 43812
rect 23164 43800 23170 43852
rect 24949 43843 25007 43849
rect 24949 43809 24961 43843
rect 24995 43840 25007 43843
rect 25038 43840 25044 43852
rect 24995 43812 25044 43840
rect 24995 43809 25007 43812
rect 24949 43803 25007 43809
rect 25038 43800 25044 43812
rect 25096 43800 25102 43852
rect 30444 43843 30502 43849
rect 30444 43809 30456 43843
rect 30490 43840 30502 43843
rect 30834 43840 30840 43852
rect 30490 43812 30840 43840
rect 30490 43809 30502 43812
rect 30444 43803 30502 43809
rect 30834 43800 30840 43812
rect 30892 43800 30898 43852
rect 33318 43772 33324 43784
rect 33279 43744 33324 43772
rect 33318 43732 33324 43744
rect 33376 43732 33382 43784
rect 33597 43775 33655 43781
rect 33597 43741 33609 43775
rect 33643 43741 33655 43775
rect 33597 43735 33655 43741
rect 31202 43664 31208 43716
rect 31260 43704 31266 43716
rect 33502 43704 33508 43716
rect 31260 43676 33508 43704
rect 31260 43664 31266 43676
rect 33502 43664 33508 43676
rect 33560 43704 33566 43716
rect 33612 43704 33640 43735
rect 33560 43676 33640 43704
rect 33560 43664 33566 43676
rect 23247 43639 23305 43645
rect 23247 43605 23259 43639
rect 23293 43636 23305 43639
rect 23566 43636 23572 43648
rect 23293 43608 23572 43636
rect 23293 43605 23305 43608
rect 23247 43599 23305 43605
rect 23566 43596 23572 43608
rect 23624 43596 23630 43648
rect 23753 43639 23811 43645
rect 23753 43605 23765 43639
rect 23799 43636 23811 43639
rect 23842 43636 23848 43648
rect 23799 43608 23848 43636
rect 23799 43605 23811 43608
rect 23753 43599 23811 43605
rect 23842 43596 23848 43608
rect 23900 43596 23906 43648
rect 24026 43636 24032 43648
rect 23987 43608 24032 43636
rect 24026 43596 24032 43608
rect 24084 43596 24090 43648
rect 25179 43639 25237 43645
rect 25179 43605 25191 43639
rect 25225 43636 25237 43639
rect 25406 43636 25412 43648
rect 25225 43608 25412 43636
rect 25225 43605 25237 43608
rect 25179 43599 25237 43605
rect 25406 43596 25412 43608
rect 25464 43596 25470 43648
rect 25590 43636 25596 43648
rect 25551 43608 25596 43636
rect 25590 43596 25596 43608
rect 25648 43596 25654 43648
rect 30374 43596 30380 43648
rect 30432 43636 30438 43648
rect 30515 43639 30573 43645
rect 30515 43636 30527 43639
rect 30432 43608 30527 43636
rect 30432 43596 30438 43608
rect 30515 43605 30527 43608
rect 30561 43605 30573 43639
rect 31018 43636 31024 43648
rect 30979 43608 31024 43636
rect 30515 43599 30573 43605
rect 31018 43596 31024 43608
rect 31076 43596 31082 43648
rect 31294 43636 31300 43648
rect 31255 43608 31300 43636
rect 31294 43596 31300 43608
rect 31352 43596 31358 43648
rect 1104 43546 48852 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 48852 43546
rect 1104 43472 48852 43494
rect 22370 43392 22376 43444
rect 22428 43432 22434 43444
rect 23106 43432 23112 43444
rect 22428 43404 23112 43432
rect 22428 43392 22434 43404
rect 23106 43392 23112 43404
rect 23164 43392 23170 43444
rect 25038 43432 25044 43444
rect 24999 43404 25044 43432
rect 25038 43392 25044 43404
rect 25096 43432 25102 43444
rect 30377 43435 30435 43441
rect 30377 43432 30389 43435
rect 25096 43404 30389 43432
rect 25096 43392 25102 43404
rect 23198 43324 23204 43376
rect 23256 43364 23262 43376
rect 24305 43367 24363 43373
rect 24305 43364 24317 43367
rect 23256 43336 24317 43364
rect 23256 43324 23262 43336
rect 24305 43333 24317 43336
rect 24351 43364 24363 43367
rect 26602 43364 26608 43376
rect 24351 43336 26608 43364
rect 24351 43333 24363 43336
rect 24305 43327 24363 43333
rect 26602 43324 26608 43336
rect 26660 43324 26666 43376
rect 23474 43256 23480 43308
rect 23532 43296 23538 43308
rect 23753 43299 23811 43305
rect 23753 43296 23765 43299
rect 23532 43268 23765 43296
rect 23532 43256 23538 43268
rect 23753 43265 23765 43268
rect 23799 43296 23811 43299
rect 24026 43296 24032 43308
rect 23799 43268 24032 43296
rect 23799 43265 23811 43268
rect 23753 43259 23811 43265
rect 24026 43256 24032 43268
rect 24084 43256 24090 43308
rect 24210 43256 24216 43308
rect 24268 43296 24274 43308
rect 25777 43299 25835 43305
rect 25777 43296 25789 43299
rect 24268 43268 25789 43296
rect 24268 43256 24274 43268
rect 25777 43265 25789 43268
rect 25823 43265 25835 43299
rect 25777 43259 25835 43265
rect 22592 43231 22650 43237
rect 22592 43228 22604 43231
rect 22388 43200 22604 43228
rect 21634 43052 21640 43104
rect 21692 43092 21698 43104
rect 22388 43101 22416 43200
rect 22592 43197 22604 43200
rect 22638 43197 22650 43231
rect 22592 43191 22650 43197
rect 27433 43231 27491 43237
rect 27433 43197 27445 43231
rect 27479 43228 27491 43231
rect 27522 43228 27528 43240
rect 27479 43200 27528 43228
rect 27479 43197 27491 43200
rect 27433 43191 27491 43197
rect 27522 43188 27528 43200
rect 27580 43188 27586 43240
rect 27982 43228 27988 43240
rect 27943 43200 27988 43228
rect 27982 43188 27988 43200
rect 28040 43188 28046 43240
rect 29983 43237 30011 43404
rect 30377 43401 30389 43404
rect 30423 43432 30435 43435
rect 30466 43432 30472 43444
rect 30423 43404 30472 43432
rect 30423 43401 30435 43404
rect 30377 43395 30435 43401
rect 30466 43392 30472 43404
rect 30524 43392 30530 43444
rect 30834 43432 30840 43444
rect 30747 43404 30840 43432
rect 30834 43392 30840 43404
rect 30892 43432 30898 43444
rect 30892 43404 33134 43432
rect 30892 43392 30898 43404
rect 30558 43324 30564 43376
rect 30616 43364 30622 43376
rect 33106 43364 33134 43404
rect 33318 43392 33324 43444
rect 33376 43432 33382 43444
rect 33870 43432 33876 43444
rect 33376 43404 33876 43432
rect 33376 43392 33382 43404
rect 33870 43392 33876 43404
rect 33928 43392 33934 43444
rect 37090 43364 37096 43376
rect 30616 43336 32720 43364
rect 33106 43336 37096 43364
rect 30616 43324 30622 43336
rect 30055 43299 30113 43305
rect 30055 43265 30067 43299
rect 30101 43296 30113 43299
rect 31021 43299 31079 43305
rect 31021 43296 31033 43299
rect 30101 43268 31033 43296
rect 30101 43265 30113 43268
rect 30055 43259 30113 43265
rect 31021 43265 31033 43268
rect 31067 43296 31079 43299
rect 31294 43296 31300 43308
rect 31067 43268 31300 43296
rect 31067 43265 31079 43268
rect 31021 43259 31079 43265
rect 31294 43256 31300 43268
rect 31352 43256 31358 43308
rect 32582 43296 32588 43308
rect 32543 43268 32588 43296
rect 32582 43256 32588 43268
rect 32640 43256 32646 43308
rect 32692 43296 32720 43336
rect 37090 43324 37096 43336
rect 37148 43324 37154 43376
rect 32861 43299 32919 43305
rect 32861 43296 32873 43299
rect 32692 43268 32873 43296
rect 32861 43265 32873 43268
rect 32907 43265 32919 43299
rect 32861 43259 32919 43265
rect 29968 43231 30026 43237
rect 29968 43197 29980 43231
rect 30014 43197 30026 43231
rect 29968 43191 30026 43197
rect 34952 43231 35010 43237
rect 34952 43197 34964 43231
rect 34998 43228 35010 43231
rect 34998 43200 35480 43228
rect 34998 43197 35010 43200
rect 34952 43191 35010 43197
rect 23842 43120 23848 43172
rect 23900 43160 23906 43172
rect 24765 43163 24823 43169
rect 23900 43132 23945 43160
rect 23900 43120 23906 43132
rect 24765 43129 24777 43163
rect 24811 43160 24823 43163
rect 25498 43160 25504 43172
rect 24811 43132 25504 43160
rect 24811 43129 24823 43132
rect 24765 43123 24823 43129
rect 25498 43120 25504 43132
rect 25556 43120 25562 43172
rect 25590 43120 25596 43172
rect 25648 43160 25654 43172
rect 25648 43132 25693 43160
rect 25648 43120 25654 43132
rect 31018 43120 31024 43172
rect 31076 43160 31082 43172
rect 31113 43163 31171 43169
rect 31113 43160 31125 43163
rect 31076 43132 31125 43160
rect 31076 43120 31082 43132
rect 31113 43129 31125 43132
rect 31159 43129 31171 43163
rect 31662 43160 31668 43172
rect 31623 43132 31668 43160
rect 31113 43123 31171 43129
rect 22373 43095 22431 43101
rect 22373 43092 22385 43095
rect 21692 43064 22385 43092
rect 21692 43052 21698 43064
rect 22373 43061 22385 43064
rect 22419 43061 22431 43095
rect 22373 43055 22431 43061
rect 22695 43095 22753 43101
rect 22695 43061 22707 43095
rect 22741 43092 22753 43095
rect 23014 43092 23020 43104
rect 22741 43064 23020 43092
rect 22741 43061 22753 43064
rect 22695 43055 22753 43061
rect 23014 43052 23020 43064
rect 23072 43052 23078 43104
rect 27614 43092 27620 43104
rect 27575 43064 27620 43092
rect 27614 43052 27620 43064
rect 27672 43052 27678 43104
rect 31128 43092 31156 43123
rect 31662 43120 31668 43132
rect 31720 43120 31726 43172
rect 32677 43163 32735 43169
rect 32677 43160 32689 43163
rect 32324 43132 32689 43160
rect 32324 43101 32352 43132
rect 32677 43129 32689 43132
rect 32723 43129 32735 43163
rect 32677 43123 32735 43129
rect 35452 43104 35480 43200
rect 32309 43095 32367 43101
rect 32309 43092 32321 43095
rect 31128 43064 32321 43092
rect 32309 43061 32321 43064
rect 32355 43061 32367 43095
rect 32309 43055 32367 43061
rect 33597 43095 33655 43101
rect 33597 43061 33609 43095
rect 33643 43092 33655 43095
rect 33686 43092 33692 43104
rect 33643 43064 33692 43092
rect 33643 43061 33655 43064
rect 33597 43055 33655 43061
rect 33686 43052 33692 43064
rect 33744 43052 33750 43104
rect 34238 43052 34244 43104
rect 34296 43092 34302 43104
rect 35023 43095 35081 43101
rect 35023 43092 35035 43095
rect 34296 43064 35035 43092
rect 34296 43052 34302 43064
rect 35023 43061 35035 43064
rect 35069 43061 35081 43095
rect 35434 43092 35440 43104
rect 35395 43064 35440 43092
rect 35023 43055 35081 43061
rect 35434 43052 35440 43064
rect 35492 43052 35498 43104
rect 1104 43002 48852 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 48852 43002
rect 1104 42928 48852 42950
rect 27617 42891 27675 42897
rect 27617 42857 27629 42891
rect 27663 42888 27675 42891
rect 27982 42888 27988 42900
rect 27663 42860 27988 42888
rect 27663 42857 27675 42860
rect 27617 42851 27675 42857
rect 27982 42848 27988 42860
rect 28040 42848 28046 42900
rect 33686 42888 33692 42900
rect 33612 42860 33692 42888
rect 23566 42820 23572 42832
rect 23527 42792 23572 42820
rect 23566 42780 23572 42792
rect 23624 42780 23630 42832
rect 23658 42780 23664 42832
rect 23716 42820 23722 42832
rect 24210 42820 24216 42832
rect 23716 42792 23761 42820
rect 24171 42792 24216 42820
rect 23716 42780 23722 42792
rect 24210 42780 24216 42792
rect 24268 42780 24274 42832
rect 25406 42780 25412 42832
rect 25464 42820 25470 42832
rect 26234 42820 26240 42832
rect 25464 42792 26240 42820
rect 25464 42780 25470 42792
rect 26234 42780 26240 42792
rect 26292 42820 26298 42832
rect 26605 42823 26663 42829
rect 26605 42820 26617 42823
rect 26292 42792 26617 42820
rect 26292 42780 26298 42792
rect 26605 42789 26617 42792
rect 26651 42789 26663 42823
rect 26605 42783 26663 42789
rect 26694 42780 26700 42832
rect 26752 42820 26758 42832
rect 26752 42792 26797 42820
rect 26752 42780 26758 42792
rect 30374 42780 30380 42832
rect 30432 42820 30438 42832
rect 30561 42823 30619 42829
rect 30561 42820 30573 42823
rect 30432 42792 30573 42820
rect 30432 42780 30438 42792
rect 30561 42789 30573 42792
rect 30607 42789 30619 42823
rect 30561 42783 30619 42789
rect 30653 42823 30711 42829
rect 30653 42789 30665 42823
rect 30699 42820 30711 42823
rect 31018 42820 31024 42832
rect 30699 42792 31024 42820
rect 30699 42789 30711 42792
rect 30653 42783 30711 42789
rect 31018 42780 31024 42792
rect 31076 42780 31082 42832
rect 31202 42820 31208 42832
rect 31163 42792 31208 42820
rect 31202 42780 31208 42792
rect 31260 42780 31266 42832
rect 33612 42829 33640 42860
rect 33686 42848 33692 42860
rect 33744 42888 33750 42900
rect 33744 42860 35204 42888
rect 33744 42848 33750 42860
rect 33597 42823 33655 42829
rect 33597 42789 33609 42823
rect 33643 42789 33655 42823
rect 33597 42783 33655 42789
rect 34790 42780 34796 42832
rect 34848 42820 34854 42832
rect 35176 42829 35204 42860
rect 35069 42823 35127 42829
rect 35069 42820 35081 42823
rect 34848 42792 35081 42820
rect 34848 42780 34854 42792
rect 35069 42789 35081 42792
rect 35115 42789 35127 42823
rect 35069 42783 35127 42789
rect 35161 42823 35219 42829
rect 35161 42789 35173 42823
rect 35207 42820 35219 42823
rect 35710 42820 35716 42832
rect 35207 42792 35716 42820
rect 35207 42789 35219 42792
rect 35161 42783 35219 42789
rect 35710 42780 35716 42792
rect 35768 42780 35774 42832
rect 22440 42755 22498 42761
rect 22440 42721 22452 42755
rect 22486 42752 22498 42755
rect 23106 42752 23112 42764
rect 22486 42724 23112 42752
rect 22486 42721 22498 42724
rect 22440 42715 22498 42721
rect 23106 42712 23112 42724
rect 23164 42712 23170 42764
rect 25225 42755 25283 42761
rect 25225 42721 25237 42755
rect 25271 42752 25283 42755
rect 25314 42752 25320 42764
rect 25271 42724 25320 42752
rect 25271 42721 25283 42724
rect 25225 42715 25283 42721
rect 25314 42712 25320 42724
rect 25372 42712 25378 42764
rect 27522 42712 27528 42764
rect 27580 42752 27586 42764
rect 29178 42752 29184 42764
rect 27580 42724 29184 42752
rect 27580 42712 27586 42724
rect 29178 42712 29184 42724
rect 29236 42712 29242 42764
rect 29457 42755 29515 42761
rect 29457 42721 29469 42755
rect 29503 42752 29515 42755
rect 29546 42752 29552 42764
rect 29503 42724 29552 42752
rect 29503 42721 29515 42724
rect 29457 42715 29515 42721
rect 29546 42712 29552 42724
rect 29604 42712 29610 42764
rect 32401 42755 32459 42761
rect 32401 42721 32413 42755
rect 32447 42752 32459 42755
rect 32490 42752 32496 42764
rect 32447 42724 32496 42752
rect 32447 42721 32459 42724
rect 32401 42715 32459 42721
rect 32490 42712 32496 42724
rect 32548 42712 32554 42764
rect 37090 42712 37096 42764
rect 37148 42752 37154 42764
rect 38105 42755 38163 42761
rect 38105 42752 38117 42755
rect 37148 42724 38117 42752
rect 37148 42712 37154 42724
rect 38105 42721 38117 42724
rect 38151 42752 38163 42755
rect 38194 42752 38200 42764
rect 38151 42724 38200 42752
rect 38151 42721 38163 42724
rect 38105 42715 38163 42721
rect 38194 42712 38200 42724
rect 38252 42712 38258 42764
rect 39850 42752 39856 42764
rect 39811 42724 39856 42752
rect 39850 42712 39856 42724
rect 39908 42712 39914 42764
rect 24394 42644 24400 42696
rect 24452 42684 24458 42696
rect 26881 42687 26939 42693
rect 26881 42684 26893 42687
rect 24452 42656 26893 42684
rect 24452 42644 24458 42656
rect 26881 42653 26893 42656
rect 26927 42653 26939 42687
rect 29638 42684 29644 42696
rect 29599 42656 29644 42684
rect 26881 42647 26939 42653
rect 29638 42644 29644 42656
rect 29696 42644 29702 42696
rect 33505 42687 33563 42693
rect 33505 42653 33517 42687
rect 33551 42684 33563 42687
rect 34238 42684 34244 42696
rect 33551 42656 34244 42684
rect 33551 42653 33563 42656
rect 33505 42647 33563 42653
rect 34238 42644 34244 42656
rect 34296 42644 34302 42696
rect 35526 42684 35532 42696
rect 35487 42656 35532 42684
rect 35526 42644 35532 42656
rect 35584 42644 35590 42696
rect 31662 42576 31668 42628
rect 31720 42616 31726 42628
rect 34054 42616 34060 42628
rect 31720 42588 34060 42616
rect 31720 42576 31726 42588
rect 34054 42576 34060 42588
rect 34112 42576 34118 42628
rect 35434 42576 35440 42628
rect 35492 42616 35498 42628
rect 39758 42616 39764 42628
rect 35492 42588 39764 42616
rect 35492 42576 35498 42588
rect 39758 42576 39764 42588
rect 39816 42616 39822 42628
rect 41414 42616 41420 42628
rect 39816 42588 41420 42616
rect 39816 42576 39822 42588
rect 41414 42576 41420 42588
rect 41472 42576 41478 42628
rect 22094 42508 22100 42560
rect 22152 42548 22158 42560
rect 22511 42551 22569 42557
rect 22511 42548 22523 42551
rect 22152 42520 22523 42548
rect 22152 42508 22158 42520
rect 22511 42517 22523 42520
rect 22557 42517 22569 42551
rect 22511 42511 22569 42517
rect 23750 42508 23756 42560
rect 23808 42548 23814 42560
rect 24489 42551 24547 42557
rect 24489 42548 24501 42551
rect 23808 42520 24501 42548
rect 23808 42508 23814 42520
rect 24489 42517 24501 42520
rect 24535 42517 24547 42551
rect 24489 42511 24547 42517
rect 25363 42551 25421 42557
rect 25363 42517 25375 42551
rect 25409 42548 25421 42551
rect 25590 42548 25596 42560
rect 25409 42520 25596 42548
rect 25409 42517 25421 42520
rect 25363 42511 25421 42517
rect 25590 42508 25596 42520
rect 25648 42548 25654 42560
rect 25685 42551 25743 42557
rect 25685 42548 25697 42551
rect 25648 42520 25697 42548
rect 25648 42508 25654 42520
rect 25685 42517 25697 42520
rect 25731 42517 25743 42551
rect 25685 42511 25743 42517
rect 32539 42551 32597 42557
rect 32539 42517 32551 42551
rect 32585 42548 32597 42551
rect 34698 42548 34704 42560
rect 32585 42520 34704 42548
rect 32585 42517 32597 42520
rect 32539 42511 32597 42517
rect 34698 42508 34704 42520
rect 34756 42508 34762 42560
rect 38243 42551 38301 42557
rect 38243 42517 38255 42551
rect 38289 42548 38301 42551
rect 38470 42548 38476 42560
rect 38289 42520 38476 42548
rect 38289 42517 38301 42520
rect 38243 42511 38301 42517
rect 38470 42508 38476 42520
rect 38528 42508 38534 42560
rect 38562 42508 38568 42560
rect 38620 42548 38626 42560
rect 39991 42551 40049 42557
rect 38620 42520 38665 42548
rect 38620 42508 38626 42520
rect 39991 42517 40003 42551
rect 40037 42548 40049 42551
rect 40310 42548 40316 42560
rect 40037 42520 40316 42548
rect 40037 42517 40049 42520
rect 39991 42511 40049 42517
rect 40310 42508 40316 42520
rect 40368 42508 40374 42560
rect 1104 42458 48852 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 48852 42458
rect 1104 42384 48852 42406
rect 18506 42304 18512 42356
rect 18564 42344 18570 42356
rect 19334 42344 19340 42356
rect 18564 42316 19340 42344
rect 18564 42304 18570 42316
rect 19334 42304 19340 42316
rect 19392 42344 19398 42356
rect 25314 42344 25320 42356
rect 19392 42316 25320 42344
rect 19392 42304 19398 42316
rect 25314 42304 25320 42316
rect 25372 42344 25378 42356
rect 30653 42347 30711 42353
rect 25372 42316 30236 42344
rect 25372 42304 25378 42316
rect 21913 42279 21971 42285
rect 21913 42245 21925 42279
rect 21959 42276 21971 42279
rect 23658 42276 23664 42288
rect 21959 42248 23664 42276
rect 21959 42245 21971 42248
rect 21913 42239 21971 42245
rect 21060 42143 21118 42149
rect 21060 42109 21072 42143
rect 21106 42140 21118 42143
rect 21453 42143 21511 42149
rect 21453 42140 21465 42143
rect 21106 42112 21465 42140
rect 21106 42109 21118 42112
rect 21060 42103 21118 42109
rect 21453 42109 21465 42112
rect 21499 42109 21511 42143
rect 21453 42103 21511 42109
rect 21131 42007 21189 42013
rect 21131 41973 21143 42007
rect 21177 42004 21189 42007
rect 21358 42004 21364 42016
rect 21177 41976 21364 42004
rect 21177 41973 21189 41976
rect 21131 41967 21189 41973
rect 21358 41964 21364 41976
rect 21416 41964 21422 42016
rect 21468 42004 21496 42103
rect 21928 42072 21956 42239
rect 23658 42236 23664 42248
rect 23716 42236 23722 42288
rect 26605 42279 26663 42285
rect 26605 42245 26617 42279
rect 26651 42276 26663 42279
rect 26694 42276 26700 42288
rect 26651 42248 26700 42276
rect 26651 42245 26663 42248
rect 26605 42239 26663 42245
rect 26694 42236 26700 42248
rect 26752 42276 26758 42288
rect 28353 42279 28411 42285
rect 28353 42276 28365 42279
rect 26752 42248 28365 42276
rect 26752 42236 26758 42248
rect 28353 42245 28365 42248
rect 28399 42245 28411 42279
rect 28353 42239 28411 42245
rect 22094 42208 22100 42220
rect 22055 42180 22100 42208
rect 22094 42168 22100 42180
rect 22152 42168 22158 42220
rect 23014 42168 23020 42220
rect 23072 42208 23078 42220
rect 23750 42208 23756 42220
rect 23072 42180 23756 42208
rect 23072 42168 23078 42180
rect 23750 42168 23756 42180
rect 23808 42168 23814 42220
rect 24394 42208 24400 42220
rect 24355 42180 24400 42208
rect 24394 42168 24400 42180
rect 24452 42168 24458 42220
rect 25590 42208 25596 42220
rect 25551 42180 25596 42208
rect 25590 42168 25596 42180
rect 25648 42168 25654 42220
rect 26973 42211 27031 42217
rect 26973 42177 26985 42211
rect 27019 42208 27031 42211
rect 27433 42211 27491 42217
rect 27433 42208 27445 42211
rect 27019 42180 27445 42208
rect 27019 42177 27031 42180
rect 26973 42171 27031 42177
rect 27433 42177 27445 42180
rect 27479 42208 27491 42211
rect 27614 42208 27620 42220
rect 27479 42180 27620 42208
rect 27479 42177 27491 42180
rect 27433 42171 27491 42177
rect 27614 42168 27620 42180
rect 27672 42168 27678 42220
rect 29638 42168 29644 42220
rect 29696 42208 29702 42220
rect 29733 42211 29791 42217
rect 29733 42208 29745 42211
rect 29696 42180 29745 42208
rect 29696 42168 29702 42180
rect 29733 42177 29745 42180
rect 29779 42177 29791 42211
rect 29733 42171 29791 42177
rect 29454 42100 29460 42152
rect 29512 42140 29518 42152
rect 30208 42140 30236 42316
rect 30653 42313 30665 42347
rect 30699 42344 30711 42347
rect 31018 42344 31024 42356
rect 30699 42316 31024 42344
rect 30699 42313 30711 42316
rect 30653 42307 30711 42313
rect 31018 42304 31024 42316
rect 31076 42304 31082 42356
rect 33091 42347 33149 42353
rect 33091 42313 33103 42347
rect 33137 42344 33149 42347
rect 33870 42344 33876 42356
rect 33137 42316 33876 42344
rect 33137 42313 33149 42316
rect 33091 42307 33149 42313
rect 33870 42304 33876 42316
rect 33928 42304 33934 42356
rect 34238 42344 34244 42356
rect 34199 42316 34244 42344
rect 34238 42304 34244 42316
rect 34296 42304 34302 42356
rect 34701 42347 34759 42353
rect 34701 42313 34713 42347
rect 34747 42344 34759 42347
rect 34790 42344 34796 42356
rect 34747 42316 34796 42344
rect 34747 42313 34759 42316
rect 34701 42307 34759 42313
rect 34790 42304 34796 42316
rect 34848 42304 34854 42356
rect 35710 42344 35716 42356
rect 35671 42316 35716 42344
rect 35710 42304 35716 42316
rect 35768 42304 35774 42356
rect 39850 42344 39856 42356
rect 35820 42316 39856 42344
rect 30374 42236 30380 42288
rect 30432 42276 30438 42288
rect 31297 42279 31355 42285
rect 31297 42276 31309 42279
rect 30432 42248 31309 42276
rect 30432 42236 30438 42248
rect 31297 42245 31309 42248
rect 31343 42245 31355 42279
rect 31297 42239 31355 42245
rect 32079 42279 32137 42285
rect 32079 42245 32091 42279
rect 32125 42276 32137 42279
rect 32125 42248 33640 42276
rect 32125 42245 32137 42248
rect 32079 42239 32137 42245
rect 30282 42168 30288 42220
rect 30340 42208 30346 42220
rect 33413 42211 33471 42217
rect 33413 42208 33425 42211
rect 30340 42180 33425 42208
rect 30340 42168 30346 42180
rect 30742 42140 30748 42152
rect 29512 42112 30097 42140
rect 30208 42112 30748 42140
rect 29512 42100 29518 42112
rect 22189 42075 22247 42081
rect 22189 42072 22201 42075
rect 21928 42044 22201 42072
rect 22189 42041 22201 42044
rect 22235 42041 22247 42075
rect 22738 42072 22744 42084
rect 22699 42044 22744 42072
rect 22189 42035 22247 42041
rect 22738 42032 22744 42044
rect 22796 42072 22802 42084
rect 23198 42072 23204 42084
rect 22796 42044 23204 42072
rect 22796 42032 22802 42044
rect 23198 42032 23204 42044
rect 23256 42032 23262 42084
rect 23845 42075 23903 42081
rect 23845 42041 23857 42075
rect 23891 42041 23903 42075
rect 25682 42072 25688 42084
rect 25595 42044 25688 42072
rect 23845 42035 23903 42041
rect 22646 42004 22652 42016
rect 21468 41976 22652 42004
rect 22646 41964 22652 41976
rect 22704 41964 22710 42016
rect 23106 42004 23112 42016
rect 23067 41976 23112 42004
rect 23106 41964 23112 41976
rect 23164 41964 23170 42016
rect 23477 42007 23535 42013
rect 23477 41973 23489 42007
rect 23523 42004 23535 42007
rect 23750 42004 23756 42016
rect 23523 41976 23756 42004
rect 23523 41973 23535 41976
rect 23477 41967 23535 41973
rect 23750 41964 23756 41976
rect 23808 42004 23814 42016
rect 23860 42004 23888 42035
rect 25682 42032 25688 42044
rect 25740 42032 25746 42084
rect 26237 42075 26295 42081
rect 26237 42041 26249 42075
rect 26283 42072 26295 42075
rect 26602 42072 26608 42084
rect 26283 42044 26608 42072
rect 26283 42041 26295 42044
rect 26237 42035 26295 42041
rect 26602 42032 26608 42044
rect 26660 42032 26666 42084
rect 27754 42075 27812 42081
rect 27754 42041 27766 42075
rect 27800 42041 27812 42075
rect 27754 42035 27812 42041
rect 28997 42075 29055 42081
rect 28997 42041 29009 42075
rect 29043 42072 29055 42075
rect 29178 42072 29184 42084
rect 29043 42044 29184 42072
rect 29043 42041 29055 42044
rect 28997 42035 29055 42041
rect 24673 42007 24731 42013
rect 24673 42004 24685 42007
rect 23808 41976 24685 42004
rect 23808 41964 23814 41976
rect 24673 41973 24685 41976
rect 24719 41973 24731 42007
rect 25700 42004 25728 42032
rect 26694 42004 26700 42016
rect 25700 41976 26700 42004
rect 24673 41967 24731 41973
rect 26694 41964 26700 41976
rect 26752 41964 26758 42016
rect 27246 42004 27252 42016
rect 27207 41976 27252 42004
rect 27246 41964 27252 41976
rect 27304 42004 27310 42016
rect 27769 42004 27797 42035
rect 29178 42032 29184 42044
rect 29236 42072 29242 42084
rect 30069 42081 30097 42112
rect 30742 42100 30748 42112
rect 30800 42100 30806 42152
rect 33035 42149 33063 42180
rect 33413 42177 33425 42180
rect 33459 42177 33471 42211
rect 33612 42208 33640 42248
rect 33686 42236 33692 42288
rect 33744 42276 33750 42288
rect 33781 42279 33839 42285
rect 33781 42276 33793 42279
rect 33744 42248 33793 42276
rect 33744 42236 33750 42248
rect 33781 42245 33793 42248
rect 33827 42245 33839 42279
rect 33781 42239 33839 42245
rect 34057 42279 34115 42285
rect 34057 42245 34069 42279
rect 34103 42276 34115 42279
rect 35618 42276 35624 42288
rect 34103 42248 35624 42276
rect 34103 42245 34115 42248
rect 34057 42239 34115 42245
rect 35618 42236 35624 42248
rect 35676 42276 35682 42288
rect 35820 42276 35848 42316
rect 39850 42304 39856 42316
rect 39908 42304 39914 42356
rect 35676 42248 35848 42276
rect 35676 42236 35682 42248
rect 35894 42236 35900 42288
rect 35952 42276 35958 42288
rect 35952 42248 39528 42276
rect 35952 42236 35958 42248
rect 35250 42208 35256 42220
rect 33612 42180 35256 42208
rect 33413 42171 33471 42177
rect 32008 42143 32066 42149
rect 32008 42109 32020 42143
rect 32054 42140 32066 42143
rect 33020 42143 33078 42149
rect 33020 42140 33032 42143
rect 32054 42112 32904 42140
rect 32998 42112 33032 42140
rect 32054 42109 32066 42112
rect 32008 42103 32066 42109
rect 30054 42075 30112 42081
rect 29236 42044 29684 42072
rect 29236 42032 29242 42044
rect 29454 42004 29460 42016
rect 27304 41976 29460 42004
rect 27304 41964 27310 41976
rect 29454 41964 29460 41976
rect 29512 42004 29518 42016
rect 29549 42007 29607 42013
rect 29549 42004 29561 42007
rect 29512 41976 29561 42004
rect 29512 41964 29518 41976
rect 29549 41973 29561 41976
rect 29595 41973 29607 42007
rect 29656 42004 29684 42044
rect 30054 42041 30066 42075
rect 30100 42041 30112 42075
rect 30054 42035 30112 42041
rect 32030 42004 32036 42016
rect 29656 41976 32036 42004
rect 29549 41967 29607 41973
rect 32030 41964 32036 41976
rect 32088 41964 32094 42016
rect 32490 42004 32496 42016
rect 32451 41976 32496 42004
rect 32490 41964 32496 41976
rect 32548 41964 32554 42016
rect 32876 42013 32904 42112
rect 33020 42109 33032 42112
rect 33066 42109 33078 42143
rect 33428 42140 33456 42171
rect 35250 42168 35256 42180
rect 35308 42168 35314 42220
rect 36357 42211 36415 42217
rect 36357 42208 36369 42211
rect 35947 42180 36369 42208
rect 34057 42143 34115 42149
rect 34057 42140 34069 42143
rect 33428 42112 34069 42140
rect 33020 42103 33078 42109
rect 34057 42109 34069 42112
rect 34103 42109 34115 42143
rect 34057 42103 34115 42109
rect 34952 42143 35010 42149
rect 34952 42109 34964 42143
rect 34998 42140 35010 42143
rect 35434 42140 35440 42152
rect 34998 42112 35440 42140
rect 34998 42109 35010 42112
rect 34952 42103 35010 42109
rect 35434 42100 35440 42112
rect 35492 42100 35498 42152
rect 35802 42100 35808 42152
rect 35860 42140 35866 42152
rect 35947 42149 35975 42180
rect 36357 42177 36369 42180
rect 36403 42177 36415 42211
rect 38470 42208 38476 42220
rect 38431 42180 38476 42208
rect 36357 42171 36415 42177
rect 38470 42168 38476 42180
rect 38528 42208 38534 42220
rect 39393 42211 39451 42217
rect 39393 42208 39405 42211
rect 38528 42180 39405 42208
rect 38528 42168 38534 42180
rect 39393 42177 39405 42180
rect 39439 42177 39451 42211
rect 39393 42171 39451 42177
rect 35932 42143 35990 42149
rect 35932 42140 35944 42143
rect 35860 42112 35944 42140
rect 35860 42100 35866 42112
rect 35932 42109 35944 42112
rect 35978 42109 35990 42143
rect 35932 42103 35990 42109
rect 36170 42100 36176 42152
rect 36228 42140 36234 42152
rect 37436 42143 37494 42149
rect 37436 42140 37448 42143
rect 36228 42112 37448 42140
rect 36228 42100 36234 42112
rect 37436 42109 37448 42112
rect 37482 42140 37494 42143
rect 39500 42140 39528 42248
rect 40532 42143 40590 42149
rect 40532 42140 40544 42143
rect 37482 42112 37964 42140
rect 39500 42112 40544 42140
rect 37482 42109 37494 42112
rect 37436 42103 37494 42109
rect 33686 42032 33692 42084
rect 33744 42072 33750 42084
rect 37936 42081 37964 42112
rect 40532 42109 40544 42112
rect 40578 42140 40590 42143
rect 40957 42143 41015 42149
rect 40957 42140 40969 42143
rect 40578 42112 40969 42140
rect 40578 42109 40590 42112
rect 40532 42103 40590 42109
rect 40957 42109 40969 42112
rect 41003 42109 41015 42143
rect 40957 42103 41015 42109
rect 36035 42075 36093 42081
rect 36035 42072 36047 42075
rect 33744 42044 36047 42072
rect 33744 42032 33750 42044
rect 36035 42041 36047 42044
rect 36081 42041 36093 42075
rect 36035 42035 36093 42041
rect 37921 42075 37979 42081
rect 37921 42041 37933 42075
rect 37967 42072 37979 42075
rect 38286 42072 38292 42084
rect 37967 42044 38292 42072
rect 37967 42041 37979 42044
rect 37921 42035 37979 42041
rect 38286 42032 38292 42044
rect 38344 42032 38350 42084
rect 38562 42072 38568 42084
rect 38523 42044 38568 42072
rect 38562 42032 38568 42044
rect 38620 42032 38626 42084
rect 39117 42075 39175 42081
rect 39117 42041 39129 42075
rect 39163 42072 39175 42075
rect 40126 42072 40132 42084
rect 39163 42044 40132 42072
rect 39163 42041 39175 42044
rect 39117 42035 39175 42041
rect 40126 42032 40132 42044
rect 40184 42032 40190 42084
rect 32861 42007 32919 42013
rect 32861 41973 32873 42007
rect 32907 42004 32919 42007
rect 32950 42004 32956 42016
rect 32907 41976 32956 42004
rect 32907 41973 32919 41976
rect 32861 41967 32919 41973
rect 32950 41964 32956 41976
rect 33008 41964 33014 42016
rect 33962 41964 33968 42016
rect 34020 42004 34026 42016
rect 35023 42007 35081 42013
rect 35023 42004 35035 42007
rect 34020 41976 35035 42004
rect 34020 41964 34026 41976
rect 35023 41973 35035 41976
rect 35069 41973 35081 42007
rect 35434 42004 35440 42016
rect 35395 41976 35440 42004
rect 35023 41967 35081 41973
rect 35434 41964 35440 41976
rect 35492 41964 35498 42016
rect 37507 42007 37565 42013
rect 37507 41973 37519 42007
rect 37553 42004 37565 42007
rect 37734 42004 37740 42016
rect 37553 41976 37740 42004
rect 37553 41973 37565 41976
rect 37507 41967 37565 41973
rect 37734 41964 37740 41976
rect 37792 41964 37798 42016
rect 38194 42004 38200 42016
rect 38155 41976 38200 42004
rect 38194 41964 38200 41976
rect 38252 41964 38258 42016
rect 40635 42007 40693 42013
rect 40635 41973 40647 42007
rect 40681 42004 40693 42007
rect 40770 42004 40776 42016
rect 40681 41976 40776 42004
rect 40681 41973 40693 41976
rect 40635 41967 40693 41973
rect 40770 41964 40776 41976
rect 40828 41964 40834 42016
rect 1104 41914 48852 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 48852 41914
rect 1104 41840 48852 41862
rect 22094 41800 22100 41812
rect 22055 41772 22100 41800
rect 22094 41760 22100 41772
rect 22152 41760 22158 41812
rect 22327 41803 22385 41809
rect 22327 41769 22339 41803
rect 22373 41800 22385 41803
rect 23474 41800 23480 41812
rect 22373 41772 23480 41800
rect 22373 41769 22385 41772
rect 22327 41763 22385 41769
rect 23474 41760 23480 41772
rect 23532 41760 23538 41812
rect 23566 41760 23572 41812
rect 23624 41800 23630 41812
rect 24213 41803 24271 41809
rect 24213 41800 24225 41803
rect 23624 41772 24225 41800
rect 23624 41760 23630 41772
rect 24213 41769 24225 41772
rect 24259 41769 24271 41803
rect 24213 41763 24271 41769
rect 25271 41803 25329 41809
rect 25271 41769 25283 41803
rect 25317 41800 25329 41803
rect 25498 41800 25504 41812
rect 25317 41772 25504 41800
rect 25317 41769 25329 41772
rect 25271 41763 25329 41769
rect 25498 41760 25504 41772
rect 25556 41760 25562 41812
rect 25682 41800 25688 41812
rect 25643 41772 25688 41800
rect 25682 41760 25688 41772
rect 25740 41760 25746 41812
rect 26234 41800 26240 41812
rect 26195 41772 26240 41800
rect 26234 41760 26240 41772
rect 26292 41760 26298 41812
rect 29638 41760 29644 41812
rect 29696 41800 29702 41812
rect 29917 41803 29975 41809
rect 29917 41800 29929 41803
rect 29696 41772 29929 41800
rect 29696 41760 29702 41772
rect 29917 41769 29929 41772
rect 29963 41769 29975 41803
rect 29917 41763 29975 41769
rect 34698 41760 34704 41812
rect 34756 41800 34762 41812
rect 34885 41803 34943 41809
rect 34885 41800 34897 41803
rect 34756 41772 34897 41800
rect 34756 41760 34762 41772
rect 34885 41769 34897 41772
rect 34931 41769 34943 41803
rect 34885 41763 34943 41769
rect 35084 41772 35388 41800
rect 21358 41692 21364 41744
rect 21416 41732 21422 41744
rect 23290 41732 23296 41744
rect 21416 41704 23296 41732
rect 21416 41692 21422 41704
rect 23290 41692 23296 41704
rect 23348 41692 23354 41744
rect 23385 41735 23443 41741
rect 23385 41701 23397 41735
rect 23431 41732 23443 41735
rect 23658 41732 23664 41744
rect 23431 41704 23664 41732
rect 23431 41701 23443 41704
rect 23385 41695 23443 41701
rect 23658 41692 23664 41704
rect 23716 41692 23722 41744
rect 23937 41735 23995 41741
rect 23937 41701 23949 41735
rect 23983 41732 23995 41735
rect 24394 41732 24400 41744
rect 23983 41704 24400 41732
rect 23983 41701 23995 41704
rect 23937 41695 23995 41701
rect 24394 41692 24400 41704
rect 24452 41692 24458 41744
rect 26694 41732 26700 41744
rect 26655 41704 26700 41732
rect 26694 41692 26700 41704
rect 26752 41692 26758 41744
rect 30650 41732 30656 41744
rect 30611 41704 30656 41732
rect 30650 41692 30656 41704
rect 30708 41692 30714 41744
rect 33686 41732 33692 41744
rect 33647 41704 33692 41732
rect 33686 41692 33692 41704
rect 33744 41692 33750 41744
rect 33781 41735 33839 41741
rect 33781 41701 33793 41735
rect 33827 41732 33839 41735
rect 34606 41732 34612 41744
rect 33827 41704 34612 41732
rect 33827 41701 33839 41704
rect 33781 41695 33839 41701
rect 34606 41692 34612 41704
rect 34664 41732 34670 41744
rect 35084 41732 35112 41772
rect 35250 41732 35256 41744
rect 34664 41704 35112 41732
rect 35211 41704 35256 41732
rect 34664 41692 34670 41704
rect 35250 41692 35256 41704
rect 35308 41692 35314 41744
rect 35360 41741 35388 41772
rect 35345 41735 35403 41741
rect 35345 41701 35357 41735
rect 35391 41701 35403 41735
rect 35345 41695 35403 41701
rect 38562 41692 38568 41744
rect 38620 41732 38626 41744
rect 38657 41735 38715 41741
rect 38657 41732 38669 41735
rect 38620 41704 38669 41732
rect 38620 41692 38626 41704
rect 38657 41701 38669 41704
rect 38703 41701 38715 41735
rect 40310 41732 40316 41744
rect 40271 41704 40316 41732
rect 38657 41695 38715 41701
rect 40310 41692 40316 41704
rect 40368 41692 40374 41744
rect 40402 41692 40408 41744
rect 40460 41732 40466 41744
rect 42242 41732 42248 41744
rect 40460 41704 42248 41732
rect 40460 41692 40466 41704
rect 42242 41692 42248 41704
rect 42300 41692 42306 41744
rect 22094 41624 22100 41676
rect 22152 41664 22158 41676
rect 22224 41667 22282 41673
rect 22224 41664 22236 41667
rect 22152 41636 22236 41664
rect 22152 41624 22158 41636
rect 22224 41633 22236 41636
rect 22270 41633 22282 41667
rect 22224 41627 22282 41633
rect 24762 41624 24768 41676
rect 24820 41664 24826 41676
rect 25200 41667 25258 41673
rect 25200 41664 25212 41667
rect 24820 41636 25212 41664
rect 24820 41624 24826 41636
rect 25200 41633 25212 41636
rect 25246 41664 25258 41667
rect 29181 41667 29239 41673
rect 25246 41636 26096 41664
rect 25246 41633 25258 41636
rect 25200 41627 25258 41633
rect 26068 41528 26096 41636
rect 29181 41633 29193 41667
rect 29227 41664 29239 41667
rect 29270 41664 29276 41676
rect 29227 41636 29276 41664
rect 29227 41633 29239 41636
rect 29181 41627 29239 41633
rect 29270 41624 29276 41636
rect 29328 41624 29334 41676
rect 29457 41667 29515 41673
rect 29457 41633 29469 41667
rect 29503 41664 29515 41667
rect 29546 41664 29552 41676
rect 29503 41636 29552 41664
rect 29503 41633 29515 41636
rect 29457 41627 29515 41633
rect 26602 41596 26608 41608
rect 26563 41568 26608 41596
rect 26602 41556 26608 41568
rect 26660 41556 26666 41608
rect 26878 41596 26884 41608
rect 26839 41568 26884 41596
rect 26878 41556 26884 41568
rect 26936 41556 26942 41608
rect 28813 41599 28871 41605
rect 28813 41565 28825 41599
rect 28859 41596 28871 41599
rect 29472 41596 29500 41627
rect 29546 41624 29552 41636
rect 29604 41624 29610 41676
rect 32306 41624 32312 41676
rect 32364 41664 32370 41676
rect 32620 41667 32678 41673
rect 32620 41664 32632 41667
rect 32364 41636 32632 41664
rect 32364 41624 32370 41636
rect 32620 41633 32632 41636
rect 32666 41633 32678 41667
rect 32620 41627 32678 41633
rect 41852 41667 41910 41673
rect 41852 41633 41864 41667
rect 41898 41664 41910 41667
rect 42058 41664 42064 41676
rect 41898 41636 42064 41664
rect 41898 41633 41910 41636
rect 41852 41627 41910 41633
rect 42058 41624 42064 41636
rect 42116 41664 42122 41676
rect 46934 41664 46940 41676
rect 42116 41636 46940 41664
rect 42116 41624 42122 41636
rect 46934 41624 46940 41636
rect 46992 41624 46998 41676
rect 28859 41568 29500 41596
rect 29641 41599 29699 41605
rect 28859 41565 28871 41568
rect 28813 41559 28871 41565
rect 29641 41565 29653 41599
rect 29687 41596 29699 41599
rect 30098 41596 30104 41608
rect 29687 41568 30104 41596
rect 29687 41565 29699 41568
rect 29641 41559 29699 41565
rect 30098 41556 30104 41568
rect 30156 41596 30162 41608
rect 30285 41599 30343 41605
rect 30285 41596 30297 41599
rect 30156 41568 30297 41596
rect 30156 41556 30162 41568
rect 30285 41565 30297 41568
rect 30331 41565 30343 41599
rect 30558 41596 30564 41608
rect 30519 41568 30564 41596
rect 30285 41559 30343 41565
rect 30558 41556 30564 41568
rect 30616 41556 30622 41608
rect 31205 41599 31263 41605
rect 31205 41565 31217 41599
rect 31251 41596 31263 41599
rect 32214 41596 32220 41608
rect 31251 41568 32220 41596
rect 31251 41565 31263 41568
rect 31205 41559 31263 41565
rect 32214 41556 32220 41568
rect 32272 41556 32278 41608
rect 34054 41596 34060 41608
rect 34015 41568 34060 41596
rect 34054 41556 34060 41568
rect 34112 41556 34118 41608
rect 35526 41596 35532 41608
rect 35487 41568 35532 41596
rect 35526 41556 35532 41568
rect 35584 41556 35590 41608
rect 38562 41596 38568 41608
rect 38523 41568 38568 41596
rect 38562 41556 38568 41568
rect 38620 41556 38626 41608
rect 40126 41556 40132 41608
rect 40184 41596 40190 41608
rect 40589 41599 40647 41605
rect 40589 41596 40601 41599
rect 40184 41568 40601 41596
rect 40184 41556 40190 41568
rect 40589 41565 40601 41568
rect 40635 41565 40647 41599
rect 40589 41559 40647 41565
rect 30834 41528 30840 41540
rect 26068 41500 30840 41528
rect 30834 41488 30840 41500
rect 30892 41488 30898 41540
rect 38654 41488 38660 41540
rect 38712 41528 38718 41540
rect 39117 41531 39175 41537
rect 39117 41528 39129 41531
rect 38712 41500 39129 41528
rect 38712 41488 38718 41500
rect 39117 41497 39129 41500
rect 39163 41528 39175 41531
rect 40862 41528 40868 41540
rect 39163 41500 40868 41528
rect 39163 41497 39175 41500
rect 39117 41491 39175 41497
rect 40862 41488 40868 41500
rect 40920 41488 40926 41540
rect 32723 41463 32781 41469
rect 32723 41429 32735 41463
rect 32769 41460 32781 41463
rect 33410 41460 33416 41472
rect 32769 41432 33416 41460
rect 32769 41429 32781 41432
rect 32723 41423 32781 41429
rect 33410 41420 33416 41432
rect 33468 41420 33474 41472
rect 36630 41460 36636 41472
rect 36591 41432 36636 41460
rect 36630 41420 36636 41432
rect 36688 41420 36694 41472
rect 41923 41463 41981 41469
rect 41923 41429 41935 41463
rect 41969 41460 41981 41463
rect 42150 41460 42156 41472
rect 41969 41432 42156 41460
rect 41969 41429 41981 41432
rect 41923 41423 41981 41429
rect 42150 41420 42156 41432
rect 42208 41420 42214 41472
rect 1104 41370 48852 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 48852 41370
rect 1104 41296 48852 41318
rect 23293 41259 23351 41265
rect 23293 41225 23305 41259
rect 23339 41256 23351 41259
rect 23474 41256 23480 41268
rect 23339 41228 23480 41256
rect 23339 41225 23351 41228
rect 23293 41219 23351 41225
rect 23474 41216 23480 41228
rect 23532 41256 23538 41268
rect 23658 41256 23664 41268
rect 23532 41228 23664 41256
rect 23532 41216 23538 41228
rect 23658 41216 23664 41228
rect 23716 41256 23722 41268
rect 23842 41256 23848 41268
rect 23716 41228 23848 41256
rect 23716 41216 23722 41228
rect 23842 41216 23848 41228
rect 23900 41216 23906 41268
rect 24762 41256 24768 41268
rect 24723 41228 24768 41256
rect 24762 41216 24768 41228
rect 24820 41216 24826 41268
rect 26602 41216 26608 41268
rect 26660 41256 26666 41268
rect 28169 41259 28227 41265
rect 28169 41256 28181 41259
rect 26660 41228 28181 41256
rect 26660 41216 26666 41228
rect 28169 41225 28181 41228
rect 28215 41225 28227 41259
rect 28169 41219 28227 41225
rect 29454 41216 29460 41268
rect 29512 41256 29518 41268
rect 29917 41259 29975 41265
rect 29917 41256 29929 41259
rect 29512 41228 29929 41256
rect 29512 41216 29518 41228
rect 29917 41225 29929 41228
rect 29963 41256 29975 41259
rect 29963 41228 30512 41256
rect 29963 41225 29975 41228
rect 29917 41219 29975 41225
rect 19242 41148 19248 41200
rect 19300 41188 19306 41200
rect 24780 41188 24808 41216
rect 19300 41160 24808 41188
rect 26513 41191 26571 41197
rect 19300 41148 19306 41160
rect 23124 41064 23152 41160
rect 26513 41157 26525 41191
rect 26559 41188 26571 41191
rect 26694 41188 26700 41200
rect 26559 41160 26700 41188
rect 26559 41157 26571 41160
rect 26513 41151 26571 41157
rect 26694 41148 26700 41160
rect 26752 41188 26758 41200
rect 27893 41191 27951 41197
rect 27893 41188 27905 41191
rect 26752 41160 27905 41188
rect 26752 41148 26758 41160
rect 27893 41157 27905 41160
rect 27939 41157 27951 41191
rect 27893 41151 27951 41157
rect 23842 41080 23848 41132
rect 23900 41120 23906 41132
rect 25041 41123 25099 41129
rect 25041 41120 25053 41123
rect 23900 41092 25053 41120
rect 23900 41080 23906 41092
rect 25041 41089 25053 41092
rect 25087 41089 25099 41123
rect 25041 41083 25099 41089
rect 26973 41123 27031 41129
rect 26973 41089 26985 41123
rect 27019 41120 27031 41123
rect 27338 41120 27344 41132
rect 27019 41092 27344 41120
rect 27019 41089 27031 41092
rect 26973 41083 27031 41089
rect 19058 41012 19064 41064
rect 19116 41052 19122 41064
rect 21856 41055 21914 41061
rect 21856 41052 21868 41055
rect 19116 41024 21868 41052
rect 19116 41012 19122 41024
rect 21856 41021 21868 41024
rect 21902 41052 21914 41055
rect 22281 41055 22339 41061
rect 22281 41052 22293 41055
rect 21902 41024 22293 41052
rect 21902 41021 21914 41024
rect 21856 41015 21914 41021
rect 22281 41021 22293 41024
rect 22327 41052 22339 41055
rect 22327 41024 22876 41052
rect 22327 41021 22339 41024
rect 22281 41015 22339 41021
rect 21959 40987 22017 40993
rect 21959 40953 21971 40987
rect 22005 40984 22017 40987
rect 22462 40984 22468 40996
rect 22005 40956 22468 40984
rect 22005 40953 22017 40956
rect 21959 40947 22017 40953
rect 22462 40944 22468 40956
rect 22520 40944 22526 40996
rect 22094 40876 22100 40928
rect 22152 40916 22158 40928
rect 22649 40919 22707 40925
rect 22649 40916 22661 40919
rect 22152 40888 22661 40916
rect 22152 40876 22158 40888
rect 22649 40885 22661 40888
rect 22695 40885 22707 40919
rect 22848 40916 22876 41024
rect 23106 41012 23112 41064
rect 23164 41012 23170 41064
rect 23198 41012 23204 41064
rect 23256 41052 23262 41064
rect 23728 41055 23786 41061
rect 23728 41052 23740 41055
rect 23256 41024 23740 41052
rect 23256 41012 23262 41024
rect 23728 41021 23740 41024
rect 23774 41052 23786 41055
rect 24121 41055 24179 41061
rect 24121 41052 24133 41055
rect 23774 41024 24133 41052
rect 23774 41021 23786 41024
rect 23728 41015 23786 41021
rect 24121 41021 24133 41024
rect 24167 41021 24179 41055
rect 24121 41015 24179 41021
rect 23934 40984 23940 40996
rect 23446 40956 23940 40984
rect 23446 40916 23474 40956
rect 23934 40944 23940 40956
rect 23992 40944 23998 40996
rect 25056 40984 25084 41083
rect 27338 41080 27344 41092
rect 27396 41080 27402 41132
rect 30098 41120 30104 41132
rect 30059 41092 30104 41120
rect 30098 41080 30104 41092
rect 30156 41080 30162 41132
rect 25222 41052 25228 41064
rect 25183 41024 25228 41052
rect 25222 41012 25228 41024
rect 25280 41012 25286 41064
rect 30484 40996 30512 41228
rect 30650 41216 30656 41268
rect 30708 41256 30714 41268
rect 31021 41259 31079 41265
rect 31021 41256 31033 41259
rect 30708 41228 31033 41256
rect 30708 41216 30714 41228
rect 31021 41225 31033 41228
rect 31067 41256 31079 41259
rect 31297 41259 31355 41265
rect 31297 41256 31309 41259
rect 31067 41228 31309 41256
rect 31067 41225 31079 41228
rect 31021 41219 31079 41225
rect 31297 41225 31309 41228
rect 31343 41225 31355 41259
rect 31297 41219 31355 41225
rect 33321 41259 33379 41265
rect 33321 41225 33333 41259
rect 33367 41256 33379 41259
rect 33686 41256 33692 41268
rect 33367 41228 33692 41256
rect 33367 41225 33379 41228
rect 33321 41219 33379 41225
rect 33686 41216 33692 41228
rect 33744 41216 33750 41268
rect 37734 41216 37740 41268
rect 37792 41256 37798 41268
rect 37829 41259 37887 41265
rect 37829 41256 37841 41259
rect 37792 41228 37841 41256
rect 37792 41216 37798 41228
rect 37829 41225 37841 41228
rect 37875 41256 37887 41259
rect 37875 41228 38516 41256
rect 37875 41225 37887 41228
rect 37829 41219 37887 41225
rect 30558 41148 30564 41200
rect 30616 41188 30622 41200
rect 35526 41188 35532 41200
rect 30616 41160 35532 41188
rect 30616 41148 30622 41160
rect 31662 41080 31668 41132
rect 31720 41120 31726 41132
rect 31938 41120 31944 41132
rect 31720 41092 31944 41120
rect 31720 41080 31726 41092
rect 31938 41080 31944 41092
rect 31996 41080 32002 41132
rect 32214 41120 32220 41132
rect 32175 41092 32220 41120
rect 32214 41080 32220 41092
rect 32272 41080 32278 41132
rect 34698 41080 34704 41132
rect 34756 41120 34762 41132
rect 35268 41129 35296 41160
rect 35526 41148 35532 41160
rect 35584 41148 35590 41200
rect 38488 41129 38516 41228
rect 34977 41123 35035 41129
rect 34977 41120 34989 41123
rect 34756 41092 34989 41120
rect 34756 41080 34762 41092
rect 34977 41089 34989 41092
rect 35023 41089 35035 41123
rect 34977 41083 35035 41089
rect 35253 41123 35311 41129
rect 35253 41089 35265 41123
rect 35299 41089 35311 41123
rect 35253 41083 35311 41089
rect 38473 41123 38531 41129
rect 38473 41089 38485 41123
rect 38519 41089 38531 41123
rect 38473 41083 38531 41089
rect 38562 41080 38568 41132
rect 38620 41120 38626 41132
rect 39393 41123 39451 41129
rect 39393 41120 39405 41123
rect 38620 41092 39405 41120
rect 38620 41080 38626 41092
rect 39393 41089 39405 41092
rect 39439 41089 39451 41123
rect 39393 41083 39451 41089
rect 40589 41123 40647 41129
rect 40589 41089 40601 41123
rect 40635 41120 40647 41123
rect 40770 41120 40776 41132
rect 40635 41092 40776 41120
rect 40635 41089 40647 41092
rect 40589 41083 40647 41089
rect 40770 41080 40776 41092
rect 40828 41080 40834 41132
rect 40862 41080 40868 41132
rect 40920 41120 40926 41132
rect 42426 41120 42432 41132
rect 40920 41092 40965 41120
rect 42387 41092 42432 41120
rect 40920 41080 40926 41092
rect 42426 41080 42432 41092
rect 42484 41080 42490 41132
rect 32766 41012 32772 41064
rect 32824 41052 32830 41064
rect 33480 41055 33538 41061
rect 33480 41052 33492 41055
rect 32824 41024 33492 41052
rect 32824 41012 32830 41024
rect 33480 41021 33492 41024
rect 33526 41052 33538 41055
rect 33873 41055 33931 41061
rect 33873 41052 33885 41055
rect 33526 41024 33885 41052
rect 33526 41021 33538 41024
rect 33480 41015 33538 41021
rect 33873 41021 33885 41024
rect 33919 41021 33931 41055
rect 36630 41052 36636 41064
rect 36591 41024 36636 41052
rect 33873 41015 33931 41021
rect 36630 41012 36636 41024
rect 36688 41012 36694 41064
rect 37553 41055 37611 41061
rect 36924 41024 37044 41052
rect 25546 40987 25604 40993
rect 25546 40984 25558 40987
rect 25056 40956 25558 40984
rect 25546 40953 25558 40956
rect 25592 40984 25604 40987
rect 26789 40987 26847 40993
rect 26789 40984 26801 40987
rect 25592 40956 26801 40984
rect 25592 40953 25604 40956
rect 25546 40947 25604 40953
rect 26789 40953 26801 40956
rect 26835 40984 26847 40987
rect 27246 40984 27252 40996
rect 26835 40956 27252 40984
rect 26835 40953 26847 40956
rect 26789 40947 26847 40953
rect 27246 40944 27252 40956
rect 27304 40993 27310 40996
rect 30466 40993 30472 40996
rect 27304 40987 27352 40993
rect 27304 40953 27306 40987
rect 27340 40953 27352 40987
rect 27304 40947 27352 40953
rect 30423 40987 30472 40993
rect 30423 40953 30435 40987
rect 30469 40953 30472 40987
rect 30423 40947 30472 40953
rect 27304 40944 27310 40947
rect 30466 40944 30472 40947
rect 30524 40984 30530 40996
rect 32033 40987 32091 40993
rect 30524 40956 30617 40984
rect 30524 40944 30530 40956
rect 32033 40953 32045 40987
rect 32079 40953 32091 40987
rect 32033 40947 32091 40953
rect 22848 40888 23474 40916
rect 23799 40919 23857 40925
rect 22649 40879 22707 40885
rect 23799 40885 23811 40919
rect 23845 40916 23857 40919
rect 24578 40916 24584 40928
rect 23845 40888 24584 40916
rect 23845 40885 23857 40888
rect 23799 40879 23857 40885
rect 24578 40876 24584 40888
rect 24636 40876 24642 40928
rect 25682 40876 25688 40928
rect 25740 40916 25746 40928
rect 26145 40919 26203 40925
rect 26145 40916 26157 40919
rect 25740 40888 26157 40916
rect 25740 40876 25746 40888
rect 26145 40885 26157 40888
rect 26191 40885 26203 40919
rect 26145 40879 26203 40885
rect 28997 40919 29055 40925
rect 28997 40885 29009 40919
rect 29043 40916 29055 40919
rect 29270 40916 29276 40928
rect 29043 40888 29276 40916
rect 29043 40885 29055 40888
rect 28997 40879 29055 40885
rect 29270 40876 29276 40888
rect 29328 40876 29334 40928
rect 29546 40916 29552 40928
rect 29507 40888 29552 40916
rect 29546 40876 29552 40888
rect 29604 40876 29610 40928
rect 31662 40916 31668 40928
rect 31623 40888 31668 40916
rect 31662 40876 31668 40888
rect 31720 40916 31726 40928
rect 32048 40916 32076 40947
rect 33686 40944 33692 40996
rect 33744 40984 33750 40996
rect 34701 40987 34759 40993
rect 34701 40984 34713 40987
rect 33744 40956 34713 40984
rect 33744 40944 33750 40956
rect 34701 40953 34713 40956
rect 34747 40984 34759 40987
rect 35069 40987 35127 40993
rect 35069 40984 35081 40987
rect 34747 40956 35081 40984
rect 34747 40953 34759 40956
rect 34701 40947 34759 40953
rect 35069 40953 35081 40956
rect 35115 40953 35127 40987
rect 35069 40947 35127 40953
rect 31720 40888 32076 40916
rect 31720 40876 31726 40888
rect 32306 40876 32312 40928
rect 32364 40916 32370 40928
rect 32861 40919 32919 40925
rect 32861 40916 32873 40919
rect 32364 40888 32873 40916
rect 32364 40876 32370 40888
rect 32861 40885 32873 40888
rect 32907 40885 32919 40919
rect 32861 40879 32919 40885
rect 33318 40876 33324 40928
rect 33376 40916 33382 40928
rect 33551 40919 33609 40925
rect 33551 40916 33563 40919
rect 33376 40888 33563 40916
rect 33376 40876 33382 40888
rect 33551 40885 33563 40888
rect 33597 40885 33609 40919
rect 33551 40879 33609 40885
rect 34333 40919 34391 40925
rect 34333 40885 34345 40919
rect 34379 40916 34391 40919
rect 34606 40916 34612 40928
rect 34379 40888 34612 40916
rect 34379 40885 34391 40888
rect 34333 40879 34391 40885
rect 34606 40876 34612 40888
rect 34664 40916 34670 40928
rect 35897 40919 35955 40925
rect 35897 40916 35909 40919
rect 34664 40888 35909 40916
rect 34664 40876 34670 40888
rect 35897 40885 35909 40888
rect 35943 40885 35955 40919
rect 36538 40916 36544 40928
rect 36499 40888 36544 40916
rect 35897 40879 35955 40885
rect 36538 40876 36544 40888
rect 36596 40916 36602 40928
rect 36924 40916 36952 41024
rect 37016 40993 37044 41024
rect 37553 41021 37565 41055
rect 37599 41052 37611 41055
rect 37599 41024 38332 41052
rect 37599 41021 37611 41024
rect 37553 41015 37611 41021
rect 38304 40993 38332 41024
rect 36995 40987 37053 40993
rect 36995 40953 37007 40987
rect 37041 40953 37053 40987
rect 36995 40947 37053 40953
rect 38289 40987 38347 40993
rect 38289 40953 38301 40987
rect 38335 40984 38347 40987
rect 38470 40984 38476 40996
rect 38335 40956 38476 40984
rect 38335 40953 38347 40956
rect 38289 40947 38347 40953
rect 38470 40944 38476 40956
rect 38528 40984 38534 40996
rect 38565 40987 38623 40993
rect 38565 40984 38577 40987
rect 38528 40956 38577 40984
rect 38528 40944 38534 40956
rect 38565 40953 38577 40956
rect 38611 40953 38623 40987
rect 39114 40984 39120 40996
rect 39075 40956 39120 40984
rect 38565 40947 38623 40953
rect 39114 40944 39120 40956
rect 39172 40944 39178 40996
rect 40681 40987 40739 40993
rect 40681 40953 40693 40987
rect 40727 40953 40739 40987
rect 40681 40947 40739 40953
rect 39942 40916 39948 40928
rect 36596 40888 36952 40916
rect 39903 40888 39948 40916
rect 36596 40876 36602 40888
rect 39942 40876 39948 40888
rect 40000 40916 40006 40928
rect 40221 40919 40279 40925
rect 40221 40916 40233 40919
rect 40000 40888 40233 40916
rect 40000 40876 40006 40888
rect 40221 40885 40233 40888
rect 40267 40916 40279 40919
rect 40402 40916 40408 40928
rect 40267 40888 40408 40916
rect 40267 40885 40279 40888
rect 40221 40879 40279 40885
rect 40402 40876 40408 40888
rect 40460 40916 40466 40928
rect 40696 40916 40724 40947
rect 41690 40944 41696 40996
rect 41748 40984 41754 40996
rect 42153 40987 42211 40993
rect 42153 40984 42165 40987
rect 41748 40956 42165 40984
rect 41748 40944 41754 40956
rect 42153 40953 42165 40956
rect 42199 40953 42211 40987
rect 42153 40947 42211 40953
rect 40460 40888 40724 40916
rect 41877 40919 41935 40925
rect 40460 40876 40466 40888
rect 41877 40885 41889 40919
rect 41923 40916 41935 40919
rect 42058 40916 42064 40928
rect 41923 40888 42064 40916
rect 41923 40885 41935 40888
rect 41877 40879 41935 40885
rect 42058 40876 42064 40888
rect 42116 40876 42122 40928
rect 42168 40916 42196 40947
rect 42242 40944 42248 40996
rect 42300 40984 42306 40996
rect 42300 40956 42345 40984
rect 42300 40944 42306 40956
rect 43073 40919 43131 40925
rect 43073 40916 43085 40919
rect 42168 40888 43085 40916
rect 43073 40885 43085 40888
rect 43119 40885 43131 40919
rect 43073 40879 43131 40885
rect 1104 40826 48852 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 48852 40826
rect 1104 40752 48852 40774
rect 23290 40672 23296 40724
rect 23348 40712 23354 40724
rect 23385 40715 23443 40721
rect 23385 40712 23397 40715
rect 23348 40684 23397 40712
rect 23348 40672 23354 40684
rect 23385 40681 23397 40684
rect 23431 40681 23443 40715
rect 23385 40675 23443 40681
rect 25222 40672 25228 40724
rect 25280 40712 25286 40724
rect 25317 40715 25375 40721
rect 25317 40712 25329 40715
rect 25280 40684 25329 40712
rect 25280 40672 25286 40684
rect 25317 40681 25329 40684
rect 25363 40712 25375 40715
rect 27433 40715 27491 40721
rect 27433 40712 27445 40715
rect 25363 40684 27445 40712
rect 25363 40681 25375 40684
rect 25317 40675 25375 40681
rect 27433 40681 27445 40684
rect 27479 40681 27491 40715
rect 27433 40675 27491 40681
rect 29917 40715 29975 40721
rect 29917 40681 29929 40715
rect 29963 40712 29975 40715
rect 30558 40712 30564 40724
rect 29963 40684 30564 40712
rect 29963 40681 29975 40684
rect 29917 40675 29975 40681
rect 30558 40672 30564 40684
rect 30616 40672 30622 40724
rect 30929 40715 30987 40721
rect 30929 40681 30941 40715
rect 30975 40712 30987 40715
rect 31662 40712 31668 40724
rect 30975 40684 31668 40712
rect 30975 40681 30987 40684
rect 30929 40675 30987 40681
rect 31662 40672 31668 40684
rect 31720 40672 31726 40724
rect 31938 40712 31944 40724
rect 31899 40684 31944 40712
rect 31938 40672 31944 40684
rect 31996 40672 32002 40724
rect 32030 40672 32036 40724
rect 32088 40712 32094 40724
rect 32088 40684 35204 40712
rect 32088 40672 32094 40684
rect 22557 40647 22615 40653
rect 22557 40613 22569 40647
rect 22603 40644 22615 40647
rect 22922 40644 22928 40656
rect 22603 40616 22928 40644
rect 22603 40613 22615 40616
rect 22557 40607 22615 40613
rect 22922 40604 22928 40616
rect 22980 40604 22986 40656
rect 24121 40647 24179 40653
rect 24121 40613 24133 40647
rect 24167 40644 24179 40647
rect 24486 40644 24492 40656
rect 24167 40616 24492 40644
rect 24167 40613 24179 40616
rect 24121 40607 24179 40613
rect 24486 40604 24492 40616
rect 24544 40604 24550 40656
rect 30371 40647 30429 40653
rect 30371 40613 30383 40647
rect 30417 40644 30429 40647
rect 30466 40644 30472 40656
rect 30417 40616 30472 40644
rect 30417 40613 30429 40616
rect 30371 40607 30429 40613
rect 30466 40604 30472 40616
rect 30524 40604 30530 40656
rect 33410 40644 33416 40656
rect 33371 40616 33416 40644
rect 33410 40604 33416 40616
rect 33468 40604 33474 40656
rect 33505 40647 33563 40653
rect 33505 40613 33517 40647
rect 33551 40644 33563 40647
rect 33686 40644 33692 40656
rect 33551 40616 33692 40644
rect 33551 40613 33563 40616
rect 33505 40607 33563 40613
rect 33686 40604 33692 40616
rect 33744 40604 33750 40656
rect 34054 40644 34060 40656
rect 34015 40616 34060 40644
rect 34054 40604 34060 40616
rect 34112 40604 34118 40656
rect 21174 40536 21180 40588
rect 21232 40576 21238 40588
rect 21396 40579 21454 40585
rect 21396 40576 21408 40579
rect 21232 40548 21408 40576
rect 21232 40536 21238 40548
rect 21396 40545 21408 40548
rect 21442 40545 21454 40579
rect 27614 40576 27620 40588
rect 27575 40548 27620 40576
rect 21396 40539 21454 40545
rect 27614 40536 27620 40548
rect 27672 40536 27678 40588
rect 27893 40579 27951 40585
rect 27893 40545 27905 40579
rect 27939 40576 27951 40579
rect 27982 40576 27988 40588
rect 27939 40548 27988 40576
rect 27939 40545 27951 40548
rect 27893 40539 27951 40545
rect 27982 40536 27988 40548
rect 28040 40536 28046 40588
rect 28718 40536 28724 40588
rect 28776 40576 28782 40588
rect 28997 40579 29055 40585
rect 28997 40576 29009 40579
rect 28776 40548 29009 40576
rect 28776 40536 28782 40548
rect 28997 40545 29009 40548
rect 29043 40545 29055 40579
rect 32122 40576 32128 40588
rect 28997 40539 29055 40545
rect 29196 40548 32128 40576
rect 22462 40508 22468 40520
rect 22423 40480 22468 40508
rect 22462 40468 22468 40480
rect 22520 40468 22526 40520
rect 22738 40508 22744 40520
rect 22699 40480 22744 40508
rect 22738 40468 22744 40480
rect 22796 40468 22802 40520
rect 24029 40511 24087 40517
rect 24029 40508 24041 40511
rect 23446 40480 24041 40508
rect 21499 40443 21557 40449
rect 21499 40409 21511 40443
rect 21545 40440 21557 40443
rect 23290 40440 23296 40452
rect 21545 40412 23296 40440
rect 21545 40409 21557 40412
rect 21499 40403 21557 40409
rect 23290 40400 23296 40412
rect 23348 40440 23354 40452
rect 23446 40440 23474 40480
rect 24029 40477 24041 40480
rect 24075 40477 24087 40511
rect 24394 40508 24400 40520
rect 24355 40480 24400 40508
rect 24029 40471 24087 40477
rect 24394 40468 24400 40480
rect 24452 40468 24458 40520
rect 29196 40449 29224 40548
rect 32122 40536 32128 40548
rect 32180 40536 32186 40588
rect 34790 40536 34796 40588
rect 34848 40576 34854 40588
rect 34920 40579 34978 40585
rect 34920 40576 34932 40579
rect 34848 40548 34932 40576
rect 34848 40536 34854 40548
rect 34920 40545 34932 40548
rect 34966 40545 34978 40579
rect 35176 40576 35204 40684
rect 35250 40672 35256 40724
rect 35308 40712 35314 40724
rect 35713 40715 35771 40721
rect 35713 40712 35725 40715
rect 35308 40684 35725 40712
rect 35308 40672 35314 40684
rect 35713 40681 35725 40684
rect 35759 40681 35771 40715
rect 35713 40675 35771 40681
rect 38243 40715 38301 40721
rect 38243 40681 38255 40715
rect 38289 40712 38301 40715
rect 38562 40712 38568 40724
rect 38289 40684 38568 40712
rect 38289 40681 38301 40684
rect 38243 40675 38301 40681
rect 38562 40672 38568 40684
rect 38620 40672 38626 40724
rect 40310 40672 40316 40724
rect 40368 40712 40374 40724
rect 40405 40715 40463 40721
rect 40405 40712 40417 40715
rect 40368 40684 40417 40712
rect 40368 40672 40374 40684
rect 40405 40681 40417 40684
rect 40451 40681 40463 40715
rect 40770 40712 40776 40724
rect 40731 40684 40776 40712
rect 40405 40675 40463 40681
rect 40770 40672 40776 40684
rect 40828 40672 40834 40724
rect 42150 40672 42156 40724
rect 42208 40712 42214 40724
rect 43254 40712 43260 40724
rect 42208 40684 43260 40712
rect 42208 40672 42214 40684
rect 43254 40672 43260 40684
rect 43312 40712 43318 40724
rect 43533 40715 43591 40721
rect 43533 40712 43545 40715
rect 43312 40684 43545 40712
rect 43312 40672 43318 40684
rect 43533 40681 43545 40684
rect 43579 40681 43591 40715
rect 43533 40675 43591 40681
rect 36630 40644 36636 40656
rect 36591 40616 36636 40644
rect 36630 40604 36636 40616
rect 36688 40604 36694 40656
rect 40083 40647 40141 40653
rect 40083 40613 40095 40647
rect 40129 40644 40141 40647
rect 41690 40644 41696 40656
rect 40129 40616 41696 40644
rect 40129 40613 40141 40616
rect 40083 40607 40141 40613
rect 41690 40604 41696 40616
rect 41748 40604 41754 40656
rect 41782 40604 41788 40656
rect 41840 40644 41846 40656
rect 42337 40647 42395 40653
rect 41840 40616 41885 40644
rect 41840 40604 41846 40616
rect 42337 40613 42349 40647
rect 42383 40644 42395 40647
rect 42426 40644 42432 40656
rect 42383 40616 42432 40644
rect 42383 40613 42395 40616
rect 42337 40607 42395 40613
rect 42426 40604 42432 40616
rect 42484 40604 42490 40656
rect 35897 40579 35955 40585
rect 35897 40576 35909 40579
rect 35176 40548 35909 40576
rect 34920 40539 34978 40545
rect 35897 40545 35909 40548
rect 35943 40576 35955 40579
rect 36262 40576 36268 40588
rect 35943 40548 36268 40576
rect 35943 40545 35955 40548
rect 35897 40539 35955 40545
rect 36262 40536 36268 40548
rect 36320 40536 36326 40588
rect 36357 40579 36415 40585
rect 36357 40545 36369 40579
rect 36403 40545 36415 40579
rect 36357 40539 36415 40545
rect 30006 40508 30012 40520
rect 29967 40480 30012 40508
rect 30006 40468 30012 40480
rect 30064 40468 30070 40520
rect 35437 40511 35495 40517
rect 35437 40477 35449 40511
rect 35483 40508 35495 40511
rect 35710 40508 35716 40520
rect 35483 40480 35716 40508
rect 35483 40477 35495 40480
rect 35437 40471 35495 40477
rect 35710 40468 35716 40480
rect 35768 40508 35774 40520
rect 36372 40508 36400 40539
rect 38010 40536 38016 40588
rect 38068 40576 38074 40588
rect 38140 40579 38198 40585
rect 38140 40576 38152 40579
rect 38068 40548 38152 40576
rect 38068 40536 38074 40548
rect 38140 40545 38152 40548
rect 38186 40545 38198 40579
rect 38140 40539 38198 40545
rect 38470 40536 38476 40588
rect 38528 40576 38534 40588
rect 38565 40579 38623 40585
rect 38565 40576 38577 40579
rect 38528 40548 38577 40576
rect 38528 40536 38534 40548
rect 38565 40545 38577 40548
rect 38611 40545 38623 40579
rect 38565 40539 38623 40545
rect 39758 40536 39764 40588
rect 39816 40576 39822 40588
rect 39980 40579 40038 40585
rect 39980 40576 39992 40579
rect 39816 40548 39992 40576
rect 39816 40536 39822 40548
rect 39980 40545 39992 40548
rect 40026 40545 40038 40579
rect 39980 40539 40038 40545
rect 41693 40511 41751 40517
rect 41693 40508 41705 40511
rect 35768 40480 36400 40508
rect 41616 40480 41705 40508
rect 35768 40468 35774 40480
rect 41616 40452 41644 40480
rect 41693 40477 41705 40480
rect 41739 40477 41751 40511
rect 41693 40471 41751 40477
rect 23348 40412 23474 40440
rect 29181 40443 29239 40449
rect 23348 40400 23354 40412
rect 29181 40409 29193 40443
rect 29227 40409 29239 40443
rect 29181 40403 29239 40409
rect 29270 40400 29276 40452
rect 29328 40440 29334 40452
rect 33134 40440 33140 40452
rect 29328 40412 33140 40440
rect 29328 40400 29334 40412
rect 33134 40400 33140 40412
rect 33192 40400 33198 40452
rect 41598 40400 41604 40452
rect 41656 40400 41662 40452
rect 27065 40375 27123 40381
rect 27065 40341 27077 40375
rect 27111 40372 27123 40375
rect 27338 40372 27344 40384
rect 27111 40344 27344 40372
rect 27111 40341 27123 40344
rect 27065 40335 27123 40341
rect 27338 40332 27344 40344
rect 27396 40332 27402 40384
rect 29546 40372 29552 40384
rect 29507 40344 29552 40372
rect 29546 40332 29552 40344
rect 29604 40372 29610 40384
rect 31205 40375 31263 40381
rect 31205 40372 31217 40375
rect 29604 40344 31217 40372
rect 29604 40332 29610 40344
rect 31205 40341 31217 40344
rect 31251 40372 31263 40375
rect 31294 40372 31300 40384
rect 31251 40344 31300 40372
rect 31251 40341 31263 40344
rect 31205 40335 31263 40341
rect 31294 40332 31300 40344
rect 31352 40372 31358 40384
rect 32309 40375 32367 40381
rect 32309 40372 32321 40375
rect 31352 40344 32321 40372
rect 31352 40332 31358 40344
rect 32309 40341 32321 40344
rect 32355 40341 32367 40375
rect 32309 40335 32367 40341
rect 33686 40332 33692 40384
rect 33744 40372 33750 40384
rect 35023 40375 35081 40381
rect 35023 40372 35035 40375
rect 33744 40344 35035 40372
rect 33744 40332 33750 40344
rect 35023 40341 35035 40344
rect 35069 40341 35081 40375
rect 35023 40335 35081 40341
rect 38746 40332 38752 40384
rect 38804 40372 38810 40384
rect 38933 40375 38991 40381
rect 38933 40372 38945 40375
rect 38804 40344 38945 40372
rect 38804 40332 38810 40344
rect 38933 40341 38945 40344
rect 38979 40341 38991 40375
rect 38933 40335 38991 40341
rect 41509 40375 41567 40381
rect 41509 40341 41521 40375
rect 41555 40372 41567 40375
rect 41690 40372 41696 40384
rect 41555 40344 41696 40372
rect 41555 40341 41567 40344
rect 41509 40335 41567 40341
rect 41690 40332 41696 40344
rect 41748 40332 41754 40384
rect 1104 40282 48852 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 48852 40282
rect 1104 40208 48852 40230
rect 23290 40128 23296 40180
rect 23348 40168 23354 40180
rect 23385 40171 23443 40177
rect 23385 40168 23397 40171
rect 23348 40140 23397 40168
rect 23348 40128 23354 40140
rect 23385 40137 23397 40140
rect 23431 40137 23443 40171
rect 23385 40131 23443 40137
rect 24394 40128 24400 40180
rect 24452 40168 24458 40180
rect 24857 40171 24915 40177
rect 24857 40168 24869 40171
rect 24452 40140 24869 40168
rect 24452 40128 24458 40140
rect 24857 40137 24869 40140
rect 24903 40168 24915 40171
rect 32122 40168 32128 40180
rect 24903 40140 25544 40168
rect 32083 40140 32128 40168
rect 24903 40137 24915 40140
rect 24857 40131 24915 40137
rect 21407 40103 21465 40109
rect 21407 40069 21419 40103
rect 21453 40100 21465 40103
rect 23566 40100 23572 40112
rect 21453 40072 23572 40100
rect 21453 40069 21465 40072
rect 21407 40063 21465 40069
rect 23566 40060 23572 40072
rect 23624 40060 23630 40112
rect 25516 40041 25544 40140
rect 32122 40128 32128 40140
rect 32180 40128 32186 40180
rect 34514 40128 34520 40180
rect 34572 40168 34578 40180
rect 34790 40168 34796 40180
rect 34572 40140 34796 40168
rect 34572 40128 34578 40140
rect 34790 40128 34796 40140
rect 34848 40168 34854 40180
rect 35069 40171 35127 40177
rect 35069 40168 35081 40171
rect 34848 40140 35081 40168
rect 34848 40128 34854 40140
rect 35069 40137 35081 40140
rect 35115 40137 35127 40171
rect 36262 40168 36268 40180
rect 36223 40140 36268 40168
rect 35069 40131 35127 40137
rect 36262 40128 36268 40140
rect 36320 40128 36326 40180
rect 38010 40128 38016 40180
rect 38068 40168 38074 40180
rect 38105 40171 38163 40177
rect 38105 40168 38117 40171
rect 38068 40140 38117 40168
rect 38068 40128 38074 40140
rect 38105 40137 38117 40140
rect 38151 40137 38163 40171
rect 38105 40131 38163 40137
rect 39114 40128 39120 40180
rect 39172 40168 39178 40180
rect 39669 40171 39727 40177
rect 39669 40168 39681 40171
rect 39172 40140 39681 40168
rect 39172 40128 39178 40140
rect 39669 40137 39681 40140
rect 39715 40168 39727 40171
rect 42426 40168 42432 40180
rect 39715 40140 42432 40168
rect 39715 40137 39727 40140
rect 39669 40131 39727 40137
rect 42426 40128 42432 40140
rect 42484 40128 42490 40180
rect 26786 40060 26792 40112
rect 26844 40100 26850 40112
rect 30653 40103 30711 40109
rect 30653 40100 30665 40103
rect 26844 40072 30665 40100
rect 26844 40060 26850 40072
rect 30653 40069 30665 40072
rect 30699 40069 30711 40103
rect 30653 40063 30711 40069
rect 25501 40035 25559 40041
rect 25501 40001 25513 40035
rect 25547 40001 25559 40035
rect 25774 40032 25780 40044
rect 25735 40004 25780 40032
rect 25501 39995 25559 40001
rect 25774 39992 25780 40004
rect 25832 39992 25838 40044
rect 29270 40032 29276 40044
rect 27540 40004 29276 40032
rect 12504 39967 12562 39973
rect 12504 39933 12516 39967
rect 12550 39964 12562 39967
rect 21336 39967 21394 39973
rect 12550 39936 13032 39964
rect 12550 39933 12562 39936
rect 12504 39927 12562 39933
rect 13004 39840 13032 39936
rect 21336 39933 21348 39967
rect 21382 39964 21394 39967
rect 21382 39936 22232 39964
rect 21382 39933 21394 39936
rect 21336 39927 21394 39933
rect 22204 39905 22232 39936
rect 23014 39924 23020 39976
rect 23072 39964 23078 39976
rect 27540 39973 27568 40004
rect 29270 39992 29276 40004
rect 29328 39992 29334 40044
rect 30006 40032 30012 40044
rect 29967 40004 30012 40032
rect 30006 39992 30012 40004
rect 30064 39992 30070 40044
rect 23728 39967 23786 39973
rect 23728 39964 23740 39967
rect 23072 39936 23740 39964
rect 23072 39924 23078 39936
rect 23728 39933 23740 39936
rect 23774 39964 23786 39967
rect 24121 39967 24179 39973
rect 24121 39964 24133 39967
rect 23774 39936 24133 39964
rect 23774 39933 23786 39936
rect 23728 39927 23786 39933
rect 24121 39933 24133 39936
rect 24167 39933 24179 39967
rect 24121 39927 24179 39933
rect 26789 39967 26847 39973
rect 26789 39933 26801 39967
rect 26835 39964 26847 39967
rect 27525 39967 27583 39973
rect 27525 39964 27537 39967
rect 26835 39936 27537 39964
rect 26835 39933 26847 39936
rect 26789 39927 26847 39933
rect 27525 39933 27537 39936
rect 27571 39933 27583 39967
rect 27525 39927 27583 39933
rect 27801 39967 27859 39973
rect 27801 39933 27813 39967
rect 27847 39964 27859 39967
rect 27982 39964 27988 39976
rect 27847 39936 27988 39964
rect 27847 39933 27859 39936
rect 27801 39927 27859 39933
rect 27982 39924 27988 39936
rect 28040 39964 28046 39976
rect 28261 39967 28319 39973
rect 28261 39964 28273 39967
rect 28040 39936 28273 39964
rect 28040 39924 28046 39936
rect 28261 39933 28273 39936
rect 28307 39933 28319 39967
rect 28261 39927 28319 39933
rect 29457 39967 29515 39973
rect 29457 39933 29469 39967
rect 29503 39933 29515 39967
rect 29457 39927 29515 39933
rect 22189 39899 22247 39905
rect 22189 39865 22201 39899
rect 22235 39896 22247 39899
rect 22554 39896 22560 39908
rect 22235 39868 22560 39896
rect 22235 39865 22247 39868
rect 22189 39859 22247 39865
rect 22554 39856 22560 39868
rect 22612 39856 22618 39908
rect 25593 39899 25651 39905
rect 25593 39865 25605 39899
rect 25639 39896 25651 39899
rect 25682 39896 25688 39908
rect 25639 39868 25688 39896
rect 25639 39865 25651 39868
rect 25593 39859 25651 39865
rect 12575 39831 12633 39837
rect 12575 39797 12587 39831
rect 12621 39828 12633 39831
rect 12802 39828 12808 39840
rect 12621 39800 12808 39828
rect 12621 39797 12633 39800
rect 12575 39791 12633 39797
rect 12802 39788 12808 39800
rect 12860 39788 12866 39840
rect 12986 39828 12992 39840
rect 12947 39800 12992 39828
rect 12986 39788 12992 39800
rect 13044 39788 13050 39840
rect 21174 39788 21180 39840
rect 21232 39828 21238 39840
rect 21729 39831 21787 39837
rect 21729 39828 21741 39831
rect 21232 39800 21741 39828
rect 21232 39788 21238 39800
rect 21729 39797 21741 39800
rect 21775 39797 21787 39831
rect 22278 39828 22284 39840
rect 22239 39800 22284 39828
rect 21729 39791 21787 39797
rect 22278 39788 22284 39800
rect 22336 39788 22342 39840
rect 22833 39831 22891 39837
rect 22833 39797 22845 39831
rect 22879 39828 22891 39831
rect 22922 39828 22928 39840
rect 22879 39800 22928 39828
rect 22879 39797 22891 39800
rect 22833 39791 22891 39797
rect 22922 39788 22928 39800
rect 22980 39788 22986 39840
rect 23658 39788 23664 39840
rect 23716 39828 23722 39840
rect 23799 39831 23857 39837
rect 23799 39828 23811 39831
rect 23716 39800 23811 39828
rect 23716 39788 23722 39800
rect 23799 39797 23811 39800
rect 23845 39797 23857 39831
rect 24486 39828 24492 39840
rect 24447 39800 24492 39828
rect 23799 39791 23857 39797
rect 24486 39788 24492 39800
rect 24544 39788 24550 39840
rect 25317 39831 25375 39837
rect 25317 39797 25329 39831
rect 25363 39828 25375 39831
rect 25608 39828 25636 39859
rect 25682 39856 25688 39868
rect 25740 39856 25746 39908
rect 27157 39899 27215 39905
rect 27157 39865 27169 39899
rect 27203 39896 27215 39899
rect 27614 39896 27620 39908
rect 27203 39868 27620 39896
rect 27203 39865 27215 39868
rect 27157 39859 27215 39865
rect 27614 39856 27620 39868
rect 27672 39896 27678 39908
rect 29089 39899 29147 39905
rect 29089 39896 29101 39899
rect 27672 39868 29101 39896
rect 27672 39856 27678 39868
rect 29089 39865 29101 39868
rect 29135 39896 29147 39899
rect 29472 39896 29500 39927
rect 29546 39924 29552 39976
rect 29604 39964 29610 39976
rect 29733 39967 29791 39973
rect 29733 39964 29745 39967
rect 29604 39936 29745 39964
rect 29604 39924 29610 39936
rect 29733 39933 29745 39936
rect 29779 39933 29791 39967
rect 30668 39964 30696 40063
rect 33318 40032 33324 40044
rect 33279 40004 33324 40032
rect 33318 39992 33324 40004
rect 33376 39992 33382 40044
rect 33502 39992 33508 40044
rect 33560 40032 33566 40044
rect 33597 40035 33655 40041
rect 33597 40032 33609 40035
rect 33560 40004 33609 40032
rect 33560 39992 33566 40004
rect 33597 40001 33609 40004
rect 33643 40001 33655 40035
rect 33597 39995 33655 40001
rect 35802 39992 35808 40044
rect 35860 40032 35866 40044
rect 38657 40035 38715 40041
rect 35860 40004 38516 40032
rect 35860 39992 35866 40004
rect 30834 39964 30840 39976
rect 30668 39936 30840 39964
rect 29733 39927 29791 39933
rect 30834 39924 30840 39936
rect 30892 39924 30898 39976
rect 31294 39964 31300 39976
rect 31255 39936 31300 39964
rect 31294 39924 31300 39936
rect 31352 39924 31358 39976
rect 35250 39964 35256 39976
rect 35211 39936 35256 39964
rect 35250 39924 35256 39936
rect 35308 39924 35314 39976
rect 35710 39964 35716 39976
rect 35671 39936 35716 39964
rect 35710 39924 35716 39936
rect 35768 39924 35774 39976
rect 35989 39967 36047 39973
rect 35989 39933 36001 39967
rect 36035 39964 36047 39967
rect 36817 39967 36875 39973
rect 36817 39964 36829 39967
rect 36035 39936 36829 39964
rect 36035 39933 36047 39936
rect 35989 39927 36047 39933
rect 36817 39933 36829 39936
rect 36863 39964 36875 39967
rect 36906 39964 36912 39976
rect 36863 39936 36912 39964
rect 36863 39933 36875 39936
rect 36817 39927 36875 39933
rect 36906 39924 36912 39936
rect 36964 39924 36970 39976
rect 30374 39896 30380 39908
rect 29135 39868 30380 39896
rect 29135 39865 29147 39868
rect 29089 39859 29147 39865
rect 30374 39856 30380 39868
rect 30432 39856 30438 39908
rect 31570 39896 31576 39908
rect 31531 39868 31576 39896
rect 31570 39856 31576 39868
rect 31628 39856 31634 39908
rect 32769 39899 32827 39905
rect 32769 39865 32781 39899
rect 32815 39896 32827 39899
rect 33042 39896 33048 39908
rect 32815 39868 33048 39896
rect 32815 39865 32827 39868
rect 32769 39859 32827 39865
rect 33042 39856 33048 39868
rect 33100 39896 33106 39908
rect 33137 39899 33195 39905
rect 33137 39896 33149 39899
rect 33100 39868 33149 39896
rect 33100 39856 33106 39868
rect 33137 39865 33149 39868
rect 33183 39896 33195 39899
rect 33413 39899 33471 39905
rect 33413 39896 33425 39899
rect 33183 39868 33425 39896
rect 33183 39865 33195 39868
rect 33137 39859 33195 39865
rect 33413 39865 33425 39868
rect 33459 39896 33471 39899
rect 33594 39896 33600 39908
rect 33459 39868 33600 39896
rect 33459 39865 33471 39868
rect 33413 39859 33471 39865
rect 33594 39856 33600 39868
rect 33652 39856 33658 39908
rect 37138 39899 37196 39905
rect 37138 39865 37150 39899
rect 37184 39865 37196 39899
rect 37138 39859 37196 39865
rect 27338 39828 27344 39840
rect 25363 39800 25636 39828
rect 27299 39800 27344 39828
rect 25363 39797 25375 39800
rect 25317 39791 25375 39797
rect 27338 39788 27344 39800
rect 27396 39788 27402 39840
rect 28718 39828 28724 39840
rect 28679 39800 28724 39828
rect 28718 39788 28724 39800
rect 28776 39788 28782 39840
rect 29454 39788 29460 39840
rect 29512 39828 29518 39840
rect 30285 39831 30343 39837
rect 30285 39828 30297 39831
rect 29512 39800 30297 39828
rect 29512 39788 29518 39800
rect 30285 39797 30297 39800
rect 30331 39797 30343 39831
rect 30285 39791 30343 39797
rect 36538 39788 36544 39840
rect 36596 39828 36602 39840
rect 36725 39831 36783 39837
rect 36725 39828 36737 39831
rect 36596 39800 36737 39828
rect 36596 39788 36602 39800
rect 36725 39797 36737 39800
rect 36771 39828 36783 39831
rect 36998 39828 37004 39840
rect 36771 39800 37004 39828
rect 36771 39797 36783 39800
rect 36725 39791 36783 39797
rect 36998 39788 37004 39800
rect 37056 39828 37062 39840
rect 37153 39828 37181 39859
rect 37734 39828 37740 39840
rect 37056 39800 37181 39828
rect 37695 39800 37740 39828
rect 37056 39788 37062 39800
rect 37734 39788 37740 39800
rect 37792 39788 37798 39840
rect 38488 39828 38516 40004
rect 38657 40001 38669 40035
rect 38703 40032 38715 40035
rect 39132 40032 39160 40128
rect 39758 40060 39764 40112
rect 39816 40100 39822 40112
rect 39945 40103 40003 40109
rect 39945 40100 39957 40103
rect 39816 40072 39957 40100
rect 39816 40060 39822 40072
rect 39945 40069 39957 40072
rect 39991 40100 40003 40103
rect 41322 40100 41328 40112
rect 39991 40072 41328 40100
rect 39991 40069 40003 40072
rect 39945 40063 40003 40069
rect 41322 40060 41328 40072
rect 41380 40060 41386 40112
rect 41984 40072 43576 40100
rect 38703 40004 39160 40032
rect 38703 40001 38715 40004
rect 38657 39995 38715 40001
rect 40862 39992 40868 40044
rect 40920 40032 40926 40044
rect 41984 40041 42012 40072
rect 41969 40035 42027 40041
rect 41969 40032 41981 40035
rect 40920 40004 41981 40032
rect 40920 39992 40926 40004
rect 41969 40001 41981 40004
rect 42015 40001 42027 40035
rect 43254 40032 43260 40044
rect 43215 40004 43260 40032
rect 41969 39995 42027 40001
rect 43254 39992 43260 40004
rect 43312 39992 43318 40044
rect 43548 40041 43576 40072
rect 43533 40035 43591 40041
rect 43533 40001 43545 40035
rect 43579 40001 43591 40035
rect 43533 39995 43591 40001
rect 40624 39967 40682 39973
rect 40624 39964 40636 39967
rect 40420 39936 40636 39964
rect 38746 39856 38752 39908
rect 38804 39896 38810 39908
rect 39298 39896 39304 39908
rect 38804 39868 38849 39896
rect 39259 39868 39304 39896
rect 38804 39856 38810 39868
rect 39298 39856 39304 39868
rect 39356 39856 39362 39908
rect 40420 39828 40448 39936
rect 40624 39933 40636 39936
rect 40670 39964 40682 39967
rect 41049 39967 41107 39973
rect 41049 39964 41061 39967
rect 40670 39936 41061 39964
rect 40670 39933 40682 39936
rect 40624 39927 40682 39933
rect 41049 39933 41061 39936
rect 41095 39964 41107 39967
rect 41138 39964 41144 39976
rect 41095 39936 41144 39964
rect 41095 39933 41107 39936
rect 41049 39927 41107 39933
rect 41138 39924 41144 39936
rect 41196 39924 41202 39976
rect 41690 39896 41696 39908
rect 41651 39868 41696 39896
rect 41690 39856 41696 39868
rect 41748 39856 41754 39908
rect 41782 39856 41788 39908
rect 41840 39896 41846 39908
rect 43070 39896 43076 39908
rect 41840 39868 41933 39896
rect 42983 39868 43076 39896
rect 41840 39856 41846 39868
rect 43070 39856 43076 39868
rect 43128 39896 43134 39908
rect 43349 39899 43407 39905
rect 43349 39896 43361 39899
rect 43128 39868 43361 39896
rect 43128 39856 43134 39868
rect 43349 39865 43361 39868
rect 43395 39865 43407 39899
rect 43349 39859 43407 39865
rect 38488 39800 40448 39828
rect 40727 39831 40785 39837
rect 40727 39797 40739 39831
rect 40773 39828 40785 39831
rect 40954 39828 40960 39840
rect 40773 39800 40960 39828
rect 40773 39797 40785 39800
rect 40727 39791 40785 39797
rect 40954 39788 40960 39800
rect 41012 39788 41018 39840
rect 41509 39831 41567 39837
rect 41509 39797 41521 39831
rect 41555 39828 41567 39831
rect 41800 39828 41828 39856
rect 42613 39831 42671 39837
rect 42613 39828 42625 39831
rect 41555 39800 42625 39828
rect 41555 39797 41567 39800
rect 41509 39791 41567 39797
rect 42613 39797 42625 39800
rect 42659 39797 42671 39831
rect 42613 39791 42671 39797
rect 1104 39738 48852 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 48852 39738
rect 1104 39664 48852 39686
rect 22186 39624 22192 39636
rect 22147 39596 22192 39624
rect 22186 39584 22192 39596
rect 22244 39584 22250 39636
rect 22462 39584 22468 39636
rect 22520 39624 22526 39636
rect 23017 39627 23075 39633
rect 23017 39624 23029 39627
rect 22520 39596 23029 39624
rect 22520 39584 22526 39596
rect 23017 39593 23029 39596
rect 23063 39593 23075 39627
rect 23017 39587 23075 39593
rect 27617 39627 27675 39633
rect 27617 39593 27629 39627
rect 27663 39624 27675 39627
rect 27982 39624 27988 39636
rect 27663 39596 27988 39624
rect 27663 39593 27675 39596
rect 27617 39587 27675 39593
rect 27982 39584 27988 39596
rect 28040 39584 28046 39636
rect 28166 39624 28172 39636
rect 28127 39596 28172 39624
rect 28166 39584 28172 39596
rect 28224 39584 28230 39636
rect 30006 39624 30012 39636
rect 29967 39596 30012 39624
rect 30006 39584 30012 39596
rect 30064 39584 30070 39636
rect 32398 39584 32404 39636
rect 32456 39624 32462 39636
rect 32493 39627 32551 39633
rect 32493 39624 32505 39627
rect 32456 39596 32505 39624
rect 32456 39584 32462 39596
rect 32493 39593 32505 39596
rect 32539 39593 32551 39627
rect 33042 39624 33048 39636
rect 33003 39596 33048 39624
rect 32493 39587 32551 39593
rect 33042 39584 33048 39596
rect 33100 39584 33106 39636
rect 33318 39584 33324 39636
rect 33376 39624 33382 39636
rect 33689 39627 33747 39633
rect 33689 39624 33701 39627
rect 33376 39596 33701 39624
rect 33376 39584 33382 39596
rect 33689 39593 33701 39596
rect 33735 39593 33747 39627
rect 36906 39624 36912 39636
rect 36867 39596 36912 39624
rect 33689 39587 33747 39593
rect 36906 39584 36912 39596
rect 36964 39584 36970 39636
rect 41598 39624 41604 39636
rect 41559 39596 41604 39624
rect 41598 39584 41604 39596
rect 41656 39624 41662 39636
rect 43487 39627 43545 39633
rect 43487 39624 43499 39627
rect 41656 39596 43499 39624
rect 41656 39584 41662 39596
rect 43487 39593 43499 39596
rect 43533 39593 43545 39627
rect 43487 39587 43545 39593
rect 22922 39516 22928 39568
rect 22980 39556 22986 39568
rect 23753 39559 23811 39565
rect 23753 39556 23765 39559
rect 22980 39528 23765 39556
rect 22980 39516 22986 39528
rect 23753 39525 23765 39528
rect 23799 39556 23811 39559
rect 24486 39556 24492 39568
rect 23799 39528 24492 39556
rect 23799 39525 23811 39528
rect 23753 39519 23811 39525
rect 24486 39516 24492 39528
rect 24544 39516 24550 39568
rect 26694 39556 26700 39568
rect 26655 39528 26700 39556
rect 26694 39516 26700 39528
rect 26752 39516 26758 39568
rect 28000 39556 28028 39584
rect 30650 39556 30656 39568
rect 28000 39528 28580 39556
rect 30611 39528 30656 39556
rect 11974 39488 11980 39500
rect 11935 39460 11980 39488
rect 11974 39448 11980 39460
rect 12032 39448 12038 39500
rect 14001 39491 14059 39497
rect 14001 39457 14013 39491
rect 14047 39488 14059 39491
rect 14826 39488 14832 39500
rect 14047 39460 14832 39488
rect 14047 39457 14059 39460
rect 14001 39451 14059 39457
rect 14826 39448 14832 39460
rect 14884 39448 14890 39500
rect 15356 39491 15414 39497
rect 15356 39457 15368 39491
rect 15402 39488 15414 39491
rect 16114 39488 16120 39500
rect 15402 39460 16120 39488
rect 15402 39457 15414 39460
rect 15356 39451 15414 39457
rect 16114 39448 16120 39460
rect 16172 39448 16178 39500
rect 25130 39488 25136 39500
rect 25091 39460 25136 39488
rect 25130 39448 25136 39460
rect 25188 39448 25194 39500
rect 28350 39488 28356 39500
rect 28311 39460 28356 39488
rect 28350 39448 28356 39460
rect 28408 39448 28414 39500
rect 28552 39497 28580 39528
rect 30650 39516 30656 39528
rect 30708 39516 30714 39568
rect 33410 39556 33416 39568
rect 33371 39528 33416 39556
rect 33410 39516 33416 39528
rect 33468 39516 33474 39568
rect 33962 39556 33968 39568
rect 33923 39528 33968 39556
rect 33962 39516 33968 39528
rect 34020 39516 34026 39568
rect 34057 39559 34115 39565
rect 34057 39525 34069 39559
rect 34103 39556 34115 39559
rect 34606 39556 34612 39568
rect 34103 39528 34612 39556
rect 34103 39525 34115 39528
rect 34057 39519 34115 39525
rect 34606 39516 34612 39528
rect 34664 39516 34670 39568
rect 37734 39516 37740 39568
rect 37792 39556 37798 39568
rect 38562 39556 38568 39568
rect 37792 39528 38568 39556
rect 37792 39516 37798 39528
rect 38562 39516 38568 39528
rect 38620 39556 38626 39568
rect 38657 39559 38715 39565
rect 38657 39556 38669 39559
rect 38620 39528 38669 39556
rect 38620 39516 38626 39528
rect 38657 39525 38669 39528
rect 38703 39525 38715 39559
rect 38657 39519 38715 39525
rect 40126 39516 40132 39568
rect 40184 39556 40190 39568
rect 40221 39559 40279 39565
rect 40221 39556 40233 39559
rect 40184 39528 40233 39556
rect 40184 39516 40190 39528
rect 40221 39525 40233 39528
rect 40267 39525 40279 39559
rect 40221 39519 40279 39525
rect 40954 39516 40960 39568
rect 41012 39556 41018 39568
rect 41506 39556 41512 39568
rect 41012 39528 41512 39556
rect 41012 39516 41018 39528
rect 41506 39516 41512 39528
rect 41564 39556 41570 39568
rect 41785 39559 41843 39565
rect 41785 39556 41797 39559
rect 41564 39528 41797 39556
rect 41564 39516 41570 39528
rect 41785 39525 41797 39528
rect 41831 39525 41843 39559
rect 41785 39519 41843 39525
rect 41877 39559 41935 39565
rect 41877 39525 41889 39559
rect 41923 39556 41935 39559
rect 43070 39556 43076 39568
rect 41923 39528 43076 39556
rect 41923 39525 41935 39528
rect 41877 39519 41935 39525
rect 43070 39516 43076 39528
rect 43128 39516 43134 39568
rect 28537 39491 28595 39497
rect 28537 39457 28549 39491
rect 28583 39457 28595 39491
rect 28537 39451 28595 39457
rect 31570 39448 31576 39500
rect 31628 39488 31634 39500
rect 32125 39491 32183 39497
rect 32125 39488 32137 39491
rect 31628 39460 32137 39488
rect 31628 39448 31634 39460
rect 32125 39457 32137 39460
rect 32171 39488 32183 39491
rect 32674 39488 32680 39500
rect 32171 39460 32680 39488
rect 32171 39457 32183 39460
rect 32125 39451 32183 39457
rect 32674 39448 32680 39460
rect 32732 39448 32738 39500
rect 36170 39488 36176 39500
rect 36131 39460 36176 39488
rect 36170 39448 36176 39460
rect 36228 39448 36234 39500
rect 36357 39491 36415 39497
rect 36357 39457 36369 39491
rect 36403 39457 36415 39491
rect 36357 39451 36415 39457
rect 10962 39380 10968 39432
rect 11020 39420 11026 39432
rect 12345 39423 12403 39429
rect 12345 39420 12357 39423
rect 11020 39392 12357 39420
rect 11020 39380 11026 39392
rect 12345 39389 12357 39392
rect 12391 39420 12403 39423
rect 12986 39420 12992 39432
rect 12391 39392 12992 39420
rect 12391 39389 12403 39392
rect 12345 39383 12403 39389
rect 12986 39380 12992 39392
rect 13044 39380 13050 39432
rect 21450 39380 21456 39432
rect 21508 39420 21514 39432
rect 21821 39423 21879 39429
rect 21821 39420 21833 39423
rect 21508 39392 21833 39420
rect 21508 39380 21514 39392
rect 21821 39389 21833 39392
rect 21867 39389 21879 39423
rect 23658 39420 23664 39432
rect 23619 39392 23664 39420
rect 21821 39383 21879 39389
rect 23658 39380 23664 39392
rect 23716 39380 23722 39432
rect 25314 39380 25320 39432
rect 25372 39420 25378 39432
rect 25593 39423 25651 39429
rect 25593 39420 25605 39423
rect 25372 39392 25605 39420
rect 25372 39380 25378 39392
rect 25593 39389 25605 39392
rect 25639 39389 25651 39423
rect 25593 39383 25651 39389
rect 26605 39423 26663 39429
rect 26605 39389 26617 39423
rect 26651 39389 26663 39423
rect 26878 39420 26884 39432
rect 26791 39392 26884 39420
rect 26605 39383 26663 39389
rect 17310 39312 17316 39364
rect 17368 39352 17374 39364
rect 24026 39352 24032 39364
rect 17368 39324 24032 39352
rect 17368 39312 17374 39324
rect 24026 39312 24032 39324
rect 24084 39312 24090 39364
rect 24210 39352 24216 39364
rect 24171 39324 24216 39352
rect 24210 39312 24216 39324
rect 24268 39352 24274 39364
rect 26234 39352 26240 39364
rect 24268 39324 26240 39352
rect 24268 39312 24274 39324
rect 26234 39312 26240 39324
rect 26292 39352 26298 39364
rect 26620 39352 26648 39383
rect 26878 39380 26884 39392
rect 26936 39380 26942 39432
rect 30561 39423 30619 39429
rect 30561 39389 30573 39423
rect 30607 39420 30619 39423
rect 30607 39392 31616 39420
rect 30607 39389 30619 39392
rect 30561 39383 30619 39389
rect 26292 39324 26648 39352
rect 26292 39312 26298 39324
rect 13630 39244 13636 39296
rect 13688 39284 13694 39296
rect 14185 39287 14243 39293
rect 14185 39284 14197 39287
rect 13688 39256 14197 39284
rect 13688 39244 13694 39256
rect 14185 39253 14197 39256
rect 14231 39253 14243 39287
rect 14185 39247 14243 39253
rect 15010 39244 15016 39296
rect 15068 39284 15074 39296
rect 15427 39287 15485 39293
rect 15427 39284 15439 39287
rect 15068 39256 15439 39284
rect 15068 39244 15074 39256
rect 15427 39253 15439 39256
rect 15473 39253 15485 39287
rect 15427 39247 15485 39253
rect 22741 39287 22799 39293
rect 22741 39253 22753 39287
rect 22787 39284 22799 39287
rect 22922 39284 22928 39296
rect 22787 39256 22928 39284
rect 22787 39253 22799 39256
rect 22741 39247 22799 39253
rect 22922 39244 22928 39256
rect 22980 39244 22986 39296
rect 24394 39244 24400 39296
rect 24452 39284 24458 39296
rect 25271 39287 25329 39293
rect 25271 39284 25283 39287
rect 24452 39256 25283 39284
rect 24452 39244 24458 39256
rect 25271 39253 25283 39256
rect 25317 39253 25329 39287
rect 25271 39247 25329 39253
rect 25774 39244 25780 39296
rect 25832 39284 25838 39296
rect 26896 39284 26924 39380
rect 31110 39352 31116 39364
rect 31071 39324 31116 39352
rect 31110 39312 31116 39324
rect 31168 39312 31174 39364
rect 31588 39361 31616 39392
rect 33134 39380 33140 39432
rect 33192 39420 33198 39432
rect 35250 39420 35256 39432
rect 33192 39392 35256 39420
rect 33192 39380 33198 39392
rect 35250 39380 35256 39392
rect 35308 39380 35314 39432
rect 36372 39420 36400 39451
rect 42426 39448 42432 39500
rect 42484 39488 42490 39500
rect 42484 39460 42529 39488
rect 42484 39448 42490 39460
rect 43162 39448 43168 39500
rect 43220 39488 43226 39500
rect 43384 39491 43442 39497
rect 43384 39488 43396 39491
rect 43220 39460 43396 39488
rect 43220 39448 43226 39460
rect 43384 39457 43396 39460
rect 43430 39457 43442 39491
rect 43384 39451 43442 39457
rect 36630 39420 36636 39432
rect 35728 39392 36400 39420
rect 36591 39392 36636 39420
rect 31573 39355 31631 39361
rect 31573 39321 31585 39355
rect 31619 39352 31631 39355
rect 33502 39352 33508 39364
rect 31619 39324 33508 39352
rect 31619 39321 31631 39324
rect 31573 39315 31631 39321
rect 33502 39312 33508 39324
rect 33560 39352 33566 39364
rect 34517 39355 34575 39361
rect 34517 39352 34529 39355
rect 33560 39324 34529 39352
rect 33560 39312 33566 39324
rect 34517 39321 34529 39324
rect 34563 39321 34575 39355
rect 34517 39315 34575 39321
rect 35728 39296 35756 39392
rect 36630 39380 36636 39392
rect 36688 39380 36694 39432
rect 38565 39423 38623 39429
rect 38565 39389 38577 39423
rect 38611 39420 38623 39423
rect 38654 39420 38660 39432
rect 38611 39392 38660 39420
rect 38611 39389 38623 39392
rect 38565 39383 38623 39389
rect 38654 39380 38660 39392
rect 38712 39380 38718 39432
rect 40129 39423 40187 39429
rect 40129 39389 40141 39423
rect 40175 39420 40187 39423
rect 40218 39420 40224 39432
rect 40175 39392 40224 39420
rect 40175 39389 40187 39392
rect 40129 39383 40187 39389
rect 40218 39380 40224 39392
rect 40276 39380 40282 39432
rect 40405 39423 40463 39429
rect 40405 39389 40417 39423
rect 40451 39389 40463 39423
rect 40405 39383 40463 39389
rect 39117 39355 39175 39361
rect 39117 39321 39129 39355
rect 39163 39352 39175 39355
rect 39298 39352 39304 39364
rect 39163 39324 39304 39352
rect 39163 39321 39175 39324
rect 39117 39315 39175 39321
rect 39298 39312 39304 39324
rect 39356 39352 39362 39364
rect 40420 39352 40448 39383
rect 39356 39324 40448 39352
rect 39356 39312 39362 39324
rect 25832 39256 26924 39284
rect 25832 39244 25838 39256
rect 29454 39244 29460 39296
rect 29512 39284 29518 39296
rect 29549 39287 29607 39293
rect 29549 39284 29561 39287
rect 29512 39256 29561 39284
rect 29512 39244 29518 39256
rect 29549 39253 29561 39256
rect 29595 39253 29607 39287
rect 35710 39284 35716 39296
rect 35671 39256 35716 39284
rect 29549 39247 29607 39253
rect 35710 39244 35716 39256
rect 35768 39244 35774 39296
rect 1104 39194 48852 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 48852 39194
rect 1104 39120 48852 39142
rect 22186 39080 22192 39092
rect 22147 39052 22192 39080
rect 22186 39040 22192 39052
rect 22244 39040 22250 39092
rect 23474 39040 23480 39092
rect 23532 39080 23538 39092
rect 23532 39052 23577 39080
rect 23532 39040 23538 39052
rect 23658 39040 23664 39092
rect 23716 39080 23722 39092
rect 24673 39083 24731 39089
rect 24673 39080 24685 39083
rect 23716 39052 24685 39080
rect 23716 39040 23722 39052
rect 24673 39049 24685 39052
rect 24719 39049 24731 39083
rect 24673 39043 24731 39049
rect 30469 39083 30527 39089
rect 30469 39049 30481 39083
rect 30515 39080 30527 39083
rect 30650 39080 30656 39092
rect 30515 39052 30656 39080
rect 30515 39049 30527 39052
rect 30469 39043 30527 39049
rect 30650 39040 30656 39052
rect 30708 39080 30714 39092
rect 30745 39083 30803 39089
rect 30745 39080 30757 39083
rect 30708 39052 30757 39080
rect 30708 39040 30714 39052
rect 30745 39049 30757 39052
rect 30791 39049 30803 39083
rect 32674 39080 32680 39092
rect 32635 39052 32680 39080
rect 30745 39043 30803 39049
rect 32674 39040 32680 39052
rect 32732 39040 32738 39092
rect 38562 39080 38568 39092
rect 38523 39052 38568 39080
rect 38562 39040 38568 39052
rect 38620 39040 38626 39092
rect 39761 39083 39819 39089
rect 39761 39049 39773 39083
rect 39807 39080 39819 39083
rect 40218 39080 40224 39092
rect 39807 39052 40224 39080
rect 39807 39049 39819 39052
rect 39761 39043 39819 39049
rect 40218 39040 40224 39052
rect 40276 39040 40282 39092
rect 40819 39083 40877 39089
rect 40819 39049 40831 39083
rect 40865 39080 40877 39083
rect 41690 39080 41696 39092
rect 40865 39052 41696 39080
rect 40865 39049 40877 39052
rect 40819 39043 40877 39049
rect 41690 39040 41696 39052
rect 41748 39040 41754 39092
rect 42702 39040 42708 39092
rect 42760 39080 42766 39092
rect 43162 39080 43168 39092
rect 42760 39052 43168 39080
rect 42760 39040 42766 39052
rect 43162 39040 43168 39052
rect 43220 39040 43226 39092
rect 26605 39015 26663 39021
rect 26605 38981 26617 39015
rect 26651 39012 26663 39015
rect 26694 39012 26700 39024
rect 26651 38984 26700 39012
rect 26651 38981 26663 38984
rect 26605 38975 26663 38981
rect 26694 38972 26700 38984
rect 26752 39012 26758 39024
rect 28353 39015 28411 39021
rect 28353 39012 28365 39015
rect 26752 38984 28365 39012
rect 26752 38972 26758 38984
rect 28353 38981 28365 38984
rect 28399 38981 28411 39015
rect 28353 38975 28411 38981
rect 31110 38972 31116 39024
rect 31168 39012 31174 39024
rect 31941 39015 31999 39021
rect 31941 39012 31953 39015
rect 31168 38984 31953 39012
rect 31168 38972 31174 38984
rect 31941 38981 31953 38984
rect 31987 39012 31999 39015
rect 32214 39012 32220 39024
rect 31987 38984 32220 39012
rect 31987 38981 31999 38984
rect 31941 38975 31999 38981
rect 32214 38972 32220 38984
rect 32272 38972 32278 39024
rect 37645 39015 37703 39021
rect 37645 38981 37657 39015
rect 37691 39012 37703 39015
rect 38746 39012 38752 39024
rect 37691 38984 38752 39012
rect 37691 38981 37703 38984
rect 37645 38975 37703 38981
rect 38746 38972 38752 38984
rect 38804 38972 38810 39024
rect 39298 39012 39304 39024
rect 39259 38984 39304 39012
rect 39298 38972 39304 38984
rect 39356 38972 39362 39024
rect 8294 38904 8300 38956
rect 8352 38944 8358 38956
rect 11146 38944 11152 38956
rect 8352 38916 11152 38944
rect 8352 38904 8358 38916
rect 11146 38904 11152 38916
rect 11204 38904 11210 38956
rect 21174 38944 21180 38956
rect 21135 38916 21180 38944
rect 21174 38904 21180 38916
rect 21232 38904 21238 38956
rect 24210 38944 24216 38956
rect 24171 38916 24216 38944
rect 24210 38904 24216 38916
rect 24268 38904 24274 38956
rect 25774 38944 25780 38956
rect 25735 38916 25780 38944
rect 25774 38904 25780 38916
rect 25832 38904 25838 38956
rect 26973 38947 27031 38953
rect 26973 38913 26985 38947
rect 27019 38944 27031 38947
rect 27433 38947 27491 38953
rect 27433 38944 27445 38947
rect 27019 38916 27445 38944
rect 27019 38913 27031 38916
rect 26973 38907 27031 38913
rect 27433 38913 27445 38916
rect 27479 38944 27491 38947
rect 28166 38944 28172 38956
rect 27479 38916 28172 38944
rect 27479 38913 27491 38916
rect 27433 38907 27491 38913
rect 28166 38904 28172 38916
rect 28224 38904 28230 38956
rect 31389 38947 31447 38953
rect 31389 38913 31401 38947
rect 31435 38944 31447 38947
rect 34333 38947 34391 38953
rect 31435 38916 34008 38944
rect 31435 38913 31447 38916
rect 31389 38907 31447 38913
rect 11885 38879 11943 38885
rect 11885 38845 11897 38879
rect 11931 38876 11943 38879
rect 11974 38876 11980 38888
rect 11931 38848 11980 38876
rect 11931 38845 11943 38848
rect 11885 38839 11943 38845
rect 11974 38836 11980 38848
rect 12032 38836 12038 38888
rect 12504 38879 12562 38885
rect 12504 38845 12516 38879
rect 12550 38876 12562 38879
rect 12802 38876 12808 38888
rect 12550 38848 12808 38876
rect 12550 38845 12562 38848
rect 12504 38839 12562 38845
rect 12802 38836 12808 38848
rect 12860 38876 12866 38888
rect 12897 38879 12955 38885
rect 12897 38876 12909 38879
rect 12860 38848 12909 38876
rect 12860 38836 12866 38848
rect 12897 38845 12909 38848
rect 12943 38845 12955 38879
rect 12897 38839 12955 38845
rect 13633 38879 13691 38885
rect 13633 38845 13645 38879
rect 13679 38876 13691 38879
rect 14369 38879 14427 38885
rect 14369 38876 14381 38879
rect 13679 38848 14381 38876
rect 13679 38845 13691 38848
rect 13633 38839 13691 38845
rect 14369 38845 14381 38848
rect 14415 38845 14427 38879
rect 14826 38876 14832 38888
rect 14739 38848 14832 38876
rect 14369 38839 14427 38845
rect 10870 38808 10876 38820
rect 10831 38780 10876 38808
rect 10870 38768 10876 38780
rect 10928 38768 10934 38820
rect 10962 38768 10968 38820
rect 11020 38808 11026 38820
rect 13722 38808 13728 38820
rect 11020 38780 11065 38808
rect 13683 38780 13728 38808
rect 11020 38768 11026 38780
rect 13722 38768 13728 38780
rect 13780 38768 13786 38820
rect 14384 38808 14412 38839
rect 14826 38836 14832 38848
rect 14884 38876 14890 38888
rect 15340 38879 15398 38885
rect 15340 38876 15352 38879
rect 14884 38848 15352 38876
rect 14884 38836 14890 38848
rect 15340 38845 15352 38848
rect 15386 38876 15398 38879
rect 16368 38879 16426 38885
rect 15386 38848 15884 38876
rect 15386 38845 15398 38848
rect 15340 38839 15398 38845
rect 15427 38811 15485 38817
rect 15427 38808 15439 38811
rect 14384 38780 15439 38808
rect 15427 38777 15439 38780
rect 15473 38777 15485 38811
rect 15427 38771 15485 38777
rect 10689 38743 10747 38749
rect 10689 38709 10701 38743
rect 10735 38740 10747 38743
rect 10980 38740 11008 38768
rect 15856 38752 15884 38848
rect 16368 38845 16380 38879
rect 16414 38876 16426 38879
rect 20692 38879 20750 38885
rect 16414 38848 16896 38876
rect 16414 38845 16426 38848
rect 16368 38839 16426 38845
rect 16868 38752 16896 38848
rect 20692 38845 20704 38879
rect 20738 38876 20750 38879
rect 21192 38876 21220 38904
rect 20738 38848 21220 38876
rect 21704 38879 21762 38885
rect 20738 38845 20750 38848
rect 20692 38839 20750 38845
rect 21704 38845 21716 38879
rect 21750 38876 21762 38879
rect 22094 38876 22100 38888
rect 21750 38848 22100 38876
rect 21750 38845 21762 38848
rect 21704 38839 21762 38845
rect 22094 38836 22100 38848
rect 22152 38876 22158 38888
rect 29089 38879 29147 38885
rect 22152 38848 22508 38876
rect 22152 38836 22158 38848
rect 22480 38752 22508 38848
rect 29089 38845 29101 38879
rect 29135 38876 29147 38879
rect 29270 38876 29276 38888
rect 29135 38848 29276 38876
rect 29135 38845 29147 38848
rect 29089 38839 29147 38845
rect 29270 38836 29276 38848
rect 29328 38876 29334 38888
rect 29549 38879 29607 38885
rect 29549 38876 29561 38879
rect 29328 38848 29561 38876
rect 29328 38836 29334 38848
rect 29549 38845 29561 38848
rect 29595 38845 29607 38879
rect 29549 38839 29607 38845
rect 23382 38768 23388 38820
rect 23440 38808 23446 38820
rect 23566 38808 23572 38820
rect 23440 38780 23572 38808
rect 23440 38768 23446 38780
rect 23566 38768 23572 38780
rect 23624 38808 23630 38820
rect 23753 38811 23811 38817
rect 23753 38808 23765 38811
rect 23624 38780 23765 38808
rect 23624 38768 23630 38780
rect 23753 38777 23765 38780
rect 23799 38777 23811 38811
rect 23753 38771 23811 38777
rect 23845 38811 23903 38817
rect 23845 38777 23857 38811
rect 23891 38777 23903 38811
rect 23845 38771 23903 38777
rect 10735 38712 11008 38740
rect 10735 38709 10747 38712
rect 10689 38703 10747 38709
rect 11882 38700 11888 38752
rect 11940 38740 11946 38752
rect 12575 38743 12633 38749
rect 12575 38740 12587 38743
rect 11940 38712 12587 38740
rect 11940 38700 11946 38712
rect 12575 38709 12587 38712
rect 12621 38709 12633 38743
rect 15838 38740 15844 38752
rect 15799 38712 15844 38740
rect 12575 38703 12633 38709
rect 15838 38700 15844 38712
rect 15896 38700 15902 38752
rect 16114 38740 16120 38752
rect 16075 38712 16120 38740
rect 16114 38700 16120 38712
rect 16172 38700 16178 38752
rect 16298 38700 16304 38752
rect 16356 38740 16362 38752
rect 16439 38743 16497 38749
rect 16439 38740 16451 38743
rect 16356 38712 16451 38740
rect 16356 38700 16362 38712
rect 16439 38709 16451 38712
rect 16485 38709 16497 38743
rect 16850 38740 16856 38752
rect 16811 38712 16856 38740
rect 16439 38703 16497 38709
rect 16850 38700 16856 38712
rect 16908 38700 16914 38752
rect 20763 38743 20821 38749
rect 20763 38709 20775 38743
rect 20809 38740 20821 38743
rect 20990 38740 20996 38752
rect 20809 38712 20996 38740
rect 20809 38709 20821 38712
rect 20763 38703 20821 38709
rect 20990 38700 20996 38712
rect 21048 38700 21054 38752
rect 21450 38740 21456 38752
rect 21411 38712 21456 38740
rect 21450 38700 21456 38712
rect 21508 38700 21514 38752
rect 21542 38700 21548 38752
rect 21600 38740 21606 38752
rect 21775 38743 21833 38749
rect 21775 38740 21787 38743
rect 21600 38712 21787 38740
rect 21600 38700 21606 38712
rect 21775 38709 21787 38712
rect 21821 38709 21833 38743
rect 22462 38740 22468 38752
rect 22423 38712 22468 38740
rect 21775 38703 21833 38709
rect 22462 38700 22468 38712
rect 22520 38700 22526 38752
rect 22922 38700 22928 38752
rect 22980 38740 22986 38752
rect 23017 38743 23075 38749
rect 23017 38740 23029 38743
rect 22980 38712 23029 38740
rect 22980 38700 22986 38712
rect 23017 38709 23029 38712
rect 23063 38709 23075 38743
rect 23017 38703 23075 38709
rect 23474 38700 23480 38752
rect 23532 38740 23538 38752
rect 23860 38740 23888 38771
rect 25314 38768 25320 38820
rect 25372 38808 25378 38820
rect 25501 38811 25559 38817
rect 25501 38808 25513 38811
rect 25372 38780 25513 38808
rect 25372 38768 25378 38780
rect 25501 38777 25513 38780
rect 25547 38777 25559 38811
rect 25501 38771 25559 38777
rect 25590 38768 25596 38820
rect 25648 38808 25654 38820
rect 27754 38811 27812 38817
rect 25648 38780 25693 38808
rect 25648 38768 25654 38780
rect 27754 38777 27766 38811
rect 27800 38808 27812 38811
rect 29454 38808 29460 38820
rect 27800 38780 29460 38808
rect 27800 38777 27812 38780
rect 27754 38771 27812 38777
rect 23532 38712 23888 38740
rect 23532 38700 23538 38712
rect 24026 38700 24032 38752
rect 24084 38740 24090 38752
rect 25130 38740 25136 38752
rect 24084 38712 25136 38740
rect 24084 38700 24090 38712
rect 25130 38700 25136 38712
rect 25188 38740 25194 38752
rect 25225 38743 25283 38749
rect 25225 38740 25237 38743
rect 25188 38712 25237 38740
rect 25188 38700 25194 38712
rect 25225 38709 25237 38712
rect 25271 38740 25283 38743
rect 25682 38740 25688 38752
rect 25271 38712 25688 38740
rect 25271 38709 25283 38712
rect 25225 38703 25283 38709
rect 25682 38700 25688 38712
rect 25740 38700 25746 38752
rect 27246 38740 27252 38752
rect 27207 38712 27252 38740
rect 27246 38700 27252 38712
rect 27304 38740 27310 38752
rect 27769 38740 27797 38771
rect 29454 38768 29460 38780
rect 29512 38808 29518 38820
rect 29914 38817 29920 38820
rect 29870 38811 29920 38817
rect 29870 38808 29882 38811
rect 29512 38780 29882 38808
rect 29512 38768 29518 38780
rect 29870 38777 29882 38780
rect 29916 38777 29920 38811
rect 29870 38771 29920 38777
rect 29914 38768 29920 38771
rect 29972 38768 29978 38820
rect 31481 38811 31539 38817
rect 31481 38777 31493 38811
rect 31527 38777 31539 38811
rect 33321 38811 33379 38817
rect 33321 38808 33333 38811
rect 31481 38771 31539 38777
rect 33106 38780 33333 38808
rect 27304 38712 27797 38740
rect 27304 38700 27310 38712
rect 28350 38700 28356 38752
rect 28408 38740 28414 38752
rect 28721 38743 28779 38749
rect 28721 38740 28733 38743
rect 28408 38712 28733 38740
rect 28408 38700 28414 38712
rect 28721 38709 28733 38712
rect 28767 38740 28779 38743
rect 29086 38740 29092 38752
rect 28767 38712 29092 38740
rect 28767 38709 28779 38712
rect 28721 38703 28779 38709
rect 29086 38700 29092 38712
rect 29144 38700 29150 38752
rect 31110 38740 31116 38752
rect 31071 38712 31116 38740
rect 31110 38700 31116 38712
rect 31168 38740 31174 38752
rect 31496 38740 31524 38771
rect 33106 38752 33134 38780
rect 33321 38777 33333 38780
rect 33367 38777 33379 38811
rect 33321 38771 33379 38777
rect 33413 38811 33471 38817
rect 33413 38777 33425 38811
rect 33459 38808 33471 38811
rect 33594 38808 33600 38820
rect 33459 38780 33600 38808
rect 33459 38777 33471 38780
rect 33413 38771 33471 38777
rect 33594 38768 33600 38780
rect 33652 38768 33658 38820
rect 33980 38817 34008 38916
rect 34333 38913 34345 38947
rect 34379 38944 34391 38947
rect 34606 38944 34612 38956
rect 34379 38916 34612 38944
rect 34379 38913 34391 38916
rect 34333 38907 34391 38913
rect 34606 38904 34612 38916
rect 34664 38904 34670 38956
rect 36630 38904 36636 38956
rect 36688 38944 36694 38956
rect 36725 38947 36783 38953
rect 36725 38944 36737 38947
rect 36688 38916 36737 38944
rect 36688 38904 36694 38916
rect 36725 38913 36737 38916
rect 36771 38913 36783 38947
rect 40236 38944 40264 39040
rect 42797 39015 42855 39021
rect 42797 38981 42809 39015
rect 42843 39012 42855 39015
rect 42889 39015 42947 39021
rect 42889 39012 42901 39015
rect 42843 38984 42901 39012
rect 42843 38981 42855 38984
rect 42797 38975 42855 38981
rect 42889 38981 42901 38984
rect 42935 39012 42947 39015
rect 43070 39012 43076 39024
rect 42935 38984 43076 39012
rect 42935 38981 42947 38984
rect 42889 38975 42947 38981
rect 43070 38972 43076 38984
rect 43128 39012 43134 39024
rect 43438 39012 43444 39024
rect 43128 38984 43444 39012
rect 43128 38972 43134 38984
rect 43438 38972 43444 38984
rect 43496 38972 43502 39024
rect 42061 38947 42119 38953
rect 42061 38944 42073 38947
rect 40236 38916 42073 38944
rect 36725 38907 36783 38913
rect 42061 38913 42073 38916
rect 42107 38944 42119 38947
rect 43625 38947 43683 38953
rect 43625 38944 43637 38947
rect 42107 38916 43637 38944
rect 42107 38913 42119 38916
rect 42061 38907 42119 38913
rect 43625 38913 43637 38916
rect 43671 38913 43683 38947
rect 43625 38907 43683 38913
rect 35250 38876 35256 38888
rect 35211 38848 35256 38876
rect 35250 38836 35256 38848
rect 35308 38836 35314 38888
rect 35710 38876 35716 38888
rect 35671 38848 35716 38876
rect 35710 38836 35716 38848
rect 35768 38836 35774 38888
rect 40748 38879 40806 38885
rect 40748 38845 40760 38879
rect 40794 38876 40806 38879
rect 40794 38848 41184 38876
rect 40794 38845 40806 38848
rect 40748 38839 40806 38845
rect 33965 38811 34023 38817
rect 33965 38777 33977 38811
rect 34011 38808 34023 38811
rect 34330 38808 34336 38820
rect 34011 38780 34336 38808
rect 34011 38777 34023 38780
rect 33965 38771 34023 38777
rect 34330 38768 34336 38780
rect 34388 38768 34394 38820
rect 34701 38811 34759 38817
rect 34701 38777 34713 38811
rect 34747 38808 34759 38811
rect 35728 38808 35756 38836
rect 35894 38808 35900 38820
rect 34747 38780 35756 38808
rect 35855 38780 35900 38808
rect 34747 38777 34759 38780
rect 34701 38771 34759 38777
rect 35894 38768 35900 38780
rect 35952 38768 35958 38820
rect 38746 38808 38752 38820
rect 38707 38780 38752 38808
rect 38746 38768 38752 38780
rect 38804 38768 38810 38820
rect 38841 38811 38899 38817
rect 38841 38777 38853 38811
rect 38887 38777 38899 38811
rect 38841 38771 38899 38777
rect 32306 38740 32312 38752
rect 31168 38712 31524 38740
rect 32267 38712 32312 38740
rect 31168 38700 31174 38712
rect 32306 38700 32312 38712
rect 32364 38700 32370 38752
rect 33042 38740 33048 38752
rect 33003 38712 33048 38740
rect 33042 38700 33048 38712
rect 33100 38712 33134 38752
rect 33100 38700 33106 38712
rect 36170 38700 36176 38752
rect 36228 38740 36234 38752
rect 36265 38743 36323 38749
rect 36265 38740 36277 38743
rect 36228 38712 36277 38740
rect 36228 38700 36234 38712
rect 36265 38709 36277 38712
rect 36311 38740 36323 38743
rect 36354 38740 36360 38752
rect 36311 38712 36360 38740
rect 36311 38709 36323 38712
rect 36265 38703 36323 38709
rect 36354 38700 36360 38712
rect 36412 38700 36418 38752
rect 36633 38743 36691 38749
rect 36633 38709 36645 38743
rect 36679 38740 36691 38743
rect 36906 38740 36912 38752
rect 36679 38712 36912 38740
rect 36679 38709 36691 38712
rect 36633 38703 36691 38709
rect 36906 38700 36912 38712
rect 36964 38700 36970 38752
rect 37090 38740 37096 38752
rect 37051 38712 37096 38740
rect 37090 38700 37096 38712
rect 37148 38700 37154 38752
rect 38102 38740 38108 38752
rect 38063 38712 38108 38740
rect 38102 38700 38108 38712
rect 38160 38740 38166 38752
rect 38856 38740 38884 38771
rect 41156 38752 41184 38848
rect 41414 38768 41420 38820
rect 41472 38808 41478 38820
rect 41785 38811 41843 38817
rect 41785 38808 41797 38811
rect 41472 38780 41797 38808
rect 41472 38768 41478 38780
rect 41785 38777 41797 38780
rect 41831 38777 41843 38811
rect 41785 38771 41843 38777
rect 41874 38768 41880 38820
rect 41932 38808 41938 38820
rect 43349 38811 43407 38817
rect 41932 38780 41977 38808
rect 41932 38768 41938 38780
rect 43349 38777 43361 38811
rect 43395 38777 43407 38811
rect 43349 38771 43407 38777
rect 40034 38740 40040 38752
rect 38160 38712 38884 38740
rect 39995 38712 40040 38740
rect 38160 38700 38166 38712
rect 40034 38700 40040 38712
rect 40092 38700 40098 38752
rect 41138 38740 41144 38752
rect 41099 38712 41144 38740
rect 41138 38700 41144 38712
rect 41196 38700 41202 38752
rect 41598 38740 41604 38752
rect 41511 38712 41604 38740
rect 41598 38700 41604 38712
rect 41656 38740 41662 38752
rect 42889 38743 42947 38749
rect 42889 38740 42901 38743
rect 41656 38712 42901 38740
rect 41656 38700 41662 38712
rect 42889 38709 42901 38712
rect 42935 38709 42947 38743
rect 43364 38740 43392 38771
rect 43438 38768 43444 38820
rect 43496 38808 43502 38820
rect 43496 38780 43541 38808
rect 43496 38768 43502 38780
rect 43530 38740 43536 38752
rect 43364 38712 43536 38740
rect 42889 38703 42947 38709
rect 43530 38700 43536 38712
rect 43588 38740 43594 38752
rect 44269 38743 44327 38749
rect 44269 38740 44281 38743
rect 43588 38712 44281 38740
rect 43588 38700 43594 38712
rect 44269 38709 44281 38712
rect 44315 38709 44327 38743
rect 44269 38703 44327 38709
rect 1104 38650 48852 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 48852 38650
rect 1104 38576 48852 38598
rect 13722 38536 13728 38548
rect 13642 38508 13728 38536
rect 9861 38471 9919 38477
rect 9861 38437 9873 38471
rect 9907 38468 9919 38471
rect 10226 38468 10232 38480
rect 9907 38440 10232 38468
rect 9907 38437 9919 38440
rect 9861 38431 9919 38437
rect 10226 38428 10232 38440
rect 10284 38428 10290 38480
rect 13642 38468 13670 38508
rect 13722 38496 13728 38508
rect 13780 38496 13786 38548
rect 23382 38496 23388 38548
rect 23440 38536 23446 38548
rect 23753 38539 23811 38545
rect 23753 38536 23765 38539
rect 23440 38508 23765 38536
rect 23440 38496 23446 38508
rect 23753 38505 23765 38508
rect 23799 38505 23811 38539
rect 23753 38499 23811 38505
rect 24578 38496 24584 38548
rect 24636 38536 24642 38548
rect 26234 38536 26240 38548
rect 24636 38508 25589 38536
rect 26195 38508 26240 38536
rect 24636 38496 24642 38508
rect 13814 38468 13820 38480
rect 13642 38440 13820 38468
rect 13814 38428 13820 38440
rect 13872 38468 13878 38480
rect 15470 38468 15476 38480
rect 13872 38440 13965 38468
rect 15431 38440 15476 38468
rect 13872 38428 13878 38440
rect 15470 38428 15476 38440
rect 15528 38428 15534 38480
rect 20990 38468 20996 38480
rect 20951 38440 20996 38468
rect 20990 38428 20996 38440
rect 21048 38428 21054 38480
rect 21082 38428 21088 38480
rect 21140 38468 21146 38480
rect 21140 38440 21185 38468
rect 21140 38428 21146 38440
rect 22278 38428 22284 38480
rect 22336 38468 22342 38480
rect 22830 38468 22836 38480
rect 22336 38440 22836 38468
rect 22336 38428 22342 38440
rect 22830 38428 22836 38440
rect 22888 38428 22894 38480
rect 22922 38428 22928 38480
rect 22980 38468 22986 38480
rect 24213 38471 24271 38477
rect 22980 38440 23025 38468
rect 22980 38428 22986 38440
rect 24213 38437 24225 38471
rect 24259 38468 24271 38471
rect 24394 38468 24400 38480
rect 24259 38440 24400 38468
rect 24259 38437 24271 38440
rect 24213 38431 24271 38437
rect 24394 38428 24400 38440
rect 24452 38428 24458 38480
rect 24489 38471 24547 38477
rect 24489 38437 24501 38471
rect 24535 38468 24547 38471
rect 25130 38468 25136 38480
rect 24535 38440 25136 38468
rect 24535 38437 24547 38440
rect 24489 38431 24547 38437
rect 25130 38428 25136 38440
rect 25188 38428 25194 38480
rect 25561 38468 25589 38508
rect 26234 38496 26240 38508
rect 26292 38496 26298 38548
rect 27982 38496 27988 38548
rect 28040 38536 28046 38548
rect 28077 38539 28135 38545
rect 28077 38536 28089 38539
rect 28040 38508 28089 38536
rect 28040 38496 28046 38508
rect 28077 38505 28089 38508
rect 28123 38505 28135 38539
rect 29270 38536 29276 38548
rect 29231 38508 29276 38536
rect 28077 38499 28135 38505
rect 26602 38468 26608 38480
rect 25561 38440 26608 38468
rect 26602 38428 26608 38440
rect 26660 38428 26666 38480
rect 26694 38428 26700 38480
rect 26752 38468 26758 38480
rect 28092 38468 28120 38499
rect 29270 38496 29276 38508
rect 29328 38496 29334 38548
rect 30745 38539 30803 38545
rect 30745 38505 30757 38539
rect 30791 38505 30803 38539
rect 30745 38499 30803 38505
rect 32585 38539 32643 38545
rect 32585 38505 32597 38539
rect 32631 38536 32643 38539
rect 33042 38536 33048 38548
rect 32631 38508 33048 38536
rect 32631 38505 32643 38508
rect 32585 38499 32643 38505
rect 30760 38468 30788 38499
rect 33042 38496 33048 38508
rect 33100 38496 33106 38548
rect 33321 38539 33379 38545
rect 33321 38505 33333 38539
rect 33367 38536 33379 38539
rect 33594 38536 33600 38548
rect 33367 38508 33600 38536
rect 33367 38505 33379 38508
rect 33321 38499 33379 38505
rect 33594 38496 33600 38508
rect 33652 38496 33658 38548
rect 33962 38496 33968 38548
rect 34020 38536 34026 38548
rect 34609 38539 34667 38545
rect 34609 38536 34621 38539
rect 34020 38508 34621 38536
rect 34020 38496 34026 38508
rect 34609 38505 34621 38508
rect 34655 38505 34667 38539
rect 34609 38499 34667 38505
rect 36630 38496 36636 38548
rect 36688 38536 36694 38548
rect 37093 38539 37151 38545
rect 37093 38536 37105 38539
rect 36688 38508 37105 38536
rect 36688 38496 36694 38508
rect 37093 38505 37105 38508
rect 37139 38505 37151 38539
rect 37093 38499 37151 38505
rect 38657 38539 38715 38545
rect 38657 38505 38669 38539
rect 38703 38536 38715 38539
rect 40034 38536 40040 38548
rect 38703 38508 40040 38536
rect 38703 38505 38715 38508
rect 38657 38499 38715 38505
rect 40034 38496 40040 38508
rect 40092 38496 40098 38548
rect 41506 38536 41512 38548
rect 41467 38508 41512 38536
rect 41506 38496 41512 38508
rect 41564 38496 41570 38548
rect 41874 38496 41880 38548
rect 41932 38536 41938 38548
rect 42153 38539 42211 38545
rect 42153 38536 42165 38539
rect 41932 38508 42165 38536
rect 41932 38496 41938 38508
rect 42153 38505 42165 38508
rect 42199 38505 42211 38539
rect 43530 38536 43536 38548
rect 43491 38508 43536 38536
rect 42153 38499 42211 38505
rect 43530 38496 43536 38508
rect 43588 38496 43594 38548
rect 33686 38468 33692 38480
rect 26752 38440 26797 38468
rect 28092 38440 30788 38468
rect 33647 38440 33692 38468
rect 26752 38428 26758 38440
rect 33686 38428 33692 38440
rect 33744 38428 33750 38480
rect 33778 38428 33784 38480
rect 33836 38468 33842 38480
rect 33836 38440 33881 38468
rect 33836 38428 33842 38440
rect 35710 38428 35716 38480
rect 35768 38468 35774 38480
rect 35989 38471 36047 38477
rect 35989 38468 36001 38471
rect 35768 38440 36001 38468
rect 35768 38428 35774 38440
rect 35989 38437 36001 38440
rect 36035 38468 36047 38471
rect 36035 38440 36584 38468
rect 36035 38437 36047 38440
rect 35989 38431 36047 38437
rect 36556 38412 36584 38440
rect 36998 38428 37004 38480
rect 37056 38468 37062 38480
rect 38058 38471 38116 38477
rect 38058 38468 38070 38471
rect 37056 38440 38070 38468
rect 37056 38428 37062 38440
rect 38058 38437 38070 38440
rect 38104 38437 38116 38471
rect 38058 38431 38116 38437
rect 38746 38428 38752 38480
rect 38804 38468 38810 38480
rect 38933 38471 38991 38477
rect 38933 38468 38945 38471
rect 38804 38440 38945 38468
rect 38804 38428 38810 38440
rect 38933 38437 38945 38440
rect 38979 38437 38991 38471
rect 38933 38431 38991 38437
rect 39114 38428 39120 38480
rect 39172 38468 39178 38480
rect 39806 38471 39864 38477
rect 39806 38468 39818 38471
rect 39172 38440 39818 38468
rect 39172 38428 39178 38440
rect 39806 38437 39818 38440
rect 39852 38437 39864 38471
rect 39806 38431 39864 38437
rect 11882 38400 11888 38412
rect 11843 38372 11888 38400
rect 11882 38360 11888 38372
rect 11940 38360 11946 38412
rect 16920 38403 16978 38409
rect 16920 38369 16932 38403
rect 16966 38400 16978 38403
rect 17770 38400 17776 38412
rect 16966 38372 17776 38400
rect 16966 38369 16978 38372
rect 16920 38363 16978 38369
rect 17770 38360 17776 38372
rect 17828 38360 17834 38412
rect 18969 38403 19027 38409
rect 18969 38369 18981 38403
rect 19015 38400 19027 38403
rect 19058 38400 19064 38412
rect 19015 38372 19064 38400
rect 19015 38369 19027 38372
rect 18969 38363 19027 38369
rect 19058 38360 19064 38372
rect 19116 38360 19122 38412
rect 29273 38403 29331 38409
rect 29273 38369 29285 38403
rect 29319 38369 29331 38403
rect 29546 38400 29552 38412
rect 29507 38372 29552 38400
rect 29273 38363 29331 38369
rect 9769 38335 9827 38341
rect 9769 38301 9781 38335
rect 9815 38301 9827 38335
rect 10042 38332 10048 38344
rect 10003 38304 10048 38332
rect 9769 38295 9827 38301
rect 7190 38224 7196 38276
rect 7248 38264 7254 38276
rect 9401 38267 9459 38273
rect 9401 38264 9413 38267
rect 7248 38236 9413 38264
rect 7248 38224 7254 38236
rect 9401 38233 9413 38236
rect 9447 38264 9459 38267
rect 9784 38264 9812 38295
rect 10042 38292 10048 38304
rect 10100 38332 10106 38344
rect 10781 38335 10839 38341
rect 10781 38332 10793 38335
rect 10100 38304 10793 38332
rect 10100 38292 10106 38304
rect 10781 38301 10793 38304
rect 10827 38332 10839 38335
rect 10870 38332 10876 38344
rect 10827 38304 10876 38332
rect 10827 38301 10839 38304
rect 10781 38295 10839 38301
rect 10870 38292 10876 38304
rect 10928 38292 10934 38344
rect 11238 38332 11244 38344
rect 11199 38304 11244 38332
rect 11238 38292 11244 38304
rect 11296 38292 11302 38344
rect 13170 38292 13176 38344
rect 13228 38332 13234 38344
rect 13725 38335 13783 38341
rect 13725 38332 13737 38335
rect 13228 38304 13737 38332
rect 13228 38292 13234 38304
rect 13725 38301 13737 38304
rect 13771 38301 13783 38335
rect 15378 38332 15384 38344
rect 13725 38295 13783 38301
rect 14200 38304 15384 38332
rect 9447 38236 9812 38264
rect 9447 38233 9459 38236
rect 9401 38227 9459 38233
rect 11146 38224 11152 38276
rect 11204 38264 11210 38276
rect 14200 38264 14228 38304
rect 15378 38292 15384 38304
rect 15436 38292 15442 38344
rect 15657 38335 15715 38341
rect 15657 38301 15669 38335
rect 15703 38332 15715 38335
rect 16114 38332 16120 38344
rect 15703 38304 16120 38332
rect 15703 38301 15715 38304
rect 15657 38295 15715 38301
rect 11204 38236 14228 38264
rect 14277 38267 14335 38273
rect 11204 38224 11210 38236
rect 14277 38233 14289 38267
rect 14323 38264 14335 38267
rect 15672 38264 15700 38295
rect 16114 38292 16120 38304
rect 16172 38292 16178 38344
rect 21637 38335 21695 38341
rect 21637 38301 21649 38335
rect 21683 38332 21695 38335
rect 21910 38332 21916 38344
rect 21683 38304 21916 38332
rect 21683 38301 21695 38304
rect 21637 38295 21695 38301
rect 21910 38292 21916 38304
rect 21968 38292 21974 38344
rect 24673 38335 24731 38341
rect 24673 38301 24685 38335
rect 24719 38332 24731 38335
rect 25314 38332 25320 38344
rect 24719 38304 25320 38332
rect 24719 38301 24731 38304
rect 24673 38295 24731 38301
rect 14323 38236 15700 38264
rect 14323 38233 14335 38236
rect 14277 38227 14335 38233
rect 16850 38224 16856 38276
rect 16908 38264 16914 38276
rect 16991 38267 17049 38273
rect 16991 38264 17003 38267
rect 16908 38236 17003 38264
rect 16908 38224 16914 38236
rect 16991 38233 17003 38236
rect 17037 38233 17049 38267
rect 16991 38227 17049 38233
rect 23385 38267 23443 38273
rect 23385 38233 23397 38267
rect 23431 38264 23443 38267
rect 24688 38264 24716 38295
rect 25314 38292 25320 38304
rect 25372 38292 25378 38344
rect 26881 38335 26939 38341
rect 26881 38301 26893 38335
rect 26927 38301 26939 38335
rect 26881 38295 26939 38301
rect 23431 38236 24716 38264
rect 25332 38264 25360 38292
rect 26896 38264 26924 38295
rect 29086 38292 29092 38344
rect 29144 38332 29150 38344
rect 29288 38332 29316 38363
rect 29546 38360 29552 38372
rect 29604 38360 29610 38412
rect 30558 38400 30564 38412
rect 30519 38372 30564 38400
rect 30558 38360 30564 38372
rect 30616 38360 30622 38412
rect 32858 38360 32864 38412
rect 32916 38400 32922 38412
rect 33042 38400 33048 38412
rect 32916 38372 33048 38400
rect 32916 38360 32922 38372
rect 33042 38360 33048 38372
rect 33100 38360 33106 38412
rect 36078 38400 36084 38412
rect 36039 38372 36084 38400
rect 36078 38360 36084 38372
rect 36136 38360 36142 38412
rect 36538 38400 36544 38412
rect 36499 38372 36544 38400
rect 36538 38360 36544 38372
rect 36596 38360 36602 38412
rect 36817 38403 36875 38409
rect 36817 38369 36829 38403
rect 36863 38400 36875 38403
rect 39482 38400 39488 38412
rect 36863 38372 39488 38400
rect 36863 38369 36875 38372
rect 36817 38363 36875 38369
rect 39482 38360 39488 38372
rect 39540 38360 39546 38412
rect 40405 38403 40463 38409
rect 40405 38369 40417 38403
rect 40451 38400 40463 38403
rect 41874 38400 41880 38412
rect 40451 38372 41880 38400
rect 40451 38369 40463 38372
rect 40405 38363 40463 38369
rect 41874 38360 41880 38372
rect 41932 38360 41938 38412
rect 43416 38403 43474 38409
rect 43416 38369 43428 38403
rect 43462 38400 43474 38403
rect 43806 38400 43812 38412
rect 43462 38372 43812 38400
rect 43462 38369 43474 38372
rect 43416 38363 43474 38369
rect 43806 38360 43812 38372
rect 43864 38360 43870 38412
rect 34330 38332 34336 38344
rect 29144 38304 30880 38332
rect 29144 38292 29150 38304
rect 25332 38236 26924 38264
rect 23431 38233 23443 38236
rect 23385 38227 23443 38233
rect 7650 38196 7656 38208
rect 7611 38168 7656 38196
rect 7650 38156 7656 38168
rect 7708 38156 7714 38208
rect 19199 38199 19257 38205
rect 19199 38165 19211 38199
rect 19245 38196 19257 38199
rect 19334 38196 19340 38208
rect 19245 38168 19340 38196
rect 19245 38165 19257 38168
rect 19199 38159 19257 38165
rect 19334 38156 19340 38168
rect 19392 38156 19398 38208
rect 19610 38196 19616 38208
rect 19523 38168 19616 38196
rect 19610 38156 19616 38168
rect 19668 38196 19674 38208
rect 21082 38196 21088 38208
rect 19668 38168 21088 38196
rect 19668 38156 19674 38168
rect 21082 38156 21088 38168
rect 21140 38156 21146 38208
rect 21726 38156 21732 38208
rect 21784 38196 21790 38208
rect 21913 38199 21971 38205
rect 21913 38196 21925 38199
rect 21784 38168 21925 38196
rect 21784 38156 21790 38168
rect 21913 38165 21925 38168
rect 21959 38165 21971 38199
rect 25498 38196 25504 38208
rect 25459 38168 25504 38196
rect 21913 38159 21971 38165
rect 25498 38156 25504 38168
rect 25556 38156 25562 38208
rect 30190 38196 30196 38208
rect 30151 38168 30196 38196
rect 30190 38156 30196 38168
rect 30248 38156 30254 38208
rect 30852 38196 30880 38304
rect 33106 38304 34336 38332
rect 31389 38267 31447 38273
rect 31389 38233 31401 38267
rect 31435 38264 31447 38267
rect 33106 38264 33134 38304
rect 34330 38292 34336 38304
rect 34388 38292 34394 38344
rect 35894 38292 35900 38344
rect 35952 38332 35958 38344
rect 37737 38335 37795 38341
rect 37737 38332 37749 38335
rect 35952 38304 37749 38332
rect 35952 38292 35958 38304
rect 37737 38301 37749 38304
rect 37783 38332 37795 38335
rect 37918 38332 37924 38344
rect 37783 38304 37924 38332
rect 37783 38301 37795 38304
rect 37737 38295 37795 38301
rect 37918 38292 37924 38304
rect 37976 38292 37982 38344
rect 38654 38292 38660 38344
rect 38712 38332 38718 38344
rect 39301 38335 39359 38341
rect 39301 38332 39313 38335
rect 38712 38304 39313 38332
rect 38712 38292 38718 38304
rect 39301 38301 39313 38304
rect 39347 38301 39359 38335
rect 41690 38332 41696 38344
rect 41651 38304 41696 38332
rect 39301 38295 39359 38301
rect 41690 38292 41696 38304
rect 41748 38292 41754 38344
rect 31435 38236 33134 38264
rect 31435 38233 31447 38236
rect 31389 38227 31447 38233
rect 41414 38224 41420 38276
rect 41472 38264 41478 38276
rect 42521 38267 42579 38273
rect 42521 38264 42533 38267
rect 41472 38236 42533 38264
rect 41472 38224 41478 38236
rect 42521 38233 42533 38236
rect 42567 38233 42579 38267
rect 42521 38227 42579 38233
rect 35250 38196 35256 38208
rect 30852 38168 35256 38196
rect 35250 38156 35256 38168
rect 35308 38156 35314 38208
rect 1104 38106 48852 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 48852 38106
rect 1104 38032 48852 38054
rect 11882 37992 11888 38004
rect 11843 37964 11888 37992
rect 11882 37952 11888 37964
rect 11940 37952 11946 38004
rect 11974 37952 11980 38004
rect 12032 37992 12038 38004
rect 12621 37995 12679 38001
rect 12621 37992 12633 37995
rect 12032 37964 12633 37992
rect 12032 37952 12038 37964
rect 12621 37961 12633 37964
rect 12667 37961 12679 37995
rect 12621 37955 12679 37961
rect 12802 37952 12808 38004
rect 12860 37992 12866 38004
rect 12897 37995 12955 38001
rect 12897 37992 12909 37995
rect 12860 37964 12909 37992
rect 12860 37952 12866 37964
rect 12897 37961 12909 37964
rect 12943 37961 12955 37995
rect 12897 37955 12955 37961
rect 13633 37995 13691 38001
rect 13633 37961 13645 37995
rect 13679 37992 13691 37995
rect 13814 37992 13820 38004
rect 13679 37964 13820 37992
rect 13679 37961 13691 37964
rect 13633 37955 13691 37961
rect 13814 37952 13820 37964
rect 13872 37952 13878 38004
rect 14185 37995 14243 38001
rect 14185 37961 14197 37995
rect 14231 37992 14243 37995
rect 15197 37995 15255 38001
rect 15197 37992 15209 37995
rect 14231 37964 15209 37992
rect 14231 37961 14243 37964
rect 14185 37955 14243 37961
rect 15197 37961 15209 37964
rect 15243 37992 15255 37995
rect 15470 37992 15476 38004
rect 15243 37964 15476 37992
rect 15243 37961 15255 37964
rect 15197 37955 15255 37961
rect 15470 37952 15476 37964
rect 15528 37952 15534 38004
rect 17770 37992 17776 38004
rect 17731 37964 17776 37992
rect 17770 37952 17776 37964
rect 17828 37952 17834 38004
rect 19058 37992 19064 38004
rect 19019 37964 19064 37992
rect 19058 37952 19064 37964
rect 19116 37952 19122 38004
rect 20625 37995 20683 38001
rect 20625 37961 20637 37995
rect 20671 37992 20683 37995
rect 20990 37992 20996 38004
rect 20671 37964 20996 37992
rect 20671 37961 20683 37964
rect 20625 37955 20683 37961
rect 20990 37952 20996 37964
rect 21048 37952 21054 38004
rect 22830 37992 22836 38004
rect 22791 37964 22836 37992
rect 22830 37952 22836 37964
rect 22888 37952 22894 38004
rect 23477 37995 23535 38001
rect 23477 37961 23489 37995
rect 23523 37992 23535 37995
rect 23750 37992 23756 38004
rect 23523 37964 23756 37992
rect 23523 37961 23535 37964
rect 23477 37955 23535 37961
rect 23750 37952 23756 37964
rect 23808 37992 23814 38004
rect 25130 37992 25136 38004
rect 23808 37964 25136 37992
rect 23808 37952 23814 37964
rect 25130 37952 25136 37964
rect 25188 37952 25194 38004
rect 25498 37952 25504 38004
rect 25556 37992 25562 38004
rect 27433 37995 27491 38001
rect 27433 37992 27445 37995
rect 25556 37964 27445 37992
rect 25556 37952 25562 37964
rect 27433 37961 27445 37964
rect 27479 37961 27491 37995
rect 29086 37992 29092 38004
rect 29047 37964 29092 37992
rect 27433 37955 27491 37961
rect 29086 37952 29092 37964
rect 29144 37952 29150 38004
rect 29914 37992 29920 38004
rect 29875 37964 29920 37992
rect 29914 37952 29920 37964
rect 29972 37952 29978 38004
rect 31021 37995 31079 38001
rect 31021 37961 31033 37995
rect 31067 37992 31079 37995
rect 31110 37992 31116 38004
rect 31067 37964 31116 37992
rect 31067 37961 31079 37964
rect 31021 37955 31079 37961
rect 31110 37952 31116 37964
rect 31168 37952 31174 38004
rect 33686 37952 33692 38004
rect 33744 37992 33750 38004
rect 34057 37995 34115 38001
rect 34057 37992 34069 37995
rect 33744 37964 34069 37992
rect 33744 37952 33750 37964
rect 34057 37961 34069 37964
rect 34103 37961 34115 37995
rect 36998 37992 37004 38004
rect 36959 37964 37004 37992
rect 34057 37955 34115 37961
rect 36998 37952 37004 37964
rect 37056 37952 37062 38004
rect 38102 37992 38108 38004
rect 38063 37964 38108 37992
rect 38102 37952 38108 37964
rect 38160 37952 38166 38004
rect 38841 37995 38899 38001
rect 38841 37961 38853 37995
rect 38887 37992 38899 37995
rect 39298 37992 39304 38004
rect 38887 37964 39304 37992
rect 38887 37961 38899 37964
rect 38841 37955 38899 37961
rect 10226 37924 10232 37936
rect 10139 37896 10232 37924
rect 10226 37884 10232 37896
rect 10284 37924 10290 37936
rect 10284 37896 13814 37924
rect 10284 37884 10290 37896
rect 8294 37856 8300 37868
rect 8255 37828 8300 37856
rect 8294 37816 8300 37828
rect 8352 37816 8358 37868
rect 9490 37856 9496 37868
rect 8404 37828 9496 37856
rect 7650 37720 7656 37732
rect 7611 37692 7656 37720
rect 7650 37680 7656 37692
rect 7708 37680 7714 37732
rect 7745 37723 7803 37729
rect 7745 37689 7757 37723
rect 7791 37720 7803 37723
rect 8404 37720 8432 37828
rect 9490 37816 9496 37828
rect 9548 37816 9554 37868
rect 9861 37859 9919 37865
rect 9861 37825 9873 37859
rect 9907 37856 9919 37859
rect 10042 37856 10048 37868
rect 9907 37828 10048 37856
rect 9907 37825 9919 37828
rect 9861 37819 9919 37825
rect 10042 37816 10048 37828
rect 10100 37816 10106 37868
rect 13786 37856 13814 37896
rect 13998 37884 14004 37936
rect 14056 37924 14062 37936
rect 14056 37896 17769 37924
rect 14056 37884 14062 37896
rect 13906 37856 13912 37868
rect 13786 37828 13912 37856
rect 13906 37816 13912 37828
rect 13964 37856 13970 37868
rect 15289 37859 15347 37865
rect 15289 37856 15301 37859
rect 13964 37828 15301 37856
rect 13964 37816 13970 37828
rect 15289 37825 15301 37828
rect 15335 37825 15347 37859
rect 15289 37819 15347 37825
rect 12437 37791 12495 37797
rect 12437 37757 12449 37791
rect 12483 37788 12495 37791
rect 12802 37788 12808 37800
rect 12483 37760 12808 37788
rect 12483 37757 12495 37760
rect 12437 37751 12495 37757
rect 12802 37748 12808 37760
rect 12860 37748 12866 37800
rect 13630 37748 13636 37800
rect 13688 37788 13694 37800
rect 13817 37791 13875 37797
rect 13817 37788 13829 37791
rect 13688 37760 13829 37788
rect 13688 37748 13694 37760
rect 13817 37757 13829 37760
rect 13863 37757 13875 37791
rect 13817 37751 13875 37757
rect 15933 37791 15991 37797
rect 15933 37757 15945 37791
rect 15979 37757 15991 37791
rect 16850 37788 16856 37800
rect 16763 37760 16856 37788
rect 15933 37751 15991 37757
rect 9030 37720 9036 37732
rect 7791 37692 8432 37720
rect 8991 37692 9036 37720
rect 7791 37689 7803 37692
rect 7745 37683 7803 37689
rect 7469 37655 7527 37661
rect 7469 37621 7481 37655
rect 7515 37652 7527 37655
rect 7760 37652 7788 37683
rect 9030 37680 9036 37692
rect 9088 37680 9094 37732
rect 9214 37720 9220 37732
rect 9175 37692 9220 37720
rect 9214 37680 9220 37692
rect 9272 37680 9278 37732
rect 9318 37723 9376 37729
rect 9318 37689 9330 37723
rect 9364 37689 9376 37723
rect 9318 37683 9376 37689
rect 7515 37624 7788 37652
rect 9048 37652 9076 37680
rect 9324 37652 9352 37683
rect 9490 37680 9496 37732
rect 9548 37720 9554 37732
rect 10870 37720 10876 37732
rect 9548 37692 10732 37720
rect 10831 37692 10876 37720
rect 9548 37680 9554 37692
rect 10704 37661 10732 37692
rect 10870 37680 10876 37692
rect 10928 37680 10934 37732
rect 10965 37723 11023 37729
rect 10965 37689 10977 37723
rect 11011 37720 11023 37723
rect 11238 37720 11244 37732
rect 11011 37692 11244 37720
rect 11011 37689 11023 37692
rect 10965 37683 11023 37689
rect 9048 37624 9352 37652
rect 10689 37655 10747 37661
rect 7515 37621 7527 37624
rect 7469 37615 7527 37621
rect 10689 37621 10701 37655
rect 10735 37652 10747 37655
rect 10980 37652 11008 37683
rect 11238 37680 11244 37692
rect 11296 37680 11302 37732
rect 11517 37723 11575 37729
rect 11517 37689 11529 37723
rect 11563 37720 11575 37723
rect 13170 37720 13176 37732
rect 11563 37692 13176 37720
rect 11563 37689 11575 37692
rect 11517 37683 11575 37689
rect 13170 37680 13176 37692
rect 13228 37680 13234 37732
rect 14829 37723 14887 37729
rect 14829 37689 14841 37723
rect 14875 37720 14887 37723
rect 15948 37720 15976 37751
rect 16850 37748 16856 37760
rect 16908 37788 16914 37800
rect 17313 37791 17371 37797
rect 17313 37788 17325 37791
rect 16908 37760 17325 37788
rect 16908 37748 16914 37760
rect 17313 37757 17325 37760
rect 17359 37757 17371 37791
rect 17741 37788 17769 37896
rect 26602 37884 26608 37936
rect 26660 37924 26666 37936
rect 28077 37927 28135 37933
rect 28077 37924 28089 37927
rect 26660 37896 28089 37924
rect 26660 37884 26666 37896
rect 28077 37893 28089 37896
rect 28123 37893 28135 37927
rect 28077 37887 28135 37893
rect 30834 37884 30840 37936
rect 30892 37924 30898 37936
rect 33413 37927 33471 37933
rect 30892 37896 33134 37924
rect 30892 37884 30898 37896
rect 19334 37816 19340 37868
rect 19392 37856 19398 37868
rect 19521 37859 19579 37865
rect 19521 37856 19533 37859
rect 19392 37828 19533 37856
rect 19392 37816 19398 37828
rect 19521 37825 19533 37828
rect 19567 37825 19579 37859
rect 19521 37819 19579 37825
rect 20993 37859 21051 37865
rect 20993 37825 21005 37859
rect 21039 37856 21051 37859
rect 21082 37856 21088 37868
rect 21039 37828 21088 37856
rect 21039 37825 21051 37828
rect 20993 37819 21051 37825
rect 21082 37816 21088 37828
rect 21140 37816 21146 37868
rect 21637 37859 21695 37865
rect 21637 37825 21649 37859
rect 21683 37856 21695 37859
rect 21726 37856 21732 37868
rect 21683 37828 21732 37856
rect 21683 37825 21695 37828
rect 21637 37819 21695 37825
rect 21726 37816 21732 37828
rect 21784 37816 21790 37868
rect 21910 37856 21916 37868
rect 21871 37828 21916 37856
rect 21910 37816 21916 37828
rect 21968 37816 21974 37868
rect 25317 37859 25375 37865
rect 25317 37825 25329 37859
rect 25363 37856 25375 37859
rect 26329 37859 26387 37865
rect 26329 37856 26341 37859
rect 25363 37828 26341 37856
rect 25363 37825 25375 37828
rect 25317 37819 25375 37825
rect 26329 37825 26341 37828
rect 26375 37825 26387 37859
rect 26329 37819 26387 37825
rect 29730 37816 29736 37868
rect 29788 37856 29794 37868
rect 30558 37856 30564 37868
rect 29788 37828 30564 37856
rect 29788 37816 29794 37828
rect 30558 37816 30564 37828
rect 30616 37856 30622 37868
rect 31297 37859 31355 37865
rect 31297 37856 31309 37859
rect 30616 37828 31309 37856
rect 30616 37816 30622 37828
rect 31297 37825 31309 37828
rect 31343 37825 31355 37859
rect 33106 37856 33134 37896
rect 33413 37893 33425 37927
rect 33459 37924 33471 37927
rect 33778 37924 33784 37936
rect 33459 37896 33784 37924
rect 33459 37893 33471 37896
rect 33413 37887 33471 37893
rect 33778 37884 33784 37896
rect 33836 37884 33842 37936
rect 36078 37924 36084 37936
rect 33888 37896 36084 37924
rect 33888 37856 33916 37896
rect 36078 37884 36084 37896
rect 36136 37884 36142 37936
rect 33106 37828 33916 37856
rect 31297 37819 31355 37825
rect 34330 37816 34336 37868
rect 34388 37856 34394 37868
rect 35253 37859 35311 37865
rect 35253 37856 35265 37859
rect 34388 37828 35265 37856
rect 34388 37816 34394 37828
rect 35253 37825 35265 37828
rect 35299 37825 35311 37859
rect 35253 37819 35311 37825
rect 37185 37859 37243 37865
rect 37185 37825 37197 37859
rect 37231 37856 37243 37859
rect 37550 37856 37556 37868
rect 37231 37828 37556 37856
rect 37231 37825 37243 37828
rect 37185 37819 37243 37825
rect 37550 37816 37556 37828
rect 37608 37816 37614 37868
rect 37826 37816 37832 37868
rect 37884 37856 37890 37868
rect 39071 37859 39129 37865
rect 39071 37856 39083 37859
rect 37884 37828 39083 37856
rect 37884 37816 37890 37828
rect 39071 37825 39083 37828
rect 39117 37825 39129 37859
rect 39071 37819 39129 37825
rect 18084 37791 18142 37797
rect 18084 37788 18096 37791
rect 17741 37760 18096 37788
rect 17313 37751 17371 37757
rect 18084 37757 18096 37760
rect 18130 37788 18142 37791
rect 18509 37791 18567 37797
rect 18509 37788 18521 37791
rect 18130 37760 18521 37788
rect 18130 37757 18142 37760
rect 18084 37751 18142 37757
rect 18509 37757 18521 37760
rect 18555 37788 18567 37791
rect 19242 37788 19248 37800
rect 18555 37760 19248 37788
rect 18555 37757 18567 37760
rect 18509 37751 18567 37757
rect 19242 37748 19248 37760
rect 19300 37748 19306 37800
rect 24213 37791 24271 37797
rect 24213 37757 24225 37791
rect 24259 37788 24271 37791
rect 26510 37788 26516 37800
rect 24259 37760 25544 37788
rect 26471 37760 26516 37788
rect 24259 37757 24271 37760
rect 24213 37751 24271 37757
rect 19610 37720 19616 37732
rect 14875 37692 15976 37720
rect 19571 37692 19616 37720
rect 14875 37689 14887 37692
rect 14829 37683 14887 37689
rect 10735 37624 11008 37652
rect 15948 37652 15976 37692
rect 19610 37680 19616 37692
rect 19668 37680 19674 37732
rect 20162 37720 20168 37732
rect 20123 37692 20168 37720
rect 20162 37680 20168 37692
rect 20220 37680 20226 37732
rect 21729 37723 21787 37729
rect 21729 37689 21741 37723
rect 21775 37689 21787 37723
rect 24534 37723 24592 37729
rect 24534 37720 24546 37723
rect 21729 37683 21787 37689
rect 24044 37692 24546 37720
rect 17037 37655 17095 37661
rect 17037 37652 17049 37655
rect 15948 37624 17049 37652
rect 10735 37621 10747 37624
rect 10689 37615 10747 37621
rect 17037 37621 17049 37624
rect 17083 37621 17095 37655
rect 17037 37615 17095 37621
rect 18187 37655 18245 37661
rect 18187 37621 18199 37655
rect 18233 37652 18245 37655
rect 18322 37652 18328 37664
rect 18233 37624 18328 37652
rect 18233 37621 18245 37624
rect 18187 37615 18245 37621
rect 18322 37612 18328 37624
rect 18380 37612 18386 37664
rect 21453 37655 21511 37661
rect 21453 37621 21465 37655
rect 21499 37652 21511 37655
rect 21744 37652 21772 37683
rect 21818 37652 21824 37664
rect 21499 37624 21824 37652
rect 21499 37621 21511 37624
rect 21453 37615 21511 37621
rect 21818 37612 21824 37624
rect 21876 37612 21882 37664
rect 23842 37612 23848 37664
rect 23900 37652 23906 37664
rect 24044 37661 24072 37692
rect 24534 37689 24546 37692
rect 24580 37720 24592 37723
rect 25317 37723 25375 37729
rect 25317 37720 25329 37723
rect 24580 37692 25329 37720
rect 24580 37689 24592 37692
rect 24534 37683 24592 37689
rect 25317 37689 25329 37692
rect 25363 37689 25375 37723
rect 25317 37683 25375 37689
rect 25516 37661 25544 37760
rect 26510 37748 26516 37760
rect 26568 37788 26574 37800
rect 27709 37791 27767 37797
rect 27709 37788 27721 37791
rect 26568 37760 27721 37788
rect 26568 37748 26574 37760
rect 27709 37757 27721 37760
rect 27755 37757 27767 37791
rect 29546 37788 29552 37800
rect 29459 37760 29552 37788
rect 27709 37751 27767 37757
rect 29546 37748 29552 37760
rect 29604 37788 29610 37800
rect 29914 37788 29920 37800
rect 29604 37760 29920 37788
rect 29604 37748 29610 37760
rect 29914 37748 29920 37760
rect 29972 37748 29978 37800
rect 30101 37791 30159 37797
rect 30101 37757 30113 37791
rect 30147 37788 30159 37791
rect 30190 37788 30196 37800
rect 30147 37760 30196 37788
rect 30147 37757 30159 37760
rect 30101 37751 30159 37757
rect 30190 37748 30196 37760
rect 30248 37748 30254 37800
rect 32398 37748 32404 37800
rect 32456 37788 32462 37800
rect 32493 37791 32551 37797
rect 32493 37788 32505 37791
rect 32456 37760 32505 37788
rect 32456 37748 32462 37760
rect 32493 37757 32505 37760
rect 32539 37757 32551 37791
rect 32493 37751 32551 37757
rect 36998 37748 37004 37800
rect 37056 37788 37062 37800
rect 38381 37791 38439 37797
rect 38381 37788 38393 37791
rect 37056 37760 38393 37788
rect 37056 37748 37062 37760
rect 26694 37720 26700 37732
rect 25976 37692 26700 37720
rect 25976 37664 26004 37692
rect 26694 37680 26700 37692
rect 26752 37680 26758 37732
rect 30006 37680 30012 37732
rect 30064 37720 30070 37732
rect 30422 37723 30480 37729
rect 30422 37720 30434 37723
rect 30064 37692 30434 37720
rect 30064 37680 30070 37692
rect 30422 37689 30434 37692
rect 30468 37720 30480 37723
rect 32306 37720 32312 37732
rect 30468 37692 32312 37720
rect 30468 37689 30480 37692
rect 30422 37683 30480 37689
rect 32306 37680 32312 37692
rect 32364 37720 32370 37732
rect 32814 37723 32872 37729
rect 32814 37720 32826 37723
rect 32364 37692 32826 37720
rect 32364 37680 32370 37692
rect 32814 37689 32826 37692
rect 32860 37689 32872 37723
rect 32814 37683 32872 37689
rect 34790 37680 34796 37732
rect 34848 37720 34854 37732
rect 34977 37723 35035 37729
rect 34977 37720 34989 37723
rect 34848 37692 34989 37720
rect 34848 37680 34854 37692
rect 34977 37689 34989 37692
rect 35023 37689 35035 37723
rect 34977 37683 35035 37689
rect 35069 37723 35127 37729
rect 35069 37689 35081 37723
rect 35115 37689 35127 37723
rect 36538 37720 36544 37732
rect 36451 37692 36544 37720
rect 35069 37683 35127 37689
rect 24029 37655 24087 37661
rect 24029 37652 24041 37655
rect 23900 37624 24041 37652
rect 23900 37612 23906 37624
rect 24029 37621 24041 37624
rect 24075 37621 24087 37655
rect 24029 37615 24087 37621
rect 25501 37655 25559 37661
rect 25501 37621 25513 37655
rect 25547 37652 25559 37655
rect 25682 37652 25688 37664
rect 25547 37624 25688 37652
rect 25547 37621 25559 37624
rect 25501 37615 25559 37621
rect 25682 37612 25688 37624
rect 25740 37612 25746 37664
rect 25958 37652 25964 37664
rect 25919 37624 25964 37652
rect 25958 37612 25964 37624
rect 26016 37612 26022 37664
rect 26881 37655 26939 37661
rect 26881 37621 26893 37655
rect 26927 37652 26939 37655
rect 27246 37652 27252 37664
rect 26927 37624 27252 37652
rect 26927 37621 26939 37624
rect 26881 37615 26939 37621
rect 27246 37612 27252 37624
rect 27304 37612 27310 37664
rect 34606 37652 34612 37664
rect 34567 37624 34612 37652
rect 34606 37612 34612 37624
rect 34664 37652 34670 37664
rect 35084 37652 35112 37683
rect 36538 37680 36544 37692
rect 36596 37720 36602 37732
rect 37090 37720 37096 37732
rect 36596 37692 37096 37720
rect 36596 37680 36602 37692
rect 37090 37680 37096 37692
rect 37148 37680 37154 37732
rect 37522 37729 37550 37760
rect 38381 37757 38393 37760
rect 38427 37757 38439 37791
rect 38381 37751 38439 37757
rect 38984 37791 39042 37797
rect 38984 37757 38996 37791
rect 39030 37788 39042 37791
rect 39178 37788 39206 37964
rect 39298 37952 39304 37964
rect 39356 37952 39362 38004
rect 39482 37952 39488 38004
rect 39540 37992 39546 38004
rect 39853 37995 39911 38001
rect 39853 37992 39865 37995
rect 39540 37964 39865 37992
rect 39540 37952 39546 37964
rect 39853 37961 39865 37964
rect 39899 37961 39911 37995
rect 39853 37955 39911 37961
rect 40911 37995 40969 38001
rect 40911 37961 40923 37995
rect 40957 37992 40969 37995
rect 41414 37992 41420 38004
rect 40957 37964 41420 37992
rect 40957 37961 40969 37964
rect 40911 37955 40969 37961
rect 41414 37952 41420 37964
rect 41472 37952 41478 38004
rect 41690 37992 41696 38004
rect 41651 37964 41696 37992
rect 41690 37952 41696 37964
rect 41748 37952 41754 38004
rect 41708 37856 41736 37952
rect 41782 37884 41788 37936
rect 41840 37924 41846 37936
rect 41840 37896 42196 37924
rect 41840 37884 41846 37896
rect 42168 37865 42196 37896
rect 41877 37859 41935 37865
rect 41877 37856 41889 37859
rect 41708 37828 41889 37856
rect 41877 37825 41889 37828
rect 41923 37825 41935 37859
rect 41877 37819 41935 37825
rect 42153 37859 42211 37865
rect 42153 37825 42165 37859
rect 42199 37825 42211 37859
rect 42153 37819 42211 37825
rect 39030 37760 39206 37788
rect 39030 37757 39042 37760
rect 38984 37751 39042 37757
rect 37507 37723 37565 37729
rect 37507 37689 37519 37723
rect 37553 37689 37565 37723
rect 38396 37720 38424 37751
rect 40402 37748 40408 37800
rect 40460 37788 40466 37800
rect 40808 37791 40866 37797
rect 40808 37788 40820 37791
rect 40460 37760 40820 37788
rect 40460 37748 40466 37760
rect 40808 37757 40820 37760
rect 40854 37788 40866 37791
rect 41233 37791 41291 37797
rect 41233 37788 41245 37791
rect 40854 37760 41245 37788
rect 40854 37757 40866 37760
rect 40808 37751 40866 37757
rect 41233 37757 41245 37760
rect 41279 37757 41291 37791
rect 41233 37751 41291 37757
rect 43416 37791 43474 37797
rect 43416 37757 43428 37791
rect 43462 37788 43474 37791
rect 43622 37788 43628 37800
rect 43462 37760 43628 37788
rect 43462 37757 43474 37760
rect 43416 37751 43474 37757
rect 43622 37748 43628 37760
rect 43680 37788 43686 37800
rect 44177 37791 44235 37797
rect 44177 37788 44189 37791
rect 43680 37760 44189 37788
rect 43680 37748 43686 37760
rect 44177 37757 44189 37760
rect 44223 37757 44235 37791
rect 44177 37751 44235 37757
rect 39114 37720 39120 37732
rect 38396 37692 39120 37720
rect 37507 37683 37565 37689
rect 39114 37680 39120 37692
rect 39172 37720 39178 37732
rect 39485 37723 39543 37729
rect 39485 37720 39497 37723
rect 39172 37692 39497 37720
rect 39172 37680 39178 37692
rect 39485 37689 39497 37692
rect 39531 37689 39543 37723
rect 39485 37683 39543 37689
rect 41874 37680 41880 37732
rect 41932 37720 41938 37732
rect 41969 37723 42027 37729
rect 41969 37720 41981 37723
rect 41932 37692 41981 37720
rect 41932 37680 41938 37692
rect 41969 37689 41981 37692
rect 42015 37689 42027 37723
rect 41969 37683 42027 37689
rect 36078 37652 36084 37664
rect 34664 37624 35112 37652
rect 36039 37624 36084 37652
rect 34664 37612 34670 37624
rect 36078 37612 36084 37624
rect 36136 37612 36142 37664
rect 42426 37612 42432 37664
rect 42484 37652 42490 37664
rect 43487 37655 43545 37661
rect 43487 37652 43499 37655
rect 42484 37624 43499 37652
rect 42484 37612 42490 37624
rect 43487 37621 43499 37624
rect 43533 37621 43545 37655
rect 43806 37652 43812 37664
rect 43767 37624 43812 37652
rect 43487 37615 43545 37621
rect 43806 37612 43812 37624
rect 43864 37612 43870 37664
rect 1104 37562 48852 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 48852 37562
rect 1104 37488 48852 37510
rect 9214 37448 9220 37460
rect 9175 37420 9220 37448
rect 9214 37408 9220 37420
rect 9272 37408 9278 37460
rect 10870 37448 10876 37460
rect 10831 37420 10876 37448
rect 10870 37408 10876 37420
rect 10928 37408 10934 37460
rect 13630 37408 13636 37460
rect 13688 37448 13694 37460
rect 13817 37451 13875 37457
rect 13817 37448 13829 37451
rect 13688 37420 13829 37448
rect 13688 37408 13694 37420
rect 13817 37417 13829 37420
rect 13863 37417 13875 37451
rect 13817 37411 13875 37417
rect 15378 37408 15384 37460
rect 15436 37448 15442 37460
rect 15473 37451 15531 37457
rect 15473 37448 15485 37451
rect 15436 37420 15485 37448
rect 15436 37408 15442 37420
rect 15473 37417 15485 37420
rect 15519 37417 15531 37451
rect 15473 37411 15531 37417
rect 19334 37408 19340 37460
rect 19392 37448 19398 37460
rect 19889 37451 19947 37457
rect 19889 37448 19901 37451
rect 19392 37420 19901 37448
rect 19392 37408 19398 37420
rect 19889 37417 19901 37420
rect 19935 37417 19947 37451
rect 19889 37411 19947 37417
rect 21726 37408 21732 37460
rect 21784 37448 21790 37460
rect 23155 37451 23213 37457
rect 23155 37448 23167 37451
rect 21784 37420 23167 37448
rect 21784 37408 21790 37420
rect 23155 37417 23167 37420
rect 23201 37417 23213 37451
rect 23155 37411 23213 37417
rect 23474 37408 23480 37460
rect 23532 37448 23538 37460
rect 25041 37451 25099 37457
rect 25041 37448 25053 37451
rect 23532 37420 25053 37448
rect 23532 37408 23538 37420
rect 25041 37417 25053 37420
rect 25087 37448 25099 37451
rect 25958 37448 25964 37460
rect 25087 37420 25964 37448
rect 25087 37417 25099 37420
rect 25041 37411 25099 37417
rect 25958 37408 25964 37420
rect 26016 37408 26022 37460
rect 26510 37408 26516 37460
rect 26568 37448 26574 37460
rect 26881 37451 26939 37457
rect 26881 37448 26893 37451
rect 26568 37420 26893 37448
rect 26568 37408 26574 37420
rect 26881 37417 26893 37420
rect 26927 37417 26939 37451
rect 26881 37411 26939 37417
rect 33781 37451 33839 37457
rect 33781 37417 33793 37451
rect 33827 37448 33839 37451
rect 34606 37448 34612 37460
rect 33827 37420 34612 37448
rect 33827 37417 33839 37420
rect 33781 37411 33839 37417
rect 34606 37408 34612 37420
rect 34664 37408 34670 37460
rect 37918 37448 37924 37460
rect 37879 37420 37924 37448
rect 37918 37408 37924 37420
rect 37976 37408 37982 37460
rect 39577 37451 39635 37457
rect 39577 37417 39589 37451
rect 39623 37448 39635 37451
rect 39942 37448 39948 37460
rect 39623 37420 39948 37448
rect 39623 37417 39635 37420
rect 39577 37411 39635 37417
rect 39942 37408 39948 37420
rect 40000 37448 40006 37460
rect 40497 37451 40555 37457
rect 40497 37448 40509 37451
rect 40000 37420 40509 37448
rect 40000 37408 40006 37420
rect 40497 37417 40509 37420
rect 40543 37448 40555 37451
rect 40678 37448 40684 37460
rect 40543 37420 40684 37448
rect 40543 37417 40555 37420
rect 40497 37411 40555 37417
rect 40678 37408 40684 37420
rect 40736 37408 40742 37460
rect 41598 37408 41604 37460
rect 41656 37448 41662 37460
rect 41693 37451 41751 37457
rect 41693 37448 41705 37451
rect 41656 37420 41705 37448
rect 41656 37408 41662 37420
rect 41693 37417 41705 37420
rect 41739 37417 41751 37451
rect 41693 37411 41751 37417
rect 41874 37408 41880 37460
rect 41932 37448 41938 37460
rect 41969 37451 42027 37457
rect 41969 37448 41981 37451
rect 41932 37420 41981 37448
rect 41932 37408 41938 37420
rect 41969 37417 41981 37420
rect 42015 37417 42027 37451
rect 42426 37448 42432 37460
rect 42387 37420 42432 37448
rect 41969 37411 42027 37417
rect 42426 37408 42432 37420
rect 42484 37408 42490 37460
rect 7009 37383 7067 37389
rect 7009 37349 7021 37383
rect 7055 37380 7067 37383
rect 7098 37380 7104 37392
rect 7055 37352 7104 37380
rect 7055 37349 7067 37352
rect 7009 37343 7067 37349
rect 7098 37340 7104 37352
rect 7156 37340 7162 37392
rect 9861 37383 9919 37389
rect 9861 37349 9873 37383
rect 9907 37380 9919 37383
rect 10226 37380 10232 37392
rect 9907 37352 10232 37380
rect 9907 37349 9919 37352
rect 9861 37343 9919 37349
rect 10226 37340 10232 37352
rect 10284 37340 10290 37392
rect 11422 37380 11428 37392
rect 11383 37352 11428 37380
rect 11422 37340 11428 37352
rect 11480 37340 11486 37392
rect 12986 37380 12992 37392
rect 12947 37352 12992 37380
rect 12986 37340 12992 37352
rect 13044 37340 13050 37392
rect 18414 37340 18420 37392
rect 18472 37380 18478 37392
rect 19061 37383 19119 37389
rect 19061 37380 19073 37383
rect 18472 37352 19073 37380
rect 18472 37340 18478 37352
rect 19061 37349 19073 37352
rect 19107 37349 19119 37383
rect 19061 37343 19119 37349
rect 21361 37383 21419 37389
rect 21361 37349 21373 37383
rect 21407 37380 21419 37383
rect 21542 37380 21548 37392
rect 21407 37352 21548 37380
rect 21407 37349 21419 37352
rect 21361 37343 21419 37349
rect 21542 37340 21548 37352
rect 21600 37340 21606 37392
rect 21637 37383 21695 37389
rect 21637 37349 21649 37383
rect 21683 37380 21695 37383
rect 21818 37380 21824 37392
rect 21683 37352 21824 37380
rect 21683 37349 21695 37352
rect 21637 37343 21695 37349
rect 21818 37340 21824 37352
rect 21876 37340 21882 37392
rect 22833 37383 22891 37389
rect 22833 37349 22845 37383
rect 22879 37380 22891 37383
rect 22922 37380 22928 37392
rect 22879 37352 22928 37380
rect 22879 37349 22891 37352
rect 22833 37343 22891 37349
rect 22922 37340 22928 37352
rect 22980 37340 22986 37392
rect 23842 37340 23848 37392
rect 23900 37380 23906 37392
rect 24442 37383 24500 37389
rect 24442 37380 24454 37383
rect 23900 37352 24454 37380
rect 23900 37340 23906 37352
rect 24442 37349 24454 37352
rect 24488 37349 24500 37383
rect 30190 37380 30196 37392
rect 24442 37343 24500 37349
rect 27080 37352 29500 37380
rect 30151 37352 30196 37380
rect 16298 37312 16304 37324
rect 16259 37284 16304 37312
rect 16298 37272 16304 37284
rect 16356 37272 16362 37324
rect 17862 37312 17868 37324
rect 17826 37284 17868 37312
rect 17862 37272 17868 37284
rect 17920 37321 17926 37324
rect 17920 37315 17974 37321
rect 17920 37281 17928 37315
rect 17962 37312 17974 37315
rect 18506 37312 18512 37324
rect 17962 37284 18512 37312
rect 17962 37281 17974 37284
rect 17920 37275 17974 37281
rect 17920 37272 17926 37275
rect 18506 37272 18512 37284
rect 18564 37272 18570 37324
rect 22646 37272 22652 37324
rect 22704 37312 22710 37324
rect 23052 37315 23110 37321
rect 23052 37312 23064 37315
rect 22704 37284 23064 37312
rect 22704 37272 22710 37284
rect 23052 37281 23064 37284
rect 23098 37281 23110 37315
rect 23052 37275 23110 37281
rect 26602 37272 26608 37324
rect 26660 37312 26666 37324
rect 27080 37321 27108 37352
rect 29472 37324 29500 37352
rect 30190 37340 30196 37352
rect 30248 37340 30254 37392
rect 32306 37340 32312 37392
rect 32364 37380 32370 37392
rect 33226 37389 33232 37392
rect 33223 37380 33232 37389
rect 32364 37352 33232 37380
rect 32364 37340 32370 37352
rect 33223 37343 33232 37352
rect 33226 37340 33232 37343
rect 33284 37340 33290 37392
rect 39019 37383 39077 37389
rect 39019 37349 39031 37383
rect 39065 37380 39077 37383
rect 39114 37380 39120 37392
rect 39065 37352 39120 37380
rect 39065 37349 39077 37352
rect 39019 37343 39077 37349
rect 39114 37340 39120 37352
rect 39172 37380 39178 37392
rect 41094 37383 41152 37389
rect 41094 37380 41106 37383
rect 39172 37352 41106 37380
rect 39172 37340 39178 37352
rect 41094 37349 41106 37352
rect 41140 37380 41152 37383
rect 41506 37380 41512 37392
rect 41140 37352 41512 37380
rect 41140 37349 41152 37352
rect 41094 37343 41152 37349
rect 41506 37340 41512 37352
rect 41564 37340 41570 37392
rect 27065 37315 27123 37321
rect 27065 37312 27077 37315
rect 26660 37284 27077 37312
rect 26660 37272 26666 37284
rect 27065 37281 27077 37284
rect 27111 37281 27123 37315
rect 27065 37275 27123 37281
rect 27341 37315 27399 37321
rect 27341 37281 27353 37315
rect 27387 37312 27399 37315
rect 27982 37312 27988 37324
rect 27387 37284 27988 37312
rect 27387 37281 27399 37284
rect 27341 37275 27399 37281
rect 27982 37272 27988 37284
rect 28040 37272 28046 37324
rect 28350 37312 28356 37324
rect 28311 37284 28356 37312
rect 28350 37272 28356 37284
rect 28408 37272 28414 37324
rect 29454 37312 29460 37324
rect 29415 37284 29460 37312
rect 29454 37272 29460 37284
rect 29512 37272 29518 37324
rect 29914 37312 29920 37324
rect 29875 37284 29920 37312
rect 29914 37272 29920 37284
rect 29972 37272 29978 37324
rect 31110 37321 31116 37324
rect 31088 37315 31116 37321
rect 31088 37312 31100 37315
rect 31023 37284 31100 37312
rect 31088 37281 31100 37284
rect 31168 37312 31174 37324
rect 35713 37315 35771 37321
rect 31168 37284 33134 37312
rect 31088 37275 31116 37281
rect 31110 37272 31116 37275
rect 31168 37272 31174 37284
rect 6914 37244 6920 37256
rect 6875 37216 6920 37244
rect 6914 37204 6920 37216
rect 6972 37204 6978 37256
rect 7190 37244 7196 37256
rect 7151 37216 7196 37244
rect 7190 37204 7196 37216
rect 7248 37204 7254 37256
rect 8938 37204 8944 37256
rect 8996 37244 9002 37256
rect 9769 37247 9827 37253
rect 9769 37244 9781 37247
rect 8996 37216 9781 37244
rect 8996 37204 9002 37216
rect 9769 37213 9781 37216
rect 9815 37213 9827 37247
rect 11330 37244 11336 37256
rect 11291 37216 11336 37244
rect 9769 37207 9827 37213
rect 11330 37204 11336 37216
rect 11388 37204 11394 37256
rect 11609 37247 11667 37253
rect 11609 37244 11621 37247
rect 11440 37216 11621 37244
rect 7650 37136 7656 37188
rect 7708 37176 7714 37188
rect 10321 37179 10379 37185
rect 10321 37176 10333 37179
rect 7708 37148 10333 37176
rect 7708 37136 7714 37148
rect 10321 37145 10333 37148
rect 10367 37176 10379 37179
rect 11440 37176 11468 37216
rect 11609 37213 11621 37216
rect 11655 37213 11667 37247
rect 12894 37244 12900 37256
rect 12855 37216 12900 37244
rect 11609 37207 11667 37213
rect 12894 37204 12900 37216
rect 12952 37204 12958 37256
rect 13170 37244 13176 37256
rect 13131 37216 13176 37244
rect 13170 37204 13176 37216
rect 13228 37244 13234 37256
rect 14185 37247 14243 37253
rect 14185 37244 14197 37247
rect 13228 37216 14197 37244
rect 13228 37204 13234 37216
rect 14185 37213 14197 37216
rect 14231 37213 14243 37247
rect 15746 37244 15752 37256
rect 15707 37216 15752 37244
rect 14185 37207 14243 37213
rect 15746 37204 15752 37216
rect 15804 37204 15810 37256
rect 18003 37247 18061 37253
rect 18003 37213 18015 37247
rect 18049 37244 18061 37247
rect 18966 37244 18972 37256
rect 18049 37216 18972 37244
rect 18049 37213 18061 37216
rect 18003 37207 18061 37213
rect 18966 37204 18972 37216
rect 19024 37204 19030 37256
rect 19334 37244 19340 37256
rect 19295 37216 19340 37244
rect 19334 37204 19340 37216
rect 19392 37244 19398 37256
rect 20162 37244 20168 37256
rect 19392 37216 20168 37244
rect 19392 37204 19398 37216
rect 20162 37204 20168 37216
rect 20220 37244 20226 37256
rect 21821 37247 21879 37253
rect 21821 37244 21833 37247
rect 20220 37216 21833 37244
rect 20220 37204 20226 37216
rect 21821 37213 21833 37216
rect 21867 37213 21879 37247
rect 21821 37207 21879 37213
rect 24026 37204 24032 37256
rect 24084 37244 24090 37256
rect 24121 37247 24179 37253
rect 24121 37244 24133 37247
rect 24084 37216 24133 37244
rect 24084 37204 24090 37216
rect 24121 37213 24133 37216
rect 24167 37244 24179 37247
rect 29362 37244 29368 37256
rect 24167 37216 29368 37244
rect 24167 37213 24179 37216
rect 24121 37207 24179 37213
rect 29362 37204 29368 37216
rect 29420 37204 29426 37256
rect 32858 37244 32864 37256
rect 32819 37216 32864 37244
rect 32858 37204 32864 37216
rect 32916 37204 32922 37256
rect 33106 37244 33134 37284
rect 35713 37281 35725 37315
rect 35759 37312 35771 37315
rect 35802 37312 35808 37324
rect 35759 37284 35808 37312
rect 35759 37281 35771 37284
rect 35713 37275 35771 37281
rect 35802 37272 35808 37284
rect 35860 37272 35866 37324
rect 35986 37312 35992 37324
rect 35947 37284 35992 37312
rect 35986 37272 35992 37284
rect 36044 37272 36050 37324
rect 43257 37315 43315 37321
rect 43257 37281 43269 37315
rect 43303 37312 43315 37315
rect 43346 37312 43352 37324
rect 43303 37284 43352 37312
rect 43303 37281 43315 37284
rect 43257 37275 43315 37281
rect 43346 37272 43352 37284
rect 43404 37272 43410 37324
rect 35434 37244 35440 37256
rect 33106 37216 35440 37244
rect 35434 37204 35440 37216
rect 35492 37244 35498 37256
rect 35894 37244 35900 37256
rect 35492 37216 35900 37244
rect 35492 37204 35498 37216
rect 35894 37204 35900 37216
rect 35952 37204 35958 37256
rect 36170 37244 36176 37256
rect 36131 37216 36176 37244
rect 36170 37204 36176 37216
rect 36228 37204 36234 37256
rect 38654 37244 38660 37256
rect 38615 37216 38660 37244
rect 38654 37204 38660 37216
rect 38712 37204 38718 37256
rect 40770 37244 40776 37256
rect 40731 37216 40776 37244
rect 40770 37204 40776 37216
rect 40828 37204 40834 37256
rect 10367 37148 11468 37176
rect 10367 37145 10379 37148
rect 10321 37139 10379 37145
rect 40586 37136 40592 37188
rect 40644 37176 40650 37188
rect 43487 37179 43545 37185
rect 43487 37176 43499 37179
rect 40644 37148 43499 37176
rect 40644 37136 40650 37148
rect 43487 37145 43499 37148
rect 43533 37145 43545 37179
rect 43487 37139 43545 37145
rect 18414 37108 18420 37120
rect 18375 37080 18420 37108
rect 18414 37068 18420 37080
rect 18472 37068 18478 37120
rect 25222 37068 25228 37120
rect 25280 37108 25286 37120
rect 28537 37111 28595 37117
rect 28537 37108 28549 37111
rect 25280 37080 28549 37108
rect 25280 37068 25286 37080
rect 28537 37077 28549 37080
rect 28583 37108 28595 37111
rect 29273 37111 29331 37117
rect 29273 37108 29285 37111
rect 28583 37080 29285 37108
rect 28583 37077 28595 37080
rect 28537 37071 28595 37077
rect 29273 37077 29285 37080
rect 29319 37108 29331 37111
rect 29730 37108 29736 37120
rect 29319 37080 29736 37108
rect 29319 37077 29331 37080
rect 29273 37071 29331 37077
rect 29730 37068 29736 37080
rect 29788 37068 29794 37120
rect 31159 37111 31217 37117
rect 31159 37077 31171 37111
rect 31205 37108 31217 37111
rect 31294 37108 31300 37120
rect 31205 37080 31300 37108
rect 31205 37077 31217 37080
rect 31159 37071 31217 37077
rect 31294 37068 31300 37080
rect 31352 37068 31358 37120
rect 32398 37068 32404 37120
rect 32456 37108 32462 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32456 37080 32505 37108
rect 32456 37068 32462 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 34790 37068 34796 37120
rect 34848 37108 34854 37120
rect 34885 37111 34943 37117
rect 34885 37108 34897 37111
rect 34848 37080 34897 37108
rect 34848 37068 34854 37080
rect 34885 37077 34897 37080
rect 34931 37077 34943 37111
rect 37090 37108 37096 37120
rect 37051 37080 37096 37108
rect 34885 37071 34943 37077
rect 37090 37068 37096 37080
rect 37148 37068 37154 37120
rect 37461 37111 37519 37117
rect 37461 37077 37473 37111
rect 37507 37108 37519 37111
rect 37550 37108 37556 37120
rect 37507 37080 37556 37108
rect 37507 37077 37519 37080
rect 37461 37071 37519 37077
rect 37550 37068 37556 37080
rect 37608 37068 37614 37120
rect 1104 37018 48852 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 48852 37018
rect 1104 36944 48852 36966
rect 5767 36907 5825 36913
rect 5767 36873 5779 36907
rect 5813 36904 5825 36907
rect 6914 36904 6920 36916
rect 5813 36876 6920 36904
rect 5813 36873 5825 36876
rect 5767 36867 5825 36873
rect 6914 36864 6920 36876
rect 6972 36904 6978 36916
rect 8113 36907 8171 36913
rect 8113 36904 8125 36907
rect 6972 36876 8125 36904
rect 6972 36864 6978 36876
rect 8113 36873 8125 36876
rect 8159 36873 8171 36907
rect 8938 36904 8944 36916
rect 8899 36876 8944 36904
rect 8113 36867 8171 36873
rect 8938 36864 8944 36876
rect 8996 36864 9002 36916
rect 9309 36907 9367 36913
rect 9309 36873 9321 36907
rect 9355 36904 9367 36907
rect 9677 36907 9735 36913
rect 9677 36904 9689 36907
rect 9355 36876 9689 36904
rect 9355 36873 9367 36876
rect 9309 36867 9367 36873
rect 9677 36873 9689 36876
rect 9723 36904 9735 36907
rect 10226 36904 10232 36916
rect 9723 36876 10232 36904
rect 9723 36873 9735 36876
rect 9677 36867 9735 36873
rect 10226 36864 10232 36876
rect 10284 36864 10290 36916
rect 11330 36864 11336 36916
rect 11388 36904 11394 36916
rect 11609 36907 11667 36913
rect 11609 36904 11621 36907
rect 11388 36876 11621 36904
rect 11388 36864 11394 36876
rect 11609 36873 11621 36876
rect 11655 36904 11667 36907
rect 11974 36904 11980 36916
rect 11655 36876 11980 36904
rect 11655 36873 11667 36876
rect 11609 36867 11667 36873
rect 11974 36864 11980 36876
rect 12032 36864 12038 36916
rect 12897 36907 12955 36913
rect 12897 36873 12909 36907
rect 12943 36904 12955 36907
rect 12986 36904 12992 36916
rect 12943 36876 12992 36904
rect 12943 36873 12955 36876
rect 12897 36867 12955 36873
rect 12986 36864 12992 36876
rect 13044 36864 13050 36916
rect 13817 36907 13875 36913
rect 13817 36873 13829 36907
rect 13863 36904 13875 36907
rect 13906 36904 13912 36916
rect 13863 36876 13912 36904
rect 13863 36873 13875 36876
rect 13817 36867 13875 36873
rect 13906 36864 13912 36876
rect 13964 36864 13970 36916
rect 16298 36864 16304 36916
rect 16356 36904 16362 36916
rect 16485 36907 16543 36913
rect 16485 36904 16497 36907
rect 16356 36876 16497 36904
rect 16356 36864 16362 36876
rect 16485 36873 16497 36876
rect 16531 36873 16543 36907
rect 17862 36904 17868 36916
rect 17823 36876 17868 36904
rect 16485 36867 16543 36873
rect 17862 36864 17868 36876
rect 17920 36864 17926 36916
rect 21450 36864 21456 36916
rect 21508 36904 21514 36916
rect 27801 36907 27859 36913
rect 21508 36876 27292 36904
rect 21508 36864 21514 36876
rect 22554 36796 22560 36848
rect 22612 36836 22618 36848
rect 26602 36836 26608 36848
rect 22612 36808 23474 36836
rect 26563 36808 26608 36836
rect 22612 36796 22618 36808
rect 7837 36771 7895 36777
rect 7837 36737 7849 36771
rect 7883 36768 7895 36771
rect 8202 36768 8208 36780
rect 7883 36740 8208 36768
rect 7883 36737 7895 36740
rect 7837 36731 7895 36737
rect 8202 36728 8208 36740
rect 8260 36768 8266 36780
rect 9214 36768 9220 36780
rect 8260 36740 9220 36768
rect 8260 36728 8266 36740
rect 9214 36728 9220 36740
rect 9272 36728 9278 36780
rect 10505 36771 10563 36777
rect 10505 36737 10517 36771
rect 10551 36768 10563 36771
rect 10870 36768 10876 36780
rect 10551 36740 10876 36768
rect 10551 36737 10563 36740
rect 10505 36731 10563 36737
rect 10870 36728 10876 36740
rect 10928 36728 10934 36780
rect 13449 36771 13507 36777
rect 13449 36737 13461 36771
rect 13495 36768 13507 36771
rect 14001 36771 14059 36777
rect 14001 36768 14013 36771
rect 13495 36740 14013 36768
rect 13495 36737 13507 36740
rect 13449 36731 13507 36737
rect 14001 36737 14013 36740
rect 14047 36768 14059 36771
rect 14274 36768 14280 36780
rect 14047 36740 14280 36768
rect 14047 36737 14059 36740
rect 14001 36731 14059 36737
rect 14274 36728 14280 36740
rect 14332 36728 14338 36780
rect 14642 36768 14648 36780
rect 14555 36740 14648 36768
rect 14642 36728 14648 36740
rect 14700 36768 14706 36780
rect 15841 36771 15899 36777
rect 15841 36768 15853 36771
rect 14700 36740 15853 36768
rect 14700 36728 14706 36740
rect 15841 36737 15853 36740
rect 15887 36737 15899 36771
rect 15841 36731 15899 36737
rect 17497 36771 17555 36777
rect 17497 36737 17509 36771
rect 17543 36768 17555 36771
rect 18322 36768 18328 36780
rect 17543 36740 18328 36768
rect 17543 36737 17555 36740
rect 17497 36731 17555 36737
rect 18322 36728 18328 36740
rect 18380 36728 18386 36780
rect 21910 36768 21916 36780
rect 21744 36740 21916 36768
rect 5664 36703 5722 36709
rect 5664 36700 5676 36703
rect 5552 36672 5676 36700
rect 5552 36576 5580 36672
rect 5664 36669 5676 36672
rect 5710 36669 5722 36703
rect 5664 36663 5722 36669
rect 21744 36644 21772 36740
rect 21910 36728 21916 36740
rect 21968 36728 21974 36780
rect 22002 36728 22008 36780
rect 22060 36768 22066 36780
rect 22189 36771 22247 36777
rect 22189 36768 22201 36771
rect 22060 36740 22201 36768
rect 22060 36728 22066 36740
rect 22189 36737 22201 36740
rect 22235 36737 22247 36771
rect 22189 36731 22247 36737
rect 22646 36728 22652 36780
rect 22704 36768 22710 36780
rect 23017 36771 23075 36777
rect 23017 36768 23029 36771
rect 22704 36740 23029 36768
rect 22704 36728 22710 36740
rect 23017 36737 23029 36740
rect 23063 36737 23075 36771
rect 23017 36731 23075 36737
rect 23446 36700 23474 36808
rect 26602 36796 26608 36808
rect 26660 36796 26666 36848
rect 23842 36728 23848 36780
rect 23900 36768 23906 36780
rect 24121 36771 24179 36777
rect 24121 36768 24133 36771
rect 23900 36740 24133 36768
rect 23900 36728 23906 36740
rect 24121 36737 24133 36740
rect 24167 36737 24179 36771
rect 25682 36768 25688 36780
rect 25643 36740 25688 36768
rect 24121 36731 24179 36737
rect 25682 36728 25688 36740
rect 25740 36728 25746 36780
rect 27264 36777 27292 36876
rect 27801 36873 27813 36907
rect 27847 36904 27859 36907
rect 27982 36904 27988 36916
rect 27847 36876 27988 36904
rect 27847 36873 27859 36876
rect 27801 36867 27859 36873
rect 27249 36771 27307 36777
rect 27249 36737 27261 36771
rect 27295 36737 27307 36771
rect 27249 36731 27307 36737
rect 23728 36703 23786 36709
rect 23728 36700 23740 36703
rect 23446 36672 23740 36700
rect 23728 36669 23740 36672
rect 23774 36700 23786 36703
rect 25041 36703 25099 36709
rect 23774 36672 24624 36700
rect 23774 36669 23786 36672
rect 23728 36663 23786 36669
rect 7193 36635 7251 36641
rect 7193 36632 7205 36635
rect 6196 36604 7205 36632
rect 6196 36576 6224 36604
rect 7193 36601 7205 36604
rect 7239 36601 7251 36635
rect 7193 36595 7251 36601
rect 7285 36635 7343 36641
rect 7285 36601 7297 36635
rect 7331 36601 7343 36635
rect 9858 36632 9864 36644
rect 9819 36604 9864 36632
rect 7285 36595 7343 36601
rect 5534 36564 5540 36576
rect 5495 36536 5540 36564
rect 5534 36524 5540 36536
rect 5592 36524 5598 36576
rect 6178 36564 6184 36576
rect 6139 36536 6184 36564
rect 6178 36524 6184 36536
rect 6236 36524 6242 36576
rect 6641 36567 6699 36573
rect 6641 36533 6653 36567
rect 6687 36564 6699 36567
rect 7098 36564 7104 36576
rect 6687 36536 7104 36564
rect 6687 36533 6699 36536
rect 6641 36527 6699 36533
rect 7098 36524 7104 36536
rect 7156 36564 7162 36576
rect 7300 36564 7328 36595
rect 9858 36592 9864 36604
rect 9916 36592 9922 36644
rect 9953 36635 10011 36641
rect 9953 36601 9965 36635
rect 9999 36632 10011 36635
rect 10226 36632 10232 36644
rect 9999 36604 10232 36632
rect 9999 36601 10011 36604
rect 9953 36595 10011 36601
rect 10226 36592 10232 36604
rect 10284 36592 10290 36644
rect 13786 36604 13952 36632
rect 7156 36536 7328 36564
rect 11333 36567 11391 36573
rect 7156 36524 7162 36536
rect 11333 36533 11345 36567
rect 11379 36564 11391 36567
rect 11422 36564 11428 36576
rect 11379 36536 11428 36564
rect 11379 36533 11391 36536
rect 11333 36527 11391 36533
rect 11422 36524 11428 36536
rect 11480 36564 11486 36576
rect 13786 36564 13814 36604
rect 11480 36536 13814 36564
rect 13924 36564 13952 36604
rect 13998 36592 14004 36644
rect 14056 36632 14062 36644
rect 14093 36635 14151 36641
rect 14093 36632 14105 36635
rect 14056 36604 14105 36632
rect 14056 36592 14062 36604
rect 14093 36601 14105 36604
rect 14139 36601 14151 36635
rect 15562 36632 15568 36644
rect 15523 36604 15568 36632
rect 14093 36595 14151 36601
rect 15562 36592 15568 36604
rect 15620 36592 15626 36644
rect 15657 36635 15715 36641
rect 15657 36601 15669 36635
rect 15703 36632 15715 36635
rect 15746 36632 15752 36644
rect 15703 36604 15752 36632
rect 15703 36601 15715 36604
rect 15657 36595 15715 36601
rect 15381 36567 15439 36573
rect 15381 36564 15393 36567
rect 13924 36536 15393 36564
rect 11480 36524 11486 36536
rect 15381 36533 15393 36536
rect 15427 36564 15439 36567
rect 15672 36564 15700 36595
rect 15746 36592 15752 36604
rect 15804 36592 15810 36644
rect 18414 36632 18420 36644
rect 18375 36604 18420 36632
rect 18414 36592 18420 36604
rect 18472 36592 18478 36644
rect 18969 36635 19027 36641
rect 18969 36601 18981 36635
rect 19015 36632 19027 36635
rect 19058 36632 19064 36644
rect 19015 36604 19064 36632
rect 19015 36601 19027 36604
rect 18969 36595 19027 36601
rect 19058 36592 19064 36604
rect 19116 36592 19122 36644
rect 19886 36632 19892 36644
rect 19847 36604 19892 36632
rect 19886 36592 19892 36604
rect 19944 36592 19950 36644
rect 19981 36635 20039 36641
rect 19981 36601 19993 36635
rect 20027 36601 20039 36635
rect 19981 36595 20039 36601
rect 20533 36635 20591 36641
rect 20533 36601 20545 36635
rect 20579 36632 20591 36635
rect 21726 36632 21732 36644
rect 20579 36604 21732 36632
rect 20579 36601 20591 36604
rect 20533 36595 20591 36601
rect 15427 36536 15700 36564
rect 18432 36564 18460 36592
rect 19245 36567 19303 36573
rect 19245 36564 19257 36567
rect 18432 36536 19257 36564
rect 15427 36533 15439 36536
rect 15381 36527 15439 36533
rect 19245 36533 19257 36536
rect 19291 36564 19303 36567
rect 19613 36567 19671 36573
rect 19613 36564 19625 36567
rect 19291 36536 19625 36564
rect 19291 36533 19303 36536
rect 19245 36527 19303 36533
rect 19613 36533 19625 36536
rect 19659 36564 19671 36567
rect 19996 36564 20024 36595
rect 21726 36592 21732 36604
rect 21784 36592 21790 36644
rect 21910 36632 21916 36644
rect 21871 36604 21916 36632
rect 21910 36592 21916 36604
rect 21968 36592 21974 36644
rect 22005 36635 22063 36641
rect 22005 36601 22017 36635
rect 22051 36601 22063 36635
rect 22005 36595 22063 36601
rect 23385 36635 23443 36641
rect 23385 36601 23397 36635
rect 23431 36632 23443 36635
rect 24026 36632 24032 36644
rect 23431 36604 24032 36632
rect 23431 36601 23443 36604
rect 23385 36595 23443 36601
rect 19659 36536 20024 36564
rect 21177 36567 21235 36573
rect 19659 36533 19671 36536
rect 19613 36527 19671 36533
rect 21177 36533 21189 36567
rect 21223 36564 21235 36567
rect 21358 36564 21364 36576
rect 21223 36536 21364 36564
rect 21223 36533 21235 36536
rect 21177 36527 21235 36533
rect 21358 36524 21364 36536
rect 21416 36564 21422 36576
rect 21453 36567 21511 36573
rect 21453 36564 21465 36567
rect 21416 36536 21465 36564
rect 21416 36524 21422 36536
rect 21453 36533 21465 36536
rect 21499 36564 21511 36567
rect 21818 36564 21824 36576
rect 21499 36536 21824 36564
rect 21499 36533 21511 36536
rect 21453 36527 21511 36533
rect 21818 36524 21824 36536
rect 21876 36564 21882 36576
rect 22020 36564 22048 36595
rect 24026 36592 24032 36604
rect 24084 36592 24090 36644
rect 21876 36536 22048 36564
rect 21876 36524 21882 36536
rect 23566 36524 23572 36576
rect 23624 36564 23630 36576
rect 24596 36573 24624 36672
rect 25041 36669 25053 36703
rect 25087 36700 25099 36703
rect 25133 36703 25191 36709
rect 25133 36700 25145 36703
rect 25087 36672 25145 36700
rect 25087 36669 25099 36672
rect 25041 36663 25099 36669
rect 25133 36669 25145 36672
rect 25179 36669 25191 36703
rect 25133 36663 25191 36669
rect 25148 36632 25176 36663
rect 25222 36660 25228 36712
rect 25280 36700 25286 36712
rect 25593 36703 25651 36709
rect 25593 36700 25605 36703
rect 25280 36672 25605 36700
rect 25280 36660 25286 36672
rect 25593 36669 25605 36672
rect 25639 36669 25651 36703
rect 25593 36663 25651 36669
rect 26237 36703 26295 36709
rect 26237 36669 26249 36703
rect 26283 36700 26295 36703
rect 26786 36700 26792 36712
rect 26283 36672 26792 36700
rect 26283 36669 26295 36672
rect 26237 36663 26295 36669
rect 26786 36660 26792 36672
rect 26844 36660 26850 36712
rect 27157 36703 27215 36709
rect 27157 36669 27169 36703
rect 27203 36700 27215 36703
rect 27614 36700 27620 36712
rect 27203 36672 27620 36700
rect 27203 36669 27215 36672
rect 27157 36663 27215 36669
rect 27614 36660 27620 36672
rect 27672 36700 27678 36712
rect 27816 36700 27844 36867
rect 27982 36864 27988 36876
rect 28040 36864 28046 36916
rect 29638 36864 29644 36916
rect 29696 36904 29702 36916
rect 31110 36904 31116 36916
rect 29696 36876 31116 36904
rect 29696 36864 29702 36876
rect 31110 36864 31116 36876
rect 31168 36864 31174 36916
rect 32306 36864 32312 36916
rect 32364 36904 32370 36916
rect 32861 36907 32919 36913
rect 32861 36904 32873 36907
rect 32364 36876 32873 36904
rect 32364 36864 32370 36876
rect 32861 36873 32873 36876
rect 32907 36873 32919 36907
rect 33778 36904 33784 36916
rect 33739 36876 33784 36904
rect 32861 36867 32919 36873
rect 33778 36864 33784 36876
rect 33836 36864 33842 36916
rect 34701 36907 34759 36913
rect 34701 36873 34713 36907
rect 34747 36904 34759 36907
rect 35802 36904 35808 36916
rect 34747 36876 35808 36904
rect 34747 36873 34759 36876
rect 34701 36867 34759 36873
rect 35802 36864 35808 36876
rect 35860 36864 35866 36916
rect 36170 36864 36176 36916
rect 36228 36904 36234 36916
rect 40221 36907 40279 36913
rect 40221 36904 40233 36907
rect 36228 36876 40233 36904
rect 36228 36864 36234 36876
rect 40221 36873 40233 36876
rect 40267 36904 40279 36907
rect 40770 36904 40776 36916
rect 40267 36876 40776 36904
rect 40267 36873 40279 36876
rect 40221 36867 40279 36873
rect 40770 36864 40776 36876
rect 40828 36864 40834 36916
rect 41506 36904 41512 36916
rect 41467 36876 41512 36904
rect 41506 36864 41512 36876
rect 41564 36864 41570 36916
rect 41598 36864 41604 36916
rect 41656 36904 41662 36916
rect 41877 36907 41935 36913
rect 41877 36904 41889 36907
rect 41656 36876 41889 36904
rect 41656 36864 41662 36876
rect 41877 36873 41889 36876
rect 41923 36873 41935 36907
rect 41877 36867 41935 36873
rect 38473 36839 38531 36845
rect 38473 36836 38485 36839
rect 31496 36808 35480 36836
rect 31496 36777 31524 36808
rect 31481 36771 31539 36777
rect 31481 36768 31493 36771
rect 27672 36672 27844 36700
rect 28552 36740 31493 36768
rect 27672 36660 27678 36672
rect 28552 36644 28580 36740
rect 31481 36737 31493 36740
rect 31527 36737 31539 36771
rect 32398 36768 32404 36780
rect 32359 36740 32404 36768
rect 31481 36731 31539 36737
rect 29549 36703 29607 36709
rect 29549 36669 29561 36703
rect 29595 36669 29607 36703
rect 29730 36700 29736 36712
rect 29691 36672 29736 36700
rect 29549 36663 29607 36669
rect 28534 36632 28540 36644
rect 25148 36604 28540 36632
rect 28534 36592 28540 36604
rect 28592 36592 28598 36644
rect 28902 36592 28908 36644
rect 28960 36632 28966 36644
rect 29089 36635 29147 36641
rect 29089 36632 29101 36635
rect 28960 36604 29101 36632
rect 28960 36592 28966 36604
rect 29089 36601 29101 36604
rect 29135 36632 29147 36635
rect 29564 36632 29592 36663
rect 29730 36660 29736 36672
rect 29788 36660 29794 36712
rect 31496 36700 31524 36731
rect 32398 36728 32404 36740
rect 32456 36728 32462 36780
rect 31665 36703 31723 36709
rect 31665 36700 31677 36703
rect 31496 36672 31677 36700
rect 31665 36669 31677 36672
rect 31711 36669 31723 36703
rect 32122 36700 32128 36712
rect 32083 36672 32128 36700
rect 31665 36663 31723 36669
rect 32122 36660 32128 36672
rect 32180 36660 32186 36712
rect 32950 36660 32956 36712
rect 33008 36700 33014 36712
rect 33280 36703 33338 36709
rect 33280 36700 33292 36703
rect 33008 36672 33292 36700
rect 33008 36660 33014 36672
rect 33280 36669 33292 36672
rect 33326 36700 33338 36703
rect 33778 36700 33784 36712
rect 33326 36672 33784 36700
rect 33326 36669 33338 36672
rect 33280 36663 33338 36669
rect 33778 36660 33784 36672
rect 33836 36660 33842 36712
rect 35452 36709 35480 36808
rect 37153 36808 38485 36836
rect 36173 36771 36231 36777
rect 36173 36737 36185 36771
rect 36219 36768 36231 36771
rect 37153 36768 37181 36808
rect 38473 36805 38485 36808
rect 38519 36836 38531 36839
rect 38654 36836 38660 36848
rect 38519 36808 38660 36836
rect 38519 36805 38531 36808
rect 38473 36799 38531 36805
rect 38654 36796 38660 36808
rect 38712 36796 38718 36848
rect 38746 36796 38752 36848
rect 38804 36836 38810 36848
rect 41782 36836 41788 36848
rect 38804 36808 41788 36836
rect 38804 36796 38810 36808
rect 37550 36768 37556 36780
rect 36219 36740 37181 36768
rect 37511 36740 37556 36768
rect 36219 36737 36231 36740
rect 36173 36731 36231 36737
rect 37550 36728 37556 36740
rect 37608 36728 37614 36780
rect 39114 36768 39120 36780
rect 39075 36740 39120 36768
rect 39114 36728 39120 36740
rect 39172 36728 39178 36780
rect 39945 36771 40003 36777
rect 39945 36737 39957 36771
rect 39991 36768 40003 36771
rect 40586 36768 40592 36780
rect 39991 36740 40592 36768
rect 39991 36737 40003 36740
rect 39945 36731 40003 36737
rect 40586 36728 40592 36740
rect 40644 36728 40650 36780
rect 40880 36777 40908 36808
rect 41782 36796 41788 36808
rect 41840 36796 41846 36848
rect 40865 36771 40923 36777
rect 40865 36737 40877 36771
rect 40911 36737 40923 36771
rect 40865 36731 40923 36737
rect 35437 36703 35495 36709
rect 35437 36669 35449 36703
rect 35483 36669 35495 36703
rect 35986 36700 35992 36712
rect 35899 36672 35992 36700
rect 35437 36663 35495 36669
rect 32398 36632 32404 36644
rect 29135 36604 32404 36632
rect 29135 36601 29147 36604
rect 29089 36595 29147 36601
rect 32398 36592 32404 36604
rect 32456 36592 32462 36644
rect 32674 36592 32680 36644
rect 32732 36632 32738 36644
rect 33367 36635 33425 36641
rect 33367 36632 33379 36635
rect 32732 36604 33379 36632
rect 32732 36592 32738 36604
rect 33367 36601 33379 36604
rect 33413 36601 33425 36635
rect 33367 36595 33425 36601
rect 35452 36576 35480 36663
rect 35986 36660 35992 36672
rect 36044 36700 36050 36712
rect 37001 36703 37059 36709
rect 37001 36700 37013 36703
rect 36044 36672 36584 36700
rect 36044 36660 36050 36672
rect 23799 36567 23857 36573
rect 23799 36564 23811 36567
rect 23624 36536 23811 36564
rect 23624 36524 23630 36536
rect 23799 36533 23811 36536
rect 23845 36533 23857 36567
rect 23799 36527 23857 36533
rect 24581 36567 24639 36573
rect 24581 36533 24593 36567
rect 24627 36564 24639 36567
rect 24670 36564 24676 36576
rect 24627 36536 24676 36564
rect 24627 36533 24639 36536
rect 24581 36527 24639 36533
rect 24670 36524 24676 36536
rect 24728 36524 24734 36576
rect 27890 36524 27896 36576
rect 27948 36564 27954 36576
rect 28350 36564 28356 36576
rect 27948 36536 28356 36564
rect 27948 36524 27954 36536
rect 28350 36524 28356 36536
rect 28408 36524 28414 36576
rect 29362 36564 29368 36576
rect 29323 36536 29368 36564
rect 29362 36524 29368 36536
rect 29420 36524 29426 36576
rect 29454 36524 29460 36576
rect 29512 36564 29518 36576
rect 30285 36567 30343 36573
rect 30285 36564 30297 36567
rect 29512 36536 30297 36564
rect 29512 36524 29518 36536
rect 30285 36533 30297 36536
rect 30331 36533 30343 36567
rect 30285 36527 30343 36533
rect 35345 36567 35403 36573
rect 35345 36533 35357 36567
rect 35391 36564 35403 36567
rect 35434 36564 35440 36576
rect 35391 36536 35440 36564
rect 35391 36533 35403 36536
rect 35345 36527 35403 36533
rect 35434 36524 35440 36536
rect 35492 36524 35498 36576
rect 36556 36573 36584 36672
rect 36832 36672 37013 36700
rect 36541 36567 36599 36573
rect 36541 36533 36553 36567
rect 36587 36564 36599 36567
rect 36630 36564 36636 36576
rect 36587 36536 36636 36564
rect 36587 36533 36599 36536
rect 36541 36527 36599 36533
rect 36630 36524 36636 36536
rect 36688 36524 36694 36576
rect 36722 36524 36728 36576
rect 36780 36564 36786 36576
rect 36832 36573 36860 36672
rect 37001 36669 37013 36672
rect 37047 36669 37059 36703
rect 37001 36663 37059 36669
rect 37090 36660 37096 36712
rect 37148 36700 37154 36712
rect 37461 36703 37519 36709
rect 37461 36700 37473 36703
rect 37148 36672 37473 36700
rect 37148 36660 37154 36672
rect 37461 36669 37473 36672
rect 37507 36700 37519 36703
rect 37918 36700 37924 36712
rect 37507 36672 37924 36700
rect 37507 36669 37519 36672
rect 37461 36663 37519 36669
rect 37918 36660 37924 36672
rect 37976 36660 37982 36712
rect 38286 36660 38292 36712
rect 38344 36700 38350 36712
rect 38724 36703 38782 36709
rect 38724 36700 38736 36703
rect 38344 36672 38736 36700
rect 38344 36660 38350 36672
rect 38724 36669 38736 36672
rect 38770 36700 38782 36703
rect 38770 36672 39620 36700
rect 38770 36669 38782 36672
rect 38724 36663 38782 36669
rect 39592 36576 39620 36672
rect 40678 36632 40684 36644
rect 40639 36604 40684 36632
rect 40678 36592 40684 36604
rect 40736 36592 40742 36644
rect 41892 36632 41920 36867
rect 41966 36796 41972 36848
rect 42024 36836 42030 36848
rect 42024 36808 42472 36836
rect 42024 36796 42030 36808
rect 42153 36771 42211 36777
rect 42153 36737 42165 36771
rect 42199 36768 42211 36771
rect 42334 36768 42340 36780
rect 42199 36740 42340 36768
rect 42199 36737 42211 36740
rect 42153 36731 42211 36737
rect 42334 36728 42340 36740
rect 42392 36728 42398 36780
rect 42444 36777 42472 36808
rect 42429 36771 42487 36777
rect 42429 36737 42441 36771
rect 42475 36737 42487 36771
rect 42429 36731 42487 36737
rect 42245 36635 42303 36641
rect 42245 36632 42257 36635
rect 41892 36604 42257 36632
rect 42245 36601 42257 36604
rect 42291 36601 42303 36635
rect 42245 36595 42303 36601
rect 36817 36567 36875 36573
rect 36817 36564 36829 36567
rect 36780 36536 36829 36564
rect 36780 36524 36786 36536
rect 36817 36533 36829 36536
rect 36863 36533 36875 36567
rect 36817 36527 36875 36533
rect 38795 36567 38853 36573
rect 38795 36533 38807 36567
rect 38841 36564 38853 36567
rect 38930 36564 38936 36576
rect 38841 36536 38936 36564
rect 38841 36533 38853 36536
rect 38795 36527 38853 36533
rect 38930 36524 38936 36536
rect 38988 36524 38994 36576
rect 39574 36564 39580 36576
rect 39535 36536 39580 36564
rect 39574 36524 39580 36536
rect 39632 36524 39638 36576
rect 43346 36564 43352 36576
rect 43307 36536 43352 36564
rect 43346 36524 43352 36536
rect 43404 36524 43410 36576
rect 1104 36474 48852 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 48852 36474
rect 1104 36400 48852 36422
rect 11422 36360 11428 36372
rect 6104 36332 7696 36360
rect 6104 36304 6132 36332
rect 6086 36292 6092 36304
rect 5999 36264 6092 36292
rect 6086 36252 6092 36264
rect 6144 36252 6150 36304
rect 6641 36295 6699 36301
rect 6641 36261 6653 36295
rect 6687 36292 6699 36295
rect 7190 36292 7196 36304
rect 6687 36264 7196 36292
rect 6687 36261 6699 36264
rect 6641 36255 6699 36261
rect 7190 36252 7196 36264
rect 7248 36252 7254 36304
rect 7668 36301 7696 36332
rect 10244 36332 11428 36360
rect 7653 36295 7711 36301
rect 7653 36261 7665 36295
rect 7699 36292 7711 36295
rect 7834 36292 7840 36304
rect 7699 36264 7840 36292
rect 7699 36261 7711 36264
rect 7653 36255 7711 36261
rect 7834 36252 7840 36264
rect 7892 36252 7898 36304
rect 8202 36292 8208 36304
rect 8163 36264 8208 36292
rect 8202 36252 8208 36264
rect 8260 36252 8266 36304
rect 9030 36252 9036 36304
rect 9088 36292 9094 36304
rect 10134 36292 10140 36304
rect 9088 36264 10140 36292
rect 9088 36252 9094 36264
rect 10134 36252 10140 36264
rect 10192 36292 10198 36304
rect 10244 36301 10272 36332
rect 11422 36320 11428 36332
rect 11480 36320 11486 36372
rect 12894 36360 12900 36372
rect 12855 36332 12900 36360
rect 12894 36320 12900 36332
rect 12952 36360 12958 36372
rect 14642 36360 14648 36372
rect 12952 36332 14648 36360
rect 12952 36320 12958 36332
rect 14642 36320 14648 36332
rect 14700 36320 14706 36372
rect 18414 36320 18420 36372
rect 18472 36360 18478 36372
rect 18509 36363 18567 36369
rect 18509 36360 18521 36363
rect 18472 36332 18521 36360
rect 18472 36320 18478 36332
rect 18509 36329 18521 36332
rect 18555 36329 18567 36363
rect 18966 36360 18972 36372
rect 18927 36332 18972 36360
rect 18509 36323 18567 36329
rect 18966 36320 18972 36332
rect 19024 36320 19030 36372
rect 20254 36360 20260 36372
rect 19403 36332 20260 36360
rect 10229 36295 10287 36301
rect 10229 36292 10241 36295
rect 10192 36264 10241 36292
rect 10192 36252 10198 36264
rect 10229 36261 10241 36264
rect 10275 36261 10287 36295
rect 10229 36255 10287 36261
rect 10781 36295 10839 36301
rect 10781 36261 10793 36295
rect 10827 36292 10839 36295
rect 10870 36292 10876 36304
rect 10827 36264 10876 36292
rect 10827 36261 10839 36264
rect 10781 36255 10839 36261
rect 10870 36252 10876 36264
rect 10928 36252 10934 36304
rect 11790 36292 11796 36304
rect 11751 36264 11796 36292
rect 11790 36252 11796 36264
rect 11848 36252 11854 36304
rect 17678 36252 17684 36304
rect 17736 36292 17742 36304
rect 17910 36295 17968 36301
rect 17910 36292 17922 36295
rect 17736 36264 17922 36292
rect 17736 36252 17742 36264
rect 17910 36261 17922 36264
rect 17956 36261 17968 36295
rect 17910 36255 17968 36261
rect 4960 36227 5018 36233
rect 4960 36193 4972 36227
rect 5006 36224 5018 36227
rect 5258 36224 5264 36236
rect 5006 36196 5264 36224
rect 5006 36193 5018 36196
rect 4960 36187 5018 36193
rect 5258 36184 5264 36196
rect 5316 36224 5322 36236
rect 5353 36227 5411 36233
rect 5353 36224 5365 36227
rect 5316 36196 5365 36224
rect 5316 36184 5322 36196
rect 5353 36193 5365 36196
rect 5399 36193 5411 36227
rect 5353 36187 5411 36193
rect 13884 36227 13942 36233
rect 13884 36193 13896 36227
rect 13930 36224 13942 36227
rect 13998 36224 14004 36236
rect 13930 36196 14004 36224
rect 13930 36193 13942 36196
rect 13884 36187 13942 36193
rect 13998 36184 14004 36196
rect 14056 36184 14062 36236
rect 16206 36224 16212 36236
rect 16167 36196 16212 36224
rect 16206 36184 16212 36196
rect 16264 36184 16270 36236
rect 19242 36184 19248 36236
rect 19300 36224 19306 36236
rect 19403 36233 19431 36332
rect 20254 36320 20260 36332
rect 20312 36360 20318 36372
rect 20312 36332 21496 36360
rect 20312 36320 20318 36332
rect 19475 36295 19533 36301
rect 19475 36261 19487 36295
rect 19521 36292 19533 36295
rect 19886 36292 19892 36304
rect 19521 36264 19892 36292
rect 19521 36261 19533 36264
rect 19475 36255 19533 36261
rect 19886 36252 19892 36264
rect 19944 36252 19950 36304
rect 21082 36252 21088 36304
rect 21140 36292 21146 36304
rect 21361 36295 21419 36301
rect 21361 36292 21373 36295
rect 21140 36264 21373 36292
rect 21140 36252 21146 36264
rect 21361 36261 21373 36264
rect 21407 36261 21419 36295
rect 21468 36292 21496 36332
rect 21910 36320 21916 36372
rect 21968 36360 21974 36372
rect 22189 36363 22247 36369
rect 22189 36360 22201 36363
rect 21968 36332 22201 36360
rect 21968 36320 21974 36332
rect 22189 36329 22201 36332
rect 22235 36360 22247 36363
rect 23566 36360 23572 36372
rect 22235 36332 23572 36360
rect 22235 36329 22247 36332
rect 22189 36323 22247 36329
rect 23566 36320 23572 36332
rect 23624 36320 23630 36372
rect 25038 36360 25044 36372
rect 23998 36332 25044 36360
rect 23998 36292 24026 36332
rect 25038 36320 25044 36332
rect 25096 36320 25102 36372
rect 25222 36360 25228 36372
rect 25183 36332 25228 36360
rect 25222 36320 25228 36332
rect 25280 36320 25286 36372
rect 27614 36360 27620 36372
rect 27575 36332 27620 36360
rect 27614 36320 27620 36332
rect 27672 36320 27678 36372
rect 29733 36363 29791 36369
rect 29733 36329 29745 36363
rect 29779 36360 29791 36363
rect 29914 36360 29920 36372
rect 29779 36332 29920 36360
rect 29779 36329 29791 36332
rect 29733 36323 29791 36329
rect 29914 36320 29920 36332
rect 29972 36320 29978 36372
rect 31570 36320 31576 36372
rect 31628 36360 31634 36372
rect 31757 36363 31815 36369
rect 31757 36360 31769 36363
rect 31628 36332 31769 36360
rect 31628 36320 31634 36332
rect 31757 36329 31769 36332
rect 31803 36360 31815 36363
rect 32122 36360 32128 36372
rect 31803 36332 32128 36360
rect 31803 36329 31815 36332
rect 31757 36323 31815 36329
rect 32122 36320 32128 36332
rect 32180 36320 32186 36372
rect 34885 36363 34943 36369
rect 34885 36329 34897 36363
rect 34931 36360 34943 36363
rect 35805 36363 35863 36369
rect 34931 36332 35480 36360
rect 34931 36329 34943 36332
rect 34885 36323 34943 36329
rect 24302 36292 24308 36304
rect 21468 36264 24026 36292
rect 24263 36264 24308 36292
rect 21361 36255 21419 36261
rect 24302 36252 24308 36264
rect 24360 36252 24366 36304
rect 26418 36252 26424 36304
rect 26476 36292 26482 36304
rect 26697 36295 26755 36301
rect 26697 36292 26709 36295
rect 26476 36264 26709 36292
rect 26476 36252 26482 36264
rect 26697 36261 26709 36264
rect 26743 36261 26755 36295
rect 30558 36292 30564 36304
rect 30519 36264 30564 36292
rect 26697 36255 26755 36261
rect 30558 36252 30564 36264
rect 30616 36252 30622 36304
rect 32140 36292 32168 36320
rect 32858 36292 32864 36304
rect 32140 36264 32628 36292
rect 32771 36264 32864 36292
rect 19388 36227 19446 36233
rect 19388 36224 19400 36227
rect 19300 36196 19400 36224
rect 19300 36184 19306 36196
rect 19388 36193 19400 36196
rect 19434 36193 19446 36227
rect 19388 36187 19446 36193
rect 22792 36227 22850 36233
rect 22792 36193 22804 36227
rect 22838 36224 22850 36227
rect 23014 36224 23020 36236
rect 22838 36196 23020 36224
rect 22838 36193 22850 36196
rect 22792 36187 22850 36193
rect 23014 36184 23020 36196
rect 23072 36184 23078 36236
rect 28902 36224 28908 36236
rect 28863 36196 28908 36224
rect 28902 36184 28908 36196
rect 28960 36184 28966 36236
rect 29086 36224 29092 36236
rect 29047 36196 29092 36224
rect 29086 36184 29092 36196
rect 29144 36184 29150 36236
rect 32398 36224 32404 36236
rect 32359 36196 32404 36224
rect 32398 36184 32404 36196
rect 32456 36184 32462 36236
rect 32600 36233 32628 36264
rect 32858 36252 32864 36264
rect 32916 36292 32922 36304
rect 35452 36301 35480 36332
rect 35805 36329 35817 36363
rect 35851 36360 35863 36363
rect 35894 36360 35900 36372
rect 35851 36332 35900 36360
rect 35851 36329 35863 36332
rect 35805 36323 35863 36329
rect 35894 36320 35900 36332
rect 35952 36360 35958 36372
rect 36262 36360 36268 36372
rect 35952 36332 36268 36360
rect 35952 36320 35958 36332
rect 36262 36320 36268 36332
rect 36320 36320 36326 36372
rect 37918 36360 37924 36372
rect 37879 36332 37924 36360
rect 37918 36320 37924 36332
rect 37976 36320 37982 36372
rect 33137 36295 33195 36301
rect 33137 36292 33149 36295
rect 32916 36264 33149 36292
rect 32916 36252 32922 36264
rect 33137 36261 33149 36264
rect 33183 36261 33195 36295
rect 33137 36255 33195 36261
rect 35437 36295 35495 36301
rect 35437 36261 35449 36295
rect 35483 36292 35495 36295
rect 35483 36264 36676 36292
rect 35483 36261 35495 36264
rect 35437 36255 35495 36261
rect 36648 36236 36676 36264
rect 38930 36252 38936 36304
rect 38988 36292 38994 36304
rect 39117 36295 39175 36301
rect 39117 36292 39129 36295
rect 38988 36264 39129 36292
rect 38988 36252 38994 36264
rect 39117 36261 39129 36264
rect 39163 36261 39175 36295
rect 39117 36255 39175 36261
rect 39206 36252 39212 36304
rect 39264 36292 39270 36304
rect 40770 36292 40776 36304
rect 39264 36264 40776 36292
rect 39264 36252 39270 36264
rect 40770 36252 40776 36264
rect 40828 36252 40834 36304
rect 32585 36227 32643 36233
rect 32585 36193 32597 36227
rect 32631 36193 32643 36227
rect 32585 36187 32643 36193
rect 33042 36184 33048 36236
rect 33100 36224 33106 36236
rect 33226 36224 33232 36236
rect 33100 36196 33232 36224
rect 33100 36184 33106 36196
rect 33226 36184 33232 36196
rect 33284 36224 33290 36236
rect 33724 36227 33782 36233
rect 33724 36224 33736 36227
rect 33284 36196 33736 36224
rect 33284 36184 33290 36196
rect 33724 36193 33736 36196
rect 33770 36193 33782 36227
rect 33724 36187 33782 36193
rect 34606 36184 34612 36236
rect 34664 36224 34670 36236
rect 34701 36227 34759 36233
rect 34701 36224 34713 36227
rect 34664 36196 34713 36224
rect 34664 36184 34670 36196
rect 34701 36193 34713 36196
rect 34747 36193 34759 36227
rect 36078 36224 36084 36236
rect 36039 36196 36084 36224
rect 34701 36187 34759 36193
rect 36078 36184 36084 36196
rect 36136 36184 36142 36236
rect 36538 36224 36544 36236
rect 36499 36196 36544 36224
rect 36538 36184 36544 36196
rect 36596 36184 36602 36236
rect 36630 36184 36636 36236
rect 36688 36224 36694 36236
rect 37737 36227 37795 36233
rect 37737 36224 37749 36227
rect 36688 36196 37749 36224
rect 36688 36184 36694 36196
rect 37737 36193 37749 36196
rect 37783 36224 37795 36227
rect 38470 36224 38476 36236
rect 37783 36196 38476 36224
rect 37783 36193 37795 36196
rect 37737 36187 37795 36193
rect 38470 36184 38476 36196
rect 38528 36184 38534 36236
rect 41690 36184 41696 36236
rect 41748 36224 41754 36236
rect 42188 36227 42246 36233
rect 42188 36224 42200 36227
rect 41748 36196 42200 36224
rect 41748 36184 41754 36196
rect 42188 36193 42200 36196
rect 42234 36193 42246 36227
rect 42188 36187 42246 36193
rect 42702 36184 42708 36236
rect 42760 36224 42766 36236
rect 43416 36227 43474 36233
rect 43416 36224 43428 36227
rect 42760 36196 43428 36224
rect 42760 36184 42766 36196
rect 43416 36193 43428 36196
rect 43462 36224 43474 36227
rect 43898 36224 43904 36236
rect 43462 36196 43904 36224
rect 43462 36193 43474 36196
rect 43416 36187 43474 36193
rect 43898 36184 43904 36196
rect 43956 36184 43962 36236
rect 5169 36159 5227 36165
rect 5169 36125 5181 36159
rect 5215 36156 5227 36159
rect 5994 36156 6000 36168
rect 5215 36128 6000 36156
rect 5215 36125 5227 36128
rect 5169 36119 5227 36125
rect 5994 36116 6000 36128
rect 6052 36116 6058 36168
rect 7561 36159 7619 36165
rect 7561 36125 7573 36159
rect 7607 36156 7619 36159
rect 8202 36156 8208 36168
rect 7607 36128 8208 36156
rect 7607 36125 7619 36128
rect 7561 36119 7619 36125
rect 8202 36116 8208 36128
rect 8260 36116 8266 36168
rect 10137 36159 10195 36165
rect 10137 36125 10149 36159
rect 10183 36156 10195 36159
rect 10410 36156 10416 36168
rect 10183 36128 10416 36156
rect 10183 36125 10195 36128
rect 10137 36119 10195 36125
rect 10410 36116 10416 36128
rect 10468 36116 10474 36168
rect 11698 36156 11704 36168
rect 11659 36128 11704 36156
rect 11698 36116 11704 36128
rect 11756 36116 11762 36168
rect 11974 36156 11980 36168
rect 11935 36128 11980 36156
rect 11974 36116 11980 36128
rect 12032 36116 12038 36168
rect 15654 36116 15660 36168
rect 15712 36156 15718 36168
rect 16025 36159 16083 36165
rect 16025 36156 16037 36159
rect 15712 36128 16037 36156
rect 15712 36116 15718 36128
rect 16025 36125 16037 36128
rect 16071 36125 16083 36159
rect 16025 36119 16083 36125
rect 17402 36116 17408 36168
rect 17460 36156 17466 36168
rect 17589 36159 17647 36165
rect 17589 36156 17601 36159
rect 17460 36128 17601 36156
rect 17460 36116 17466 36128
rect 17589 36125 17601 36128
rect 17635 36125 17647 36159
rect 17589 36119 17647 36125
rect 20714 36116 20720 36168
rect 20772 36156 20778 36168
rect 21269 36159 21327 36165
rect 21269 36156 21281 36159
rect 20772 36128 21281 36156
rect 20772 36116 20778 36128
rect 21269 36125 21281 36128
rect 21315 36156 21327 36159
rect 22879 36159 22937 36165
rect 22879 36156 22891 36159
rect 21315 36128 22891 36156
rect 21315 36125 21327 36128
rect 21269 36119 21327 36125
rect 22879 36125 22891 36128
rect 22925 36125 22937 36159
rect 22879 36119 22937 36125
rect 24213 36159 24271 36165
rect 24213 36125 24225 36159
rect 24259 36125 24271 36159
rect 24486 36156 24492 36168
rect 24447 36128 24492 36156
rect 24213 36119 24271 36125
rect 19058 36048 19064 36100
rect 19116 36088 19122 36100
rect 21821 36091 21879 36097
rect 21821 36088 21833 36091
rect 19116 36060 21833 36088
rect 19116 36048 19122 36060
rect 21821 36057 21833 36060
rect 21867 36088 21879 36091
rect 22002 36088 22008 36100
rect 21867 36060 22008 36088
rect 21867 36057 21879 36060
rect 21821 36051 21879 36057
rect 22002 36048 22008 36060
rect 22060 36048 22066 36100
rect 24118 36048 24124 36100
rect 24176 36088 24182 36100
rect 24228 36088 24256 36119
rect 24486 36116 24492 36128
rect 24544 36116 24550 36168
rect 26605 36159 26663 36165
rect 26605 36125 26617 36159
rect 26651 36156 26663 36159
rect 27522 36156 27528 36168
rect 26651 36128 27528 36156
rect 26651 36125 26663 36128
rect 26605 36119 26663 36125
rect 27522 36116 27528 36128
rect 27580 36116 27586 36168
rect 29362 36156 29368 36168
rect 29323 36128 29368 36156
rect 29362 36116 29368 36128
rect 29420 36116 29426 36168
rect 30466 36156 30472 36168
rect 30427 36128 30472 36156
rect 30466 36116 30472 36128
rect 30524 36116 30530 36168
rect 36814 36156 36820 36168
rect 36775 36128 36820 36156
rect 36814 36116 36820 36128
rect 36872 36116 36878 36168
rect 39390 36156 39396 36168
rect 39351 36128 39396 36156
rect 39390 36116 39396 36128
rect 39448 36116 39454 36168
rect 40310 36116 40316 36168
rect 40368 36156 40374 36168
rect 40681 36159 40739 36165
rect 40681 36156 40693 36159
rect 40368 36128 40693 36156
rect 40368 36116 40374 36128
rect 40681 36125 40693 36128
rect 40727 36125 40739 36159
rect 41322 36156 41328 36168
rect 41283 36128 41328 36156
rect 40681 36119 40739 36125
rect 41322 36116 41328 36128
rect 41380 36156 41386 36168
rect 43254 36156 43260 36168
rect 41380 36128 43260 36156
rect 41380 36116 41386 36128
rect 43254 36116 43260 36128
rect 43312 36116 43318 36168
rect 24176 36060 24256 36088
rect 24504 36088 24532 36116
rect 27157 36091 27215 36097
rect 27157 36088 27169 36091
rect 24504 36060 27169 36088
rect 24176 36048 24182 36060
rect 27157 36057 27169 36060
rect 27203 36088 27215 36091
rect 27246 36088 27252 36100
rect 27203 36060 27252 36088
rect 27203 36057 27215 36060
rect 27157 36051 27215 36057
rect 27246 36048 27252 36060
rect 27304 36048 27310 36100
rect 29270 36048 29276 36100
rect 29328 36088 29334 36100
rect 30009 36091 30067 36097
rect 30009 36088 30021 36091
rect 29328 36060 30021 36088
rect 29328 36048 29334 36060
rect 30009 36057 30021 36060
rect 30055 36057 30067 36091
rect 31018 36088 31024 36100
rect 30979 36060 31024 36088
rect 30009 36051 30067 36057
rect 31018 36048 31024 36060
rect 31076 36048 31082 36100
rect 32490 36048 32496 36100
rect 32548 36088 32554 36100
rect 34054 36088 34060 36100
rect 32548 36060 34060 36088
rect 32548 36048 32554 36060
rect 34054 36048 34060 36060
rect 34112 36088 34118 36100
rect 41138 36088 41144 36100
rect 34112 36060 41144 36088
rect 34112 36048 34118 36060
rect 41138 36048 41144 36060
rect 41196 36088 41202 36100
rect 41690 36088 41696 36100
rect 41196 36060 41696 36088
rect 41196 36048 41202 36060
rect 41690 36048 41696 36060
rect 41748 36048 41754 36100
rect 41782 36048 41788 36100
rect 41840 36088 41846 36100
rect 43487 36091 43545 36097
rect 43487 36088 43499 36091
rect 41840 36060 43499 36088
rect 41840 36048 41846 36060
rect 43487 36057 43499 36060
rect 43533 36057 43545 36091
rect 43487 36051 43545 36057
rect 4614 36020 4620 36032
rect 4575 35992 4620 36020
rect 4614 35980 4620 35992
rect 4672 35980 4678 36032
rect 7098 36020 7104 36032
rect 7059 35992 7104 36020
rect 7098 35980 7104 35992
rect 7156 35980 7162 36032
rect 9858 36020 9864 36032
rect 9819 35992 9864 36020
rect 9858 35980 9864 35992
rect 9916 35980 9922 36032
rect 13630 36020 13636 36032
rect 13543 35992 13636 36020
rect 13630 35980 13636 35992
rect 13688 36020 13694 36032
rect 13955 36023 14013 36029
rect 13955 36020 13967 36023
rect 13688 35992 13967 36020
rect 13688 35980 13694 35992
rect 13955 35989 13967 35992
rect 14001 35989 14013 36023
rect 15562 36020 15568 36032
rect 15475 35992 15568 36020
rect 13955 35983 14013 35989
rect 15562 35980 15568 35992
rect 15620 36020 15626 36032
rect 16022 36020 16028 36032
rect 15620 35992 16028 36020
rect 15620 35980 15626 35992
rect 16022 35980 16028 35992
rect 16080 35980 16086 36032
rect 24026 36020 24032 36032
rect 23987 35992 24032 36020
rect 24026 35980 24032 35992
rect 24084 35980 24090 36032
rect 33827 36023 33885 36029
rect 33827 35989 33839 36023
rect 33873 36020 33885 36023
rect 34698 36020 34704 36032
rect 33873 35992 34704 36020
rect 33873 35989 33885 35992
rect 33827 35983 33885 35989
rect 34698 35980 34704 35992
rect 34756 35980 34762 36032
rect 42291 36023 42349 36029
rect 42291 35989 42303 36023
rect 42337 36020 42349 36023
rect 42981 36023 43039 36029
rect 42981 36020 42993 36023
rect 42337 35992 42993 36020
rect 42337 35989 42349 35992
rect 42291 35983 42349 35989
rect 42981 35989 42993 35992
rect 43027 36020 43039 36023
rect 43070 36020 43076 36032
rect 43027 35992 43076 36020
rect 43027 35989 43039 35992
rect 42981 35983 43039 35989
rect 43070 35980 43076 35992
rect 43128 35980 43134 36032
rect 1104 35930 48852 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 48852 35930
rect 1104 35856 48852 35878
rect 5534 35816 5540 35828
rect 5495 35788 5540 35816
rect 5534 35776 5540 35788
rect 5592 35776 5598 35828
rect 5997 35819 6055 35825
rect 5997 35785 6009 35819
rect 6043 35816 6055 35819
rect 6086 35816 6092 35828
rect 6043 35788 6092 35816
rect 6043 35785 6055 35788
rect 5997 35779 6055 35785
rect 6086 35776 6092 35788
rect 6144 35776 6150 35828
rect 10134 35816 10140 35828
rect 10095 35788 10140 35816
rect 10134 35776 10140 35788
rect 10192 35776 10198 35828
rect 11698 35776 11704 35828
rect 11756 35816 11762 35828
rect 12161 35819 12219 35825
rect 12161 35816 12173 35819
rect 11756 35788 12173 35816
rect 11756 35776 11762 35788
rect 12161 35785 12173 35788
rect 12207 35785 12219 35819
rect 16206 35816 16212 35828
rect 16167 35788 16212 35816
rect 12161 35779 12219 35785
rect 16206 35776 16212 35788
rect 16264 35816 16270 35828
rect 16853 35819 16911 35825
rect 16853 35816 16865 35819
rect 16264 35788 16865 35816
rect 16264 35776 16270 35788
rect 16853 35785 16865 35788
rect 16899 35785 16911 35819
rect 19242 35816 19248 35828
rect 19203 35788 19248 35816
rect 16853 35779 16911 35785
rect 19242 35776 19248 35788
rect 19300 35776 19306 35828
rect 20533 35819 20591 35825
rect 20533 35785 20545 35819
rect 20579 35816 20591 35819
rect 20717 35819 20775 35825
rect 20717 35816 20729 35819
rect 20579 35788 20729 35816
rect 20579 35785 20591 35788
rect 20533 35779 20591 35785
rect 20717 35785 20729 35788
rect 20763 35816 20775 35819
rect 21082 35816 21088 35828
rect 20763 35788 21088 35816
rect 20763 35785 20775 35788
rect 20717 35779 20775 35785
rect 21082 35776 21088 35788
rect 21140 35776 21146 35828
rect 22833 35819 22891 35825
rect 22833 35785 22845 35819
rect 22879 35816 22891 35819
rect 23014 35816 23020 35828
rect 22879 35788 23020 35816
rect 22879 35785 22891 35788
rect 22833 35779 22891 35785
rect 23014 35776 23020 35788
rect 23072 35776 23078 35828
rect 28307 35819 28365 35825
rect 28307 35785 28319 35819
rect 28353 35816 28365 35819
rect 30466 35816 30472 35828
rect 28353 35788 30472 35816
rect 28353 35785 28365 35788
rect 28307 35779 28365 35785
rect 30466 35776 30472 35788
rect 30524 35776 30530 35828
rect 30558 35776 30564 35828
rect 30616 35816 30622 35828
rect 31205 35819 31263 35825
rect 30616 35788 30661 35816
rect 30616 35776 30622 35788
rect 31205 35785 31217 35819
rect 31251 35816 31263 35819
rect 31294 35816 31300 35828
rect 31251 35788 31300 35816
rect 31251 35785 31263 35788
rect 31205 35779 31263 35785
rect 31294 35776 31300 35788
rect 31352 35776 31358 35828
rect 31570 35816 31576 35828
rect 31531 35788 31576 35816
rect 31570 35776 31576 35788
rect 31628 35776 31634 35828
rect 32398 35776 32404 35828
rect 32456 35816 32462 35828
rect 32769 35819 32827 35825
rect 32769 35816 32781 35819
rect 32456 35788 32781 35816
rect 32456 35776 32462 35788
rect 32769 35785 32781 35788
rect 32815 35816 32827 35819
rect 35802 35816 35808 35828
rect 32815 35788 35808 35816
rect 32815 35785 32827 35788
rect 32769 35779 32827 35785
rect 35802 35776 35808 35788
rect 35860 35776 35866 35828
rect 36998 35776 37004 35828
rect 37056 35816 37062 35828
rect 37093 35819 37151 35825
rect 37093 35816 37105 35819
rect 37056 35788 37105 35816
rect 37056 35776 37062 35788
rect 37093 35785 37105 35788
rect 37139 35785 37151 35819
rect 38470 35816 38476 35828
rect 38431 35788 38476 35816
rect 37093 35779 37151 35785
rect 38470 35776 38476 35788
rect 38528 35776 38534 35828
rect 38930 35816 38936 35828
rect 38891 35788 38936 35816
rect 38930 35776 38936 35788
rect 38988 35776 38994 35828
rect 39163 35819 39221 35825
rect 39163 35785 39175 35819
rect 39209 35816 39221 35819
rect 40310 35816 40316 35828
rect 39209 35788 40316 35816
rect 39209 35785 39221 35788
rect 39163 35779 39221 35785
rect 40310 35776 40316 35788
rect 40368 35776 40374 35828
rect 40770 35816 40776 35828
rect 40731 35788 40776 35816
rect 40770 35776 40776 35788
rect 40828 35776 40834 35828
rect 41690 35776 41696 35828
rect 41748 35816 41754 35828
rect 42429 35819 42487 35825
rect 42429 35816 42441 35819
rect 41748 35788 42441 35816
rect 41748 35776 41754 35788
rect 42429 35785 42441 35788
rect 42475 35785 42487 35819
rect 42429 35779 42487 35785
rect 3743 35751 3801 35757
rect 3743 35717 3755 35751
rect 3789 35748 3801 35751
rect 6178 35748 6184 35760
rect 3789 35720 6184 35748
rect 3789 35717 3801 35720
rect 3743 35711 3801 35717
rect 6178 35708 6184 35720
rect 6236 35708 6242 35760
rect 11790 35708 11796 35760
rect 11848 35748 11854 35760
rect 11885 35751 11943 35757
rect 11885 35748 11897 35751
rect 11848 35720 11897 35748
rect 11848 35708 11854 35720
rect 11885 35717 11897 35720
rect 11931 35748 11943 35751
rect 14921 35751 14979 35757
rect 14921 35748 14933 35751
rect 11931 35720 14933 35748
rect 11931 35717 11943 35720
rect 11885 35711 11943 35717
rect 14921 35717 14933 35720
rect 14967 35748 14979 35751
rect 15286 35748 15292 35760
rect 14967 35720 15292 35748
rect 14967 35717 14979 35720
rect 14921 35711 14979 35717
rect 15286 35708 15292 35720
rect 15344 35708 15350 35760
rect 19981 35751 20039 35757
rect 19981 35717 19993 35751
rect 20027 35748 20039 35751
rect 21634 35748 21640 35760
rect 20027 35720 21640 35748
rect 20027 35717 20039 35720
rect 19981 35711 20039 35717
rect 21634 35708 21640 35720
rect 21692 35748 21698 35760
rect 21821 35751 21879 35757
rect 21821 35748 21833 35751
rect 21692 35720 21833 35748
rect 21692 35708 21698 35720
rect 21821 35717 21833 35720
rect 21867 35717 21879 35751
rect 21821 35711 21879 35717
rect 23198 35708 23204 35760
rect 23256 35748 23262 35760
rect 28077 35751 28135 35757
rect 23256 35720 28028 35748
rect 23256 35708 23262 35720
rect 6917 35683 6975 35689
rect 6917 35649 6929 35683
rect 6963 35680 6975 35683
rect 7190 35680 7196 35692
rect 6963 35652 7196 35680
rect 6963 35649 6975 35652
rect 6917 35643 6975 35649
rect 7190 35640 7196 35652
rect 7248 35640 7254 35692
rect 7561 35683 7619 35689
rect 7561 35649 7573 35683
rect 7607 35680 7619 35683
rect 8938 35680 8944 35692
rect 7607 35652 8944 35680
rect 7607 35649 7619 35652
rect 7561 35643 7619 35649
rect 8938 35640 8944 35652
rect 8996 35640 9002 35692
rect 11517 35683 11575 35689
rect 11517 35649 11529 35683
rect 11563 35680 11575 35683
rect 11974 35680 11980 35692
rect 11563 35652 11980 35680
rect 11563 35649 11575 35652
rect 11517 35643 11575 35649
rect 11974 35640 11980 35652
rect 12032 35640 12038 35692
rect 13630 35680 13636 35692
rect 13591 35652 13636 35680
rect 13630 35640 13636 35652
rect 13688 35640 13694 35692
rect 14274 35680 14280 35692
rect 14187 35652 14280 35680
rect 14274 35640 14280 35652
rect 14332 35680 14338 35692
rect 15473 35683 15531 35689
rect 15473 35680 15485 35683
rect 14332 35652 15485 35680
rect 14332 35640 14338 35652
rect 15473 35649 15485 35652
rect 15519 35649 15531 35683
rect 15473 35643 15531 35649
rect 21269 35683 21327 35689
rect 21269 35649 21281 35683
rect 21315 35680 21327 35683
rect 22186 35680 22192 35692
rect 21315 35652 22192 35680
rect 21315 35649 21327 35652
rect 21269 35643 21327 35649
rect 22186 35640 22192 35652
rect 22244 35640 22250 35692
rect 23477 35683 23535 35689
rect 23477 35649 23489 35683
rect 23523 35680 23535 35683
rect 24121 35683 24179 35689
rect 24121 35680 24133 35683
rect 23523 35652 24133 35680
rect 23523 35649 23535 35652
rect 23477 35643 23535 35649
rect 24121 35649 24133 35652
rect 24167 35680 24179 35683
rect 24302 35680 24308 35692
rect 24167 35652 24308 35680
rect 24167 35649 24179 35652
rect 24121 35643 24179 35649
rect 24302 35640 24308 35652
rect 24360 35640 24366 35692
rect 24949 35683 25007 35689
rect 24949 35649 24961 35683
rect 24995 35680 25007 35683
rect 26878 35680 26884 35692
rect 24995 35652 26884 35680
rect 24995 35649 25007 35652
rect 24949 35643 25007 35649
rect 26878 35640 26884 35652
rect 26936 35640 26942 35692
rect 26970 35640 26976 35692
rect 27028 35680 27034 35692
rect 28000 35680 28028 35720
rect 28077 35717 28089 35751
rect 28123 35748 28135 35751
rect 28902 35748 28908 35760
rect 28123 35720 28908 35748
rect 28123 35717 28135 35720
rect 28077 35711 28135 35717
rect 28902 35708 28908 35720
rect 28960 35708 28966 35760
rect 31312 35680 31340 35776
rect 33226 35708 33232 35760
rect 33284 35748 33290 35760
rect 34241 35751 34299 35757
rect 34241 35748 34253 35751
rect 33284 35720 34253 35748
rect 33284 35708 33290 35720
rect 34241 35717 34253 35720
rect 34287 35717 34299 35751
rect 34241 35711 34299 35717
rect 39945 35751 40003 35757
rect 39945 35717 39957 35751
rect 39991 35748 40003 35751
rect 40788 35748 40816 35776
rect 39991 35720 40816 35748
rect 39991 35717 40003 35720
rect 39945 35711 40003 35717
rect 31757 35683 31815 35689
rect 31757 35680 31769 35683
rect 27028 35652 27073 35680
rect 28000 35652 28279 35680
rect 31312 35652 31769 35680
rect 27028 35640 27034 35652
rect 3672 35615 3730 35621
rect 3672 35581 3684 35615
rect 3718 35612 3730 35615
rect 4614 35612 4620 35624
rect 3718 35584 4154 35612
rect 4575 35584 4620 35612
rect 3718 35581 3730 35584
rect 3672 35575 3730 35581
rect 4126 35488 4154 35584
rect 4614 35572 4620 35584
rect 4672 35572 4678 35624
rect 28251 35621 28279 35652
rect 31757 35649 31769 35652
rect 31803 35649 31815 35683
rect 31757 35643 31815 35649
rect 32401 35683 32459 35689
rect 32401 35649 32413 35683
rect 32447 35680 32459 35683
rect 32447 35652 34008 35680
rect 32447 35649 32459 35652
rect 32401 35643 32459 35649
rect 12596 35615 12654 35621
rect 12596 35581 12608 35615
rect 12642 35612 12654 35615
rect 16669 35615 16727 35621
rect 12642 35584 13124 35612
rect 12642 35581 12654 35584
rect 12596 35575 12654 35581
rect 4938 35547 4996 35553
rect 4938 35513 4950 35547
rect 4984 35513 4996 35547
rect 4938 35507 4996 35513
rect 6641 35547 6699 35553
rect 6641 35513 6653 35547
rect 6687 35544 6699 35547
rect 7009 35547 7067 35553
rect 7009 35544 7021 35547
rect 6687 35516 7021 35544
rect 6687 35513 6699 35516
rect 6641 35507 6699 35513
rect 7009 35513 7021 35516
rect 7055 35544 7067 35547
rect 7098 35544 7104 35556
rect 7055 35516 7104 35544
rect 7055 35513 7067 35516
rect 7009 35507 7067 35513
rect 4126 35448 4160 35488
rect 4154 35436 4160 35448
rect 4212 35476 4218 35488
rect 4525 35479 4583 35485
rect 4212 35448 4257 35476
rect 4212 35436 4218 35448
rect 4525 35445 4537 35479
rect 4571 35476 4583 35479
rect 4706 35476 4712 35488
rect 4571 35448 4712 35476
rect 4571 35445 4583 35448
rect 4525 35439 4583 35445
rect 4706 35436 4712 35448
rect 4764 35476 4770 35488
rect 4953 35476 4981 35507
rect 7098 35504 7104 35516
rect 7156 35544 7162 35556
rect 9306 35544 9312 35556
rect 7156 35516 9312 35544
rect 7156 35504 7162 35516
rect 9306 35504 9312 35516
rect 9364 35504 9370 35556
rect 9769 35547 9827 35553
rect 9769 35513 9781 35547
rect 9815 35544 9827 35547
rect 10410 35544 10416 35556
rect 9815 35516 10416 35544
rect 9815 35513 9827 35516
rect 9769 35507 9827 35513
rect 10410 35504 10416 35516
rect 10468 35504 10474 35556
rect 10870 35544 10876 35556
rect 10831 35516 10876 35544
rect 10870 35504 10876 35516
rect 10928 35504 10934 35556
rect 13096 35553 13124 35584
rect 16669 35581 16681 35615
rect 16715 35612 16727 35615
rect 28236 35615 28294 35621
rect 16715 35584 17264 35612
rect 16715 35581 16727 35584
rect 16669 35575 16727 35581
rect 10965 35547 11023 35553
rect 10965 35513 10977 35547
rect 11011 35544 11023 35547
rect 13081 35547 13139 35553
rect 11011 35516 13032 35544
rect 11011 35513 11023 35516
rect 10965 35507 11023 35513
rect 7834 35476 7840 35488
rect 4764 35448 4981 35476
rect 7795 35448 7840 35476
rect 4764 35436 4770 35448
rect 7834 35436 7840 35448
rect 7892 35436 7898 35488
rect 8202 35476 8208 35488
rect 8163 35448 8208 35476
rect 8202 35436 8208 35448
rect 8260 35436 8266 35488
rect 10686 35476 10692 35488
rect 10599 35448 10692 35476
rect 10686 35436 10692 35448
rect 10744 35476 10750 35488
rect 10980 35476 11008 35507
rect 10744 35448 11008 35476
rect 12667 35479 12725 35485
rect 10744 35436 10750 35448
rect 12667 35445 12679 35479
rect 12713 35476 12725 35479
rect 12894 35476 12900 35488
rect 12713 35448 12900 35476
rect 12713 35445 12725 35448
rect 12667 35439 12725 35445
rect 12894 35436 12900 35448
rect 12952 35436 12958 35488
rect 13004 35476 13032 35516
rect 13081 35513 13093 35547
rect 13127 35544 13139 35547
rect 13446 35544 13452 35556
rect 13127 35516 13452 35544
rect 13127 35513 13139 35516
rect 13081 35507 13139 35513
rect 13446 35504 13452 35516
rect 13504 35504 13510 35556
rect 13722 35544 13728 35556
rect 13683 35516 13728 35544
rect 13722 35504 13728 35516
rect 13780 35504 13786 35556
rect 15197 35547 15255 35553
rect 15197 35544 15209 35547
rect 14568 35516 15209 35544
rect 13357 35479 13415 35485
rect 13357 35476 13369 35479
rect 13004 35448 13369 35476
rect 13357 35445 13369 35448
rect 13403 35476 13415 35479
rect 13740 35476 13768 35504
rect 14568 35488 14596 35516
rect 15197 35513 15209 35516
rect 15243 35513 15255 35547
rect 15197 35507 15255 35513
rect 15286 35504 15292 35556
rect 15344 35544 15350 35556
rect 15344 35516 15389 35544
rect 15344 35504 15350 35516
rect 17236 35488 17264 35584
rect 28236 35581 28248 35615
rect 28282 35612 28294 35615
rect 29270 35612 29276 35624
rect 28282 35581 28304 35612
rect 29231 35584 29276 35612
rect 28236 35575 28304 35581
rect 18325 35547 18383 35553
rect 18325 35513 18337 35547
rect 18371 35544 18383 35547
rect 18877 35547 18935 35553
rect 18877 35544 18889 35547
rect 18371 35516 18889 35544
rect 18371 35513 18383 35516
rect 18325 35507 18383 35513
rect 18877 35513 18889 35516
rect 18923 35544 18935 35547
rect 19429 35547 19487 35553
rect 19429 35544 19441 35547
rect 18923 35516 19441 35544
rect 18923 35513 18935 35516
rect 18877 35507 18935 35513
rect 19429 35513 19441 35516
rect 19475 35513 19487 35547
rect 19429 35507 19487 35513
rect 19521 35547 19579 35553
rect 19521 35513 19533 35547
rect 19567 35544 19579 35547
rect 19886 35544 19892 35556
rect 19567 35516 19892 35544
rect 19567 35513 19579 35516
rect 19521 35507 19579 35513
rect 19886 35504 19892 35516
rect 19944 35544 19950 35556
rect 20533 35547 20591 35553
rect 20533 35544 20545 35547
rect 19944 35516 20545 35544
rect 19944 35504 19950 35516
rect 20533 35513 20545 35516
rect 20579 35513 20591 35547
rect 20533 35507 20591 35513
rect 21085 35547 21143 35553
rect 21085 35513 21097 35547
rect 21131 35544 21143 35547
rect 21358 35544 21364 35556
rect 21131 35516 21364 35544
rect 21131 35513 21143 35516
rect 21085 35507 21143 35513
rect 21358 35504 21364 35516
rect 21416 35504 21422 35556
rect 24026 35504 24032 35556
rect 24084 35544 24090 35556
rect 24305 35547 24363 35553
rect 24305 35544 24317 35547
rect 24084 35516 24317 35544
rect 24084 35504 24090 35516
rect 24305 35513 24317 35516
rect 24351 35513 24363 35547
rect 24305 35507 24363 35513
rect 24394 35504 24400 35556
rect 24452 35544 24458 35556
rect 24452 35516 24497 35544
rect 24452 35504 24458 35516
rect 26326 35504 26332 35556
rect 26384 35544 26390 35556
rect 26513 35547 26571 35553
rect 26513 35544 26525 35547
rect 26384 35516 26525 35544
rect 26384 35504 26390 35516
rect 26513 35513 26525 35516
rect 26559 35513 26571 35547
rect 26513 35507 26571 35513
rect 26605 35547 26663 35553
rect 26605 35513 26617 35547
rect 26651 35513 26663 35547
rect 26605 35507 26663 35513
rect 14550 35476 14556 35488
rect 13403 35448 13768 35476
rect 14511 35448 14556 35476
rect 13403 35445 13415 35448
rect 13357 35439 13415 35445
rect 14550 35436 14556 35448
rect 14608 35436 14614 35488
rect 17218 35476 17224 35488
rect 17179 35448 17224 35476
rect 17218 35436 17224 35448
rect 17276 35436 17282 35488
rect 17678 35476 17684 35488
rect 17639 35448 17684 35476
rect 17678 35436 17684 35448
rect 17736 35436 17742 35488
rect 24118 35436 24124 35488
rect 24176 35476 24182 35488
rect 25225 35479 25283 35485
rect 25225 35476 25237 35479
rect 24176 35448 25237 35476
rect 24176 35436 24182 35448
rect 25225 35445 25237 35448
rect 25271 35445 25283 35479
rect 25225 35439 25283 35445
rect 25961 35479 26019 35485
rect 25961 35445 25973 35479
rect 26007 35476 26019 35479
rect 26237 35479 26295 35485
rect 26237 35476 26249 35479
rect 26007 35448 26249 35476
rect 26007 35445 26019 35448
rect 25961 35439 26019 35445
rect 26237 35445 26249 35448
rect 26283 35476 26295 35479
rect 26418 35476 26424 35488
rect 26283 35448 26424 35476
rect 26283 35445 26295 35448
rect 26237 35439 26295 35445
rect 26418 35436 26424 35448
rect 26476 35476 26482 35488
rect 26620 35476 26648 35507
rect 28276 35488 28304 35575
rect 29270 35572 29276 35584
rect 29328 35572 29334 35624
rect 29089 35547 29147 35553
rect 29089 35513 29101 35547
rect 29135 35544 29147 35547
rect 29546 35544 29552 35556
rect 29135 35516 29552 35544
rect 29135 35513 29147 35516
rect 29089 35507 29147 35513
rect 29546 35504 29552 35516
rect 29604 35553 29610 35556
rect 29604 35547 29652 35553
rect 29604 35513 29606 35547
rect 29640 35513 29652 35547
rect 31846 35544 31852 35556
rect 31807 35516 31852 35544
rect 29604 35507 29652 35513
rect 29604 35504 29610 35507
rect 31846 35504 31852 35516
rect 31904 35504 31910 35556
rect 33318 35544 33324 35556
rect 33279 35516 33324 35544
rect 33318 35504 33324 35516
rect 33376 35504 33382 35556
rect 33410 35504 33416 35556
rect 33468 35544 33474 35556
rect 33980 35553 34008 35652
rect 36814 35640 36820 35692
rect 36872 35680 36878 35692
rect 41230 35680 41236 35692
rect 36872 35652 41236 35680
rect 36872 35640 36878 35652
rect 41230 35640 41236 35652
rect 41288 35640 41294 35692
rect 43070 35680 43076 35692
rect 43031 35652 43076 35680
rect 43070 35640 43076 35652
rect 43128 35640 43134 35692
rect 43254 35640 43260 35692
rect 43312 35680 43318 35692
rect 43349 35683 43407 35689
rect 43349 35680 43361 35683
rect 43312 35652 43361 35680
rect 43312 35640 43318 35652
rect 43349 35649 43361 35652
rect 43395 35649 43407 35683
rect 43349 35643 43407 35649
rect 35894 35612 35900 35624
rect 35855 35584 35900 35612
rect 35894 35572 35900 35584
rect 35952 35572 35958 35624
rect 36265 35615 36323 35621
rect 36265 35581 36277 35615
rect 36311 35581 36323 35615
rect 36265 35575 36323 35581
rect 36449 35615 36507 35621
rect 36449 35581 36461 35615
rect 36495 35612 36507 35615
rect 37274 35612 37280 35624
rect 36495 35584 37280 35612
rect 36495 35581 36507 35584
rect 36449 35575 36507 35581
rect 33965 35547 34023 35553
rect 33468 35516 33513 35544
rect 33468 35504 33474 35516
rect 33965 35513 33977 35547
rect 34011 35544 34023 35547
rect 34238 35544 34244 35556
rect 34011 35516 34244 35544
rect 34011 35513 34023 35516
rect 33965 35507 34023 35513
rect 34238 35504 34244 35516
rect 34296 35504 34302 35556
rect 35621 35547 35679 35553
rect 35621 35513 35633 35547
rect 35667 35544 35679 35547
rect 36280 35544 36308 35575
rect 37274 35572 37280 35584
rect 37332 35572 37338 35624
rect 38010 35572 38016 35624
rect 38068 35612 38074 35624
rect 39060 35615 39118 35621
rect 39060 35612 39072 35615
rect 38068 35584 39072 35612
rect 38068 35572 38074 35584
rect 39060 35581 39072 35584
rect 39106 35612 39118 35615
rect 39485 35615 39543 35621
rect 39485 35612 39497 35615
rect 39106 35584 39497 35612
rect 39106 35581 39118 35584
rect 39060 35575 39118 35581
rect 39485 35581 39497 35584
rect 39531 35581 39543 35615
rect 39485 35575 39543 35581
rect 35667 35516 36584 35544
rect 35667 35513 35679 35516
rect 35621 35507 35679 35513
rect 27522 35476 27528 35488
rect 26476 35448 26648 35476
rect 27483 35448 27528 35476
rect 26476 35436 26482 35448
rect 27522 35436 27528 35448
rect 27580 35436 27586 35488
rect 28258 35436 28264 35488
rect 28316 35476 28322 35488
rect 28629 35479 28687 35485
rect 28629 35476 28641 35479
rect 28316 35448 28641 35476
rect 28316 35436 28322 35448
rect 28629 35445 28641 35448
rect 28675 35445 28687 35479
rect 30190 35476 30196 35488
rect 30151 35448 30196 35476
rect 28629 35439 28687 35445
rect 30190 35436 30196 35448
rect 30248 35436 30254 35488
rect 33042 35476 33048 35488
rect 32955 35448 33048 35476
rect 33042 35436 33048 35448
rect 33100 35476 33106 35488
rect 33428 35476 33456 35504
rect 36556 35488 36584 35516
rect 36998 35504 37004 35556
rect 37056 35544 37062 35556
rect 37598 35547 37656 35553
rect 37598 35544 37610 35547
rect 37056 35516 37610 35544
rect 37056 35504 37062 35516
rect 37598 35513 37610 35516
rect 37644 35513 37656 35547
rect 39206 35544 39212 35556
rect 37598 35507 37656 35513
rect 38212 35516 39212 35544
rect 33100 35448 33456 35476
rect 33100 35436 33106 35448
rect 34606 35436 34612 35488
rect 34664 35476 34670 35488
rect 35069 35479 35127 35485
rect 35069 35476 35081 35479
rect 34664 35448 35081 35476
rect 34664 35436 34670 35448
rect 35069 35445 35081 35448
rect 35115 35445 35127 35479
rect 35069 35439 35127 35445
rect 36538 35436 36544 35488
rect 36596 35476 36602 35488
rect 38212 35485 38240 35516
rect 39206 35504 39212 35516
rect 39264 35504 39270 35556
rect 41554 35547 41612 35553
rect 41554 35544 41566 35547
rect 41064 35516 41566 35544
rect 36725 35479 36783 35485
rect 36725 35476 36737 35479
rect 36596 35448 36737 35476
rect 36596 35436 36602 35448
rect 36725 35445 36737 35448
rect 36771 35445 36783 35479
rect 36725 35439 36783 35445
rect 38197 35479 38255 35485
rect 38197 35445 38209 35479
rect 38243 35445 38255 35479
rect 38197 35439 38255 35445
rect 39114 35436 39120 35488
rect 39172 35476 39178 35488
rect 41064 35485 41092 35516
rect 41554 35513 41566 35516
rect 41600 35513 41612 35547
rect 42797 35547 42855 35553
rect 42797 35544 42809 35547
rect 41554 35507 41612 35513
rect 42168 35516 42809 35544
rect 41049 35479 41107 35485
rect 41049 35476 41061 35479
rect 39172 35448 41061 35476
rect 39172 35436 39178 35448
rect 41049 35445 41061 35448
rect 41095 35445 41107 35479
rect 41049 35439 41107 35445
rect 41874 35436 41880 35488
rect 41932 35476 41938 35488
rect 42168 35485 42196 35516
rect 42797 35513 42809 35516
rect 42843 35513 42855 35547
rect 42797 35507 42855 35513
rect 43165 35547 43223 35553
rect 43165 35513 43177 35547
rect 43211 35513 43223 35547
rect 43165 35507 43223 35513
rect 42153 35479 42211 35485
rect 42153 35476 42165 35479
rect 41932 35448 42165 35476
rect 41932 35436 41938 35448
rect 42153 35445 42165 35448
rect 42199 35445 42211 35479
rect 42812 35476 42840 35507
rect 43180 35476 43208 35507
rect 42812 35448 43208 35476
rect 42153 35439 42211 35445
rect 43898 35436 43904 35488
rect 43956 35476 43962 35488
rect 43993 35479 44051 35485
rect 43993 35476 44005 35479
rect 43956 35448 44005 35476
rect 43956 35436 43962 35448
rect 43993 35445 44005 35448
rect 44039 35445 44051 35479
rect 43993 35439 44051 35445
rect 1104 35386 48852 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 48852 35386
rect 1104 35312 48852 35334
rect 4706 35272 4712 35284
rect 4667 35244 4712 35272
rect 4706 35232 4712 35244
rect 4764 35232 4770 35284
rect 5258 35272 5264 35284
rect 5219 35244 5264 35272
rect 5258 35232 5264 35244
rect 5316 35232 5322 35284
rect 5994 35272 6000 35284
rect 5955 35244 6000 35272
rect 5994 35232 6000 35244
rect 6052 35232 6058 35284
rect 13078 35272 13084 35284
rect 13039 35244 13084 35272
rect 13078 35232 13084 35244
rect 13136 35232 13142 35284
rect 13633 35275 13691 35281
rect 13633 35241 13645 35275
rect 13679 35272 13691 35275
rect 13998 35272 14004 35284
rect 13679 35244 14004 35272
rect 13679 35241 13691 35244
rect 13633 35235 13691 35241
rect 13998 35232 14004 35244
rect 14056 35232 14062 35284
rect 19337 35275 19395 35281
rect 19337 35241 19349 35275
rect 19383 35272 19395 35275
rect 20714 35272 20720 35284
rect 19383 35244 19748 35272
rect 20675 35244 20720 35272
rect 19383 35241 19395 35244
rect 19337 35235 19395 35241
rect 6086 35164 6092 35216
rect 6144 35204 6150 35216
rect 6410 35207 6468 35213
rect 6410 35204 6422 35207
rect 6144 35176 6422 35204
rect 6144 35164 6150 35176
rect 6410 35173 6422 35176
rect 6456 35173 6468 35207
rect 6410 35167 6468 35173
rect 7926 35164 7932 35216
rect 7984 35204 7990 35216
rect 8021 35207 8079 35213
rect 8021 35204 8033 35207
rect 7984 35176 8033 35204
rect 7984 35164 7990 35176
rect 8021 35173 8033 35176
rect 8067 35173 8079 35207
rect 8021 35167 8079 35173
rect 8573 35207 8631 35213
rect 8573 35173 8585 35207
rect 8619 35204 8631 35207
rect 8938 35204 8944 35216
rect 8619 35176 8944 35204
rect 8619 35173 8631 35176
rect 8573 35167 8631 35173
rect 8938 35164 8944 35176
rect 8996 35164 9002 35216
rect 9306 35164 9312 35216
rect 9364 35204 9370 35216
rect 9861 35207 9919 35213
rect 9861 35204 9873 35207
rect 9364 35176 9873 35204
rect 9364 35164 9370 35176
rect 9861 35173 9873 35176
rect 9907 35204 9919 35207
rect 10686 35204 10692 35216
rect 9907 35176 10692 35204
rect 9907 35173 9919 35176
rect 9861 35167 9919 35173
rect 10686 35164 10692 35176
rect 10744 35164 10750 35216
rect 11698 35204 11704 35216
rect 11659 35176 11704 35204
rect 11698 35164 11704 35176
rect 11756 35164 11762 35216
rect 13722 35164 13728 35216
rect 13780 35204 13786 35216
rect 15565 35207 15623 35213
rect 15565 35204 15577 35207
rect 13780 35176 15577 35204
rect 13780 35164 13786 35176
rect 15565 35173 15577 35176
rect 15611 35204 15623 35207
rect 15654 35204 15660 35216
rect 15611 35176 15660 35204
rect 15611 35173 15623 35176
rect 15565 35167 15623 35173
rect 15654 35164 15660 35176
rect 15712 35164 15718 35216
rect 17678 35164 17684 35216
rect 17736 35204 17742 35216
rect 18779 35207 18837 35213
rect 18779 35204 18791 35207
rect 17736 35176 18791 35204
rect 17736 35164 17742 35176
rect 18779 35173 18791 35176
rect 18825 35204 18837 35207
rect 19150 35204 19156 35216
rect 18825 35176 19156 35204
rect 18825 35173 18837 35176
rect 18779 35167 18837 35173
rect 19150 35164 19156 35176
rect 19208 35164 19214 35216
rect 19720 35213 19748 35244
rect 20714 35232 20720 35244
rect 20772 35232 20778 35284
rect 21266 35272 21272 35284
rect 21227 35244 21272 35272
rect 21266 35232 21272 35244
rect 21324 35232 21330 35284
rect 21358 35232 21364 35284
rect 21416 35272 21422 35284
rect 21821 35275 21879 35281
rect 21821 35272 21833 35275
rect 21416 35244 21833 35272
rect 21416 35232 21422 35244
rect 21821 35241 21833 35244
rect 21867 35241 21879 35275
rect 21821 35235 21879 35241
rect 22186 35232 22192 35284
rect 22244 35272 22250 35284
rect 22787 35275 22845 35281
rect 22787 35272 22799 35275
rect 22244 35244 22799 35272
rect 22244 35232 22250 35244
rect 22787 35241 22799 35244
rect 22833 35241 22845 35275
rect 26970 35272 26976 35284
rect 22787 35235 22845 35241
rect 25561 35244 26976 35272
rect 19705 35207 19763 35213
rect 19705 35173 19717 35207
rect 19751 35204 19763 35207
rect 19886 35204 19892 35216
rect 19751 35176 19892 35204
rect 19751 35173 19763 35176
rect 19705 35167 19763 35173
rect 19886 35164 19892 35176
rect 19944 35164 19950 35216
rect 24302 35204 24308 35216
rect 24263 35176 24308 35204
rect 24302 35164 24308 35176
rect 24360 35164 24366 35216
rect 24857 35207 24915 35213
rect 24857 35173 24869 35207
rect 24903 35204 24915 35207
rect 25561 35204 25589 35244
rect 26970 35232 26976 35244
rect 27028 35232 27034 35284
rect 28905 35275 28963 35281
rect 28905 35241 28917 35275
rect 28951 35272 28963 35275
rect 29086 35272 29092 35284
rect 28951 35244 29092 35272
rect 28951 35241 28963 35244
rect 28905 35235 28963 35241
rect 29086 35232 29092 35244
rect 29144 35232 29150 35284
rect 30466 35232 30472 35284
rect 30524 35272 30530 35284
rect 30929 35275 30987 35281
rect 30929 35272 30941 35275
rect 30524 35244 30941 35272
rect 30524 35232 30530 35244
rect 30929 35241 30941 35244
rect 30975 35241 30987 35275
rect 33042 35272 33048 35284
rect 30929 35235 30987 35241
rect 31496 35244 33048 35272
rect 24903 35176 25589 35204
rect 24903 35173 24915 35176
rect 24857 35167 24915 35173
rect 26418 35164 26424 35216
rect 26476 35204 26482 35216
rect 26697 35207 26755 35213
rect 26697 35204 26709 35207
rect 26476 35176 26709 35204
rect 26476 35164 26482 35176
rect 26697 35173 26709 35176
rect 26743 35173 26755 35207
rect 26697 35167 26755 35173
rect 29546 35164 29552 35216
rect 29604 35204 29610 35216
rect 29730 35213 29736 35216
rect 29686 35207 29736 35213
rect 29686 35204 29698 35207
rect 29604 35176 29698 35204
rect 29604 35164 29610 35176
rect 29686 35173 29698 35176
rect 29732 35173 29736 35207
rect 29686 35167 29736 35173
rect 29730 35164 29736 35167
rect 29788 35164 29794 35216
rect 30190 35164 30196 35216
rect 30248 35204 30254 35216
rect 30653 35207 30711 35213
rect 30653 35204 30665 35207
rect 30248 35176 30665 35204
rect 30248 35164 30254 35176
rect 30653 35173 30665 35176
rect 30699 35204 30711 35207
rect 31496 35204 31524 35244
rect 33042 35232 33048 35244
rect 33100 35232 33106 35284
rect 33410 35232 33416 35284
rect 33468 35272 33474 35284
rect 37274 35272 37280 35284
rect 33468 35244 35480 35272
rect 37235 35244 37280 35272
rect 33468 35232 33474 35244
rect 33888 35213 33916 35244
rect 32309 35207 32367 35213
rect 32309 35204 32321 35207
rect 30699 35176 31524 35204
rect 31864 35176 32321 35204
rect 30699 35173 30711 35176
rect 30653 35167 30711 35173
rect 31864 35148 31892 35176
rect 32309 35173 32321 35176
rect 32355 35173 32367 35207
rect 32309 35167 32367 35173
rect 33873 35207 33931 35213
rect 33873 35173 33885 35207
rect 33919 35173 33931 35207
rect 33873 35167 33931 35173
rect 34698 35164 34704 35216
rect 34756 35204 34762 35216
rect 35342 35204 35348 35216
rect 34756 35176 35348 35204
rect 34756 35164 34762 35176
rect 35342 35164 35348 35176
rect 35400 35164 35406 35216
rect 35452 35213 35480 35244
rect 37274 35232 37280 35244
rect 37332 35232 37338 35284
rect 41230 35272 41236 35284
rect 41191 35244 41236 35272
rect 41230 35232 41236 35244
rect 41288 35232 41294 35284
rect 35437 35207 35495 35213
rect 35437 35173 35449 35207
rect 35483 35204 35495 35207
rect 35710 35204 35716 35216
rect 35483 35176 35716 35204
rect 35483 35173 35495 35176
rect 35437 35167 35495 35173
rect 35710 35164 35716 35176
rect 35768 35164 35774 35216
rect 38194 35204 38200 35216
rect 38073 35176 38200 35204
rect 4154 35096 4160 35148
rect 4212 35136 4218 35148
rect 7009 35139 7067 35145
rect 7009 35136 7021 35139
rect 4212 35108 7021 35136
rect 4212 35096 4218 35108
rect 7009 35105 7021 35108
rect 7055 35105 7067 35139
rect 7009 35099 7067 35105
rect 11584 35139 11642 35145
rect 11584 35105 11596 35139
rect 11630 35136 11642 35139
rect 11882 35136 11888 35148
rect 11630 35108 11888 35136
rect 11630 35105 11642 35108
rect 11584 35099 11642 35105
rect 11882 35096 11888 35108
rect 11940 35096 11946 35148
rect 17012 35139 17070 35145
rect 17012 35105 17024 35139
rect 17058 35136 17070 35139
rect 17218 35136 17224 35148
rect 17058 35108 17224 35136
rect 17058 35105 17070 35108
rect 17012 35099 17070 35105
rect 17218 35096 17224 35108
rect 17276 35096 17282 35148
rect 22716 35139 22774 35145
rect 22716 35105 22728 35139
rect 22762 35136 22774 35139
rect 22830 35136 22836 35148
rect 22762 35108 22836 35136
rect 22762 35105 22774 35108
rect 22716 35099 22774 35105
rect 22830 35096 22836 35108
rect 22888 35136 22894 35148
rect 23198 35136 23204 35148
rect 22888 35108 23204 35136
rect 22888 35096 22894 35108
rect 23198 35096 23204 35108
rect 23256 35096 23262 35148
rect 28388 35139 28446 35145
rect 28388 35105 28400 35139
rect 28434 35105 28446 35139
rect 29362 35136 29368 35148
rect 29323 35108 29368 35136
rect 28388 35099 28446 35105
rect 4062 35028 4068 35080
rect 4120 35068 4126 35080
rect 4341 35071 4399 35077
rect 4341 35068 4353 35071
rect 4120 35040 4353 35068
rect 4120 35028 4126 35040
rect 4341 35037 4353 35040
rect 4387 35037 4399 35071
rect 4341 35031 4399 35037
rect 6089 35071 6147 35077
rect 6089 35037 6101 35071
rect 6135 35068 6147 35071
rect 6454 35068 6460 35080
rect 6135 35040 6460 35068
rect 6135 35037 6147 35040
rect 6089 35031 6147 35037
rect 6454 35028 6460 35040
rect 6512 35028 6518 35080
rect 7926 35068 7932 35080
rect 7887 35040 7932 35068
rect 7926 35028 7932 35040
rect 7984 35028 7990 35080
rect 8570 35028 8576 35080
rect 8628 35068 8634 35080
rect 9769 35071 9827 35077
rect 9769 35068 9781 35071
rect 8628 35040 9781 35068
rect 8628 35028 8634 35040
rect 9769 35037 9781 35040
rect 9815 35037 9827 35071
rect 10410 35068 10416 35080
rect 10371 35040 10416 35068
rect 9769 35031 9827 35037
rect 9784 35000 9812 35031
rect 10410 35028 10416 35040
rect 10468 35028 10474 35080
rect 12710 35068 12716 35080
rect 12671 35040 12716 35068
rect 12710 35028 12716 35040
rect 12768 35028 12774 35080
rect 15473 35071 15531 35077
rect 15473 35037 15485 35071
rect 15519 35068 15531 35071
rect 16574 35068 16580 35080
rect 15519 35040 16580 35068
rect 15519 35037 15531 35040
rect 15473 35031 15531 35037
rect 16574 35028 16580 35040
rect 16632 35028 16638 35080
rect 18414 35068 18420 35080
rect 18375 35040 18420 35068
rect 18414 35028 18420 35040
rect 18472 35028 18478 35080
rect 20530 35028 20536 35080
rect 20588 35068 20594 35080
rect 20901 35071 20959 35077
rect 20901 35068 20913 35071
rect 20588 35040 20913 35068
rect 20588 35028 20594 35040
rect 20901 35037 20913 35040
rect 20947 35037 20959 35071
rect 20901 35031 20959 35037
rect 21818 35028 21824 35080
rect 21876 35068 21882 35080
rect 22097 35071 22155 35077
rect 22097 35068 22109 35071
rect 21876 35040 22109 35068
rect 21876 35028 21882 35040
rect 22097 35037 22109 35040
rect 22143 35037 22155 35071
rect 24210 35068 24216 35080
rect 24171 35040 24216 35068
rect 22097 35031 22155 35037
rect 24210 35028 24216 35040
rect 24268 35028 24274 35080
rect 26602 35068 26608 35080
rect 26563 35040 26608 35068
rect 26602 35028 26608 35040
rect 26660 35028 26666 35080
rect 26878 35068 26884 35080
rect 26839 35040 26884 35068
rect 26878 35028 26884 35040
rect 26936 35028 26942 35080
rect 28403 35068 28431 35099
rect 29362 35096 29368 35108
rect 29420 35096 29426 35148
rect 30285 35139 30343 35145
rect 30285 35105 30297 35139
rect 30331 35136 30343 35139
rect 30558 35136 30564 35148
rect 30331 35108 30564 35136
rect 30331 35105 30343 35108
rect 30285 35099 30343 35105
rect 30558 35096 30564 35108
rect 30616 35136 30622 35148
rect 31665 35139 31723 35145
rect 31665 35136 31677 35139
rect 30616 35108 31677 35136
rect 30616 35096 30622 35108
rect 31665 35105 31677 35108
rect 31711 35136 31723 35139
rect 31846 35136 31852 35148
rect 31711 35108 31852 35136
rect 31711 35105 31723 35108
rect 31665 35099 31723 35105
rect 31846 35096 31852 35108
rect 31904 35096 31910 35148
rect 38073 35145 38101 35176
rect 38194 35164 38200 35176
rect 38252 35164 38258 35216
rect 39206 35204 39212 35216
rect 39167 35176 39212 35204
rect 39206 35164 39212 35176
rect 39264 35164 39270 35216
rect 41874 35204 41880 35216
rect 41835 35176 41880 35204
rect 41874 35164 41880 35176
rect 41932 35164 41938 35216
rect 38059 35139 38117 35145
rect 38059 35105 38071 35139
rect 38105 35105 38117 35139
rect 40586 35136 40592 35148
rect 40547 35108 40592 35136
rect 38059 35099 38117 35105
rect 40586 35096 40592 35108
rect 40644 35096 40650 35148
rect 43254 35136 43260 35148
rect 43215 35108 43260 35136
rect 43254 35096 43260 35108
rect 43312 35096 43318 35148
rect 29546 35068 29552 35080
rect 28403 35040 29552 35068
rect 11146 35000 11152 35012
rect 9784 34972 11152 35000
rect 11146 34960 11152 34972
rect 11204 34960 11210 35012
rect 16022 35000 16028 35012
rect 15983 34972 16028 35000
rect 16022 34960 16028 34972
rect 16080 34960 16086 35012
rect 25774 34960 25780 35012
rect 25832 35000 25838 35012
rect 28403 35000 28431 35040
rect 29546 35028 29552 35040
rect 29604 35028 29610 35080
rect 32214 35068 32220 35080
rect 32175 35040 32220 35068
rect 32214 35028 32220 35040
rect 32272 35028 32278 35080
rect 33778 35068 33784 35080
rect 33739 35040 33784 35068
rect 33778 35028 33784 35040
rect 33836 35028 33842 35080
rect 34057 35071 34115 35077
rect 34057 35037 34069 35071
rect 34103 35037 34115 35071
rect 35618 35068 35624 35080
rect 35579 35040 35624 35068
rect 34057 35031 34115 35037
rect 25832 34972 28431 35000
rect 32769 35003 32827 35009
rect 25832 34960 25838 34972
rect 32769 34969 32781 35003
rect 32815 35000 32827 35003
rect 32858 35000 32864 35012
rect 32815 34972 32864 35000
rect 32815 34969 32827 34972
rect 32769 34963 32827 34969
rect 32858 34960 32864 34972
rect 32916 35000 32922 35012
rect 34072 35000 34100 35031
rect 35618 35028 35624 35040
rect 35676 35028 35682 35080
rect 38151 35071 38209 35077
rect 38151 35037 38163 35071
rect 38197 35068 38209 35071
rect 39114 35068 39120 35080
rect 38197 35040 39120 35068
rect 38197 35037 38209 35040
rect 38151 35031 38209 35037
rect 39114 35028 39120 35040
rect 39172 35028 39178 35080
rect 40727 35071 40785 35077
rect 40727 35037 40739 35071
rect 40773 35068 40785 35071
rect 40862 35068 40868 35080
rect 40773 35040 40868 35068
rect 40773 35037 40785 35040
rect 40727 35031 40785 35037
rect 40862 35028 40868 35040
rect 40920 35028 40926 35080
rect 41782 35068 41788 35080
rect 41743 35040 41788 35068
rect 41782 35028 41788 35040
rect 41840 35028 41846 35080
rect 42429 35071 42487 35077
rect 42429 35037 42441 35071
rect 42475 35068 42487 35071
rect 42886 35068 42892 35080
rect 42475 35040 42892 35068
rect 42475 35037 42487 35040
rect 42429 35031 42487 35037
rect 42886 35028 42892 35040
rect 42944 35028 42950 35080
rect 38838 35000 38844 35012
rect 32916 34972 34100 35000
rect 38751 34972 38844 35000
rect 32916 34960 32922 34972
rect 38838 34960 38844 34972
rect 38896 35000 38902 35012
rect 39669 35003 39727 35009
rect 39669 35000 39681 35003
rect 38896 34972 39681 35000
rect 38896 34960 38902 34972
rect 39669 34969 39681 34972
rect 39715 35000 39727 35003
rect 41138 35000 41144 35012
rect 39715 34972 41144 35000
rect 39715 34969 39727 34972
rect 39669 34963 39727 34969
rect 41138 34960 41144 34972
rect 41196 34960 41202 35012
rect 7190 34892 7196 34944
rect 7248 34932 7254 34944
rect 7285 34935 7343 34941
rect 7285 34932 7297 34935
rect 7248 34904 7297 34932
rect 7248 34892 7254 34904
rect 7285 34901 7297 34904
rect 7331 34901 7343 34935
rect 8846 34932 8852 34944
rect 8807 34904 8852 34932
rect 7285 34895 7343 34901
rect 8846 34892 8852 34904
rect 8904 34892 8910 34944
rect 10870 34932 10876 34944
rect 10831 34904 10876 34932
rect 10870 34892 10876 34904
rect 10928 34892 10934 34944
rect 16206 34892 16212 34944
rect 16264 34932 16270 34944
rect 17083 34935 17141 34941
rect 17083 34932 17095 34935
rect 16264 34904 17095 34932
rect 16264 34892 16270 34904
rect 17083 34901 17095 34904
rect 17129 34901 17141 34935
rect 17083 34895 17141 34901
rect 17402 34892 17408 34944
rect 17460 34932 17466 34944
rect 17589 34935 17647 34941
rect 17589 34932 17601 34935
rect 17460 34904 17601 34932
rect 17460 34892 17466 34904
rect 17589 34901 17601 34904
rect 17635 34901 17647 34935
rect 17589 34895 17647 34901
rect 18141 34935 18199 34941
rect 18141 34901 18153 34935
rect 18187 34932 18199 34935
rect 18506 34932 18512 34944
rect 18187 34904 18512 34932
rect 18187 34901 18199 34904
rect 18141 34895 18199 34901
rect 18506 34892 18512 34904
rect 18564 34892 18570 34944
rect 23750 34932 23756 34944
rect 23711 34904 23756 34932
rect 23750 34892 23756 34904
rect 23808 34892 23814 34944
rect 26326 34932 26332 34944
rect 26287 34904 26332 34932
rect 26326 34892 26332 34904
rect 26384 34892 26390 34944
rect 28491 34935 28549 34941
rect 28491 34901 28503 34935
rect 28537 34932 28549 34935
rect 30006 34932 30012 34944
rect 28537 34904 30012 34932
rect 28537 34901 28549 34904
rect 28491 34895 28549 34901
rect 30006 34892 30012 34904
rect 30064 34892 30070 34944
rect 33318 34932 33324 34944
rect 33231 34904 33324 34932
rect 33318 34892 33324 34904
rect 33376 34932 33382 34944
rect 33962 34932 33968 34944
rect 33376 34904 33968 34932
rect 33376 34892 33382 34904
rect 33962 34892 33968 34904
rect 34020 34892 34026 34944
rect 36078 34892 36084 34944
rect 36136 34932 36142 34944
rect 36265 34935 36323 34941
rect 36265 34932 36277 34935
rect 36136 34904 36277 34932
rect 36136 34892 36142 34904
rect 36265 34901 36277 34904
rect 36311 34901 36323 34935
rect 36265 34895 36323 34901
rect 42518 34892 42524 34944
rect 42576 34932 42582 34944
rect 42797 34935 42855 34941
rect 42797 34932 42809 34935
rect 42576 34904 42809 34932
rect 42576 34892 42582 34904
rect 42797 34901 42809 34904
rect 42843 34932 42855 34935
rect 43487 34935 43545 34941
rect 43487 34932 43499 34935
rect 42843 34904 43499 34932
rect 42843 34901 42855 34904
rect 42797 34895 42855 34901
rect 43487 34901 43499 34904
rect 43533 34901 43545 34935
rect 43487 34895 43545 34901
rect 1104 34842 48852 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 48852 34842
rect 1104 34768 48852 34790
rect 7331 34731 7389 34737
rect 7331 34697 7343 34731
rect 7377 34728 7389 34731
rect 8202 34728 8208 34740
rect 7377 34700 8208 34728
rect 7377 34697 7389 34700
rect 7331 34691 7389 34697
rect 8202 34688 8208 34700
rect 8260 34688 8266 34740
rect 9306 34728 9312 34740
rect 9267 34700 9312 34728
rect 9306 34688 9312 34700
rect 9364 34688 9370 34740
rect 10870 34688 10876 34740
rect 10928 34728 10934 34740
rect 11471 34731 11529 34737
rect 11471 34728 11483 34731
rect 10928 34700 11483 34728
rect 10928 34688 10934 34700
rect 11471 34697 11483 34700
rect 11517 34697 11529 34731
rect 11471 34691 11529 34697
rect 12894 34688 12900 34740
rect 12952 34728 12958 34740
rect 14645 34731 14703 34737
rect 14645 34728 14657 34731
rect 12952 34700 14657 34728
rect 12952 34688 12958 34700
rect 14645 34697 14657 34700
rect 14691 34697 14703 34731
rect 14645 34691 14703 34697
rect 10410 34660 10416 34672
rect 10371 34632 10416 34660
rect 10410 34620 10416 34632
rect 10468 34620 10474 34672
rect 11146 34660 11152 34672
rect 11107 34632 11152 34660
rect 11146 34620 11152 34632
rect 11204 34620 11210 34672
rect 3559 34595 3617 34601
rect 3559 34561 3571 34595
rect 3605 34592 3617 34595
rect 7009 34595 7067 34601
rect 7009 34592 7021 34595
rect 3605 34564 7021 34592
rect 3605 34561 3617 34564
rect 3559 34555 3617 34561
rect 7009 34561 7021 34564
rect 7055 34592 7067 34595
rect 7926 34592 7932 34604
rect 7055 34564 7932 34592
rect 7055 34561 7067 34564
rect 7009 34555 7067 34561
rect 7926 34552 7932 34564
rect 7984 34552 7990 34604
rect 8297 34595 8355 34601
rect 8297 34561 8309 34595
rect 8343 34592 8355 34595
rect 8754 34592 8760 34604
rect 8343 34564 8760 34592
rect 8343 34561 8355 34564
rect 8297 34555 8355 34561
rect 8754 34552 8760 34564
rect 8812 34552 8818 34604
rect 9490 34552 9496 34604
rect 9548 34592 9554 34604
rect 9861 34595 9919 34601
rect 9861 34592 9873 34595
rect 9548 34564 9873 34592
rect 9548 34552 9554 34564
rect 9861 34561 9873 34564
rect 9907 34592 9919 34595
rect 10781 34595 10839 34601
rect 10781 34592 10793 34595
rect 9907 34564 10793 34592
rect 9907 34561 9919 34564
rect 9861 34555 9919 34561
rect 10781 34561 10793 34564
rect 10827 34561 10839 34595
rect 10781 34555 10839 34561
rect 13265 34595 13323 34601
rect 13265 34561 13277 34595
rect 13311 34592 13323 34595
rect 13630 34592 13636 34604
rect 13311 34564 13636 34592
rect 13311 34561 13323 34564
rect 13265 34555 13323 34561
rect 13630 34552 13636 34564
rect 13688 34552 13694 34604
rect 14660 34592 14688 34691
rect 15286 34688 15292 34740
rect 15344 34728 15350 34740
rect 15381 34731 15439 34737
rect 15381 34728 15393 34731
rect 15344 34700 15393 34728
rect 15344 34688 15350 34700
rect 15381 34697 15393 34700
rect 15427 34697 15439 34731
rect 16574 34728 16580 34740
rect 16535 34700 16580 34728
rect 15381 34691 15439 34697
rect 16574 34688 16580 34700
rect 16632 34688 16638 34740
rect 17037 34731 17095 34737
rect 17037 34697 17049 34731
rect 17083 34728 17095 34731
rect 17218 34728 17224 34740
rect 17083 34700 17224 34728
rect 17083 34697 17095 34700
rect 17037 34691 17095 34697
rect 17218 34688 17224 34700
rect 17276 34688 17282 34740
rect 20254 34728 20260 34740
rect 20215 34700 20260 34728
rect 20254 34688 20260 34700
rect 20312 34688 20318 34740
rect 21266 34728 21272 34740
rect 21179 34700 21272 34728
rect 21266 34688 21272 34700
rect 21324 34728 21330 34740
rect 22830 34728 22836 34740
rect 21324 34700 22508 34728
rect 22791 34700 22836 34728
rect 21324 34688 21330 34700
rect 15105 34663 15163 34669
rect 15105 34629 15117 34663
rect 15151 34660 15163 34663
rect 15562 34660 15568 34672
rect 15151 34632 15568 34660
rect 15151 34629 15163 34632
rect 15105 34623 15163 34629
rect 15562 34620 15568 34632
rect 15620 34620 15626 34672
rect 19150 34660 19156 34672
rect 19063 34632 19156 34660
rect 19150 34620 19156 34632
rect 19208 34660 19214 34672
rect 21284 34660 21312 34688
rect 19208 34632 21312 34660
rect 19208 34620 19214 34632
rect 22002 34620 22008 34672
rect 22060 34660 22066 34672
rect 22373 34663 22431 34669
rect 22373 34660 22385 34663
rect 22060 34632 22385 34660
rect 22060 34620 22066 34632
rect 22373 34629 22385 34632
rect 22419 34629 22431 34663
rect 22480 34660 22508 34700
rect 22830 34688 22836 34700
rect 22888 34688 22894 34740
rect 24302 34688 24308 34740
rect 24360 34728 24366 34740
rect 24581 34731 24639 34737
rect 24581 34728 24593 34731
rect 24360 34700 24593 34728
rect 24360 34688 24366 34700
rect 24581 34697 24593 34700
rect 24627 34728 24639 34731
rect 24857 34731 24915 34737
rect 24857 34728 24869 34731
rect 24627 34700 24869 34728
rect 24627 34697 24639 34700
rect 24581 34691 24639 34697
rect 24857 34697 24869 34700
rect 24903 34697 24915 34731
rect 28307 34731 28365 34737
rect 28307 34728 28319 34731
rect 24857 34691 24915 34697
rect 25562 34700 28319 34728
rect 23290 34660 23296 34672
rect 22480 34632 23296 34660
rect 22373 34623 22431 34629
rect 23290 34620 23296 34632
rect 23348 34660 23354 34672
rect 23477 34663 23535 34669
rect 23477 34660 23489 34663
rect 23348 34632 23489 34660
rect 23348 34620 23354 34632
rect 23477 34629 23489 34632
rect 23523 34660 23535 34663
rect 23842 34660 23848 34672
rect 23523 34632 23848 34660
rect 23523 34629 23535 34632
rect 23477 34623 23535 34629
rect 23842 34620 23848 34632
rect 23900 34620 23906 34672
rect 24026 34620 24032 34672
rect 24084 34660 24090 34672
rect 25562 34660 25590 34700
rect 28307 34697 28319 34700
rect 28353 34697 28365 34731
rect 28307 34691 28365 34697
rect 29362 34688 29368 34740
rect 29420 34728 29426 34740
rect 30101 34731 30159 34737
rect 30101 34728 30113 34731
rect 29420 34700 30113 34728
rect 29420 34688 29426 34700
rect 30101 34697 30113 34700
rect 30147 34697 30159 34731
rect 30101 34691 30159 34697
rect 31665 34731 31723 34737
rect 31665 34697 31677 34731
rect 31711 34728 31723 34731
rect 31846 34728 31852 34740
rect 31711 34700 31852 34728
rect 31711 34697 31723 34700
rect 31665 34691 31723 34697
rect 31846 34688 31852 34700
rect 31904 34728 31910 34740
rect 31941 34731 31999 34737
rect 31941 34728 31953 34731
rect 31904 34700 31953 34728
rect 31904 34688 31910 34700
rect 31941 34697 31953 34700
rect 31987 34697 31999 34731
rect 31941 34691 31999 34697
rect 33597 34731 33655 34737
rect 33597 34697 33609 34731
rect 33643 34728 33655 34731
rect 33778 34728 33784 34740
rect 33643 34700 33784 34728
rect 33643 34697 33655 34700
rect 33597 34691 33655 34697
rect 33778 34688 33784 34700
rect 33836 34737 33842 34740
rect 33836 34731 33885 34737
rect 33836 34697 33839 34731
rect 33873 34697 33885 34731
rect 33836 34691 33885 34697
rect 33836 34688 33842 34691
rect 33962 34688 33968 34740
rect 34020 34728 34026 34740
rect 35023 34731 35081 34737
rect 35023 34728 35035 34731
rect 34020 34700 35035 34728
rect 34020 34688 34026 34700
rect 35023 34697 35035 34700
rect 35069 34697 35081 34731
rect 35023 34691 35081 34697
rect 35342 34688 35348 34740
rect 35400 34728 35406 34740
rect 36081 34731 36139 34737
rect 36081 34728 36093 34731
rect 35400 34700 36093 34728
rect 35400 34688 35406 34700
rect 36081 34697 36093 34700
rect 36127 34697 36139 34731
rect 36081 34691 36139 34697
rect 36909 34731 36967 34737
rect 36909 34697 36921 34731
rect 36955 34728 36967 34731
rect 36998 34728 37004 34740
rect 36955 34700 37004 34728
rect 36955 34697 36967 34700
rect 36909 34691 36967 34697
rect 36998 34688 37004 34700
rect 37056 34688 37062 34740
rect 39206 34688 39212 34740
rect 39264 34728 39270 34740
rect 39761 34731 39819 34737
rect 39761 34728 39773 34731
rect 39264 34700 39773 34728
rect 39264 34688 39270 34700
rect 39761 34697 39773 34700
rect 39807 34697 39819 34731
rect 41414 34728 41420 34740
rect 41375 34700 41420 34728
rect 39761 34691 39819 34697
rect 41414 34688 41420 34700
rect 41472 34688 41478 34740
rect 41785 34731 41843 34737
rect 41785 34697 41797 34731
rect 41831 34728 41843 34731
rect 41874 34728 41880 34740
rect 41831 34700 41880 34728
rect 41831 34697 41843 34700
rect 41785 34691 41843 34697
rect 41874 34688 41880 34700
rect 41932 34728 41938 34740
rect 42245 34731 42303 34737
rect 42245 34728 42257 34731
rect 41932 34700 42257 34728
rect 41932 34688 41938 34700
rect 42245 34697 42257 34700
rect 42291 34697 42303 34731
rect 42245 34691 42303 34697
rect 24084 34632 25590 34660
rect 25731 34663 25789 34669
rect 24084 34620 24090 34632
rect 25731 34629 25743 34663
rect 25777 34660 25789 34663
rect 26602 34660 26608 34672
rect 25777 34632 26608 34660
rect 25777 34629 25789 34632
rect 25731 34623 25789 34629
rect 26602 34620 26608 34632
rect 26660 34620 26666 34672
rect 27246 34660 27252 34672
rect 27207 34632 27252 34660
rect 27246 34620 27252 34632
rect 27304 34620 27310 34672
rect 29089 34663 29147 34669
rect 29089 34629 29101 34663
rect 29135 34660 29147 34663
rect 29546 34660 29552 34672
rect 29135 34632 29552 34660
rect 29135 34629 29147 34632
rect 29089 34623 29147 34629
rect 29546 34620 29552 34632
rect 29604 34620 29610 34672
rect 29730 34660 29736 34672
rect 29691 34632 29736 34660
rect 29730 34620 29736 34632
rect 29788 34620 29794 34672
rect 32674 34660 32680 34672
rect 32140 34632 32680 34660
rect 15657 34595 15715 34601
rect 15657 34592 15669 34595
rect 14660 34564 15669 34592
rect 15657 34561 15669 34564
rect 15703 34561 15715 34595
rect 16022 34592 16028 34604
rect 15983 34564 16028 34592
rect 15657 34555 15715 34561
rect 16022 34552 16028 34564
rect 16080 34552 16086 34604
rect 18414 34552 18420 34604
rect 18472 34592 18478 34604
rect 18601 34595 18659 34601
rect 18601 34592 18613 34595
rect 18472 34564 18613 34592
rect 18472 34552 18478 34564
rect 18601 34561 18613 34564
rect 18647 34561 18659 34595
rect 18601 34555 18659 34561
rect 19843 34595 19901 34601
rect 19843 34561 19855 34595
rect 19889 34592 19901 34595
rect 24210 34592 24216 34604
rect 19889 34564 24216 34592
rect 19889 34561 19901 34564
rect 19843 34555 19901 34561
rect 24210 34552 24216 34564
rect 24268 34552 24274 34604
rect 25866 34552 25872 34604
rect 25924 34592 25930 34604
rect 26697 34595 26755 34601
rect 26697 34592 26709 34595
rect 25924 34564 26709 34592
rect 25924 34552 25930 34564
rect 26697 34561 26709 34564
rect 26743 34592 26755 34595
rect 27985 34595 28043 34601
rect 27985 34592 27997 34595
rect 26743 34564 27997 34592
rect 26743 34561 26755 34564
rect 26697 34555 26755 34561
rect 27985 34561 27997 34564
rect 28031 34561 28043 34595
rect 27985 34555 28043 34561
rect 30006 34552 30012 34604
rect 30064 34592 30070 34604
rect 30377 34595 30435 34601
rect 30377 34592 30389 34595
rect 30064 34564 30389 34592
rect 30064 34552 30070 34564
rect 30377 34561 30389 34564
rect 30423 34592 30435 34595
rect 30834 34592 30840 34604
rect 30423 34564 30840 34592
rect 30423 34561 30435 34564
rect 30377 34555 30435 34561
rect 30834 34552 30840 34564
rect 30892 34552 30898 34604
rect 31018 34592 31024 34604
rect 30979 34564 31024 34592
rect 31018 34552 31024 34564
rect 31076 34552 31082 34604
rect 32140 34592 32168 34632
rect 32674 34620 32680 34632
rect 32732 34620 32738 34672
rect 32769 34663 32827 34669
rect 32769 34629 32781 34663
rect 32815 34660 32827 34663
rect 32950 34660 32956 34672
rect 32815 34632 32956 34660
rect 32815 34629 32827 34632
rect 32769 34623 32827 34629
rect 32950 34620 32956 34632
rect 33008 34660 33014 34672
rect 35618 34660 35624 34672
rect 33008 34632 35624 34660
rect 33008 34620 33014 34632
rect 35618 34620 35624 34632
rect 35676 34620 35682 34672
rect 35710 34620 35716 34672
rect 35768 34660 35774 34672
rect 40586 34660 40592 34672
rect 35768 34632 35813 34660
rect 36464 34632 40592 34660
rect 35768 34620 35774 34632
rect 32048 34564 32168 34592
rect 3326 34524 3332 34536
rect 3287 34496 3332 34524
rect 3326 34484 3332 34496
rect 3384 34524 3390 34536
rect 3456 34527 3514 34533
rect 3456 34524 3468 34527
rect 3384 34496 3468 34524
rect 3384 34484 3390 34496
rect 3456 34493 3468 34496
rect 3502 34493 3514 34527
rect 3456 34487 3514 34493
rect 4433 34527 4491 34533
rect 4433 34493 4445 34527
rect 4479 34524 4491 34527
rect 4890 34524 4896 34536
rect 4479 34496 4896 34524
rect 4479 34493 4491 34496
rect 4433 34487 4491 34493
rect 4890 34484 4896 34496
rect 4948 34524 4954 34536
rect 5629 34527 5687 34533
rect 5629 34524 5641 34527
rect 4948 34496 5641 34524
rect 4948 34484 4954 34496
rect 5629 34493 5641 34496
rect 5675 34493 5687 34527
rect 5629 34487 5687 34493
rect 7193 34527 7251 34533
rect 7193 34493 7205 34527
rect 7239 34524 7251 34527
rect 7282 34524 7288 34536
rect 7239 34496 7288 34524
rect 7239 34493 7251 34496
rect 7193 34487 7251 34493
rect 7282 34484 7288 34496
rect 7340 34484 7346 34536
rect 11400 34527 11458 34533
rect 11400 34493 11412 34527
rect 11446 34524 11458 34527
rect 12161 34527 12219 34533
rect 12161 34524 12173 34527
rect 11446 34496 12173 34524
rect 11446 34493 11458 34496
rect 11400 34487 11458 34493
rect 12161 34493 12173 34496
rect 12207 34524 12219 34527
rect 12250 34524 12256 34536
rect 12207 34496 12256 34524
rect 12207 34493 12219 34496
rect 12161 34487 12219 34493
rect 12250 34484 12256 34496
rect 12308 34484 12314 34536
rect 17865 34527 17923 34533
rect 17865 34493 17877 34527
rect 17911 34524 17923 34527
rect 18230 34524 18236 34536
rect 17911 34496 18236 34524
rect 17911 34493 17923 34496
rect 17865 34487 17923 34493
rect 18230 34484 18236 34496
rect 18288 34484 18294 34536
rect 18506 34524 18512 34536
rect 18467 34496 18512 34524
rect 18506 34484 18512 34496
rect 18564 34484 18570 34536
rect 19756 34527 19814 34533
rect 19756 34493 19768 34527
rect 19802 34524 19814 34527
rect 20254 34524 20260 34536
rect 19802 34496 20260 34524
rect 19802 34493 19814 34496
rect 19756 34487 19814 34493
rect 20254 34484 20260 34496
rect 20312 34484 20318 34536
rect 20784 34527 20842 34533
rect 20784 34493 20796 34527
rect 20830 34524 20842 34527
rect 23661 34527 23719 34533
rect 20830 34496 21680 34524
rect 20830 34493 20842 34496
rect 20784 34487 20842 34493
rect 8389 34459 8447 34465
rect 4816 34428 6132 34456
rect 3973 34391 4031 34397
rect 3973 34357 3985 34391
rect 4019 34388 4031 34391
rect 4341 34391 4399 34397
rect 4341 34388 4353 34391
rect 4019 34360 4353 34388
rect 4019 34357 4031 34360
rect 3973 34351 4031 34357
rect 4341 34357 4353 34360
rect 4387 34388 4399 34391
rect 4706 34388 4712 34400
rect 4387 34360 4712 34388
rect 4387 34357 4399 34360
rect 4341 34351 4399 34357
rect 4706 34348 4712 34360
rect 4764 34388 4770 34400
rect 4816 34397 4844 34428
rect 6104 34400 6132 34428
rect 8389 34425 8401 34459
rect 8435 34425 8447 34459
rect 8389 34419 8447 34425
rect 8941 34459 8999 34465
rect 8941 34425 8953 34459
rect 8987 34456 8999 34459
rect 9858 34456 9864 34468
rect 8987 34428 9864 34456
rect 8987 34425 8999 34428
rect 8941 34419 8999 34425
rect 4801 34391 4859 34397
rect 4801 34388 4813 34391
rect 4764 34360 4813 34388
rect 4764 34348 4770 34360
rect 4801 34357 4813 34360
rect 4847 34357 4859 34391
rect 5350 34388 5356 34400
rect 5311 34360 5356 34388
rect 4801 34351 4859 34357
rect 5350 34348 5356 34360
rect 5408 34348 5414 34400
rect 6086 34388 6092 34400
rect 6047 34360 6092 34388
rect 6086 34348 6092 34360
rect 6144 34348 6150 34400
rect 6454 34388 6460 34400
rect 6415 34360 6460 34388
rect 6454 34348 6460 34360
rect 6512 34348 6518 34400
rect 7834 34348 7840 34400
rect 7892 34388 7898 34400
rect 7929 34391 7987 34397
rect 7929 34388 7941 34391
rect 7892 34360 7941 34388
rect 7892 34348 7898 34360
rect 7929 34357 7941 34360
rect 7975 34388 7987 34391
rect 8294 34388 8300 34400
rect 7975 34360 8300 34388
rect 7975 34357 7987 34360
rect 7929 34351 7987 34357
rect 8294 34348 8300 34360
rect 8352 34388 8358 34400
rect 8404 34388 8432 34419
rect 9858 34416 9864 34428
rect 9916 34416 9922 34468
rect 9953 34459 10011 34465
rect 9953 34425 9965 34459
rect 9999 34456 10011 34459
rect 11790 34456 11796 34468
rect 9999 34428 11796 34456
rect 9999 34425 10011 34428
rect 9953 34419 10011 34425
rect 9677 34391 9735 34397
rect 9677 34388 9689 34391
rect 8352 34360 9689 34388
rect 8352 34348 8358 34360
rect 9677 34357 9689 34360
rect 9723 34388 9735 34391
rect 9968 34388 9996 34419
rect 11790 34416 11796 34428
rect 11848 34416 11854 34468
rect 12805 34459 12863 34465
rect 12805 34425 12817 34459
rect 12851 34456 12863 34459
rect 13078 34456 13084 34468
rect 12851 34428 13084 34456
rect 12851 34425 12863 34428
rect 12805 34419 12863 34425
rect 13078 34416 13084 34428
rect 13136 34456 13142 34468
rect 13173 34459 13231 34465
rect 13173 34456 13185 34459
rect 13136 34428 13185 34456
rect 13136 34416 13142 34428
rect 13173 34425 13185 34428
rect 13219 34456 13231 34459
rect 13627 34459 13685 34465
rect 13627 34456 13639 34459
rect 13219 34428 13639 34456
rect 13219 34425 13231 34428
rect 13173 34419 13231 34425
rect 13627 34425 13639 34428
rect 13673 34456 13685 34459
rect 13722 34456 13728 34468
rect 13673 34428 13728 34456
rect 13673 34425 13685 34428
rect 13627 34419 13685 34425
rect 13722 34416 13728 34428
rect 13780 34416 13786 34468
rect 15286 34416 15292 34468
rect 15344 34456 15350 34468
rect 15749 34459 15807 34465
rect 15749 34456 15761 34459
rect 15344 34428 15761 34456
rect 15344 34416 15350 34428
rect 15749 34425 15761 34428
rect 15795 34425 15807 34459
rect 15749 34419 15807 34425
rect 20070 34416 20076 34468
rect 20128 34456 20134 34468
rect 20530 34456 20536 34468
rect 20128 34428 20536 34456
rect 20128 34416 20134 34428
rect 20530 34416 20536 34428
rect 20588 34416 20594 34468
rect 11882 34388 11888 34400
rect 9723 34360 9996 34388
rect 11795 34360 11888 34388
rect 9723 34357 9735 34360
rect 9677 34351 9735 34357
rect 11882 34348 11888 34360
rect 11940 34388 11946 34400
rect 12342 34388 12348 34400
rect 11940 34360 12348 34388
rect 11940 34348 11946 34360
rect 12342 34348 12348 34360
rect 12400 34348 12406 34400
rect 14182 34388 14188 34400
rect 14143 34360 14188 34388
rect 14182 34348 14188 34360
rect 14240 34348 14246 34400
rect 20855 34391 20913 34397
rect 20855 34357 20867 34391
rect 20901 34388 20913 34391
rect 21082 34388 21088 34400
rect 20901 34360 21088 34388
rect 20901 34357 20913 34360
rect 20855 34351 20913 34357
rect 21082 34348 21088 34360
rect 21140 34348 21146 34400
rect 21652 34397 21680 34496
rect 23661 34493 23673 34527
rect 23707 34524 23719 34527
rect 23750 34524 23756 34536
rect 23707 34496 23756 34524
rect 23707 34493 23719 34496
rect 23661 34487 23719 34493
rect 23750 34484 23756 34496
rect 23808 34484 23814 34536
rect 25660 34527 25718 34533
rect 25660 34493 25672 34527
rect 25706 34524 25718 34527
rect 26142 34524 26148 34536
rect 25706 34496 26148 34524
rect 25706 34493 25718 34496
rect 25660 34487 25718 34493
rect 26142 34484 26148 34496
rect 26200 34484 26206 34536
rect 28236 34527 28294 34533
rect 28236 34493 28248 34527
rect 28282 34524 28294 34527
rect 29340 34527 29398 34533
rect 28282 34496 28764 34524
rect 28282 34493 28294 34496
rect 28236 34487 28294 34493
rect 21818 34456 21824 34468
rect 21779 34428 21824 34456
rect 21818 34416 21824 34428
rect 21876 34416 21882 34468
rect 21910 34416 21916 34468
rect 21968 34456 21974 34468
rect 21968 34428 22013 34456
rect 22572 34428 23704 34456
rect 21968 34416 21974 34428
rect 21637 34391 21695 34397
rect 21637 34357 21649 34391
rect 21683 34388 21695 34391
rect 22572 34388 22600 34428
rect 21683 34360 22600 34388
rect 23676 34388 23704 34428
rect 23842 34416 23848 34468
rect 23900 34456 23906 34468
rect 23982 34459 24040 34465
rect 23982 34456 23994 34459
rect 23900 34428 23994 34456
rect 23900 34416 23906 34428
rect 23982 34425 23994 34428
rect 24028 34425 24040 34459
rect 23982 34419 24040 34425
rect 26789 34459 26847 34465
rect 26789 34425 26801 34459
rect 26835 34456 26847 34459
rect 26878 34456 26884 34468
rect 26835 34428 26884 34456
rect 26835 34425 26847 34428
rect 26789 34419 26847 34425
rect 26878 34416 26884 34428
rect 26936 34416 26942 34468
rect 25590 34388 25596 34400
rect 23676 34360 25596 34388
rect 21683 34357 21695 34360
rect 21637 34351 21695 34357
rect 25590 34348 25596 34360
rect 25648 34348 25654 34400
rect 26418 34388 26424 34400
rect 26379 34360 26424 34388
rect 26418 34348 26424 34360
rect 26476 34348 26482 34400
rect 26896 34388 26924 34416
rect 28736 34397 28764 34496
rect 29340 34493 29352 34527
rect 29386 34524 29398 34527
rect 29546 34524 29552 34536
rect 29386 34496 29552 34524
rect 29386 34493 29398 34496
rect 29340 34487 29398 34493
rect 29546 34484 29552 34496
rect 29604 34484 29610 34536
rect 30190 34416 30196 34468
rect 30248 34456 30254 34468
rect 30469 34459 30527 34465
rect 30469 34456 30481 34459
rect 30248 34428 30481 34456
rect 30248 34416 30254 34428
rect 30469 34425 30481 34428
rect 30515 34425 30527 34459
rect 32048 34456 32076 34564
rect 32214 34552 32220 34604
rect 32272 34592 32278 34604
rect 33137 34595 33195 34601
rect 33137 34592 33149 34595
rect 32272 34564 33149 34592
rect 32272 34552 32278 34564
rect 33137 34561 33149 34564
rect 33183 34561 33195 34595
rect 33137 34555 33195 34561
rect 34609 34595 34667 34601
rect 34609 34561 34621 34595
rect 34655 34592 34667 34595
rect 35728 34592 35756 34620
rect 34655 34564 35756 34592
rect 34655 34561 34667 34564
rect 34609 34555 34667 34561
rect 33756 34527 33814 34533
rect 33756 34493 33768 34527
rect 33802 34493 33814 34527
rect 33756 34487 33814 34493
rect 34952 34527 35010 34533
rect 34952 34493 34964 34527
rect 34998 34524 35010 34527
rect 35437 34527 35495 34533
rect 35437 34524 35449 34527
rect 34998 34496 35449 34524
rect 34998 34493 35010 34496
rect 34952 34487 35010 34493
rect 35437 34493 35449 34496
rect 35483 34524 35495 34527
rect 35526 34524 35532 34536
rect 35483 34496 35532 34524
rect 35483 34493 35495 34496
rect 35437 34487 35495 34493
rect 32217 34459 32275 34465
rect 32217 34456 32229 34459
rect 32048 34428 32229 34456
rect 30469 34419 30527 34425
rect 32217 34425 32229 34428
rect 32263 34425 32275 34459
rect 32217 34419 32275 34425
rect 32309 34459 32367 34465
rect 32309 34425 32321 34459
rect 32355 34425 32367 34459
rect 32309 34419 32367 34425
rect 27617 34391 27675 34397
rect 27617 34388 27629 34391
rect 26896 34360 27629 34388
rect 27617 34357 27629 34360
rect 27663 34357 27675 34391
rect 27617 34351 27675 34357
rect 28721 34391 28779 34397
rect 28721 34357 28733 34391
rect 28767 34388 28779 34391
rect 28902 34388 28908 34400
rect 28767 34360 28908 34388
rect 28767 34357 28779 34360
rect 28721 34351 28779 34357
rect 28902 34348 28908 34360
rect 28960 34348 28966 34400
rect 29178 34348 29184 34400
rect 29236 34388 29242 34400
rect 29411 34391 29469 34397
rect 29411 34388 29423 34391
rect 29236 34360 29423 34388
rect 29236 34348 29242 34360
rect 29411 34357 29423 34360
rect 29457 34357 29469 34391
rect 29411 34351 29469 34357
rect 31846 34348 31852 34400
rect 31904 34388 31910 34400
rect 32324 34388 32352 34419
rect 33594 34416 33600 34468
rect 33652 34456 33658 34468
rect 33771 34456 33799 34487
rect 35526 34484 35532 34496
rect 35584 34524 35590 34536
rect 36464 34524 36492 34632
rect 40586 34620 40592 34632
rect 40644 34660 40650 34672
rect 40957 34663 41015 34669
rect 40957 34660 40969 34663
rect 40644 34632 40969 34660
rect 40644 34620 40650 34632
rect 40957 34629 40969 34632
rect 41003 34629 41015 34663
rect 40957 34623 41015 34629
rect 38838 34592 38844 34604
rect 38799 34564 38844 34592
rect 38838 34552 38844 34564
rect 38896 34552 38902 34604
rect 38930 34552 38936 34604
rect 38988 34592 38994 34604
rect 38988 34564 39528 34592
rect 38988 34552 38994 34564
rect 35584 34496 36492 34524
rect 36541 34527 36599 34533
rect 35584 34484 35590 34496
rect 36541 34493 36553 34527
rect 36587 34524 36599 34527
rect 36814 34524 36820 34536
rect 36587 34496 36820 34524
rect 36587 34493 36599 34496
rect 36541 34487 36599 34493
rect 36814 34484 36820 34496
rect 36872 34524 36878 34536
rect 37001 34527 37059 34533
rect 37001 34524 37013 34527
rect 36872 34496 37013 34524
rect 36872 34484 36878 34496
rect 37001 34493 37013 34496
rect 37047 34493 37059 34527
rect 39500 34524 39528 34564
rect 40564 34527 40622 34533
rect 40564 34524 40576 34527
rect 37001 34487 37059 34493
rect 37108 34496 38654 34524
rect 39500 34496 40576 34524
rect 34241 34459 34299 34465
rect 34241 34456 34253 34459
rect 33652 34428 34253 34456
rect 33652 34416 33658 34428
rect 34241 34425 34253 34428
rect 34287 34456 34299 34459
rect 37108 34456 37136 34496
rect 34287 34428 37136 34456
rect 37363 34459 37421 34465
rect 34287 34425 34299 34428
rect 34241 34419 34299 34425
rect 37363 34425 37375 34459
rect 37409 34425 37421 34459
rect 38626 34456 38654 34496
rect 40564 34493 40576 34496
rect 40610 34524 40622 34527
rect 41414 34524 41420 34536
rect 40610 34496 41420 34524
rect 40610 34493 40622 34496
rect 40564 34487 40622 34493
rect 41414 34484 41420 34496
rect 41472 34484 41478 34536
rect 38838 34456 38844 34468
rect 38626 34428 38844 34456
rect 37363 34419 37421 34425
rect 31904 34360 32352 34388
rect 31904 34348 31910 34360
rect 36998 34348 37004 34400
rect 37056 34388 37062 34400
rect 37378 34388 37406 34419
rect 38838 34416 38844 34428
rect 38896 34416 38902 34468
rect 38933 34459 38991 34465
rect 38933 34425 38945 34459
rect 38979 34425 38991 34459
rect 39482 34456 39488 34468
rect 39443 34428 39488 34456
rect 38933 34419 38991 34425
rect 37918 34388 37924 34400
rect 37056 34360 37406 34388
rect 37879 34360 37924 34388
rect 37056 34348 37062 34360
rect 37918 34348 37924 34360
rect 37976 34348 37982 34400
rect 38194 34388 38200 34400
rect 38155 34360 38200 34388
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 38654 34388 38660 34400
rect 38615 34360 38660 34388
rect 38654 34348 38660 34360
rect 38712 34388 38718 34400
rect 38948 34388 38976 34419
rect 39482 34416 39488 34428
rect 39540 34416 39546 34468
rect 42260 34456 42288 34691
rect 42610 34688 42616 34740
rect 42668 34728 42674 34740
rect 43254 34728 43260 34740
rect 42668 34700 43260 34728
rect 42668 34688 42674 34700
rect 43254 34688 43260 34700
rect 43312 34728 43318 34740
rect 43441 34731 43499 34737
rect 43441 34728 43453 34731
rect 43312 34700 43453 34728
rect 43312 34688 43318 34700
rect 43441 34697 43453 34700
rect 43487 34697 43499 34731
rect 43441 34691 43499 34697
rect 42518 34592 42524 34604
rect 42479 34564 42524 34592
rect 42518 34552 42524 34564
rect 42576 34552 42582 34604
rect 42794 34552 42800 34604
rect 42852 34592 42858 34604
rect 42852 34564 42897 34592
rect 42852 34552 42858 34564
rect 42613 34459 42671 34465
rect 42613 34456 42625 34459
rect 42260 34428 42625 34456
rect 42613 34425 42625 34428
rect 42659 34456 42671 34459
rect 44358 34456 44364 34468
rect 42659 34428 44364 34456
rect 42659 34425 42671 34428
rect 42613 34419 42671 34425
rect 44358 34416 44364 34428
rect 44416 34416 44422 34468
rect 38712 34360 38976 34388
rect 40635 34391 40693 34397
rect 38712 34348 38718 34360
rect 40635 34357 40647 34391
rect 40681 34388 40693 34391
rect 40770 34388 40776 34400
rect 40681 34360 40776 34388
rect 40681 34357 40693 34360
rect 40635 34351 40693 34357
rect 40770 34348 40776 34360
rect 40828 34348 40834 34400
rect 1104 34298 48852 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 48852 34298
rect 1104 34224 48852 34246
rect 6135 34187 6193 34193
rect 6135 34153 6147 34187
rect 6181 34184 6193 34187
rect 7190 34184 7196 34196
rect 6181 34156 7196 34184
rect 6181 34153 6193 34156
rect 6135 34147 6193 34153
rect 7190 34144 7196 34156
rect 7248 34144 7254 34196
rect 7699 34187 7757 34193
rect 7699 34153 7711 34187
rect 7745 34184 7757 34187
rect 8570 34184 8576 34196
rect 7745 34156 8576 34184
rect 7745 34153 7757 34156
rect 7699 34147 7757 34153
rect 8570 34144 8576 34156
rect 8628 34144 8634 34196
rect 8711 34187 8769 34193
rect 8711 34153 8723 34187
rect 8757 34184 8769 34187
rect 8846 34184 8852 34196
rect 8757 34156 8852 34184
rect 8757 34153 8769 34156
rect 8711 34147 8769 34153
rect 8846 34144 8852 34156
rect 8904 34144 8910 34196
rect 12250 34184 12256 34196
rect 12211 34156 12256 34184
rect 12250 34144 12256 34156
rect 12308 34144 12314 34196
rect 13495 34187 13553 34193
rect 13495 34153 13507 34187
rect 13541 34184 13553 34187
rect 14550 34184 14556 34196
rect 13541 34156 14556 34184
rect 13541 34153 13553 34156
rect 13495 34147 13553 34153
rect 14550 34144 14556 34156
rect 14608 34144 14614 34196
rect 17402 34184 17408 34196
rect 17363 34156 17408 34184
rect 17402 34144 17408 34156
rect 17460 34144 17466 34196
rect 18414 34184 18420 34196
rect 18375 34156 18420 34184
rect 18414 34144 18420 34156
rect 18472 34144 18478 34196
rect 21818 34144 21824 34196
rect 21876 34184 21882 34196
rect 22603 34187 22661 34193
rect 22603 34184 22615 34187
rect 21876 34156 22615 34184
rect 21876 34144 21882 34156
rect 22603 34153 22615 34156
rect 22649 34153 22661 34187
rect 22603 34147 22661 34153
rect 23983 34187 24041 34193
rect 23983 34153 23995 34187
rect 24029 34184 24041 34187
rect 24118 34184 24124 34196
rect 24029 34156 24124 34184
rect 24029 34153 24041 34156
rect 23983 34147 24041 34153
rect 24118 34144 24124 34156
rect 24176 34144 24182 34196
rect 24210 34144 24216 34196
rect 24268 34184 24274 34196
rect 24305 34187 24363 34193
rect 24305 34184 24317 34187
rect 24268 34156 24317 34184
rect 24268 34144 24274 34156
rect 24305 34153 24317 34156
rect 24351 34153 24363 34187
rect 24305 34147 24363 34153
rect 25547 34187 25605 34193
rect 25547 34153 25559 34187
rect 25593 34184 25605 34187
rect 25866 34184 25872 34196
rect 25593 34156 25872 34184
rect 25593 34153 25605 34156
rect 25547 34147 25605 34153
rect 25866 34144 25872 34156
rect 25924 34144 25930 34196
rect 26329 34187 26387 34193
rect 26329 34153 26341 34187
rect 26375 34184 26387 34187
rect 26602 34184 26608 34196
rect 26375 34156 26608 34184
rect 26375 34153 26387 34156
rect 26329 34147 26387 34153
rect 26602 34144 26608 34156
rect 26660 34144 26666 34196
rect 26786 34144 26792 34196
rect 26844 34184 26850 34196
rect 29362 34184 29368 34196
rect 26844 34156 29368 34184
rect 26844 34144 26850 34156
rect 29362 34144 29368 34156
rect 29420 34144 29426 34196
rect 30834 34184 30840 34196
rect 30795 34156 30840 34184
rect 30834 34144 30840 34156
rect 30892 34144 30898 34196
rect 32214 34144 32220 34196
rect 32272 34184 32278 34196
rect 32401 34187 32459 34193
rect 32401 34184 32413 34187
rect 32272 34156 32413 34184
rect 32272 34144 32278 34156
rect 32401 34153 32413 34156
rect 32447 34153 32459 34187
rect 32674 34184 32680 34196
rect 32635 34156 32680 34184
rect 32401 34147 32459 34153
rect 32674 34144 32680 34156
rect 32732 34144 32738 34196
rect 32950 34184 32956 34196
rect 32911 34156 32956 34184
rect 32950 34144 32956 34156
rect 33008 34144 33014 34196
rect 34563 34187 34621 34193
rect 34563 34153 34575 34187
rect 34609 34184 34621 34187
rect 34790 34184 34796 34196
rect 34609 34156 34796 34184
rect 34609 34153 34621 34156
rect 34563 34147 34621 34153
rect 34790 34144 34796 34156
rect 34848 34144 34854 34196
rect 38654 34184 38660 34196
rect 38615 34156 38660 34184
rect 38654 34144 38660 34156
rect 38712 34144 38718 34196
rect 39114 34184 39120 34196
rect 39075 34156 39120 34184
rect 39114 34144 39120 34156
rect 39172 34144 39178 34196
rect 39390 34184 39396 34196
rect 39351 34156 39396 34184
rect 39390 34144 39396 34156
rect 39448 34144 39454 34196
rect 41782 34184 41788 34196
rect 41743 34156 41788 34184
rect 41782 34144 41788 34156
rect 41840 34144 41846 34196
rect 8294 34116 8300 34128
rect 8255 34088 8300 34116
rect 8294 34076 8300 34088
rect 8352 34076 8358 34128
rect 9306 34076 9312 34128
rect 9364 34116 9370 34128
rect 9582 34116 9588 34128
rect 9364 34088 9588 34116
rect 9364 34076 9370 34088
rect 9582 34076 9588 34088
rect 9640 34116 9646 34128
rect 9861 34119 9919 34125
rect 9861 34116 9873 34119
rect 9640 34088 9873 34116
rect 9640 34076 9646 34088
rect 9861 34085 9873 34088
rect 9907 34085 9919 34119
rect 9861 34079 9919 34085
rect 11695 34119 11753 34125
rect 11695 34085 11707 34119
rect 11741 34116 11753 34119
rect 11882 34116 11888 34128
rect 11741 34088 11888 34116
rect 11741 34085 11753 34088
rect 11695 34079 11753 34085
rect 11882 34076 11888 34088
rect 11940 34076 11946 34128
rect 15286 34076 15292 34128
rect 15344 34116 15350 34128
rect 15565 34119 15623 34125
rect 15565 34116 15577 34119
rect 15344 34088 15577 34116
rect 15344 34076 15350 34088
rect 15565 34085 15577 34088
rect 15611 34085 15623 34119
rect 19426 34116 19432 34128
rect 19387 34088 19432 34116
rect 15565 34079 15623 34085
rect 19426 34076 19432 34088
rect 19484 34076 19490 34128
rect 21085 34119 21143 34125
rect 21085 34085 21097 34119
rect 21131 34116 21143 34119
rect 21266 34116 21272 34128
rect 21131 34088 21272 34116
rect 21131 34085 21143 34088
rect 21085 34079 21143 34085
rect 21266 34076 21272 34088
rect 21324 34116 21330 34128
rect 21910 34116 21916 34128
rect 21324 34088 21916 34116
rect 21324 34076 21330 34088
rect 21910 34076 21916 34088
rect 21968 34076 21974 34128
rect 26878 34116 26884 34128
rect 26839 34088 26884 34116
rect 26878 34076 26884 34088
rect 26936 34076 26942 34128
rect 29270 34116 29276 34128
rect 29231 34088 29276 34116
rect 29270 34076 29276 34088
rect 29328 34076 29334 34128
rect 36814 34116 36820 34128
rect 36775 34088 36820 34116
rect 36814 34076 36820 34088
rect 36872 34076 36878 34128
rect 36998 34076 37004 34128
rect 37056 34116 37062 34128
rect 37826 34116 37832 34128
rect 37056 34088 37832 34116
rect 37056 34076 37062 34088
rect 37826 34076 37832 34088
rect 37884 34116 37890 34128
rect 38058 34119 38116 34125
rect 38058 34116 38070 34119
rect 37884 34088 38070 34116
rect 37884 34076 37890 34088
rect 38058 34085 38070 34088
rect 38104 34085 38116 34119
rect 40586 34116 40592 34128
rect 40547 34088 40592 34116
rect 38058 34079 38116 34085
rect 40586 34076 40592 34088
rect 40644 34076 40650 34128
rect 41138 34116 41144 34128
rect 41051 34088 41144 34116
rect 41138 34076 41144 34088
rect 41196 34116 41202 34128
rect 42794 34116 42800 34128
rect 41196 34088 42800 34116
rect 41196 34076 41202 34088
rect 42794 34076 42800 34088
rect 42852 34076 42858 34128
rect 43530 34116 43536 34128
rect 43491 34088 43536 34116
rect 43530 34076 43536 34088
rect 43588 34076 43594 34128
rect 4706 34048 4712 34060
rect 4667 34020 4712 34048
rect 4706 34008 4712 34020
rect 4764 34008 4770 34060
rect 4893 34051 4951 34057
rect 4893 34017 4905 34051
rect 4939 34048 4951 34051
rect 5166 34048 5172 34060
rect 4939 34020 5172 34048
rect 4939 34017 4951 34020
rect 4893 34011 4951 34017
rect 5166 34008 5172 34020
rect 5224 34008 5230 34060
rect 5350 34008 5356 34060
rect 5408 34048 5414 34060
rect 6032 34051 6090 34057
rect 6032 34048 6044 34051
rect 5408 34020 6044 34048
rect 5408 34008 5414 34020
rect 6032 34017 6044 34020
rect 6078 34048 6090 34051
rect 6178 34048 6184 34060
rect 6078 34020 6184 34048
rect 6078 34017 6090 34020
rect 6032 34011 6090 34017
rect 6178 34008 6184 34020
rect 6236 34008 6242 34060
rect 7628 34051 7686 34057
rect 7628 34017 7640 34051
rect 7674 34048 7686 34051
rect 8018 34048 8024 34060
rect 7674 34020 8024 34048
rect 7674 34017 7686 34020
rect 7628 34011 7686 34017
rect 8018 34008 8024 34020
rect 8076 34008 8082 34060
rect 8478 34008 8484 34060
rect 8536 34048 8542 34060
rect 8608 34051 8666 34057
rect 8608 34048 8620 34051
rect 8536 34020 8620 34048
rect 8536 34008 8542 34020
rect 8608 34017 8620 34020
rect 8654 34017 8666 34051
rect 8608 34011 8666 34017
rect 13424 34051 13482 34057
rect 13424 34017 13436 34051
rect 13470 34048 13482 34051
rect 14182 34048 14188 34060
rect 13470 34020 14188 34048
rect 13470 34017 13482 34020
rect 13424 34011 13482 34017
rect 14182 34008 14188 34020
rect 14240 34008 14246 34060
rect 16206 34048 16212 34060
rect 16167 34020 16212 34048
rect 16206 34008 16212 34020
rect 16264 34008 16270 34060
rect 17126 34048 17132 34060
rect 17087 34020 17132 34048
rect 17126 34008 17132 34020
rect 17184 34008 17190 34060
rect 17678 34048 17684 34060
rect 17639 34020 17684 34048
rect 17678 34008 17684 34020
rect 17736 34008 17742 34060
rect 21634 34008 21640 34060
rect 21692 34048 21698 34060
rect 21692 34020 21737 34048
rect 21692 34008 21698 34020
rect 22370 34008 22376 34060
rect 22428 34048 22434 34060
rect 22500 34051 22558 34057
rect 22500 34048 22512 34051
rect 22428 34020 22512 34048
rect 22428 34008 22434 34020
rect 22500 34017 22512 34020
rect 22546 34017 22558 34051
rect 22500 34011 22558 34017
rect 23106 34008 23112 34060
rect 23164 34048 23170 34060
rect 23880 34051 23938 34057
rect 23880 34048 23892 34051
rect 23164 34020 23892 34048
rect 23164 34008 23170 34020
rect 23880 34017 23892 34020
rect 23926 34048 23938 34051
rect 24670 34048 24676 34060
rect 23926 34020 24676 34048
rect 23926 34017 23938 34020
rect 23880 34011 23938 34017
rect 24670 34008 24676 34020
rect 24728 34008 24734 34060
rect 25406 34048 25412 34060
rect 25464 34057 25470 34060
rect 25464 34051 25502 34057
rect 24964 34020 25412 34048
rect 4982 33980 4988 33992
rect 4943 33952 4988 33980
rect 4982 33940 4988 33952
rect 5040 33940 5046 33992
rect 9766 33980 9772 33992
rect 9727 33952 9772 33980
rect 9766 33940 9772 33952
rect 9824 33940 9830 33992
rect 9858 33940 9864 33992
rect 9916 33980 9922 33992
rect 10045 33983 10103 33989
rect 10045 33980 10057 33983
rect 9916 33952 10057 33980
rect 9916 33940 9922 33952
rect 10045 33949 10057 33952
rect 10091 33949 10103 33983
rect 11330 33980 11336 33992
rect 11291 33952 11336 33980
rect 10045 33943 10103 33949
rect 11330 33940 11336 33952
rect 11388 33940 11394 33992
rect 19153 33983 19211 33989
rect 19153 33949 19165 33983
rect 19199 33980 19211 33983
rect 19334 33980 19340 33992
rect 19199 33952 19340 33980
rect 19199 33949 19211 33952
rect 19153 33943 19211 33949
rect 19334 33940 19340 33952
rect 19392 33940 19398 33992
rect 20990 33980 20996 33992
rect 20951 33952 20996 33980
rect 20990 33940 20996 33952
rect 21048 33940 21054 33992
rect 23014 33940 23020 33992
rect 23072 33980 23078 33992
rect 24964 33980 24992 34020
rect 25406 34008 25412 34020
rect 25490 34017 25502 34051
rect 28534 34048 28540 34060
rect 28495 34020 28540 34048
rect 25464 34011 25502 34017
rect 25464 34008 25470 34011
rect 28534 34008 28540 34020
rect 28592 34008 28598 34060
rect 28810 34008 28816 34060
rect 28868 34048 28874 34060
rect 29086 34048 29092 34060
rect 28868 34020 29092 34048
rect 28868 34008 28874 34020
rect 29086 34008 29092 34020
rect 29144 34008 29150 34060
rect 32033 34051 32091 34057
rect 32033 34017 32045 34051
rect 32079 34048 32091 34051
rect 32122 34048 32128 34060
rect 32079 34020 32128 34048
rect 32079 34017 32091 34020
rect 32033 34011 32091 34017
rect 32122 34008 32128 34020
rect 32180 34008 32186 34060
rect 33413 34051 33471 34057
rect 33413 34017 33425 34051
rect 33459 34048 33471 34051
rect 33502 34048 33508 34060
rect 33459 34020 33508 34048
rect 33459 34017 33471 34020
rect 33413 34011 33471 34017
rect 33502 34008 33508 34020
rect 33560 34008 33566 34060
rect 34422 34048 34428 34060
rect 34383 34020 34428 34048
rect 34422 34008 34428 34020
rect 34480 34008 34486 34060
rect 36354 34048 36360 34060
rect 36315 34020 36360 34048
rect 36354 34008 36360 34020
rect 36412 34008 36418 34060
rect 36538 34048 36544 34060
rect 36499 34020 36544 34048
rect 36538 34008 36544 34020
rect 36596 34008 36602 34060
rect 41230 34008 41236 34060
rect 41288 34048 41294 34060
rect 42242 34048 42248 34060
rect 42300 34057 42306 34060
rect 42300 34051 42338 34057
rect 41288 34020 42248 34048
rect 41288 34008 41294 34020
rect 42242 34008 42248 34020
rect 42326 34017 42338 34051
rect 42300 34011 42338 34017
rect 42300 34008 42306 34011
rect 26786 33980 26792 33992
rect 23072 33952 24992 33980
rect 26747 33952 26792 33980
rect 23072 33940 23078 33952
rect 26786 33940 26792 33952
rect 26844 33940 26850 33992
rect 27062 33980 27068 33992
rect 27023 33952 27068 33980
rect 27062 33940 27068 33952
rect 27120 33940 27126 33992
rect 30374 33980 30380 33992
rect 30335 33952 30380 33980
rect 30374 33940 30380 33952
rect 30432 33940 30438 33992
rect 37734 33980 37740 33992
rect 37695 33952 37740 33980
rect 37734 33940 37740 33952
rect 37792 33940 37798 33992
rect 40497 33983 40555 33989
rect 40497 33949 40509 33983
rect 40543 33980 40555 33983
rect 40862 33980 40868 33992
rect 40543 33952 40868 33980
rect 40543 33949 40555 33952
rect 40497 33943 40555 33949
rect 40862 33940 40868 33952
rect 40920 33980 40926 33992
rect 41506 33980 41512 33992
rect 40920 33952 41512 33980
rect 40920 33940 40926 33952
rect 41506 33940 41512 33952
rect 41564 33940 41570 33992
rect 42383 33983 42441 33989
rect 42383 33949 42395 33983
rect 42429 33980 42441 33983
rect 43070 33980 43076 33992
rect 42429 33952 43076 33980
rect 42429 33949 42441 33952
rect 42383 33943 42441 33949
rect 43070 33940 43076 33952
rect 43128 33980 43134 33992
rect 43441 33983 43499 33989
rect 43441 33980 43453 33983
rect 43128 33952 43453 33980
rect 43128 33940 43134 33952
rect 43441 33949 43453 33952
rect 43487 33949 43499 33983
rect 43441 33943 43499 33949
rect 43717 33983 43775 33989
rect 43717 33949 43729 33983
rect 43763 33949 43775 33983
rect 43717 33943 43775 33949
rect 19886 33912 19892 33924
rect 19847 33884 19892 33912
rect 19886 33872 19892 33884
rect 19944 33872 19950 33924
rect 42886 33872 42892 33924
rect 42944 33912 42950 33924
rect 43732 33912 43760 33943
rect 42944 33884 43760 33912
rect 42944 33872 42950 33884
rect 4062 33804 4068 33856
rect 4120 33844 4126 33856
rect 4249 33847 4307 33853
rect 4249 33844 4261 33847
rect 4120 33816 4261 33844
rect 4120 33804 4126 33816
rect 4249 33813 4261 33816
rect 4295 33813 4307 33847
rect 7282 33844 7288 33856
rect 7243 33816 7288 33844
rect 4249 33807 4307 33813
rect 7282 33804 7288 33816
rect 7340 33804 7346 33856
rect 12710 33804 12716 33856
rect 12768 33844 12774 33856
rect 12805 33847 12863 33853
rect 12805 33844 12817 33847
rect 12768 33816 12817 33844
rect 12768 33804 12774 33816
rect 12805 33813 12817 33816
rect 12851 33844 12863 33847
rect 13262 33844 13268 33856
rect 12851 33816 13268 33844
rect 12851 33813 12863 33816
rect 12805 33807 12863 33813
rect 13262 33804 13268 33816
rect 13320 33804 13326 33856
rect 13630 33804 13636 33856
rect 13688 33844 13694 33856
rect 13817 33847 13875 33853
rect 13817 33844 13829 33847
rect 13688 33816 13829 33844
rect 13688 33804 13694 33816
rect 13817 33813 13829 33816
rect 13863 33813 13875 33847
rect 13817 33807 13875 33813
rect 23753 33847 23811 33853
rect 23753 33813 23765 33847
rect 23799 33844 23811 33847
rect 23842 33844 23848 33856
rect 23799 33816 23848 33844
rect 23799 33813 23811 33816
rect 23753 33807 23811 33813
rect 23842 33804 23848 33816
rect 23900 33804 23906 33856
rect 29546 33844 29552 33856
rect 29507 33816 29552 33844
rect 29546 33804 29552 33816
rect 29604 33804 29610 33856
rect 31846 33804 31852 33856
rect 31904 33844 31910 33856
rect 33134 33844 33140 33856
rect 31904 33816 33140 33844
rect 31904 33804 31910 33816
rect 33134 33804 33140 33816
rect 33192 33804 33198 33856
rect 33551 33847 33609 33853
rect 33551 33813 33563 33847
rect 33597 33844 33609 33847
rect 35526 33844 35532 33856
rect 33597 33816 35532 33844
rect 33597 33813 33609 33816
rect 33551 33807 33609 33813
rect 35526 33804 35532 33816
rect 35584 33804 35590 33856
rect 42702 33844 42708 33856
rect 42663 33816 42708 33844
rect 42702 33804 42708 33816
rect 42760 33804 42766 33856
rect 1104 33754 48852 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 48852 33754
rect 1104 33680 48852 33702
rect 3326 33600 3332 33652
rect 3384 33640 3390 33652
rect 5905 33643 5963 33649
rect 5905 33640 5917 33643
rect 3384 33612 5917 33640
rect 3384 33600 3390 33612
rect 5905 33609 5917 33612
rect 5951 33609 5963 33643
rect 6178 33640 6184 33652
rect 6139 33612 6184 33640
rect 5905 33603 5963 33609
rect 6178 33600 6184 33612
rect 6236 33600 6242 33652
rect 7282 33600 7288 33652
rect 7340 33640 7346 33652
rect 7745 33643 7803 33649
rect 7745 33640 7757 33643
rect 7340 33612 7757 33640
rect 7340 33600 7346 33612
rect 7745 33609 7757 33612
rect 7791 33609 7803 33643
rect 8018 33640 8024 33652
rect 7979 33612 8024 33640
rect 7745 33603 7803 33609
rect 8018 33600 8024 33612
rect 8076 33640 8082 33652
rect 8386 33640 8392 33652
rect 8076 33612 8392 33640
rect 8076 33600 8082 33612
rect 8386 33600 8392 33612
rect 8444 33600 8450 33652
rect 9125 33643 9183 33649
rect 9125 33609 9137 33643
rect 9171 33640 9183 33643
rect 9766 33640 9772 33652
rect 9171 33612 9772 33640
rect 9171 33609 9183 33612
rect 9125 33603 9183 33609
rect 9766 33600 9772 33612
rect 9824 33640 9830 33652
rect 10367 33643 10425 33649
rect 10367 33640 10379 33643
rect 9824 33612 10379 33640
rect 9824 33600 9830 33612
rect 10367 33609 10379 33612
rect 10413 33609 10425 33643
rect 10367 33603 10425 33609
rect 11241 33643 11299 33649
rect 11241 33609 11253 33643
rect 11287 33640 11299 33643
rect 11330 33640 11336 33652
rect 11287 33612 11336 33640
rect 11287 33609 11299 33612
rect 11241 33603 11299 33609
rect 11330 33600 11336 33612
rect 11388 33600 11394 33652
rect 14001 33643 14059 33649
rect 14001 33609 14013 33643
rect 14047 33640 14059 33643
rect 14182 33640 14188 33652
rect 14047 33612 14188 33640
rect 14047 33609 14059 33612
rect 14001 33603 14059 33609
rect 14182 33600 14188 33612
rect 14240 33600 14246 33652
rect 15933 33643 15991 33649
rect 15933 33609 15945 33643
rect 15979 33640 15991 33643
rect 16206 33640 16212 33652
rect 15979 33612 16212 33640
rect 15979 33609 15991 33612
rect 15933 33603 15991 33609
rect 16206 33600 16212 33612
rect 16264 33600 16270 33652
rect 16574 33640 16580 33652
rect 16535 33612 16580 33640
rect 16574 33600 16580 33612
rect 16632 33600 16638 33652
rect 17126 33640 17132 33652
rect 17087 33612 17132 33640
rect 17126 33600 17132 33612
rect 17184 33600 17190 33652
rect 19426 33600 19432 33652
rect 19484 33640 19490 33652
rect 19521 33643 19579 33649
rect 19521 33640 19533 33643
rect 19484 33612 19533 33640
rect 19484 33600 19490 33612
rect 19521 33609 19533 33612
rect 19567 33640 19579 33643
rect 19797 33643 19855 33649
rect 19797 33640 19809 33643
rect 19567 33612 19809 33640
rect 19567 33609 19579 33612
rect 19521 33603 19579 33609
rect 19797 33609 19809 33612
rect 19843 33609 19855 33643
rect 19797 33603 19855 33609
rect 20257 33643 20315 33649
rect 20257 33609 20269 33643
rect 20303 33640 20315 33643
rect 20487 33643 20545 33649
rect 20487 33640 20499 33643
rect 20303 33612 20499 33640
rect 20303 33609 20315 33612
rect 20257 33603 20315 33609
rect 20487 33609 20499 33612
rect 20533 33640 20545 33643
rect 20990 33640 20996 33652
rect 20533 33612 20996 33640
rect 20533 33609 20545 33612
rect 20487 33603 20545 33609
rect 20990 33600 20996 33612
rect 21048 33600 21054 33652
rect 21266 33640 21272 33652
rect 21227 33612 21272 33640
rect 21266 33600 21272 33612
rect 21324 33600 21330 33652
rect 22370 33600 22376 33652
rect 22428 33640 22434 33652
rect 22465 33643 22523 33649
rect 22465 33640 22477 33643
rect 22428 33612 22477 33640
rect 22428 33600 22434 33612
rect 22465 33609 22477 33612
rect 22511 33609 22523 33643
rect 22465 33603 22523 33609
rect 24302 33600 24308 33652
rect 24360 33640 24366 33652
rect 24670 33640 24676 33652
rect 24360 33612 24676 33640
rect 24360 33600 24366 33612
rect 24670 33600 24676 33612
rect 24728 33600 24734 33652
rect 25406 33640 25412 33652
rect 25367 33612 25412 33640
rect 25406 33600 25412 33612
rect 25464 33600 25470 33652
rect 27522 33600 27528 33652
rect 27580 33640 27586 33652
rect 28307 33643 28365 33649
rect 28307 33640 28319 33643
rect 27580 33612 28319 33640
rect 27580 33600 27586 33612
rect 28307 33609 28319 33612
rect 28353 33609 28365 33643
rect 28307 33603 28365 33609
rect 28534 33600 28540 33652
rect 28592 33640 28598 33652
rect 28997 33643 29055 33649
rect 28997 33640 29009 33643
rect 28592 33612 29009 33640
rect 28592 33600 28598 33612
rect 28997 33609 29009 33612
rect 29043 33609 29055 33643
rect 28997 33603 29055 33609
rect 30374 33600 30380 33652
rect 30432 33640 30438 33652
rect 30469 33643 30527 33649
rect 30469 33640 30481 33643
rect 30432 33612 30481 33640
rect 30432 33600 30438 33612
rect 30469 33609 30481 33612
rect 30515 33609 30527 33643
rect 30469 33603 30527 33609
rect 31941 33643 31999 33649
rect 31941 33609 31953 33643
rect 31987 33640 31999 33643
rect 33502 33640 33508 33652
rect 31987 33612 33508 33640
rect 31987 33609 31999 33612
rect 31941 33603 31999 33609
rect 9490 33572 9496 33584
rect 9451 33544 9496 33572
rect 9490 33532 9496 33544
rect 9548 33532 9554 33584
rect 9582 33532 9588 33584
rect 9640 33572 9646 33584
rect 9677 33575 9735 33581
rect 9677 33572 9689 33575
rect 9640 33544 9689 33572
rect 9640 33532 9646 33544
rect 9677 33541 9689 33544
rect 9723 33541 9735 33575
rect 9677 33535 9735 33541
rect 19334 33532 19340 33584
rect 19392 33572 19398 33584
rect 22005 33575 22063 33581
rect 22005 33572 22017 33575
rect 19392 33544 22017 33572
rect 19392 33532 19398 33544
rect 22005 33541 22017 33544
rect 22051 33541 22063 33575
rect 22005 33535 22063 33541
rect 26970 33532 26976 33584
rect 27028 33572 27034 33584
rect 27249 33575 27307 33581
rect 27249 33572 27261 33575
rect 27028 33544 27261 33572
rect 27028 33532 27034 33544
rect 27249 33541 27261 33544
rect 27295 33541 27307 33575
rect 27249 33535 27307 33541
rect 28721 33575 28779 33581
rect 28721 33541 28733 33575
rect 28767 33572 28779 33575
rect 29638 33572 29644 33584
rect 28767 33544 29644 33572
rect 28767 33541 28779 33544
rect 28721 33535 28779 33541
rect 4982 33504 4988 33516
rect 4943 33476 4988 33504
rect 4982 33464 4988 33476
rect 5040 33464 5046 33516
rect 13630 33504 13636 33516
rect 13591 33476 13636 33504
rect 13630 33464 13636 33476
rect 13688 33464 13694 33516
rect 21082 33464 21088 33516
rect 21140 33504 21146 33516
rect 21453 33507 21511 33513
rect 21453 33504 21465 33507
rect 21140 33476 21465 33504
rect 21140 33464 21146 33476
rect 21453 33473 21465 33476
rect 21499 33504 21511 33507
rect 22833 33507 22891 33513
rect 22833 33504 22845 33507
rect 21499 33476 22845 33504
rect 21499 33473 21511 33476
rect 21453 33467 21511 33473
rect 22833 33473 22845 33476
rect 22879 33473 22891 33507
rect 22833 33467 22891 33473
rect 23934 33464 23940 33516
rect 23992 33504 23998 33516
rect 25731 33507 25789 33513
rect 23992 33476 25671 33504
rect 23992 33464 23998 33476
rect 3329 33439 3387 33445
rect 3329 33405 3341 33439
rect 3375 33436 3387 33439
rect 3694 33436 3700 33448
rect 3375 33408 3700 33436
rect 3375 33405 3387 33408
rect 3329 33399 3387 33405
rect 3694 33396 3700 33408
rect 3752 33396 3758 33448
rect 3970 33436 3976 33448
rect 3931 33408 3976 33436
rect 3970 33396 3976 33408
rect 4028 33396 4034 33448
rect 4157 33439 4215 33445
rect 4157 33405 4169 33439
rect 4203 33436 4215 33439
rect 6454 33436 6460 33448
rect 4203 33408 6460 33436
rect 4203 33405 4215 33408
rect 4157 33399 4215 33405
rect 6454 33396 6460 33408
rect 6512 33396 6518 33448
rect 6822 33436 6828 33448
rect 6783 33408 6828 33436
rect 6822 33396 6828 33408
rect 6880 33396 6886 33448
rect 9284 33439 9342 33445
rect 9284 33405 9296 33439
rect 9330 33436 9342 33439
rect 9582 33436 9588 33448
rect 9330 33408 9588 33436
rect 9330 33405 9342 33408
rect 9284 33399 9342 33405
rect 9582 33396 9588 33408
rect 9640 33436 9646 33448
rect 10045 33439 10103 33445
rect 10045 33436 10057 33439
rect 9640 33408 10057 33436
rect 9640 33396 9646 33408
rect 10045 33405 10057 33408
rect 10091 33405 10103 33439
rect 10045 33399 10103 33405
rect 10296 33439 10354 33445
rect 10296 33405 10308 33439
rect 10342 33405 10354 33439
rect 10296 33399 10354 33405
rect 11400 33439 11458 33445
rect 11400 33405 11412 33439
rect 11446 33436 11458 33439
rect 11514 33436 11520 33448
rect 11446 33408 11520 33436
rect 11446 33405 11458 33408
rect 11400 33399 11458 33405
rect 4893 33371 4951 33377
rect 4893 33337 4905 33371
rect 4939 33368 4951 33371
rect 5347 33371 5405 33377
rect 5347 33368 5359 33371
rect 4939 33340 5359 33368
rect 4939 33337 4951 33340
rect 4893 33331 4951 33337
rect 5347 33337 5359 33340
rect 5393 33368 5405 33371
rect 6086 33368 6092 33380
rect 5393 33340 6092 33368
rect 5393 33337 5405 33340
rect 5347 33331 5405 33337
rect 6086 33328 6092 33340
rect 6144 33368 6150 33380
rect 6641 33371 6699 33377
rect 6641 33368 6653 33371
rect 6144 33340 6653 33368
rect 6144 33328 6150 33340
rect 6641 33337 6653 33340
rect 6687 33368 6699 33371
rect 7187 33371 7245 33377
rect 7187 33368 7199 33371
rect 6687 33340 7199 33368
rect 6687 33337 6699 33340
rect 6641 33331 6699 33337
rect 7187 33337 7199 33340
rect 7233 33368 7245 33371
rect 7834 33368 7840 33380
rect 7233 33340 7840 33368
rect 7233 33337 7245 33340
rect 7187 33331 7245 33337
rect 7834 33328 7840 33340
rect 7892 33328 7898 33380
rect 8846 33328 8852 33380
rect 8904 33368 8910 33380
rect 10311 33368 10339 33399
rect 11514 33396 11520 33408
rect 11572 33436 11578 33448
rect 12161 33439 12219 33445
rect 12161 33436 12173 33439
rect 11572 33408 12173 33436
rect 11572 33396 11578 33408
rect 12161 33405 12173 33408
rect 12207 33405 12219 33439
rect 12161 33399 12219 33405
rect 12805 33439 12863 33445
rect 12805 33405 12817 33439
rect 12851 33436 12863 33439
rect 13173 33439 13231 33445
rect 13173 33436 13185 33439
rect 12851 33408 13185 33436
rect 12851 33405 12863 33408
rect 12805 33399 12863 33405
rect 13173 33405 13185 33408
rect 13219 33436 13231 33439
rect 13354 33436 13360 33448
rect 13219 33408 13360 33436
rect 13219 33405 13231 33408
rect 13173 33399 13231 33405
rect 13354 33396 13360 33408
rect 13412 33396 13418 33448
rect 13449 33439 13507 33445
rect 13449 33405 13461 33439
rect 13495 33436 13507 33439
rect 13538 33436 13544 33448
rect 13495 33408 13544 33436
rect 13495 33405 13507 33408
rect 13449 33399 13507 33405
rect 13538 33396 13544 33408
rect 13596 33396 13602 33448
rect 14642 33436 14648 33448
rect 14603 33408 14648 33436
rect 14642 33396 14648 33408
rect 14700 33396 14706 33448
rect 15565 33439 15623 33445
rect 15565 33405 15577 33439
rect 15611 33436 15623 33439
rect 16209 33439 16267 33445
rect 16209 33436 16221 33439
rect 15611 33408 16221 33436
rect 15611 33405 15623 33408
rect 15565 33399 15623 33405
rect 16209 33405 16221 33408
rect 16255 33436 16267 33439
rect 16428 33439 16486 33445
rect 16428 33436 16440 33439
rect 16255 33408 16440 33436
rect 16255 33405 16267 33408
rect 16209 33399 16267 33405
rect 16428 33405 16440 33408
rect 16474 33405 16486 33439
rect 18598 33436 18604 33448
rect 18559 33408 18604 33436
rect 16428 33399 16486 33405
rect 18598 33396 18604 33408
rect 18656 33396 18662 33448
rect 20416 33439 20474 33445
rect 20416 33405 20428 33439
rect 20462 33436 20474 33439
rect 20898 33436 20904 33448
rect 20462 33408 20904 33436
rect 20462 33405 20474 33408
rect 20416 33399 20474 33405
rect 20898 33396 20904 33408
rect 20956 33396 20962 33448
rect 23382 33436 23388 33448
rect 23295 33408 23388 33436
rect 23382 33396 23388 33408
rect 23440 33436 23446 33448
rect 23661 33439 23719 33445
rect 23661 33436 23673 33439
rect 23440 33408 23673 33436
rect 23440 33396 23446 33408
rect 23661 33405 23673 33408
rect 23707 33405 23719 33439
rect 23661 33399 23719 33405
rect 23842 33396 23848 33448
rect 23900 33436 23906 33448
rect 24118 33436 24124 33448
rect 23900 33408 24124 33436
rect 23900 33396 23906 33408
rect 24118 33396 24124 33408
rect 24176 33396 24182 33448
rect 25643 33445 25671 33476
rect 25731 33473 25743 33507
rect 25777 33504 25789 33507
rect 26697 33507 26755 33513
rect 26697 33504 26709 33507
rect 25777 33476 26709 33504
rect 25777 33473 25789 33476
rect 25731 33467 25789 33473
rect 26697 33473 26709 33476
rect 26743 33504 26755 33507
rect 27985 33507 28043 33513
rect 27985 33504 27997 33507
rect 26743 33476 27997 33504
rect 26743 33473 26755 33476
rect 26697 33467 26755 33473
rect 27985 33473 27997 33476
rect 28031 33473 28043 33507
rect 28736 33504 28764 33535
rect 29638 33532 29644 33544
rect 29696 33532 29702 33584
rect 29454 33504 29460 33516
rect 27985 33467 28043 33473
rect 28251 33476 28764 33504
rect 29196 33476 29460 33504
rect 25628 33439 25686 33445
rect 25628 33405 25640 33439
rect 25674 33436 25686 33439
rect 26050 33436 26056 33448
rect 25674 33408 26056 33436
rect 25674 33405 25686 33408
rect 25628 33399 25686 33405
rect 26050 33396 26056 33408
rect 26108 33396 26114 33448
rect 28251 33445 28279 33476
rect 29196 33448 29224 33476
rect 29454 33464 29460 33476
rect 29512 33464 29518 33516
rect 30484 33504 30512 33603
rect 33502 33600 33508 33612
rect 33560 33600 33566 33652
rect 34422 33640 34428 33652
rect 34383 33612 34428 33640
rect 34422 33600 34428 33612
rect 34480 33600 34486 33652
rect 36354 33600 36360 33652
rect 36412 33640 36418 33652
rect 37185 33643 37243 33649
rect 37185 33640 37197 33643
rect 36412 33612 37197 33640
rect 36412 33600 36418 33612
rect 37185 33609 37197 33612
rect 37231 33609 37243 33643
rect 37826 33640 37832 33652
rect 37787 33612 37832 33640
rect 37185 33603 37243 33609
rect 37826 33600 37832 33612
rect 37884 33600 37890 33652
rect 37918 33600 37924 33652
rect 37976 33640 37982 33652
rect 38565 33643 38623 33649
rect 38565 33640 38577 33643
rect 37976 33612 38577 33640
rect 37976 33600 37982 33612
rect 38565 33609 38577 33612
rect 38611 33640 38623 33643
rect 38930 33640 38936 33652
rect 38611 33612 38936 33640
rect 38611 33609 38623 33612
rect 38565 33603 38623 33609
rect 38930 33600 38936 33612
rect 38988 33600 38994 33652
rect 39945 33643 40003 33649
rect 39945 33609 39957 33643
rect 39991 33640 40003 33643
rect 40313 33643 40371 33649
rect 40313 33640 40325 33643
rect 39991 33612 40325 33640
rect 39991 33609 40003 33612
rect 39945 33603 40003 33609
rect 40313 33609 40325 33612
rect 40359 33640 40371 33643
rect 40586 33640 40592 33652
rect 40359 33612 40592 33640
rect 40359 33609 40371 33612
rect 40313 33603 40371 33609
rect 40586 33600 40592 33612
rect 40644 33600 40650 33652
rect 41506 33640 41512 33652
rect 41467 33612 41512 33640
rect 41506 33600 41512 33612
rect 41564 33600 41570 33652
rect 42242 33640 42248 33652
rect 42203 33612 42248 33640
rect 42242 33600 42248 33612
rect 42300 33600 42306 33652
rect 32950 33572 32956 33584
rect 32508 33544 32956 33572
rect 30745 33507 30803 33513
rect 30745 33504 30757 33507
rect 30484 33476 30757 33504
rect 30745 33473 30757 33476
rect 30791 33473 30803 33507
rect 31018 33504 31024 33516
rect 30979 33476 31024 33504
rect 30745 33467 30803 33473
rect 31018 33464 31024 33476
rect 31076 33464 31082 33516
rect 32508 33513 32536 33544
rect 32950 33532 32956 33544
rect 33008 33532 33014 33584
rect 33226 33532 33232 33584
rect 33284 33572 33290 33584
rect 34606 33572 34612 33584
rect 33284 33544 34612 33572
rect 33284 33532 33290 33544
rect 34606 33532 34612 33544
rect 34664 33532 34670 33584
rect 39390 33572 39396 33584
rect 38856 33544 39396 33572
rect 32493 33507 32551 33513
rect 32493 33473 32505 33507
rect 32539 33473 32551 33507
rect 32766 33504 32772 33516
rect 32727 33476 32772 33504
rect 32493 33467 32551 33473
rect 32766 33464 32772 33476
rect 32824 33464 32830 33516
rect 35345 33507 35403 33513
rect 35345 33504 35357 33507
rect 34935 33476 35357 33504
rect 28236 33439 28294 33445
rect 28236 33405 28248 33439
rect 28282 33405 28294 33439
rect 28236 33399 28294 33405
rect 29178 33396 29184 33448
rect 29236 33396 29242 33448
rect 29324 33439 29382 33445
rect 29324 33405 29336 33439
rect 29370 33436 29382 33439
rect 29370 33408 29868 33436
rect 29370 33405 29382 33408
rect 29324 33399 29382 33405
rect 10689 33371 10747 33377
rect 10689 33368 10701 33371
rect 8904 33340 10701 33368
rect 8904 33328 8910 33340
rect 10689 33337 10701 33340
rect 10735 33337 10747 33371
rect 11882 33368 11888 33380
rect 11795 33340 11888 33368
rect 10689 33331 10747 33337
rect 11882 33328 11888 33340
rect 11940 33368 11946 33380
rect 13722 33368 13728 33380
rect 11940 33340 13728 33368
rect 11940 33328 11946 33340
rect 13722 33328 13728 33340
rect 13780 33368 13786 33380
rect 14553 33371 14611 33377
rect 14553 33368 14565 33371
rect 13780 33340 14565 33368
rect 13780 33328 13786 33340
rect 14553 33337 14565 33340
rect 14599 33368 14611 33371
rect 15007 33371 15065 33377
rect 15007 33368 15019 33371
rect 14599 33340 15019 33368
rect 14599 33337 14611 33340
rect 14553 33331 14611 33337
rect 15007 33337 15019 33340
rect 15053 33368 15065 33371
rect 15470 33368 15476 33380
rect 15053 33340 15476 33368
rect 15053 33337 15065 33340
rect 15007 33331 15065 33337
rect 15470 33328 15476 33340
rect 15528 33328 15534 33380
rect 17589 33371 17647 33377
rect 17589 33337 17601 33371
rect 17635 33368 17647 33371
rect 17678 33368 17684 33380
rect 17635 33340 17684 33368
rect 17635 33337 17647 33340
rect 17589 33331 17647 33337
rect 17678 33328 17684 33340
rect 17736 33368 17742 33380
rect 18506 33368 18512 33380
rect 17736 33340 18512 33368
rect 17736 33328 17742 33340
rect 18506 33328 18512 33340
rect 18564 33328 18570 33380
rect 18690 33328 18696 33380
rect 18748 33368 18754 33380
rect 18963 33371 19021 33377
rect 18963 33368 18975 33371
rect 18748 33340 18975 33368
rect 18748 33328 18754 33340
rect 18963 33337 18975 33340
rect 19009 33368 19021 33371
rect 19150 33368 19156 33380
rect 19009 33340 19156 33368
rect 19009 33337 19021 33340
rect 18963 33331 19021 33337
rect 19150 33328 19156 33340
rect 19208 33328 19214 33380
rect 21545 33371 21603 33377
rect 21545 33337 21557 33371
rect 21591 33337 21603 33371
rect 21545 33331 21603 33337
rect 4525 33303 4583 33309
rect 4525 33269 4537 33303
rect 4571 33300 4583 33303
rect 4706 33300 4712 33312
rect 4571 33272 4712 33300
rect 4571 33269 4583 33272
rect 4525 33263 4583 33269
rect 4706 33260 4712 33272
rect 4764 33260 4770 33312
rect 8478 33260 8484 33312
rect 8536 33300 8542 33312
rect 8573 33303 8631 33309
rect 8573 33300 8585 33303
rect 8536 33272 8585 33300
rect 8536 33260 8542 33272
rect 8573 33269 8585 33272
rect 8619 33269 8631 33303
rect 8573 33263 8631 33269
rect 11471 33303 11529 33309
rect 11471 33269 11483 33303
rect 11517 33300 11529 33303
rect 12434 33300 12440 33312
rect 11517 33272 12440 33300
rect 11517 33269 11529 33272
rect 11471 33263 11529 33269
rect 12434 33260 12440 33272
rect 12492 33260 12498 33312
rect 18417 33303 18475 33309
rect 18417 33269 18429 33303
rect 18463 33300 18475 33303
rect 18708 33300 18736 33328
rect 20898 33300 20904 33312
rect 18463 33272 18736 33300
rect 20859 33272 20904 33300
rect 18463 33269 18475 33272
rect 18417 33263 18475 33269
rect 20898 33260 20904 33272
rect 20956 33260 20962 33312
rect 21266 33260 21272 33312
rect 21324 33300 21330 33312
rect 21560 33300 21588 33331
rect 25958 33328 25964 33380
rect 26016 33368 26022 33380
rect 26421 33371 26479 33377
rect 26421 33368 26433 33371
rect 26016 33340 26433 33368
rect 26016 33328 26022 33340
rect 26421 33337 26433 33340
rect 26467 33368 26479 33371
rect 26789 33371 26847 33377
rect 26789 33368 26801 33371
rect 26467 33340 26801 33368
rect 26467 33337 26479 33340
rect 26421 33331 26479 33337
rect 26789 33337 26801 33340
rect 26835 33368 26847 33371
rect 26878 33368 26884 33380
rect 26835 33340 26884 33368
rect 26835 33337 26847 33340
rect 26789 33331 26847 33337
rect 26878 33328 26884 33340
rect 26936 33328 26942 33380
rect 27706 33328 27712 33380
rect 27764 33368 27770 33380
rect 29411 33371 29469 33377
rect 29411 33368 29423 33371
rect 27764 33340 29423 33368
rect 27764 33328 27770 33340
rect 29411 33337 29423 33340
rect 29457 33337 29469 33371
rect 29411 33331 29469 33337
rect 23750 33300 23756 33312
rect 21324 33272 21588 33300
rect 23711 33272 23756 33300
rect 21324 33260 21330 33272
rect 23750 33260 23756 33272
rect 23808 33260 23814 33312
rect 26896 33300 26924 33328
rect 27617 33303 27675 33309
rect 27617 33300 27629 33303
rect 26896 33272 27629 33300
rect 27617 33269 27629 33272
rect 27663 33269 27675 33303
rect 27617 33263 27675 33269
rect 29730 33260 29736 33312
rect 29788 33300 29794 33312
rect 29840 33309 29868 33408
rect 34054 33396 34060 33448
rect 34112 33436 34118 33448
rect 34935 33445 34963 33476
rect 35345 33473 35357 33476
rect 35391 33473 35403 33507
rect 35345 33467 35403 33473
rect 36081 33507 36139 33513
rect 36081 33473 36093 33507
rect 36127 33504 36139 33507
rect 36909 33507 36967 33513
rect 36127 33476 36584 33504
rect 36127 33473 36139 33476
rect 36081 33467 36139 33473
rect 36556 33448 36584 33476
rect 36909 33473 36921 33507
rect 36955 33504 36967 33507
rect 37734 33504 37740 33516
rect 36955 33476 37740 33504
rect 36955 33473 36967 33476
rect 36909 33467 36967 33473
rect 37734 33464 37740 33476
rect 37792 33504 37798 33516
rect 38856 33513 38884 33544
rect 39390 33532 39396 33544
rect 39448 33572 39454 33584
rect 41141 33575 41199 33581
rect 41141 33572 41153 33575
rect 39448 33544 41153 33572
rect 39448 33532 39454 33544
rect 41141 33541 41153 33544
rect 41187 33572 41199 33575
rect 42886 33572 42892 33584
rect 41187 33544 42892 33572
rect 41187 33541 41199 33544
rect 41141 33535 41199 33541
rect 42886 33532 42892 33544
rect 42944 33532 42950 33584
rect 38105 33507 38163 33513
rect 38105 33504 38117 33507
rect 37792 33476 38117 33504
rect 37792 33464 37798 33476
rect 38105 33473 38117 33476
rect 38151 33473 38163 33507
rect 38105 33467 38163 33473
rect 38841 33507 38899 33513
rect 38841 33473 38853 33507
rect 38887 33473 38899 33507
rect 38841 33467 38899 33473
rect 39206 33464 39212 33516
rect 39264 33504 39270 33516
rect 39482 33504 39488 33516
rect 39264 33476 39488 33504
rect 39264 33464 39270 33476
rect 39482 33464 39488 33476
rect 39540 33464 39546 33516
rect 40589 33507 40647 33513
rect 40589 33473 40601 33507
rect 40635 33504 40647 33507
rect 40770 33504 40776 33516
rect 40635 33476 40776 33504
rect 40635 33473 40647 33476
rect 40589 33467 40647 33473
rect 40770 33464 40776 33476
rect 40828 33504 40834 33516
rect 41877 33507 41935 33513
rect 41877 33504 41889 33507
rect 40828 33476 41889 33504
rect 40828 33464 40834 33476
rect 41877 33473 41889 33476
rect 41923 33473 41935 33507
rect 42702 33504 42708 33516
rect 42663 33476 42708 33504
rect 41877 33467 41935 33473
rect 42702 33464 42708 33476
rect 42760 33464 42766 33516
rect 42794 33464 42800 33516
rect 42852 33504 42858 33516
rect 42981 33507 43039 33513
rect 42981 33504 42993 33507
rect 42852 33476 42993 33504
rect 42852 33464 42858 33476
rect 42981 33473 42993 33476
rect 43027 33473 43039 33507
rect 44542 33504 44548 33516
rect 44503 33476 44548 33504
rect 42981 33467 43039 33473
rect 44542 33464 44548 33476
rect 44600 33464 44606 33516
rect 34920 33439 34978 33445
rect 34920 33436 34932 33439
rect 34112 33408 34932 33436
rect 34112 33396 34118 33408
rect 34920 33405 34932 33408
rect 34966 33405 34978 33439
rect 34920 33399 34978 33405
rect 35250 33396 35256 33448
rect 35308 33436 35314 33448
rect 36449 33439 36507 33445
rect 36449 33436 36461 33439
rect 35308 33408 36461 33436
rect 35308 33396 35314 33408
rect 36449 33405 36461 33408
rect 36495 33405 36507 33439
rect 36449 33399 36507 33405
rect 30193 33371 30251 33377
rect 30193 33337 30205 33371
rect 30239 33368 30251 33371
rect 30558 33368 30564 33380
rect 30239 33340 30564 33368
rect 30239 33337 30251 33340
rect 30193 33331 30251 33337
rect 30558 33328 30564 33340
rect 30616 33368 30622 33380
rect 30837 33371 30895 33377
rect 30837 33368 30849 33371
rect 30616 33340 30849 33368
rect 30616 33328 30622 33340
rect 30837 33337 30849 33340
rect 30883 33337 30895 33371
rect 30837 33331 30895 33337
rect 31849 33371 31907 33377
rect 31849 33337 31861 33371
rect 31895 33368 31907 33371
rect 32585 33371 32643 33377
rect 31895 33340 32352 33368
rect 31895 33337 31907 33340
rect 31849 33331 31907 33337
rect 29825 33303 29883 33309
rect 29825 33300 29837 33303
rect 29788 33272 29837 33300
rect 29788 33260 29794 33272
rect 29825 33269 29837 33272
rect 29871 33300 29883 33303
rect 31941 33303 31999 33309
rect 31941 33300 31953 33303
rect 29871 33272 31953 33300
rect 29871 33269 29883 33272
rect 29825 33263 29883 33269
rect 31941 33269 31953 33272
rect 31987 33269 31999 33303
rect 32122 33300 32128 33312
rect 32083 33272 32128 33300
rect 31941 33263 31999 33269
rect 32122 33260 32128 33272
rect 32180 33260 32186 33312
rect 32324 33300 32352 33340
rect 32585 33337 32597 33371
rect 32631 33337 32643 33371
rect 35894 33368 35900 33380
rect 32585 33331 32643 33337
rect 35268 33340 35900 33368
rect 32600 33300 32628 33331
rect 35268 33312 35296 33340
rect 35894 33328 35900 33340
rect 35952 33328 35958 33380
rect 36464 33368 36492 33399
rect 36538 33396 36544 33448
rect 36596 33436 36602 33448
rect 36633 33439 36691 33445
rect 36633 33436 36645 33439
rect 36596 33408 36645 33436
rect 36596 33396 36602 33408
rect 36633 33405 36645 33408
rect 36679 33405 36691 33439
rect 36633 33399 36691 33405
rect 36906 33368 36912 33380
rect 36464 33340 36912 33368
rect 36906 33328 36912 33340
rect 36964 33328 36970 33380
rect 38930 33328 38936 33380
rect 38988 33368 38994 33380
rect 38988 33340 39033 33368
rect 38988 33328 38994 33340
rect 40678 33328 40684 33380
rect 40736 33368 40742 33380
rect 42794 33368 42800 33380
rect 40736 33340 40781 33368
rect 42707 33340 42800 33368
rect 40736 33328 40742 33340
rect 42794 33328 42800 33340
rect 42852 33368 42858 33380
rect 43530 33368 43536 33380
rect 42852 33340 43536 33368
rect 42852 33328 42858 33340
rect 43530 33328 43536 33340
rect 43588 33368 43594 33380
rect 43717 33371 43775 33377
rect 43717 33368 43729 33371
rect 43588 33340 43729 33368
rect 43588 33328 43594 33340
rect 43717 33337 43729 33340
rect 43763 33368 43775 33371
rect 44082 33368 44088 33380
rect 43763 33340 44088 33368
rect 43763 33337 43775 33340
rect 43717 33331 43775 33337
rect 44082 33328 44088 33340
rect 44140 33328 44146 33380
rect 44269 33371 44327 33377
rect 44269 33337 44281 33371
rect 44315 33337 44327 33371
rect 44269 33331 44327 33337
rect 33042 33300 33048 33312
rect 32324 33272 33048 33300
rect 33042 33260 33048 33272
rect 33100 33260 33106 33312
rect 33410 33260 33416 33312
rect 33468 33300 33474 33312
rect 35023 33303 35081 33309
rect 35023 33300 35035 33303
rect 33468 33272 35035 33300
rect 33468 33260 33474 33272
rect 35023 33269 35035 33272
rect 35069 33269 35081 33303
rect 35023 33263 35081 33269
rect 35250 33260 35256 33312
rect 35308 33260 35314 33312
rect 38102 33260 38108 33312
rect 38160 33300 38166 33312
rect 39574 33300 39580 33312
rect 38160 33272 39580 33300
rect 38160 33260 38166 33272
rect 39574 33260 39580 33272
rect 39632 33260 39638 33312
rect 43990 33300 43996 33312
rect 43951 33272 43996 33300
rect 43990 33260 43996 33272
rect 44048 33300 44054 33312
rect 44284 33300 44312 33331
rect 44358 33328 44364 33380
rect 44416 33368 44422 33380
rect 44416 33340 44461 33368
rect 44416 33328 44422 33340
rect 44048 33272 44312 33300
rect 44048 33260 44054 33272
rect 1104 33210 48852 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 48852 33210
rect 1104 33136 48852 33158
rect 4062 33056 4068 33108
rect 4120 33096 4126 33108
rect 4157 33099 4215 33105
rect 4157 33096 4169 33099
rect 4120 33068 4169 33096
rect 4120 33056 4126 33068
rect 4157 33065 4169 33068
rect 4203 33065 4215 33099
rect 4157 33059 4215 33065
rect 4982 33056 4988 33108
rect 5040 33096 5046 33108
rect 5445 33099 5503 33105
rect 5445 33096 5457 33099
rect 5040 33068 5457 33096
rect 5040 33056 5046 33068
rect 5445 33065 5457 33068
rect 5491 33065 5503 33099
rect 7834 33096 7840 33108
rect 7795 33068 7840 33096
rect 5445 33059 5503 33065
rect 7834 33056 7840 33068
rect 7892 33056 7898 33108
rect 8389 33099 8447 33105
rect 8389 33065 8401 33099
rect 8435 33096 8447 33099
rect 8478 33096 8484 33108
rect 8435 33068 8484 33096
rect 8435 33065 8447 33068
rect 8389 33059 8447 33065
rect 8478 33056 8484 33068
rect 8536 33056 8542 33108
rect 9582 33056 9588 33108
rect 9640 33096 9646 33108
rect 10597 33099 10655 33105
rect 10597 33096 10609 33099
rect 9640 33068 10609 33096
rect 9640 33056 9646 33068
rect 10597 33065 10609 33068
rect 10643 33065 10655 33099
rect 12342 33096 12348 33108
rect 12303 33068 12348 33096
rect 10597 33059 10655 33065
rect 12342 33056 12348 33068
rect 12400 33056 12406 33108
rect 13262 33096 13268 33108
rect 13223 33068 13268 33096
rect 13262 33056 13268 33068
rect 13320 33056 13326 33108
rect 13446 33056 13452 33108
rect 13504 33096 13510 33108
rect 14642 33096 14648 33108
rect 13504 33068 13814 33096
rect 14603 33068 14648 33096
rect 13504 33056 13510 33068
rect 3970 32988 3976 33040
rect 4028 33028 4034 33040
rect 10039 33031 10097 33037
rect 4028 33000 4660 33028
rect 4028 32988 4034 33000
rect 3510 32920 3516 32972
rect 3568 32960 3574 32972
rect 4632 32969 4660 33000
rect 10039 32997 10051 33031
rect 10085 33028 10097 33031
rect 11422 33028 11428 33040
rect 10085 33000 11428 33028
rect 10085 32997 10097 33000
rect 10039 32991 10097 32997
rect 11422 32988 11428 33000
rect 11480 33028 11486 33040
rect 11746 33031 11804 33037
rect 11746 33028 11758 33031
rect 11480 33000 11758 33028
rect 11480 32988 11486 33000
rect 11746 32997 11758 33000
rect 11792 33028 11804 33031
rect 11882 33028 11888 33040
rect 11792 33000 11888 33028
rect 11792 32997 11804 33000
rect 11746 32991 11804 32997
rect 11882 32988 11888 33000
rect 11940 32988 11946 33040
rect 4065 32963 4123 32969
rect 4065 32960 4077 32963
rect 3568 32932 4077 32960
rect 3568 32920 3574 32932
rect 4065 32929 4077 32932
rect 4111 32929 4123 32963
rect 4065 32923 4123 32929
rect 4617 32963 4675 32969
rect 4617 32929 4629 32963
rect 4663 32960 4675 32963
rect 5166 32960 5172 32972
rect 4663 32932 5172 32960
rect 4663 32929 4675 32932
rect 4617 32923 4675 32929
rect 5166 32920 5172 32932
rect 5224 32920 5230 32972
rect 6089 32963 6147 32969
rect 6089 32929 6101 32963
rect 6135 32929 6147 32963
rect 6362 32960 6368 32972
rect 6323 32932 6368 32960
rect 6089 32923 6147 32929
rect 6104 32892 6132 32923
rect 6362 32920 6368 32932
rect 6420 32920 6426 32972
rect 6549 32963 6607 32969
rect 6549 32929 6561 32963
rect 6595 32960 6607 32963
rect 6822 32960 6828 32972
rect 6595 32932 6828 32960
rect 6595 32929 6607 32932
rect 6549 32923 6607 32929
rect 6822 32920 6828 32932
rect 6880 32920 6886 32972
rect 13446 32960 13452 32972
rect 13407 32932 13452 32960
rect 13446 32920 13452 32932
rect 13504 32920 13510 32972
rect 13633 32963 13691 32969
rect 13633 32929 13645 32963
rect 13679 32929 13691 32963
rect 13786 32960 13814 33068
rect 14642 33056 14648 33068
rect 14700 33056 14706 33108
rect 18598 33096 18604 33108
rect 18559 33068 18604 33096
rect 18598 33056 18604 33068
rect 18656 33056 18662 33108
rect 19058 33096 19064 33108
rect 19019 33068 19064 33096
rect 19058 33056 19064 33068
rect 19116 33096 19122 33108
rect 20254 33096 20260 33108
rect 19116 33068 19288 33096
rect 20167 33068 20260 33096
rect 19116 33056 19122 33068
rect 15470 32988 15476 33040
rect 15528 33028 15534 33040
rect 15610 33031 15668 33037
rect 15610 33028 15622 33031
rect 15528 33000 15622 33028
rect 15528 32988 15534 33000
rect 15610 32997 15622 33000
rect 15656 32997 15668 33031
rect 15610 32991 15668 32997
rect 17402 32988 17408 33040
rect 17460 33028 17466 33040
rect 17726 33031 17784 33037
rect 17726 33028 17738 33031
rect 17460 33000 17738 33028
rect 17460 32988 17466 33000
rect 17726 32997 17738 33000
rect 17772 33028 17784 33031
rect 18690 33028 18696 33040
rect 17772 33000 18696 33028
rect 17772 32997 17784 33000
rect 17726 32991 17784 32997
rect 18690 32988 18696 33000
rect 18748 32988 18754 33040
rect 19260 33037 19288 33068
rect 20254 33056 20260 33068
rect 20312 33096 20318 33108
rect 21634 33096 21640 33108
rect 20312 33068 21640 33096
rect 20312 33056 20318 33068
rect 21634 33056 21640 33068
rect 21692 33056 21698 33108
rect 22370 33056 22376 33108
rect 22428 33096 22434 33108
rect 23474 33096 23480 33108
rect 22428 33068 23480 33096
rect 22428 33056 22434 33068
rect 23474 33056 23480 33068
rect 23532 33056 23538 33108
rect 23569 33099 23627 33105
rect 23569 33065 23581 33099
rect 23615 33065 23627 33099
rect 23569 33059 23627 33065
rect 19245 33031 19303 33037
rect 19245 32997 19257 33031
rect 19291 32997 19303 33031
rect 19245 32991 19303 32997
rect 19334 32988 19340 33040
rect 19392 33028 19398 33040
rect 19392 33000 19437 33028
rect 19392 32988 19398 33000
rect 23290 32988 23296 33040
rect 23348 33028 23354 33040
rect 23584 33028 23612 33059
rect 26786 33056 26792 33108
rect 26844 33096 26850 33108
rect 27433 33099 27491 33105
rect 27433 33096 27445 33099
rect 26844 33068 27445 33096
rect 26844 33056 26850 33068
rect 27433 33065 27445 33068
rect 27479 33096 27491 33099
rect 27706 33096 27712 33108
rect 27479 33068 27712 33096
rect 27479 33065 27491 33068
rect 27433 33059 27491 33065
rect 27706 33056 27712 33068
rect 27764 33056 27770 33108
rect 29546 33056 29552 33108
rect 29604 33096 29610 33108
rect 32766 33096 32772 33108
rect 29604 33068 32772 33096
rect 29604 33056 29610 33068
rect 30650 33028 30656 33040
rect 23348 33000 23612 33028
rect 30611 33000 30656 33028
rect 23348 32988 23354 33000
rect 30650 32988 30656 33000
rect 30708 32988 30714 33040
rect 31220 33037 31248 33068
rect 32766 33056 32772 33068
rect 32824 33056 32830 33108
rect 33042 33096 33048 33108
rect 33003 33068 33048 33096
rect 33042 33056 33048 33068
rect 33100 33056 33106 33108
rect 33318 33056 33324 33108
rect 33376 33096 33382 33108
rect 34146 33096 34152 33108
rect 33376 33068 34152 33096
rect 33376 33056 33382 33068
rect 34146 33056 34152 33068
rect 34204 33056 34210 33108
rect 38378 33056 38384 33108
rect 38436 33096 38442 33108
rect 39850 33096 39856 33108
rect 38436 33068 39856 33096
rect 38436 33056 38442 33068
rect 39850 33056 39856 33068
rect 39908 33056 39914 33108
rect 42702 33056 42708 33108
rect 42760 33096 42766 33108
rect 43070 33096 43076 33108
rect 42760 33068 42978 33096
rect 43031 33068 43076 33096
rect 42760 33056 42766 33068
rect 31205 33031 31263 33037
rect 31205 32997 31217 33031
rect 31251 32997 31263 33031
rect 32398 33028 32404 33040
rect 32359 33000 32404 33028
rect 31205 32991 31263 32997
rect 32398 32988 32404 33000
rect 32456 32988 32462 33040
rect 33502 32988 33508 33040
rect 33560 33028 33566 33040
rect 34057 33031 34115 33037
rect 34057 33028 34069 33031
rect 33560 33000 34069 33028
rect 33560 32988 33566 33000
rect 34057 32997 34069 33000
rect 34103 33028 34115 33031
rect 35621 33031 35679 33037
rect 35621 33028 35633 33031
rect 34103 33000 35633 33028
rect 34103 32997 34115 33000
rect 34057 32991 34115 32997
rect 35621 32997 35633 33000
rect 35667 32997 35679 33031
rect 36906 33028 36912 33040
rect 36867 33000 36912 33028
rect 35621 32991 35679 32997
rect 36906 32988 36912 33000
rect 36964 32988 36970 33040
rect 39022 33028 39028 33040
rect 38983 33000 39028 33028
rect 39022 32988 39028 33000
rect 39080 32988 39086 33040
rect 40586 33028 40592 33040
rect 40547 33000 40592 33028
rect 40586 32988 40592 33000
rect 40644 32988 40650 33040
rect 42794 33028 42800 33040
rect 42755 33000 42800 33028
rect 42794 32988 42800 33000
rect 42852 32988 42858 33040
rect 42950 33028 42978 33068
rect 43070 33056 43076 33068
rect 43128 33056 43134 33108
rect 44269 33099 44327 33105
rect 44269 33065 44281 33099
rect 44315 33096 44327 33099
rect 44358 33096 44364 33108
rect 44315 33068 44364 33096
rect 44315 33065 44327 33068
rect 44269 33059 44327 33065
rect 44358 33056 44364 33068
rect 44416 33056 44422 33108
rect 43487 33031 43545 33037
rect 43487 33028 43499 33031
rect 42950 33000 43499 33028
rect 43487 32997 43499 33000
rect 43533 32997 43545 33031
rect 43487 32991 43545 32997
rect 16209 32963 16267 32969
rect 16209 32960 16221 32963
rect 13786 32932 16221 32960
rect 13633 32923 13691 32929
rect 16209 32929 16221 32932
rect 16255 32929 16267 32963
rect 16209 32923 16267 32929
rect 21913 32963 21971 32969
rect 21913 32929 21925 32963
rect 21959 32929 21971 32963
rect 21913 32923 21971 32929
rect 6270 32892 6276 32904
rect 6104 32864 6276 32892
rect 6270 32852 6276 32864
rect 6328 32852 6334 32904
rect 7466 32892 7472 32904
rect 7427 32864 7472 32892
rect 7466 32852 7472 32864
rect 7524 32852 7530 32904
rect 9677 32895 9735 32901
rect 9677 32861 9689 32895
rect 9723 32892 9735 32895
rect 10410 32892 10416 32904
rect 9723 32864 10416 32892
rect 9723 32861 9735 32864
rect 9677 32855 9735 32861
rect 10410 32852 10416 32864
rect 10468 32852 10474 32904
rect 11425 32895 11483 32901
rect 11425 32861 11437 32895
rect 11471 32892 11483 32895
rect 11882 32892 11888 32904
rect 11471 32864 11888 32892
rect 11471 32861 11483 32864
rect 11425 32855 11483 32861
rect 11882 32852 11888 32864
rect 11940 32852 11946 32904
rect 13538 32892 13544 32904
rect 13004 32864 13544 32892
rect 13004 32768 13032 32864
rect 13538 32852 13544 32864
rect 13596 32892 13602 32904
rect 13648 32892 13676 32923
rect 15286 32892 15292 32904
rect 13596 32864 13676 32892
rect 15247 32864 15292 32892
rect 13596 32852 13602 32864
rect 15286 32852 15292 32864
rect 15344 32852 15350 32904
rect 17405 32895 17463 32901
rect 17405 32861 17417 32895
rect 17451 32861 17463 32895
rect 19886 32892 19892 32904
rect 19799 32864 19892 32892
rect 17405 32855 17463 32861
rect 3234 32716 3240 32768
rect 3292 32756 3298 32768
rect 3421 32759 3479 32765
rect 3421 32756 3433 32759
rect 3292 32728 3433 32756
rect 3292 32716 3298 32728
rect 3421 32725 3433 32728
rect 3467 32756 3479 32759
rect 3970 32756 3976 32768
rect 3467 32728 3976 32756
rect 3467 32725 3479 32728
rect 3421 32719 3479 32725
rect 3970 32716 3976 32728
rect 4028 32716 4034 32768
rect 5166 32756 5172 32768
rect 5127 32728 5172 32756
rect 5166 32716 5172 32728
rect 5224 32716 5230 32768
rect 12986 32756 12992 32768
rect 12947 32728 12992 32756
rect 12986 32716 12992 32728
rect 13044 32716 13050 32768
rect 17310 32756 17316 32768
rect 17271 32728 17316 32756
rect 17310 32716 17316 32728
rect 17368 32756 17374 32768
rect 17420 32756 17448 32855
rect 19886 32852 19892 32864
rect 19944 32892 19950 32904
rect 20438 32892 20444 32904
rect 19944 32864 20444 32892
rect 19944 32852 19950 32864
rect 20438 32852 20444 32864
rect 20496 32852 20502 32904
rect 21928 32892 21956 32923
rect 22094 32920 22100 32972
rect 22152 32960 22158 32972
rect 22189 32963 22247 32969
rect 22189 32960 22201 32963
rect 22152 32932 22201 32960
rect 22152 32920 22158 32932
rect 22189 32929 22201 32932
rect 22235 32960 22247 32963
rect 24118 32960 24124 32972
rect 22235 32932 24124 32960
rect 22235 32929 22247 32932
rect 22189 32923 22247 32929
rect 24118 32920 24124 32932
rect 24176 32920 24182 32972
rect 25476 32963 25534 32969
rect 25476 32929 25488 32963
rect 25522 32960 25534 32963
rect 25590 32960 25596 32972
rect 25522 32932 25596 32960
rect 25522 32929 25534 32932
rect 25476 32923 25534 32929
rect 25590 32920 25596 32932
rect 25648 32920 25654 32972
rect 26234 32960 26240 32972
rect 25786 32932 26240 32960
rect 22278 32892 22284 32904
rect 21928 32864 22284 32892
rect 22278 32852 22284 32864
rect 22336 32852 22342 32904
rect 22373 32895 22431 32901
rect 22373 32861 22385 32895
rect 22419 32892 22431 32895
rect 22830 32892 22836 32904
rect 22419 32864 22836 32892
rect 22419 32861 22431 32864
rect 22373 32855 22431 32861
rect 22830 32852 22836 32864
rect 22888 32892 22894 32904
rect 23201 32895 23259 32901
rect 23201 32892 23213 32895
rect 22888 32864 23213 32892
rect 22888 32852 22894 32864
rect 23201 32861 23213 32864
rect 23247 32861 23259 32895
rect 23201 32855 23259 32861
rect 23474 32852 23480 32904
rect 23532 32892 23538 32904
rect 25786 32892 25814 32932
rect 26234 32920 26240 32932
rect 26292 32960 26298 32972
rect 26548 32963 26606 32969
rect 26548 32960 26560 32963
rect 26292 32932 26560 32960
rect 26292 32920 26298 32932
rect 26548 32929 26560 32932
rect 26594 32929 26606 32963
rect 26548 32923 26606 32929
rect 27576 32963 27634 32969
rect 27576 32929 27588 32963
rect 27622 32960 27634 32963
rect 28074 32960 28080 32972
rect 27622 32932 28080 32960
rect 27622 32929 27634 32932
rect 27576 32923 27634 32929
rect 28074 32920 28080 32932
rect 28132 32920 28138 32972
rect 29178 32960 29184 32972
rect 29091 32932 29184 32960
rect 29178 32920 29184 32932
rect 29236 32920 29242 32972
rect 29362 32960 29368 32972
rect 29323 32932 29368 32960
rect 29362 32920 29368 32932
rect 29420 32920 29426 32972
rect 37734 32960 37740 32972
rect 37647 32932 37740 32960
rect 37734 32920 37740 32932
rect 37792 32960 37798 32972
rect 38746 32960 38752 32972
rect 37792 32932 38752 32960
rect 37792 32920 37798 32932
rect 38746 32920 38752 32932
rect 38804 32920 38810 32972
rect 43257 32963 43315 32969
rect 43257 32929 43269 32963
rect 43303 32960 43315 32963
rect 43346 32960 43352 32972
rect 43303 32932 43352 32960
rect 43303 32929 43315 32932
rect 43257 32923 43315 32929
rect 43346 32920 43352 32932
rect 43404 32960 43410 32972
rect 43806 32960 43812 32972
rect 43404 32932 43812 32960
rect 43404 32920 43410 32932
rect 43806 32920 43812 32932
rect 43864 32920 43870 32972
rect 23532 32864 25814 32892
rect 23532 32852 23538 32864
rect 26326 32852 26332 32904
rect 26384 32892 26390 32904
rect 27663 32895 27721 32901
rect 27663 32892 27675 32895
rect 26384 32864 27675 32892
rect 26384 32852 26390 32864
rect 27663 32861 27675 32864
rect 27709 32861 27721 32895
rect 27663 32855 27721 32861
rect 18325 32827 18383 32833
rect 18325 32793 18337 32827
rect 18371 32824 18383 32827
rect 19334 32824 19340 32836
rect 18371 32796 19340 32824
rect 18371 32793 18383 32796
rect 18325 32787 18383 32793
rect 19334 32784 19340 32796
rect 19392 32784 19398 32836
rect 26694 32784 26700 32836
rect 26752 32824 26758 32836
rect 26973 32827 27031 32833
rect 26973 32824 26985 32827
rect 26752 32796 26985 32824
rect 26752 32784 26758 32796
rect 26973 32793 26985 32796
rect 27019 32793 27031 32827
rect 26973 32787 27031 32793
rect 28994 32784 29000 32836
rect 29052 32824 29058 32836
rect 29196 32824 29224 32920
rect 29546 32892 29552 32904
rect 29507 32864 29552 32892
rect 29546 32852 29552 32864
rect 29604 32852 29610 32904
rect 30561 32895 30619 32901
rect 30561 32861 30573 32895
rect 30607 32892 30619 32895
rect 30742 32892 30748 32904
rect 30607 32864 30748 32892
rect 30607 32861 30619 32864
rect 30561 32855 30619 32861
rect 30742 32852 30748 32864
rect 30800 32852 30806 32904
rect 32125 32895 32183 32901
rect 32125 32861 32137 32895
rect 32171 32892 32183 32895
rect 32306 32892 32312 32904
rect 32171 32864 32312 32892
rect 32171 32861 32183 32864
rect 32125 32855 32183 32861
rect 32306 32852 32312 32864
rect 32364 32852 32370 32904
rect 33962 32892 33968 32904
rect 33923 32864 33968 32892
rect 33962 32852 33968 32864
rect 34020 32852 34026 32904
rect 34238 32892 34244 32904
rect 34199 32864 34244 32892
rect 34238 32852 34244 32864
rect 34296 32852 34302 32904
rect 35526 32892 35532 32904
rect 35487 32864 35532 32892
rect 35526 32852 35532 32864
rect 35584 32852 35590 32904
rect 35802 32892 35808 32904
rect 35763 32864 35808 32892
rect 35802 32852 35808 32864
rect 35860 32852 35866 32904
rect 38930 32892 38936 32904
rect 38891 32864 38936 32892
rect 38930 32852 38936 32864
rect 38988 32852 38994 32904
rect 40497 32895 40555 32901
rect 40497 32861 40509 32895
rect 40543 32892 40555 32895
rect 41230 32892 41236 32904
rect 40543 32864 41236 32892
rect 40543 32861 40555 32864
rect 40497 32855 40555 32861
rect 41230 32852 41236 32864
rect 41288 32852 41294 32904
rect 42245 32895 42303 32901
rect 42245 32861 42257 32895
rect 42291 32892 42303 32895
rect 43990 32892 43996 32904
rect 42291 32864 43996 32892
rect 42291 32861 42303 32864
rect 42245 32855 42303 32861
rect 43990 32852 43996 32864
rect 44048 32852 44054 32904
rect 29052 32796 30046 32824
rect 29052 32784 29058 32796
rect 21358 32756 21364 32768
rect 17368 32728 17448 32756
rect 21319 32728 21364 32756
rect 17368 32716 17374 32728
rect 21358 32716 21364 32728
rect 21416 32716 21422 32768
rect 24118 32756 24124 32768
rect 24079 32728 24124 32756
rect 24118 32716 24124 32728
rect 24176 32716 24182 32768
rect 25222 32756 25228 32768
rect 25183 32728 25228 32756
rect 25222 32716 25228 32728
rect 25280 32716 25286 32768
rect 25547 32759 25605 32765
rect 25547 32725 25559 32759
rect 25593 32756 25605 32759
rect 26510 32756 26516 32768
rect 25593 32728 26516 32756
rect 25593 32725 25605 32728
rect 25547 32719 25605 32725
rect 26510 32716 26516 32728
rect 26568 32716 26574 32768
rect 26602 32716 26608 32768
rect 26660 32756 26666 32768
rect 26789 32759 26847 32765
rect 26789 32756 26801 32759
rect 26660 32728 26801 32756
rect 26660 32716 26666 32728
rect 26789 32725 26801 32728
rect 26835 32725 26847 32759
rect 26789 32719 26847 32725
rect 28629 32759 28687 32765
rect 28629 32725 28641 32759
rect 28675 32756 28687 32759
rect 28810 32756 28816 32768
rect 28675 32728 28816 32756
rect 28675 32725 28687 32728
rect 28629 32719 28687 32725
rect 28810 32716 28816 32728
rect 28868 32756 28874 32768
rect 29086 32756 29092 32768
rect 28868 32728 29092 32756
rect 28868 32716 28874 32728
rect 29086 32716 29092 32728
rect 29144 32716 29150 32768
rect 29914 32756 29920 32768
rect 29875 32728 29920 32756
rect 29914 32716 29920 32728
rect 29972 32716 29978 32768
rect 30018 32756 30046 32796
rect 33134 32784 33140 32836
rect 33192 32824 33198 32836
rect 33778 32824 33784 32836
rect 33192 32796 33784 32824
rect 33192 32784 33198 32796
rect 33778 32784 33784 32796
rect 33836 32784 33842 32836
rect 36538 32824 36544 32836
rect 36451 32796 36544 32824
rect 36538 32784 36544 32796
rect 36596 32824 36602 32836
rect 37921 32827 37979 32833
rect 37921 32824 37933 32827
rect 36596 32796 37933 32824
rect 36596 32784 36602 32796
rect 37921 32793 37933 32796
rect 37967 32793 37979 32827
rect 37921 32787 37979 32793
rect 39206 32784 39212 32836
rect 39264 32824 39270 32836
rect 39485 32827 39543 32833
rect 39485 32824 39497 32827
rect 39264 32796 39497 32824
rect 39264 32784 39270 32796
rect 39485 32793 39497 32796
rect 39531 32824 39543 32827
rect 41049 32827 41107 32833
rect 41049 32824 41061 32827
rect 39531 32796 41061 32824
rect 39531 32793 39543 32796
rect 39485 32787 39543 32793
rect 41049 32793 41061 32796
rect 41095 32793 41107 32827
rect 41049 32787 41107 32793
rect 35618 32756 35624 32768
rect 30018 32728 35624 32756
rect 35618 32716 35624 32728
rect 35676 32756 35682 32768
rect 36722 32756 36728 32768
rect 35676 32728 36728 32756
rect 35676 32716 35682 32728
rect 36722 32716 36728 32728
rect 36780 32756 36786 32768
rect 38838 32756 38844 32768
rect 36780 32728 38844 32756
rect 36780 32716 36786 32728
rect 38838 32716 38844 32728
rect 38896 32716 38902 32768
rect 42058 32756 42064 32768
rect 42019 32728 42064 32756
rect 42058 32716 42064 32728
rect 42116 32716 42122 32768
rect 43901 32759 43959 32765
rect 43901 32725 43913 32759
rect 43947 32756 43959 32759
rect 44082 32756 44088 32768
rect 43947 32728 44088 32756
rect 43947 32725 43959 32728
rect 43901 32719 43959 32725
rect 44082 32716 44088 32728
rect 44140 32716 44146 32768
rect 1104 32666 48852 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 48852 32666
rect 1104 32592 48852 32614
rect 3234 32552 3240 32564
rect 3195 32524 3240 32552
rect 3234 32512 3240 32524
rect 3292 32512 3298 32564
rect 5166 32552 5172 32564
rect 5079 32524 5172 32552
rect 5166 32512 5172 32524
rect 5224 32552 5230 32564
rect 5629 32555 5687 32561
rect 5629 32552 5641 32555
rect 5224 32524 5641 32552
rect 5224 32512 5230 32524
rect 5629 32521 5641 32524
rect 5675 32552 5687 32555
rect 6362 32552 6368 32564
rect 5675 32524 6368 32552
rect 5675 32521 5687 32524
rect 5629 32515 5687 32521
rect 6362 32512 6368 32524
rect 6420 32552 6426 32564
rect 7009 32555 7067 32561
rect 7009 32552 7021 32555
rect 6420 32524 7021 32552
rect 6420 32512 6426 32524
rect 7009 32521 7021 32524
rect 7055 32521 7067 32555
rect 8846 32552 8852 32564
rect 8807 32524 8852 32552
rect 7009 32515 7067 32521
rect 8846 32512 8852 32524
rect 8904 32512 8910 32564
rect 15381 32555 15439 32561
rect 15381 32521 15393 32555
rect 15427 32552 15439 32555
rect 15470 32552 15476 32564
rect 15427 32524 15476 32552
rect 15427 32521 15439 32524
rect 15381 32515 15439 32521
rect 15470 32512 15476 32524
rect 15528 32552 15534 32564
rect 17402 32552 17408 32564
rect 15528 32524 17408 32552
rect 15528 32512 15534 32524
rect 17402 32512 17408 32524
rect 17460 32512 17466 32564
rect 19245 32555 19303 32561
rect 19245 32521 19257 32555
rect 19291 32552 19303 32555
rect 19334 32552 19340 32564
rect 19291 32524 19340 32552
rect 19291 32521 19303 32524
rect 19245 32515 19303 32521
rect 19334 32512 19340 32524
rect 19392 32512 19398 32564
rect 22278 32552 22284 32564
rect 20818 32524 22284 32552
rect 8386 32444 8392 32496
rect 8444 32484 8450 32496
rect 10597 32487 10655 32493
rect 10597 32484 10609 32487
rect 8444 32456 10609 32484
rect 8444 32444 8450 32456
rect 10597 32453 10609 32456
rect 10643 32453 10655 32487
rect 20818 32484 20846 32524
rect 22278 32512 22284 32524
rect 22336 32512 22342 32564
rect 22830 32552 22836 32564
rect 22791 32524 22836 32552
rect 22830 32512 22836 32524
rect 22888 32512 22894 32564
rect 25958 32512 25964 32564
rect 26016 32552 26022 32564
rect 26145 32555 26203 32561
rect 26145 32552 26157 32555
rect 26016 32524 26157 32552
rect 26016 32512 26022 32524
rect 26145 32521 26157 32524
rect 26191 32521 26203 32555
rect 26145 32515 26203 32521
rect 26234 32512 26240 32564
rect 26292 32552 26298 32564
rect 26513 32555 26571 32561
rect 26513 32552 26525 32555
rect 26292 32524 26525 32552
rect 26292 32512 26298 32524
rect 26513 32521 26525 32524
rect 26559 32552 26571 32555
rect 27706 32552 27712 32564
rect 26559 32524 27712 32552
rect 26559 32521 26571 32524
rect 26513 32515 26571 32521
rect 27706 32512 27712 32524
rect 27764 32512 27770 32564
rect 28994 32552 29000 32564
rect 28955 32524 29000 32552
rect 28994 32512 29000 32524
rect 29052 32512 29058 32564
rect 29638 32552 29644 32564
rect 29599 32524 29644 32552
rect 29638 32512 29644 32524
rect 29696 32512 29702 32564
rect 30558 32512 30564 32564
rect 30616 32552 30622 32564
rect 30745 32555 30803 32561
rect 30745 32552 30757 32555
rect 30616 32524 30757 32552
rect 30616 32512 30622 32524
rect 30745 32521 30757 32524
rect 30791 32552 30803 32555
rect 33045 32555 33103 32561
rect 33045 32552 33057 32555
rect 30791 32524 33057 32552
rect 30791 32521 30803 32524
rect 30745 32515 30803 32521
rect 33045 32521 33057 32524
rect 33091 32552 33103 32555
rect 33502 32552 33508 32564
rect 33091 32524 33508 32552
rect 33091 32521 33103 32524
rect 33045 32515 33103 32521
rect 33502 32512 33508 32524
rect 33560 32552 33566 32564
rect 34241 32555 34299 32561
rect 34241 32552 34253 32555
rect 33560 32524 34253 32552
rect 33560 32512 33566 32524
rect 34241 32521 34253 32524
rect 34287 32552 34299 32555
rect 34609 32555 34667 32561
rect 34609 32552 34621 32555
rect 34287 32524 34621 32552
rect 34287 32521 34299 32524
rect 34241 32515 34299 32521
rect 34609 32521 34621 32524
rect 34655 32521 34667 32555
rect 34609 32515 34667 32521
rect 35526 32512 35532 32564
rect 35584 32552 35590 32564
rect 36817 32555 36875 32561
rect 36817 32552 36829 32555
rect 35584 32524 36829 32552
rect 35584 32512 35590 32524
rect 36817 32521 36829 32524
rect 36863 32521 36875 32555
rect 36817 32515 36875 32521
rect 38289 32555 38347 32561
rect 38289 32521 38301 32555
rect 38335 32552 38347 32555
rect 39022 32552 39028 32564
rect 38335 32524 39028 32552
rect 38335 32521 38347 32524
rect 38289 32515 38347 32521
rect 39022 32512 39028 32524
rect 39080 32512 39086 32564
rect 39850 32552 39856 32564
rect 39811 32524 39856 32552
rect 39850 32512 39856 32524
rect 39908 32512 39914 32564
rect 40313 32555 40371 32561
rect 40313 32521 40325 32555
rect 40359 32552 40371 32555
rect 40402 32552 40408 32564
rect 40359 32524 40408 32552
rect 40359 32521 40371 32524
rect 40313 32515 40371 32521
rect 40402 32512 40408 32524
rect 40460 32512 40466 32564
rect 10597 32447 10655 32453
rect 18386 32456 20846 32484
rect 21177 32487 21235 32493
rect 4614 32416 4620 32428
rect 4575 32388 4620 32416
rect 4614 32376 4620 32388
rect 4672 32376 4678 32428
rect 7929 32419 7987 32425
rect 7929 32385 7941 32419
rect 7975 32416 7987 32419
rect 8294 32416 8300 32428
rect 7975 32388 8300 32416
rect 7975 32385 7987 32388
rect 7929 32379 7987 32385
rect 8294 32376 8300 32388
rect 8352 32376 8358 32428
rect 14642 32416 14648 32428
rect 14603 32388 14648 32416
rect 14642 32376 14648 32388
rect 14700 32376 14706 32428
rect 15286 32376 15292 32428
rect 15344 32416 15350 32428
rect 16393 32419 16451 32425
rect 16393 32416 16405 32419
rect 15344 32388 16405 32416
rect 15344 32376 15350 32388
rect 16393 32385 16405 32388
rect 16439 32416 16451 32419
rect 17037 32419 17095 32425
rect 17037 32416 17049 32419
rect 16439 32388 17049 32416
rect 16439 32385 16451 32388
rect 16393 32379 16451 32385
rect 17037 32385 17049 32388
rect 17083 32385 17095 32419
rect 17037 32379 17095 32385
rect 17865 32419 17923 32425
rect 17865 32385 17877 32419
rect 17911 32416 17923 32419
rect 18386 32416 18414 32456
rect 21177 32453 21189 32487
rect 21223 32484 21235 32487
rect 22094 32484 22100 32496
rect 21223 32456 22100 32484
rect 21223 32453 21235 32456
rect 21177 32447 21235 32453
rect 22094 32444 22100 32456
rect 22152 32444 22158 32496
rect 24673 32487 24731 32493
rect 24673 32484 24685 32487
rect 24038 32456 24685 32484
rect 18598 32416 18604 32428
rect 17911 32388 18414 32416
rect 18559 32388 18604 32416
rect 17911 32385 17923 32388
rect 17865 32379 17923 32385
rect 3234 32308 3240 32360
rect 3292 32348 3298 32360
rect 3973 32351 4031 32357
rect 3973 32348 3985 32351
rect 3292 32320 3985 32348
rect 3292 32308 3298 32320
rect 3973 32317 3985 32320
rect 4019 32348 4031 32351
rect 4065 32351 4123 32357
rect 4065 32348 4077 32351
rect 4019 32320 4077 32348
rect 4019 32317 4031 32320
rect 3973 32311 4031 32317
rect 4065 32317 4077 32320
rect 4111 32317 4123 32351
rect 4522 32348 4528 32360
rect 4435 32320 4528 32348
rect 4065 32311 4123 32317
rect 4522 32308 4528 32320
rect 4580 32348 4586 32360
rect 5166 32348 5172 32360
rect 4580 32320 5172 32348
rect 4580 32308 4586 32320
rect 5166 32308 5172 32320
rect 5224 32308 5230 32360
rect 5788 32351 5846 32357
rect 5788 32317 5800 32351
rect 5834 32348 5846 32351
rect 6178 32348 6184 32360
rect 5834 32320 6184 32348
rect 5834 32317 5846 32320
rect 5788 32311 5846 32317
rect 6178 32308 6184 32320
rect 6236 32308 6242 32360
rect 6641 32351 6699 32357
rect 6641 32317 6653 32351
rect 6687 32348 6699 32351
rect 6825 32351 6883 32357
rect 6825 32348 6837 32351
rect 6687 32320 6837 32348
rect 6687 32317 6699 32320
rect 6641 32311 6699 32317
rect 6825 32317 6837 32320
rect 6871 32348 6883 32351
rect 7374 32348 7380 32360
rect 6871 32320 7380 32348
rect 6871 32317 6883 32320
rect 6825 32311 6883 32317
rect 7374 32308 7380 32320
rect 7432 32308 7438 32360
rect 9674 32348 9680 32360
rect 9635 32320 9680 32348
rect 9674 32308 9680 32320
rect 9732 32308 9738 32360
rect 11146 32308 11152 32360
rect 11204 32348 11210 32360
rect 12161 32351 12219 32357
rect 12161 32348 12173 32351
rect 11204 32320 12173 32348
rect 11204 32308 11210 32320
rect 12161 32317 12173 32320
rect 12207 32348 12219 32351
rect 12437 32351 12495 32357
rect 12437 32348 12449 32351
rect 12207 32320 12449 32348
rect 12207 32317 12219 32320
rect 12161 32311 12219 32317
rect 12437 32317 12449 32320
rect 12483 32317 12495 32351
rect 12986 32348 12992 32360
rect 12947 32320 12992 32348
rect 12437 32311 12495 32317
rect 12986 32308 12992 32320
rect 13044 32308 13050 32360
rect 13998 32348 14004 32360
rect 13911 32320 14004 32348
rect 13998 32308 14004 32320
rect 14056 32348 14062 32360
rect 14093 32351 14151 32357
rect 14093 32348 14105 32351
rect 14056 32320 14105 32348
rect 14056 32308 14062 32320
rect 14093 32317 14105 32320
rect 14139 32317 14151 32351
rect 14093 32311 14151 32317
rect 14553 32351 14611 32357
rect 14553 32317 14565 32351
rect 14599 32317 14611 32351
rect 15654 32348 15660 32360
rect 15615 32320 15660 32348
rect 14553 32311 14611 32317
rect 7469 32283 7527 32289
rect 7469 32249 7481 32283
rect 7515 32280 7527 32283
rect 7834 32280 7840 32292
rect 7515 32252 7840 32280
rect 7515 32249 7527 32252
rect 7469 32243 7527 32249
rect 7834 32240 7840 32252
rect 7892 32280 7898 32292
rect 8291 32283 8349 32289
rect 8291 32280 8303 32283
rect 7892 32252 8303 32280
rect 7892 32240 7898 32252
rect 8291 32249 8303 32252
rect 8337 32280 8349 32283
rect 9217 32283 9275 32289
rect 9217 32280 9229 32283
rect 8337 32252 9229 32280
rect 8337 32249 8349 32252
rect 8291 32243 8349 32249
rect 9217 32249 9229 32252
rect 9263 32280 9275 32283
rect 9585 32283 9643 32289
rect 9585 32280 9597 32283
rect 9263 32252 9597 32280
rect 9263 32249 9275 32252
rect 9217 32243 9275 32249
rect 9585 32249 9597 32252
rect 9631 32280 9643 32283
rect 9998 32283 10056 32289
rect 9998 32280 10010 32283
rect 9631 32252 10010 32280
rect 9631 32249 9643 32252
rect 9585 32243 9643 32249
rect 9998 32249 10010 32252
rect 10044 32280 10056 32283
rect 11422 32280 11428 32292
rect 10044 32252 11428 32280
rect 10044 32249 10056 32252
rect 9998 32243 10056 32249
rect 11422 32240 11428 32252
rect 11480 32240 11486 32292
rect 11882 32280 11888 32292
rect 11795 32252 11888 32280
rect 11882 32240 11888 32252
rect 11940 32280 11946 32292
rect 11940 32252 12296 32280
rect 11940 32240 11946 32252
rect 3510 32212 3516 32224
rect 3471 32184 3516 32212
rect 3510 32172 3516 32184
rect 3568 32172 3574 32224
rect 5859 32215 5917 32221
rect 5859 32181 5871 32215
rect 5905 32212 5917 32215
rect 6086 32212 6092 32224
rect 5905 32184 6092 32212
rect 5905 32181 5917 32184
rect 5859 32175 5917 32181
rect 6086 32172 6092 32184
rect 6144 32172 6150 32224
rect 6270 32212 6276 32224
rect 6231 32184 6276 32212
rect 6270 32172 6276 32184
rect 6328 32172 6334 32224
rect 10410 32172 10416 32224
rect 10468 32212 10474 32224
rect 10873 32215 10931 32221
rect 10873 32212 10885 32215
rect 10468 32184 10885 32212
rect 10468 32172 10474 32184
rect 10873 32181 10885 32184
rect 10919 32181 10931 32215
rect 12268 32212 12296 32252
rect 14182 32240 14188 32292
rect 14240 32280 14246 32292
rect 14568 32280 14596 32311
rect 15654 32308 15660 32320
rect 15712 32308 15718 32360
rect 18340 32357 18368 32388
rect 18598 32376 18604 32388
rect 18656 32376 18662 32428
rect 19797 32419 19855 32425
rect 19797 32385 19809 32419
rect 19843 32416 19855 32419
rect 20254 32416 20260 32428
rect 19843 32388 20260 32416
rect 19843 32385 19855 32388
rect 19797 32379 19855 32385
rect 20254 32376 20260 32388
rect 20312 32376 20318 32428
rect 21726 32416 21732 32428
rect 21687 32388 21732 32416
rect 21726 32376 21732 32388
rect 21784 32376 21790 32428
rect 23753 32419 23811 32425
rect 23753 32385 23765 32419
rect 23799 32416 23811 32419
rect 24038 32416 24066 32456
rect 24673 32453 24685 32456
rect 24719 32484 24731 32487
rect 26970 32484 26976 32496
rect 24719 32456 26976 32484
rect 24719 32453 24731 32456
rect 24673 32447 24731 32453
rect 26970 32444 26976 32456
rect 27028 32484 27034 32496
rect 27617 32487 27675 32493
rect 27617 32484 27629 32487
rect 27028 32456 27629 32484
rect 27028 32444 27034 32456
rect 27617 32453 27629 32456
rect 27663 32453 27675 32487
rect 28074 32484 28080 32496
rect 27987 32456 28080 32484
rect 27617 32447 27675 32453
rect 28074 32444 28080 32456
rect 28132 32484 28138 32496
rect 32122 32484 32128 32496
rect 28132 32456 32128 32484
rect 28132 32444 28138 32456
rect 32122 32444 32128 32456
rect 32180 32444 32186 32496
rect 35618 32484 35624 32496
rect 35579 32456 35624 32484
rect 35618 32444 35624 32456
rect 35676 32444 35682 32496
rect 39531 32487 39589 32493
rect 39531 32453 39543 32487
rect 39577 32484 39589 32487
rect 42058 32484 42064 32496
rect 39577 32456 42064 32484
rect 39577 32453 39589 32456
rect 39531 32447 39589 32453
rect 42058 32444 42064 32456
rect 42116 32484 42122 32496
rect 44269 32487 44327 32493
rect 44269 32484 44281 32487
rect 42116 32456 42196 32484
rect 42116 32444 42122 32456
rect 24210 32416 24216 32428
rect 23799 32388 24066 32416
rect 24171 32388 24216 32416
rect 23799 32385 23811 32388
rect 23753 32379 23811 32385
rect 24210 32376 24216 32388
rect 24268 32376 24274 32428
rect 26510 32376 26516 32428
rect 26568 32416 26574 32428
rect 27065 32419 27123 32425
rect 27065 32416 27077 32419
rect 26568 32388 27077 32416
rect 26568 32376 26574 32388
rect 27065 32385 27077 32388
rect 27111 32416 27123 32419
rect 27522 32416 27528 32428
rect 27111 32388 27528 32416
rect 27111 32385 27123 32388
rect 27065 32379 27123 32385
rect 27522 32376 27528 32388
rect 27580 32376 27586 32428
rect 29825 32419 29883 32425
rect 29825 32385 29837 32419
rect 29871 32416 29883 32419
rect 29914 32416 29920 32428
rect 29871 32388 29920 32416
rect 29871 32385 29883 32388
rect 29825 32379 29883 32385
rect 29914 32376 29920 32388
rect 29972 32376 29978 32428
rect 32398 32416 32404 32428
rect 30392 32388 32404 32416
rect 16209 32351 16267 32357
rect 16209 32317 16221 32351
rect 16255 32348 16267 32351
rect 16669 32351 16727 32357
rect 16669 32348 16681 32351
rect 16255 32320 16681 32348
rect 16255 32317 16267 32320
rect 16209 32311 16267 32317
rect 16669 32317 16681 32320
rect 16715 32317 16727 32351
rect 16669 32311 16727 32317
rect 18325 32351 18383 32357
rect 18325 32317 18337 32351
rect 18371 32317 18383 32351
rect 18506 32348 18512 32360
rect 18419 32320 18512 32348
rect 18325 32311 18383 32317
rect 16224 32280 16252 32311
rect 18506 32308 18512 32320
rect 18564 32308 18570 32360
rect 25222 32348 25228 32360
rect 25183 32320 25228 32348
rect 25222 32308 25228 32320
rect 25280 32308 25286 32360
rect 14240 32252 16252 32280
rect 14240 32240 14246 32252
rect 17862 32240 17868 32292
rect 17920 32280 17926 32292
rect 18524 32280 18552 32308
rect 17920 32252 18552 32280
rect 17920 32240 17926 32252
rect 19886 32240 19892 32292
rect 19944 32280 19950 32292
rect 20438 32280 20444 32292
rect 19944 32252 19989 32280
rect 20399 32252 20444 32280
rect 19944 32240 19950 32252
rect 20438 32240 20444 32252
rect 20496 32240 20502 32292
rect 20809 32283 20867 32289
rect 20809 32249 20821 32283
rect 20855 32280 20867 32283
rect 21174 32280 21180 32292
rect 20855 32252 21180 32280
rect 20855 32249 20867 32252
rect 20809 32243 20867 32249
rect 21174 32240 21180 32252
rect 21232 32280 21238 32292
rect 21361 32283 21419 32289
rect 21361 32280 21373 32283
rect 21232 32252 21373 32280
rect 21232 32240 21238 32252
rect 21361 32249 21373 32252
rect 21407 32249 21419 32283
rect 21361 32243 21419 32249
rect 21450 32240 21456 32292
rect 21508 32280 21514 32292
rect 23845 32283 23903 32289
rect 21508 32252 21553 32280
rect 21508 32240 21514 32252
rect 23845 32249 23857 32283
rect 23891 32280 23903 32283
rect 24118 32280 24124 32292
rect 23891 32252 24124 32280
rect 23891 32249 23903 32252
rect 23845 32243 23903 32249
rect 24118 32240 24124 32252
rect 24176 32240 24182 32292
rect 25041 32283 25099 32289
rect 25041 32280 25053 32283
rect 24596 32252 25053 32280
rect 12529 32215 12587 32221
rect 12529 32212 12541 32215
rect 12268 32184 12541 32212
rect 10873 32175 10931 32181
rect 12529 32181 12541 32184
rect 12575 32181 12587 32215
rect 13446 32212 13452 32224
rect 13407 32184 13452 32212
rect 12529 32175 12587 32181
rect 13446 32172 13452 32184
rect 13504 32172 13510 32224
rect 19613 32215 19671 32221
rect 19613 32181 19625 32215
rect 19659 32212 19671 32215
rect 19904 32212 19932 32240
rect 22370 32212 22376 32224
rect 19659 32184 19932 32212
rect 22331 32184 22376 32212
rect 19659 32181 19671 32184
rect 19613 32175 19671 32181
rect 22370 32172 22376 32184
rect 22428 32172 22434 32224
rect 23014 32172 23020 32224
rect 23072 32212 23078 32224
rect 23201 32215 23259 32221
rect 23201 32212 23213 32215
rect 23072 32184 23213 32212
rect 23072 32172 23078 32184
rect 23201 32181 23213 32184
rect 23247 32212 23259 32215
rect 23290 32212 23296 32224
rect 23247 32184 23296 32212
rect 23247 32181 23259 32184
rect 23201 32175 23259 32181
rect 23290 32172 23296 32184
rect 23348 32212 23354 32224
rect 24596 32212 24624 32252
rect 25041 32249 25053 32252
rect 25087 32280 25099 32283
rect 25546 32283 25604 32289
rect 25546 32280 25558 32283
rect 25087 32252 25558 32280
rect 25087 32249 25099 32252
rect 25041 32243 25099 32249
rect 25546 32249 25558 32252
rect 25592 32249 25604 32283
rect 25546 32243 25604 32249
rect 26694 32240 26700 32292
rect 26752 32280 26758 32292
rect 27157 32283 27215 32289
rect 27157 32280 27169 32283
rect 26752 32252 27169 32280
rect 26752 32240 26758 32252
rect 27157 32249 27169 32252
rect 27203 32249 27215 32283
rect 27157 32243 27215 32249
rect 29638 32240 29644 32292
rect 29696 32280 29702 32292
rect 30146 32283 30204 32289
rect 30146 32280 30158 32283
rect 29696 32252 30158 32280
rect 29696 32240 29702 32252
rect 30146 32249 30158 32252
rect 30192 32280 30204 32283
rect 30392 32280 30420 32388
rect 32398 32376 32404 32388
rect 32456 32416 32462 32428
rect 32585 32419 32643 32425
rect 32585 32416 32597 32419
rect 32456 32388 32597 32416
rect 32456 32376 32462 32388
rect 32585 32385 32597 32388
rect 32631 32385 32643 32419
rect 32585 32379 32643 32385
rect 33321 32419 33379 32425
rect 33321 32385 33333 32419
rect 33367 32416 33379 32419
rect 33410 32416 33416 32428
rect 33367 32388 33416 32416
rect 33367 32385 33379 32388
rect 33321 32379 33379 32385
rect 33410 32376 33416 32388
rect 33468 32376 33474 32428
rect 33778 32376 33784 32428
rect 33836 32416 33842 32428
rect 33836 32388 33881 32416
rect 33836 32376 33842 32388
rect 31481 32351 31539 32357
rect 31481 32317 31493 32351
rect 31527 32348 31539 32351
rect 31846 32348 31852 32360
rect 31527 32320 31852 32348
rect 31527 32317 31539 32320
rect 31481 32311 31539 32317
rect 31846 32308 31852 32320
rect 31904 32308 31910 32360
rect 32030 32348 32036 32360
rect 31991 32320 32036 32348
rect 32030 32308 32036 32320
rect 32088 32308 32094 32360
rect 35636 32348 35664 32444
rect 40589 32419 40647 32425
rect 40589 32385 40601 32419
rect 40635 32416 40647 32419
rect 40770 32416 40776 32428
rect 40635 32388 40776 32416
rect 40635 32385 40647 32388
rect 40589 32379 40647 32385
rect 40770 32376 40776 32388
rect 40828 32416 40834 32428
rect 42168 32425 42196 32456
rect 42766 32456 44281 32484
rect 41509 32419 41567 32425
rect 41509 32416 41521 32419
rect 40828 32388 41521 32416
rect 40828 32376 40834 32388
rect 41509 32385 41521 32388
rect 41555 32385 41567 32419
rect 41509 32379 41567 32385
rect 42153 32419 42211 32425
rect 42153 32385 42165 32419
rect 42199 32385 42211 32419
rect 42426 32416 42432 32428
rect 42387 32388 42432 32416
rect 42153 32379 42211 32385
rect 42426 32376 42432 32388
rect 42484 32416 42490 32428
rect 42766 32416 42794 32456
rect 44269 32453 44281 32456
rect 44315 32484 44327 32487
rect 44542 32484 44548 32496
rect 44315 32456 44548 32484
rect 44315 32453 44327 32456
rect 44269 32447 44327 32453
rect 44542 32444 44548 32456
rect 44600 32444 44606 32496
rect 42484 32388 42794 32416
rect 42484 32376 42490 32388
rect 43530 32376 43536 32428
rect 43588 32416 43594 32428
rect 43717 32419 43775 32425
rect 43717 32416 43729 32419
rect 43588 32388 43729 32416
rect 43588 32376 43594 32388
rect 43717 32385 43729 32388
rect 43763 32416 43775 32419
rect 44637 32419 44695 32425
rect 44637 32416 44649 32419
rect 43763 32388 44649 32416
rect 43763 32385 43775 32388
rect 43717 32379 43775 32385
rect 44637 32385 44649 32388
rect 44683 32385 44695 32419
rect 44637 32379 44695 32385
rect 35805 32351 35863 32357
rect 35805 32348 35817 32351
rect 35636 32320 35817 32348
rect 35805 32317 35817 32320
rect 35851 32317 35863 32351
rect 35805 32311 35863 32317
rect 36357 32351 36415 32357
rect 36357 32317 36369 32351
rect 36403 32348 36415 32351
rect 36446 32348 36452 32360
rect 36403 32320 36452 32348
rect 36403 32317 36415 32320
rect 36357 32311 36415 32317
rect 30192 32252 30420 32280
rect 30192 32249 30204 32252
rect 30146 32243 30204 32249
rect 30466 32240 30472 32292
rect 30524 32280 30530 32292
rect 30650 32280 30656 32292
rect 30524 32252 30656 32280
rect 30524 32240 30530 32252
rect 30650 32240 30656 32252
rect 30708 32280 30714 32292
rect 31021 32283 31079 32289
rect 31021 32280 31033 32283
rect 30708 32252 31033 32280
rect 30708 32240 30714 32252
rect 31021 32249 31033 32252
rect 31067 32249 31079 32283
rect 31021 32243 31079 32249
rect 28626 32212 28632 32224
rect 23348 32184 24624 32212
rect 28587 32184 28632 32212
rect 23348 32172 23354 32184
rect 28626 32172 28632 32184
rect 28684 32172 28690 32224
rect 31864 32212 31892 32308
rect 32306 32280 32312 32292
rect 32267 32252 32312 32280
rect 32306 32240 32312 32252
rect 32364 32240 32370 32292
rect 33413 32283 33471 32289
rect 33413 32249 33425 32283
rect 33459 32280 33471 32283
rect 33502 32280 33508 32292
rect 33459 32252 33508 32280
rect 33459 32249 33471 32252
rect 33413 32243 33471 32249
rect 33502 32240 33508 32252
rect 33560 32240 33566 32292
rect 35345 32283 35403 32289
rect 35345 32249 35357 32283
rect 35391 32280 35403 32283
rect 36372 32280 36400 32311
rect 36446 32308 36452 32320
rect 36504 32308 36510 32360
rect 36541 32351 36599 32357
rect 36541 32317 36553 32351
rect 36587 32348 36599 32351
rect 37366 32348 37372 32360
rect 36587 32320 37372 32348
rect 36587 32317 36599 32320
rect 36541 32311 36599 32317
rect 37366 32308 37372 32320
rect 37424 32308 37430 32360
rect 39460 32351 39518 32357
rect 39460 32317 39472 32351
rect 39506 32348 39518 32351
rect 39850 32348 39856 32360
rect 39506 32320 39856 32348
rect 39506 32317 39518 32320
rect 39460 32311 39518 32317
rect 39850 32308 39856 32320
rect 39908 32308 39914 32360
rect 35391 32252 36400 32280
rect 37731 32283 37789 32289
rect 35391 32249 35403 32252
rect 35345 32243 35403 32249
rect 37731 32249 37743 32283
rect 37777 32249 37789 32283
rect 37731 32243 37789 32249
rect 33134 32212 33140 32224
rect 31864 32184 33140 32212
rect 33134 32172 33140 32184
rect 33192 32172 33198 32224
rect 37277 32215 37335 32221
rect 37277 32181 37289 32215
rect 37323 32212 37335 32215
rect 37746 32212 37774 32243
rect 40402 32240 40408 32292
rect 40460 32280 40466 32292
rect 40681 32283 40739 32289
rect 40681 32280 40693 32283
rect 40460 32252 40693 32280
rect 40460 32240 40466 32252
rect 40681 32249 40693 32252
rect 40727 32249 40739 32283
rect 41230 32280 41236 32292
rect 41191 32252 41236 32280
rect 40681 32243 40739 32249
rect 37826 32212 37832 32224
rect 37323 32184 37832 32212
rect 37323 32181 37335 32184
rect 37277 32175 37335 32181
rect 37826 32172 37832 32184
rect 37884 32172 37890 32224
rect 38657 32215 38715 32221
rect 38657 32181 38669 32215
rect 38703 32212 38715 32215
rect 38746 32212 38752 32224
rect 38703 32184 38752 32212
rect 38703 32181 38715 32184
rect 38657 32175 38715 32181
rect 38746 32172 38752 32184
rect 38804 32172 38810 32224
rect 40696 32212 40724 32243
rect 41230 32240 41236 32252
rect 41288 32240 41294 32292
rect 42245 32283 42303 32289
rect 42245 32280 42257 32283
rect 41892 32252 42257 32280
rect 41892 32221 41920 32252
rect 42245 32249 42257 32252
rect 42291 32249 42303 32283
rect 42245 32243 42303 32249
rect 43809 32283 43867 32289
rect 43809 32249 43821 32283
rect 43855 32280 43867 32283
rect 44082 32280 44088 32292
rect 43855 32252 44088 32280
rect 43855 32249 43867 32252
rect 43809 32243 43867 32249
rect 44082 32240 44088 32252
rect 44140 32240 44146 32292
rect 41877 32215 41935 32221
rect 41877 32212 41889 32215
rect 40696 32184 41889 32212
rect 41877 32181 41889 32184
rect 41923 32181 41935 32215
rect 43346 32212 43352 32224
rect 43307 32184 43352 32212
rect 41877 32175 41935 32181
rect 43346 32172 43352 32184
rect 43404 32172 43410 32224
rect 1104 32122 48852 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 48852 32122
rect 1104 32048 48852 32070
rect 9493 32011 9551 32017
rect 9493 31977 9505 32011
rect 9539 32008 9551 32011
rect 9674 32008 9680 32020
rect 9539 31980 9680 32008
rect 9539 31977 9551 31980
rect 9493 31971 9551 31977
rect 9674 31968 9680 31980
rect 9732 32008 9738 32020
rect 9769 32011 9827 32017
rect 9769 32008 9781 32011
rect 9732 31980 9781 32008
rect 9732 31968 9738 31980
rect 9769 31977 9781 31980
rect 9815 31977 9827 32011
rect 9769 31971 9827 31977
rect 11238 31968 11244 32020
rect 11296 32008 11302 32020
rect 11425 32011 11483 32017
rect 11425 32008 11437 32011
rect 11296 31980 11437 32008
rect 11296 31968 11302 31980
rect 11425 31977 11437 31980
rect 11471 31977 11483 32011
rect 14182 32008 14188 32020
rect 14143 31980 14188 32008
rect 11425 31971 11483 31977
rect 14182 31968 14188 31980
rect 14240 31968 14246 32020
rect 14826 31968 14832 32020
rect 14884 32008 14890 32020
rect 15654 32008 15660 32020
rect 14884 31980 15660 32008
rect 14884 31968 14890 31980
rect 15654 31968 15660 31980
rect 15712 31968 15718 32020
rect 17310 32008 17316 32020
rect 17271 31980 17316 32008
rect 17310 31968 17316 31980
rect 17368 31968 17374 32020
rect 22094 32008 22100 32020
rect 22055 31980 22100 32008
rect 22094 31968 22100 31980
rect 22152 31968 22158 32020
rect 23014 32008 23020 32020
rect 22975 31980 23020 32008
rect 23014 31968 23020 31980
rect 23072 31968 23078 32020
rect 23937 32011 23995 32017
rect 23937 31977 23949 32011
rect 23983 32008 23995 32011
rect 24118 32008 24124 32020
rect 23983 31980 24124 32008
rect 23983 31977 23995 31980
rect 23937 31971 23995 31977
rect 24118 31968 24124 31980
rect 24176 31968 24182 32020
rect 24486 31968 24492 32020
rect 24544 32008 24550 32020
rect 27522 32008 27528 32020
rect 24544 31980 27292 32008
rect 27483 31980 27528 32008
rect 24544 31968 24550 31980
rect 4801 31943 4859 31949
rect 4801 31909 4813 31943
rect 4847 31940 4859 31943
rect 4890 31940 4896 31952
rect 4847 31912 4896 31940
rect 4847 31909 4859 31912
rect 4801 31903 4859 31909
rect 4890 31900 4896 31912
rect 4948 31900 4954 31952
rect 8711 31943 8769 31949
rect 8711 31909 8723 31943
rect 8757 31940 8769 31943
rect 12066 31940 12072 31952
rect 8757 31912 12072 31940
rect 8757 31909 8769 31912
rect 8711 31903 8769 31909
rect 12066 31900 12072 31912
rect 12124 31900 12130 31952
rect 19426 31940 19432 31952
rect 19387 31912 19432 31940
rect 19426 31900 19432 31912
rect 19484 31900 19490 31952
rect 21174 31900 21180 31952
rect 21232 31940 21238 31952
rect 21683 31943 21741 31949
rect 21683 31940 21695 31943
rect 21232 31912 21695 31940
rect 21232 31900 21238 31912
rect 21683 31909 21695 31912
rect 21729 31909 21741 31943
rect 24578 31940 24584 31952
rect 21683 31903 21741 31909
rect 23584 31912 24584 31940
rect 3786 31832 3792 31884
rect 3844 31872 3850 31884
rect 4065 31875 4123 31881
rect 4065 31872 4077 31875
rect 3844 31844 4077 31872
rect 3844 31832 3850 31844
rect 4065 31841 4077 31844
rect 4111 31841 4123 31875
rect 4522 31872 4528 31884
rect 4483 31844 4528 31872
rect 4065 31835 4123 31841
rect 4522 31832 4528 31844
rect 4580 31832 4586 31884
rect 5696 31875 5754 31881
rect 5696 31841 5708 31875
rect 5742 31872 5754 31875
rect 5810 31872 5816 31884
rect 5742 31844 5816 31872
rect 5742 31841 5754 31844
rect 5696 31835 5754 31841
rect 5810 31832 5816 31844
rect 5868 31832 5874 31884
rect 6362 31832 6368 31884
rect 6420 31872 6426 31884
rect 6917 31875 6975 31881
rect 6917 31872 6929 31875
rect 6420 31844 6929 31872
rect 6420 31832 6426 31844
rect 6917 31841 6929 31844
rect 6963 31841 6975 31875
rect 7374 31872 7380 31884
rect 7335 31844 7380 31872
rect 6917 31835 6975 31841
rect 7374 31832 7380 31844
rect 7432 31832 7438 31884
rect 8386 31832 8392 31884
rect 8444 31872 8450 31884
rect 8608 31875 8666 31881
rect 8608 31872 8620 31875
rect 8444 31844 8620 31872
rect 8444 31832 8450 31844
rect 8608 31841 8620 31844
rect 8654 31841 8666 31875
rect 8608 31835 8666 31841
rect 9582 31832 9588 31884
rect 9640 31872 9646 31884
rect 9677 31875 9735 31881
rect 9677 31872 9689 31875
rect 9640 31844 9689 31872
rect 9640 31832 9646 31844
rect 9677 31841 9689 31844
rect 9723 31841 9735 31875
rect 10134 31872 10140 31884
rect 10095 31844 10140 31872
rect 9677 31835 9735 31841
rect 10134 31832 10140 31844
rect 10192 31832 10198 31884
rect 11422 31872 11428 31884
rect 11383 31844 11428 31872
rect 11422 31832 11428 31844
rect 11480 31832 11486 31884
rect 11885 31875 11943 31881
rect 11885 31841 11897 31875
rect 11931 31872 11943 31875
rect 12250 31872 12256 31884
rect 11931 31844 12256 31872
rect 11931 31841 11943 31844
rect 11885 31835 11943 31841
rect 12250 31832 12256 31844
rect 12308 31832 12314 31884
rect 13262 31832 13268 31884
rect 13320 31872 13326 31884
rect 13449 31875 13507 31881
rect 13449 31872 13461 31875
rect 13320 31844 13461 31872
rect 13320 31832 13326 31844
rect 13449 31841 13461 31844
rect 13495 31841 13507 31875
rect 13449 31835 13507 31841
rect 16092 31875 16150 31881
rect 16092 31841 16104 31875
rect 16138 31872 16150 31875
rect 16482 31872 16488 31884
rect 16138 31844 16488 31872
rect 16138 31841 16150 31844
rect 16092 31835 16150 31841
rect 16482 31832 16488 31844
rect 16540 31832 16546 31884
rect 17310 31872 17316 31884
rect 17271 31844 17316 31872
rect 17310 31832 17316 31844
rect 17368 31832 17374 31884
rect 17589 31875 17647 31881
rect 17589 31841 17601 31875
rect 17635 31872 17647 31875
rect 17862 31872 17868 31884
rect 17635 31844 17868 31872
rect 17635 31841 17647 31844
rect 17589 31835 17647 31841
rect 17862 31832 17868 31844
rect 17920 31832 17926 31884
rect 21453 31875 21511 31881
rect 21453 31841 21465 31875
rect 21499 31872 21511 31875
rect 21542 31872 21548 31884
rect 21499 31844 21548 31872
rect 21499 31841 21511 31844
rect 21453 31835 21511 31841
rect 21542 31832 21548 31844
rect 21600 31832 21606 31884
rect 23584 31881 23612 31912
rect 24578 31900 24584 31912
rect 24636 31900 24642 31952
rect 26694 31940 26700 31952
rect 26655 31912 26700 31940
rect 26694 31900 26700 31912
rect 26752 31900 26758 31952
rect 27264 31949 27292 31980
rect 27522 31968 27528 31980
rect 27580 31968 27586 32020
rect 29638 31968 29644 32020
rect 29696 32008 29702 32020
rect 29917 32011 29975 32017
rect 29917 32008 29929 32011
rect 29696 31980 29929 32008
rect 29696 31968 29702 31980
rect 29917 31977 29929 31980
rect 29963 31977 29975 32011
rect 30466 32008 30472 32020
rect 30427 31980 30472 32008
rect 29917 31971 29975 31977
rect 30466 31968 30472 31980
rect 30524 31968 30530 32020
rect 30742 32008 30748 32020
rect 30703 31980 30748 32008
rect 30742 31968 30748 31980
rect 30800 31968 30806 32020
rect 32306 32008 32312 32020
rect 32267 31980 32312 32008
rect 32306 31968 32312 31980
rect 32364 31968 32370 32020
rect 32999 32011 33057 32017
rect 32999 31977 33011 32011
rect 33045 32008 33057 32011
rect 33781 32011 33839 32017
rect 33781 32008 33793 32011
rect 33045 31980 33793 32008
rect 33045 31977 33057 31980
rect 32999 31971 33057 31977
rect 33781 31977 33793 31980
rect 33827 32008 33839 32011
rect 33962 32008 33968 32020
rect 33827 31980 33968 32008
rect 33827 31977 33839 31980
rect 33781 31971 33839 31977
rect 33962 31968 33968 31980
rect 34020 31968 34026 32020
rect 37366 32008 37372 32020
rect 37327 31980 37372 32008
rect 37366 31968 37372 31980
rect 37424 31968 37430 32020
rect 38657 32011 38715 32017
rect 38657 31977 38669 32011
rect 38703 32008 38715 32011
rect 40586 32008 40592 32020
rect 38703 31980 40592 32008
rect 38703 31977 38715 31980
rect 38657 31971 38715 31977
rect 40586 31968 40592 31980
rect 40644 32008 40650 32020
rect 40681 32011 40739 32017
rect 40681 32008 40693 32011
rect 40644 31980 40693 32008
rect 40644 31968 40650 31980
rect 40681 31977 40693 31980
rect 40727 31977 40739 32011
rect 40681 31971 40739 31977
rect 42429 32011 42487 32017
rect 42429 31977 42441 32011
rect 42475 31977 42487 32011
rect 42429 31971 42487 31977
rect 27249 31943 27307 31949
rect 27249 31909 27261 31943
rect 27295 31909 27307 31943
rect 33410 31940 33416 31952
rect 33371 31912 33416 31940
rect 27249 31903 27307 31909
rect 33410 31900 33416 31912
rect 33468 31900 33474 31952
rect 33502 31900 33508 31952
rect 33560 31940 33566 31952
rect 34057 31943 34115 31949
rect 34057 31940 34069 31943
rect 33560 31912 34069 31940
rect 33560 31900 33566 31912
rect 34057 31909 34069 31912
rect 34103 31909 34115 31943
rect 37734 31940 37740 31952
rect 34057 31903 34115 31909
rect 36096 31912 37740 31940
rect 23569 31875 23627 31881
rect 23569 31841 23581 31875
rect 23615 31841 23627 31875
rect 29546 31872 29552 31884
rect 29507 31844 29552 31872
rect 23569 31835 23627 31841
rect 29546 31832 29552 31844
rect 29604 31832 29610 31884
rect 32582 31832 32588 31884
rect 32640 31872 32646 31884
rect 32896 31875 32954 31881
rect 32896 31872 32908 31875
rect 32640 31844 32908 31872
rect 32640 31832 32646 31844
rect 32896 31841 32908 31844
rect 32942 31841 32954 31875
rect 32896 31835 32954 31841
rect 35342 31832 35348 31884
rect 35400 31872 35406 31884
rect 35529 31875 35587 31881
rect 35529 31872 35541 31875
rect 35400 31844 35541 31872
rect 35400 31832 35406 31844
rect 35529 31841 35541 31844
rect 35575 31872 35587 31875
rect 35710 31872 35716 31884
rect 35575 31844 35716 31872
rect 35575 31841 35587 31844
rect 35529 31835 35587 31841
rect 35710 31832 35716 31844
rect 35768 31832 35774 31884
rect 35986 31832 35992 31884
rect 36044 31872 36050 31884
rect 36096 31881 36124 31912
rect 37734 31900 37740 31912
rect 37792 31900 37798 31952
rect 37826 31900 37832 31952
rect 37884 31940 37890 31952
rect 38099 31943 38157 31949
rect 38099 31940 38111 31943
rect 37884 31912 38111 31940
rect 37884 31900 37890 31912
rect 38099 31909 38111 31912
rect 38145 31940 38157 31943
rect 38470 31940 38476 31952
rect 38145 31912 38476 31940
rect 38145 31909 38157 31912
rect 38099 31903 38157 31909
rect 38470 31900 38476 31912
rect 38528 31900 38534 31952
rect 38930 31940 38936 31952
rect 38891 31912 38936 31940
rect 38930 31900 38936 31912
rect 38988 31900 38994 31952
rect 39666 31900 39672 31952
rect 39724 31940 39730 31952
rect 39806 31943 39864 31949
rect 39806 31940 39818 31943
rect 39724 31912 39818 31940
rect 39724 31900 39730 31912
rect 39806 31909 39818 31912
rect 39852 31909 39864 31943
rect 39806 31903 39864 31909
rect 41506 31900 41512 31952
rect 41564 31940 41570 31952
rect 41830 31943 41888 31949
rect 41830 31940 41842 31943
rect 41564 31912 41842 31940
rect 41564 31900 41570 31912
rect 41830 31909 41842 31912
rect 41876 31909 41888 31943
rect 42444 31940 42472 31971
rect 43533 31943 43591 31949
rect 43533 31940 43545 31943
rect 42444 31912 43545 31940
rect 41830 31903 41888 31909
rect 43533 31909 43545 31912
rect 43579 31940 43591 31943
rect 44082 31940 44088 31952
rect 43579 31912 44088 31940
rect 43579 31909 43591 31912
rect 43533 31903 43591 31909
rect 44082 31900 44088 31912
rect 44140 31900 44146 31952
rect 36081 31875 36139 31881
rect 36081 31872 36093 31875
rect 36044 31844 36093 31872
rect 36044 31832 36050 31844
rect 36081 31841 36093 31844
rect 36127 31841 36139 31875
rect 36081 31835 36139 31841
rect 36265 31875 36323 31881
rect 36265 31841 36277 31875
rect 36311 31872 36323 31875
rect 40402 31872 40408 31884
rect 36311 31844 39849 31872
rect 40363 31844 40408 31872
rect 36311 31841 36323 31844
rect 36265 31835 36323 31841
rect 7466 31804 7472 31816
rect 7427 31776 7472 31804
rect 7466 31764 7472 31776
rect 7524 31804 7530 31816
rect 7929 31807 7987 31813
rect 7929 31804 7941 31807
rect 7524 31776 7941 31804
rect 7524 31764 7530 31776
rect 7929 31773 7941 31776
rect 7975 31773 7987 31807
rect 19334 31804 19340 31816
rect 19295 31776 19340 31804
rect 7929 31767 7987 31773
rect 19334 31764 19340 31776
rect 19392 31764 19398 31816
rect 19613 31807 19671 31813
rect 19613 31773 19625 31807
rect 19659 31804 19671 31807
rect 20438 31804 20444 31816
rect 19659 31776 20444 31804
rect 19659 31773 19671 31776
rect 19613 31767 19671 31773
rect 5767 31739 5825 31745
rect 5767 31705 5779 31739
rect 5813 31736 5825 31739
rect 7834 31736 7840 31748
rect 5813 31708 7840 31736
rect 5813 31705 5825 31708
rect 5767 31699 5825 31705
rect 7834 31696 7840 31708
rect 7892 31696 7898 31748
rect 15286 31696 15292 31748
rect 15344 31736 15350 31748
rect 16163 31739 16221 31745
rect 16163 31736 16175 31739
rect 15344 31708 16175 31736
rect 15344 31696 15350 31708
rect 16163 31705 16175 31708
rect 16209 31705 16221 31739
rect 16163 31699 16221 31705
rect 16482 31696 16488 31748
rect 16540 31736 16546 31748
rect 19628 31736 19656 31767
rect 20438 31764 20444 31776
rect 20496 31764 20502 31816
rect 22646 31804 22652 31816
rect 22607 31776 22652 31804
rect 22646 31764 22652 31776
rect 22704 31764 22710 31816
rect 24486 31804 24492 31816
rect 24447 31776 24492 31804
rect 24486 31764 24492 31776
rect 24544 31764 24550 31816
rect 24765 31807 24823 31813
rect 24765 31773 24777 31807
rect 24811 31773 24823 31807
rect 26602 31804 26608 31816
rect 26563 31776 26608 31804
rect 24765 31767 24823 31773
rect 16540 31708 19656 31736
rect 16540 31696 16546 31708
rect 24210 31696 24216 31748
rect 24268 31736 24274 31748
rect 24780 31736 24808 31767
rect 26602 31764 26608 31776
rect 26660 31764 26666 31816
rect 26878 31764 26884 31816
rect 26936 31804 26942 31816
rect 28077 31807 28135 31813
rect 28077 31804 28089 31807
rect 26936 31776 28089 31804
rect 26936 31764 26942 31776
rect 28077 31773 28089 31776
rect 28123 31773 28135 31807
rect 31754 31804 31760 31816
rect 28077 31767 28135 31773
rect 28321 31776 31760 31804
rect 24268 31708 24808 31736
rect 24268 31696 24274 31708
rect 26234 31696 26240 31748
rect 26292 31736 26298 31748
rect 28321 31736 28349 31776
rect 31754 31764 31760 31776
rect 31812 31804 31818 31816
rect 33594 31804 33600 31816
rect 31812 31776 33600 31804
rect 31812 31764 31818 31776
rect 33594 31764 33600 31776
rect 33652 31764 33658 31816
rect 33962 31804 33968 31816
rect 33923 31776 33968 31804
rect 33962 31764 33968 31776
rect 34020 31764 34026 31816
rect 34241 31807 34299 31813
rect 34241 31773 34253 31807
rect 34287 31773 34299 31807
rect 37734 31804 37740 31816
rect 37695 31776 37740 31804
rect 34241 31767 34299 31773
rect 26292 31708 28349 31736
rect 26292 31696 26298 31708
rect 33778 31696 33784 31748
rect 33836 31736 33842 31748
rect 34256 31736 34284 31767
rect 37734 31764 37740 31776
rect 37792 31764 37798 31816
rect 39482 31804 39488 31816
rect 39443 31776 39488 31804
rect 39482 31764 39488 31776
rect 39540 31764 39546 31816
rect 39821 31804 39849 31844
rect 40402 31832 40408 31844
rect 40460 31832 40466 31884
rect 41509 31807 41567 31813
rect 41509 31804 41521 31807
rect 39821 31776 41521 31804
rect 41509 31773 41521 31776
rect 41555 31804 41567 31807
rect 41874 31804 41880 31816
rect 41555 31776 41880 31804
rect 41555 31773 41567 31776
rect 41509 31767 41567 31773
rect 41874 31764 41880 31776
rect 41932 31764 41938 31816
rect 43438 31804 43444 31816
rect 43399 31776 43444 31804
rect 43438 31764 43444 31776
rect 43496 31764 43502 31816
rect 43717 31807 43775 31813
rect 43717 31804 43729 31807
rect 43548 31776 43729 31804
rect 33836 31708 34284 31736
rect 33836 31696 33842 31708
rect 34422 31696 34428 31748
rect 34480 31736 34486 31748
rect 38562 31736 38568 31748
rect 34480 31708 38568 31736
rect 34480 31696 34486 31708
rect 38562 31696 38568 31708
rect 38620 31696 38626 31748
rect 41141 31739 41199 31745
rect 41141 31705 41153 31739
rect 41187 31736 41199 31739
rect 41230 31736 41236 31748
rect 41187 31708 41236 31736
rect 41187 31705 41199 31708
rect 41141 31699 41199 31705
rect 41230 31696 41236 31708
rect 41288 31736 41294 31748
rect 43548 31736 43576 31776
rect 43717 31773 43729 31776
rect 43763 31773 43775 31807
rect 43717 31767 43775 31773
rect 41288 31708 43576 31736
rect 41288 31696 41294 31708
rect 5166 31628 5172 31680
rect 5224 31668 5230 31680
rect 5445 31671 5503 31677
rect 5445 31668 5457 31671
rect 5224 31640 5457 31668
rect 5224 31628 5230 31640
rect 5445 31637 5457 31640
rect 5491 31637 5503 31671
rect 6178 31668 6184 31680
rect 6139 31640 6184 31668
rect 5445 31631 5503 31637
rect 6178 31628 6184 31640
rect 6236 31628 6242 31680
rect 8294 31668 8300 31680
rect 8255 31640 8300 31668
rect 8294 31628 8300 31640
rect 8352 31628 8358 31680
rect 12250 31628 12256 31680
rect 12308 31668 12314 31680
rect 12437 31671 12495 31677
rect 12437 31668 12449 31671
rect 12308 31640 12449 31668
rect 12308 31628 12314 31640
rect 12437 31637 12449 31640
rect 12483 31668 12495 31671
rect 12986 31668 12992 31680
rect 12483 31640 12992 31668
rect 12483 31637 12495 31640
rect 12437 31631 12495 31637
rect 12986 31628 12992 31640
rect 13044 31668 13050 31680
rect 13173 31671 13231 31677
rect 13173 31668 13185 31671
rect 13044 31640 13185 31668
rect 13044 31628 13050 31640
rect 13173 31637 13185 31640
rect 13219 31668 13231 31671
rect 13633 31671 13691 31677
rect 13633 31668 13645 31671
rect 13219 31640 13645 31668
rect 13219 31637 13231 31640
rect 13173 31631 13231 31637
rect 13633 31637 13645 31640
rect 13679 31668 13691 31671
rect 14182 31668 14188 31680
rect 13679 31640 14188 31668
rect 13679 31637 13691 31640
rect 13633 31631 13691 31637
rect 14182 31628 14188 31640
rect 14240 31628 14246 31680
rect 17862 31628 17868 31680
rect 17920 31668 17926 31680
rect 18049 31671 18107 31677
rect 18049 31668 18061 31671
rect 17920 31640 18061 31668
rect 17920 31628 17926 31640
rect 18049 31637 18061 31640
rect 18095 31637 18107 31671
rect 18966 31668 18972 31680
rect 18927 31640 18972 31668
rect 18049 31631 18107 31637
rect 18966 31628 18972 31640
rect 19024 31628 19030 31680
rect 21358 31668 21364 31680
rect 21319 31640 21364 31668
rect 21358 31628 21364 31640
rect 21416 31628 21422 31680
rect 25501 31671 25559 31677
rect 25501 31637 25513 31671
rect 25547 31668 25559 31671
rect 25590 31668 25596 31680
rect 25547 31640 25596 31668
rect 25547 31637 25559 31640
rect 25501 31631 25559 31637
rect 25590 31628 25596 31640
rect 25648 31628 25654 31680
rect 28626 31628 28632 31680
rect 28684 31668 28690 31680
rect 29362 31668 29368 31680
rect 28684 31640 29368 31668
rect 28684 31628 28690 31640
rect 29362 31628 29368 31640
rect 29420 31668 29426 31680
rect 30466 31668 30472 31680
rect 29420 31640 30472 31668
rect 29420 31628 29426 31640
rect 30466 31628 30472 31640
rect 30524 31668 30530 31680
rect 31573 31671 31631 31677
rect 31573 31668 31585 31671
rect 30524 31640 31585 31668
rect 30524 31628 30530 31640
rect 31573 31637 31585 31640
rect 31619 31668 31631 31671
rect 32030 31668 32036 31680
rect 31619 31640 32036 31668
rect 31619 31637 31631 31640
rect 31573 31631 31631 31637
rect 32030 31628 32036 31640
rect 32088 31628 32094 31680
rect 35342 31668 35348 31680
rect 35303 31640 35348 31668
rect 35342 31628 35348 31640
rect 35400 31628 35406 31680
rect 36170 31628 36176 31680
rect 36228 31668 36234 31680
rect 39390 31668 39396 31680
rect 36228 31640 39396 31668
rect 36228 31628 36234 31640
rect 39390 31628 39396 31640
rect 39448 31628 39454 31680
rect 1104 31578 48852 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 48852 31578
rect 1104 31504 48852 31526
rect 4614 31424 4620 31476
rect 4672 31464 4678 31476
rect 4893 31467 4951 31473
rect 4893 31464 4905 31467
rect 4672 31436 4905 31464
rect 4672 31424 4678 31436
rect 4893 31433 4905 31436
rect 4939 31433 4951 31467
rect 16482 31464 16488 31476
rect 16443 31436 16488 31464
rect 4893 31427 4951 31433
rect 16482 31424 16488 31436
rect 16540 31424 16546 31476
rect 18509 31467 18567 31473
rect 18509 31433 18521 31467
rect 18555 31464 18567 31467
rect 19426 31464 19432 31476
rect 18555 31436 19432 31464
rect 18555 31433 18567 31436
rect 18509 31427 18567 31433
rect 19426 31424 19432 31436
rect 19484 31464 19490 31476
rect 19889 31467 19947 31473
rect 19889 31464 19901 31467
rect 19484 31436 19901 31464
rect 19484 31424 19490 31436
rect 19889 31433 19901 31436
rect 19935 31433 19947 31467
rect 21542 31464 21548 31476
rect 21503 31436 21548 31464
rect 19889 31427 19947 31433
rect 21542 31424 21548 31436
rect 21600 31464 21606 31476
rect 24394 31464 24400 31476
rect 21600 31436 24400 31464
rect 21600 31424 21606 31436
rect 24394 31424 24400 31436
rect 24452 31424 24458 31476
rect 24578 31424 24584 31476
rect 24636 31464 24642 31476
rect 25317 31467 25375 31473
rect 25317 31464 25329 31467
rect 24636 31436 25329 31464
rect 24636 31424 24642 31436
rect 25317 31433 25329 31436
rect 25363 31433 25375 31467
rect 25958 31464 25964 31476
rect 25919 31436 25964 31464
rect 25317 31427 25375 31433
rect 25958 31424 25964 31436
rect 26016 31424 26022 31476
rect 26602 31424 26608 31476
rect 26660 31464 26666 31476
rect 27801 31467 27859 31473
rect 27801 31464 27813 31467
rect 26660 31436 27813 31464
rect 26660 31424 26666 31436
rect 27801 31433 27813 31436
rect 27847 31433 27859 31467
rect 27801 31427 27859 31433
rect 29638 31424 29644 31476
rect 29696 31464 29702 31476
rect 30282 31464 30288 31476
rect 29696 31436 30288 31464
rect 29696 31424 29702 31436
rect 30282 31424 30288 31436
rect 30340 31424 30346 31476
rect 32582 31424 32588 31476
rect 32640 31464 32646 31476
rect 32861 31467 32919 31473
rect 32861 31464 32873 31467
rect 32640 31436 32873 31464
rect 32640 31424 32646 31436
rect 32861 31433 32873 31436
rect 32907 31433 32919 31467
rect 32861 31427 32919 31433
rect 33735 31467 33793 31473
rect 33735 31433 33747 31467
rect 33781 31464 33793 31467
rect 33962 31464 33968 31476
rect 33781 31436 33968 31464
rect 33781 31433 33793 31436
rect 33735 31427 33793 31433
rect 33962 31424 33968 31436
rect 34020 31424 34026 31476
rect 34146 31464 34152 31476
rect 34107 31436 34152 31464
rect 34146 31424 34152 31436
rect 34204 31424 34210 31476
rect 35986 31464 35992 31476
rect 35947 31436 35992 31464
rect 35986 31424 35992 31436
rect 36044 31424 36050 31476
rect 36357 31467 36415 31473
rect 36357 31433 36369 31467
rect 36403 31464 36415 31467
rect 36446 31464 36452 31476
rect 36403 31436 36452 31464
rect 36403 31433 36415 31436
rect 36357 31427 36415 31433
rect 36446 31424 36452 31436
rect 36504 31424 36510 31476
rect 37734 31424 37740 31476
rect 37792 31464 37798 31476
rect 38657 31467 38715 31473
rect 38657 31464 38669 31467
rect 37792 31436 38669 31464
rect 37792 31424 37798 31436
rect 38657 31433 38669 31436
rect 38703 31433 38715 31467
rect 39390 31464 39396 31476
rect 39351 31436 39396 31464
rect 38657 31427 38715 31433
rect 39390 31424 39396 31436
rect 39448 31424 39454 31476
rect 40770 31464 40776 31476
rect 40731 31436 40776 31464
rect 40770 31424 40776 31436
rect 40828 31424 40834 31476
rect 41874 31464 41880 31476
rect 41835 31436 41880 31464
rect 41874 31424 41880 31436
rect 41932 31424 41938 31476
rect 42383 31467 42441 31473
rect 42383 31433 42395 31467
rect 42429 31464 42441 31467
rect 43165 31467 43223 31473
rect 43165 31464 43177 31467
rect 42429 31436 43177 31464
rect 42429 31433 42441 31436
rect 42383 31427 42441 31433
rect 43165 31433 43177 31436
rect 43211 31464 43223 31467
rect 43438 31464 43444 31476
rect 43211 31436 43444 31464
rect 43211 31433 43223 31436
rect 43165 31427 43223 31433
rect 43438 31424 43444 31436
rect 43496 31424 43502 31476
rect 43622 31424 43628 31476
rect 43680 31464 43686 31476
rect 43717 31467 43775 31473
rect 43717 31464 43729 31467
rect 43680 31436 43729 31464
rect 43680 31424 43686 31436
rect 43717 31433 43729 31436
rect 43763 31433 43775 31467
rect 44082 31464 44088 31476
rect 44043 31436 44088 31464
rect 43717 31427 43775 31433
rect 44082 31424 44088 31436
rect 44140 31424 44146 31476
rect 14645 31399 14703 31405
rect 14645 31365 14657 31399
rect 14691 31396 14703 31399
rect 14691 31368 15424 31396
rect 14691 31365 14703 31368
rect 14645 31359 14703 31365
rect 6641 31331 6699 31337
rect 6641 31297 6653 31331
rect 6687 31328 6699 31331
rect 7006 31328 7012 31340
rect 6687 31300 7012 31328
rect 6687 31297 6699 31300
rect 6641 31291 6699 31297
rect 7006 31288 7012 31300
rect 7064 31288 7070 31340
rect 10134 31288 10140 31340
rect 10192 31328 10198 31340
rect 13262 31328 13268 31340
rect 10192 31300 13268 31328
rect 10192 31288 10198 31300
rect 13262 31288 13268 31300
rect 13320 31328 13326 31340
rect 13449 31331 13507 31337
rect 13449 31328 13461 31331
rect 13320 31300 13461 31328
rect 13320 31288 13326 31300
rect 13449 31297 13461 31300
rect 13495 31297 13507 31331
rect 13449 31291 13507 31297
rect 4500 31263 4558 31269
rect 4500 31229 4512 31263
rect 4546 31229 4558 31263
rect 4500 31223 4558 31229
rect 4515 31192 4543 31223
rect 5166 31220 5172 31272
rect 5224 31260 5230 31272
rect 5480 31263 5538 31269
rect 5480 31260 5492 31263
rect 5224 31232 5492 31260
rect 5224 31220 5230 31232
rect 5480 31229 5492 31232
rect 5526 31229 5538 31263
rect 5480 31223 5538 31229
rect 10689 31263 10747 31269
rect 10689 31229 10701 31263
rect 10735 31260 10747 31263
rect 10778 31260 10784 31272
rect 10735 31232 10784 31260
rect 10735 31229 10747 31232
rect 10689 31223 10747 31229
rect 10778 31220 10784 31232
rect 10836 31220 10842 31272
rect 11146 31220 11152 31272
rect 11204 31260 11210 31272
rect 11241 31263 11299 31269
rect 11241 31260 11253 31263
rect 11204 31232 11253 31260
rect 11204 31220 11210 31232
rect 11241 31229 11253 31232
rect 11287 31229 11299 31263
rect 14458 31260 14464 31272
rect 14419 31232 14464 31260
rect 11241 31223 11299 31229
rect 14458 31220 14464 31232
rect 14516 31260 14522 31272
rect 14921 31263 14979 31269
rect 14921 31260 14933 31263
rect 14516 31232 14933 31260
rect 14516 31220 14522 31232
rect 14921 31229 14933 31232
rect 14967 31260 14979 31263
rect 15286 31260 15292 31272
rect 14967 31232 15292 31260
rect 14967 31229 14979 31232
rect 14921 31223 14979 31229
rect 15286 31220 15292 31232
rect 15344 31220 15350 31272
rect 15396 31269 15424 31368
rect 18690 31356 18696 31408
rect 18748 31396 18754 31408
rect 18785 31399 18843 31405
rect 18785 31396 18797 31399
rect 18748 31368 18797 31396
rect 18748 31356 18754 31368
rect 18785 31365 18797 31368
rect 18831 31365 18843 31399
rect 18785 31359 18843 31365
rect 15381 31263 15439 31269
rect 15381 31229 15393 31263
rect 15427 31260 15439 31263
rect 15565 31263 15623 31269
rect 15565 31260 15577 31263
rect 15427 31232 15577 31260
rect 15427 31229 15439 31232
rect 15381 31223 15439 31229
rect 15565 31229 15577 31232
rect 15611 31229 15623 31263
rect 15565 31223 15623 31229
rect 5583 31195 5641 31201
rect 4515 31164 5396 31192
rect 5368 31136 5396 31164
rect 5583 31161 5595 31195
rect 5629 31192 5641 31195
rect 6917 31195 6975 31201
rect 6917 31192 6929 31195
rect 5629 31164 6929 31192
rect 5629 31161 5641 31164
rect 5583 31155 5641 31161
rect 6917 31161 6929 31164
rect 6963 31161 6975 31195
rect 6917 31155 6975 31161
rect 3786 31084 3792 31136
rect 3844 31124 3850 31136
rect 4065 31127 4123 31133
rect 4065 31124 4077 31127
rect 3844 31096 4077 31124
rect 3844 31084 3850 31096
rect 4065 31093 4077 31096
rect 4111 31093 4123 31127
rect 4065 31087 4123 31093
rect 4571 31127 4629 31133
rect 4571 31093 4583 31127
rect 4617 31124 4629 31127
rect 4982 31124 4988 31136
rect 4617 31096 4988 31124
rect 4617 31093 4629 31096
rect 4571 31087 4629 31093
rect 4982 31084 4988 31096
rect 5040 31084 5046 31136
rect 5350 31124 5356 31136
rect 5311 31096 5356 31124
rect 5350 31084 5356 31096
rect 5408 31084 5414 31136
rect 6273 31127 6331 31133
rect 6273 31093 6285 31127
rect 6319 31124 6331 31127
rect 6362 31124 6368 31136
rect 6319 31096 6368 31124
rect 6319 31093 6331 31096
rect 6273 31087 6331 31093
rect 6362 31084 6368 31096
rect 6420 31084 6426 31136
rect 6932 31124 6960 31155
rect 7006 31152 7012 31204
rect 7064 31192 7070 31204
rect 7561 31195 7619 31201
rect 7064 31164 7109 31192
rect 7064 31152 7070 31164
rect 7561 31161 7573 31195
rect 7607 31192 7619 31195
rect 8846 31192 8852 31204
rect 7607 31164 8852 31192
rect 7607 31161 7619 31164
rect 7561 31155 7619 31161
rect 8846 31152 8852 31164
rect 8904 31152 8910 31204
rect 8938 31152 8944 31204
rect 8996 31192 9002 31204
rect 9493 31195 9551 31201
rect 8996 31164 9041 31192
rect 8996 31152 9002 31164
rect 9493 31161 9505 31195
rect 9539 31192 9551 31195
rect 9674 31192 9680 31204
rect 9539 31164 9680 31192
rect 9539 31161 9551 31164
rect 9493 31155 9551 31161
rect 9674 31152 9680 31164
rect 9732 31152 9738 31204
rect 12526 31192 12532 31204
rect 12487 31164 12532 31192
rect 12526 31152 12532 31164
rect 12584 31152 12590 31204
rect 12621 31195 12679 31201
rect 12621 31161 12633 31195
rect 12667 31161 12679 31195
rect 13170 31192 13176 31204
rect 13131 31164 13176 31192
rect 12621 31155 12679 31161
rect 7837 31127 7895 31133
rect 7837 31124 7849 31127
rect 6932 31096 7849 31124
rect 7837 31093 7849 31096
rect 7883 31093 7895 31127
rect 7837 31087 7895 31093
rect 8297 31127 8355 31133
rect 8297 31093 8309 31127
rect 8343 31124 8355 31127
rect 8386 31124 8392 31136
rect 8343 31096 8392 31124
rect 8343 31093 8355 31096
rect 8297 31087 8355 31093
rect 8386 31084 8392 31096
rect 8444 31084 8450 31136
rect 8665 31127 8723 31133
rect 8665 31093 8677 31127
rect 8711 31124 8723 31127
rect 8956 31124 8984 31152
rect 8711 31096 8984 31124
rect 8711 31093 8723 31096
rect 8665 31087 8723 31093
rect 9582 31084 9588 31136
rect 9640 31124 9646 31136
rect 9769 31127 9827 31133
rect 9769 31124 9781 31127
rect 9640 31096 9781 31124
rect 9640 31084 9646 31096
rect 9769 31093 9781 31096
rect 9815 31093 9827 31127
rect 10134 31124 10140 31136
rect 10095 31096 10140 31124
rect 9769 31087 9827 31093
rect 10134 31084 10140 31096
rect 10192 31084 10198 31136
rect 10870 31124 10876 31136
rect 10831 31096 10876 31124
rect 10870 31084 10876 31096
rect 10928 31084 10934 31136
rect 11422 31084 11428 31136
rect 11480 31124 11486 31136
rect 11793 31127 11851 31133
rect 11793 31124 11805 31127
rect 11480 31096 11805 31124
rect 11480 31084 11486 31096
rect 11793 31093 11805 31096
rect 11839 31093 11851 31127
rect 11793 31087 11851 31093
rect 12253 31127 12311 31133
rect 12253 31093 12265 31127
rect 12299 31124 12311 31127
rect 12636 31124 12664 31155
rect 13170 31152 13176 31164
rect 13228 31152 13234 31204
rect 13906 31192 13912 31204
rect 13280 31164 13912 31192
rect 12894 31124 12900 31136
rect 12299 31096 12900 31124
rect 12299 31093 12311 31096
rect 12253 31087 12311 31093
rect 12894 31084 12900 31096
rect 12952 31124 12958 31136
rect 13280 31124 13308 31164
rect 13906 31152 13912 31164
rect 13964 31192 13970 31204
rect 15473 31195 15531 31201
rect 15473 31192 15485 31195
rect 13964 31164 15485 31192
rect 13964 31152 13970 31164
rect 15473 31161 15485 31164
rect 15519 31161 15531 31195
rect 15473 31155 15531 31161
rect 17129 31195 17187 31201
rect 17129 31161 17141 31195
rect 17175 31192 17187 31195
rect 17310 31192 17316 31204
rect 17175 31164 17316 31192
rect 17175 31161 17187 31164
rect 17129 31155 17187 31161
rect 17310 31152 17316 31164
rect 17368 31192 17374 31204
rect 17770 31192 17776 31204
rect 17368 31164 17776 31192
rect 17368 31152 17374 31164
rect 17770 31152 17776 31164
rect 17828 31152 17834 31204
rect 18800 31192 18828 31359
rect 19334 31356 19340 31408
rect 19392 31396 19398 31408
rect 20257 31399 20315 31405
rect 20257 31396 20269 31399
rect 19392 31368 20269 31396
rect 19392 31356 19398 31368
rect 20257 31365 20269 31368
rect 20303 31396 20315 31399
rect 21726 31396 21732 31408
rect 20303 31368 21732 31396
rect 20303 31365 20315 31368
rect 20257 31359 20315 31365
rect 21726 31356 21732 31368
rect 21784 31356 21790 31408
rect 32493 31399 32551 31405
rect 32493 31365 32505 31399
rect 32539 31396 32551 31399
rect 32766 31396 32772 31408
rect 32539 31368 32772 31396
rect 32539 31365 32551 31368
rect 32493 31359 32551 31365
rect 32766 31356 32772 31368
rect 32824 31356 32830 31408
rect 33134 31356 33140 31408
rect 33192 31396 33198 31408
rect 33192 31368 36302 31396
rect 33192 31356 33198 31368
rect 22646 31328 22652 31340
rect 22559 31300 22652 31328
rect 22646 31288 22652 31300
rect 22704 31328 22710 31340
rect 23293 31331 23351 31337
rect 23293 31328 23305 31331
rect 22704 31300 23305 31328
rect 22704 31288 22710 31300
rect 23293 31297 23305 31300
rect 23339 31297 23351 31331
rect 23293 31291 23351 31297
rect 25041 31331 25099 31337
rect 25041 31297 25053 31331
rect 25087 31328 25099 31331
rect 25222 31328 25228 31340
rect 25087 31300 25228 31328
rect 25087 31297 25099 31300
rect 25041 31291 25099 31297
rect 25222 31288 25228 31300
rect 25280 31288 25286 31340
rect 26697 31331 26755 31337
rect 26697 31297 26709 31331
rect 26743 31328 26755 31331
rect 26878 31328 26884 31340
rect 26743 31300 26884 31328
rect 26743 31297 26755 31300
rect 26697 31291 26755 31297
rect 26878 31288 26884 31300
rect 26936 31288 26942 31340
rect 27154 31328 27160 31340
rect 27115 31300 27160 31328
rect 27154 31288 27160 31300
rect 27212 31288 27218 31340
rect 29914 31328 29920 31340
rect 29875 31300 29920 31328
rect 29914 31288 29920 31300
rect 29972 31288 29978 31340
rect 30374 31288 30380 31340
rect 30432 31328 30438 31340
rect 31938 31328 31944 31340
rect 30432 31300 30880 31328
rect 31851 31300 31944 31328
rect 30432 31288 30438 31300
rect 18966 31260 18972 31272
rect 18927 31232 18972 31260
rect 18966 31220 18972 31232
rect 19024 31220 19030 31272
rect 20717 31263 20775 31269
rect 20717 31229 20729 31263
rect 20763 31260 20775 31263
rect 21910 31260 21916 31272
rect 20763 31232 21312 31260
rect 21871 31232 21916 31260
rect 20763 31229 20775 31232
rect 20717 31223 20775 31229
rect 19242 31192 19248 31204
rect 18800 31164 19248 31192
rect 19242 31152 19248 31164
rect 19300 31201 19306 31204
rect 19300 31195 19348 31201
rect 19300 31161 19302 31195
rect 19336 31161 19348 31195
rect 19300 31155 19348 31161
rect 19300 31152 19306 31155
rect 12952 31096 13308 31124
rect 17497 31127 17555 31133
rect 12952 31084 12958 31096
rect 17497 31093 17509 31127
rect 17543 31124 17555 31127
rect 17862 31124 17868 31136
rect 17543 31096 17868 31124
rect 17543 31093 17555 31096
rect 17497 31087 17555 31093
rect 17862 31084 17868 31096
rect 17920 31084 17926 31136
rect 20898 31124 20904 31136
rect 20859 31096 20904 31124
rect 20898 31084 20904 31096
rect 20956 31084 20962 31136
rect 21284 31133 21312 31232
rect 21910 31220 21916 31232
rect 21968 31220 21974 31272
rect 22094 31220 22100 31272
rect 22152 31260 22158 31272
rect 22373 31263 22431 31269
rect 22373 31260 22385 31263
rect 22152 31232 22385 31260
rect 22152 31220 22158 31232
rect 22373 31229 22385 31232
rect 22419 31229 22431 31263
rect 22373 31223 22431 31229
rect 24029 31263 24087 31269
rect 24029 31229 24041 31263
rect 24075 31260 24087 31263
rect 24305 31263 24363 31269
rect 24305 31260 24317 31263
rect 24075 31232 24317 31260
rect 24075 31229 24087 31232
rect 24029 31223 24087 31229
rect 24305 31229 24317 31232
rect 24351 31229 24363 31263
rect 24305 31223 24363 31229
rect 22388 31192 22416 31223
rect 24578 31220 24584 31272
rect 24636 31260 24642 31272
rect 24765 31263 24823 31269
rect 24765 31260 24777 31263
rect 24636 31232 24777 31260
rect 24636 31220 24642 31232
rect 24765 31229 24777 31232
rect 24811 31229 24823 31263
rect 24765 31223 24823 31229
rect 29089 31263 29147 31269
rect 29089 31229 29101 31263
rect 29135 31260 29147 31263
rect 29454 31260 29460 31272
rect 29135 31232 29460 31260
rect 29135 31229 29147 31232
rect 29089 31223 29147 31229
rect 29454 31220 29460 31232
rect 29512 31220 29518 31272
rect 29825 31263 29883 31269
rect 29825 31229 29837 31263
rect 29871 31260 29883 31263
rect 30466 31260 30472 31272
rect 29871 31232 30472 31260
rect 29871 31229 29883 31232
rect 29825 31223 29883 31229
rect 30466 31220 30472 31232
rect 30524 31220 30530 31272
rect 30852 31269 30880 31300
rect 31938 31288 31944 31300
rect 31996 31328 32002 31340
rect 34238 31328 34244 31340
rect 31996 31300 34244 31328
rect 31996 31288 32002 31300
rect 34238 31288 34244 31300
rect 34296 31288 34302 31340
rect 35434 31328 35440 31340
rect 35176 31300 35440 31328
rect 30837 31263 30895 31269
rect 30837 31229 30849 31263
rect 30883 31260 30895 31263
rect 31297 31263 31355 31269
rect 31297 31260 31309 31263
rect 30883 31232 31309 31260
rect 30883 31229 30895 31232
rect 30837 31223 30895 31229
rect 31297 31229 31309 31232
rect 31343 31229 31355 31263
rect 31297 31223 31355 31229
rect 33410 31220 33416 31272
rect 33468 31260 33474 31272
rect 33664 31263 33722 31269
rect 33664 31260 33676 31263
rect 33468 31232 33676 31260
rect 33468 31220 33474 31232
rect 33664 31229 33676 31232
rect 33710 31260 33722 31263
rect 34146 31260 34152 31272
rect 33710 31232 34152 31260
rect 33710 31229 33722 31232
rect 33664 31223 33722 31229
rect 34146 31220 34152 31232
rect 34204 31220 34210 31272
rect 35176 31269 35204 31300
rect 35434 31288 35440 31300
rect 35492 31288 35498 31340
rect 35161 31263 35219 31269
rect 35161 31229 35173 31263
rect 35207 31229 35219 31263
rect 35161 31223 35219 31229
rect 35345 31263 35403 31269
rect 35345 31229 35357 31263
rect 35391 31260 35403 31263
rect 35986 31260 35992 31272
rect 35391 31232 35992 31260
rect 35391 31229 35403 31232
rect 35345 31223 35403 31229
rect 24596 31192 24624 31220
rect 22388 31164 24624 31192
rect 25958 31152 25964 31204
rect 26016 31192 26022 31204
rect 26973 31195 27031 31201
rect 26973 31192 26985 31195
rect 26016 31164 26985 31192
rect 26016 31152 26022 31164
rect 26973 31161 26985 31164
rect 27019 31161 27031 31195
rect 26973 31155 27031 31161
rect 32033 31195 32091 31201
rect 32033 31161 32045 31195
rect 32079 31161 32091 31195
rect 32033 31155 32091 31161
rect 34701 31195 34759 31201
rect 34701 31161 34713 31195
rect 34747 31192 34759 31195
rect 35360 31192 35388 31223
rect 35986 31220 35992 31232
rect 36044 31220 36050 31272
rect 36274 31260 36302 31368
rect 36464 31328 36492 31424
rect 37185 31331 37243 31337
rect 36464 31300 36952 31328
rect 36446 31260 36452 31272
rect 36274 31232 36452 31260
rect 36446 31220 36452 31232
rect 36504 31220 36510 31272
rect 36924 31269 36952 31300
rect 37185 31297 37197 31331
rect 37231 31328 37243 31331
rect 37752 31328 37780 31424
rect 39666 31396 39672 31408
rect 38488 31368 39672 31396
rect 38488 31340 38516 31368
rect 39666 31356 39672 31368
rect 39724 31396 39730 31408
rect 41506 31396 41512 31408
rect 39724 31368 41512 31396
rect 39724 31356 39730 31368
rect 41506 31356 41512 31368
rect 41564 31356 41570 31408
rect 37231 31300 37780 31328
rect 37829 31331 37887 31337
rect 37231 31297 37243 31300
rect 37185 31291 37243 31297
rect 37829 31297 37841 31331
rect 37875 31328 37887 31331
rect 38470 31328 38476 31340
rect 37875 31300 38476 31328
rect 37875 31297 37887 31300
rect 37829 31291 37887 31297
rect 38470 31288 38476 31300
rect 38528 31288 38534 31340
rect 38562 31288 38568 31340
rect 38620 31328 38626 31340
rect 43395 31331 43453 31337
rect 38620 31300 43346 31328
rect 38620 31288 38626 31300
rect 36909 31263 36967 31269
rect 36909 31229 36921 31263
rect 36955 31229 36967 31263
rect 36909 31223 36967 31229
rect 38197 31263 38255 31269
rect 38197 31229 38209 31263
rect 38243 31260 38255 31263
rect 38286 31260 38292 31272
rect 38243 31232 38292 31260
rect 38243 31229 38255 31232
rect 38197 31223 38255 31229
rect 38286 31220 38292 31232
rect 38344 31220 38350 31272
rect 39114 31220 39120 31272
rect 39172 31260 39178 31272
rect 39209 31263 39267 31269
rect 39209 31260 39221 31263
rect 39172 31232 39221 31260
rect 39172 31220 39178 31232
rect 39209 31229 39221 31232
rect 39255 31260 39267 31263
rect 40037 31263 40095 31269
rect 40037 31260 40049 31263
rect 39255 31232 40049 31260
rect 39255 31229 39267 31232
rect 39209 31223 39267 31229
rect 40037 31229 40049 31232
rect 40083 31229 40095 31263
rect 40037 31223 40095 31229
rect 40564 31263 40622 31269
rect 40564 31229 40576 31263
rect 40610 31260 40622 31263
rect 40610 31232 41092 31260
rect 40610 31229 40622 31232
rect 40564 31223 40622 31229
rect 34747 31164 35388 31192
rect 35621 31195 35679 31201
rect 34747 31161 34759 31164
rect 34701 31155 34759 31161
rect 35621 31161 35633 31195
rect 35667 31192 35679 31195
rect 39025 31195 39083 31201
rect 39025 31192 39037 31195
rect 35667 31164 39037 31192
rect 35667 31161 35679 31164
rect 35621 31155 35679 31161
rect 39025 31161 39037 31164
rect 39071 31192 39083 31195
rect 39482 31192 39488 31204
rect 39071 31164 39488 31192
rect 39071 31161 39083 31164
rect 39025 31155 39083 31161
rect 21269 31127 21327 31133
rect 21269 31093 21281 31127
rect 21315 31124 21327 31127
rect 21634 31124 21640 31136
rect 21315 31096 21640 31124
rect 21315 31093 21327 31096
rect 21269 31087 21327 31093
rect 21634 31084 21640 31096
rect 21692 31084 21698 31136
rect 22278 31084 22284 31136
rect 22336 31124 22342 31136
rect 22925 31127 22983 31133
rect 22925 31124 22937 31127
rect 22336 31096 22937 31124
rect 22336 31084 22342 31096
rect 22925 31093 22937 31096
rect 22971 31124 22983 31127
rect 23014 31124 23020 31136
rect 22971 31096 23020 31124
rect 22971 31093 22983 31096
rect 22925 31087 22983 31093
rect 23014 31084 23020 31096
rect 23072 31084 23078 31136
rect 23750 31084 23756 31136
rect 23808 31124 23814 31136
rect 24029 31127 24087 31133
rect 24029 31124 24041 31127
rect 23808 31096 24041 31124
rect 23808 31084 23814 31096
rect 24029 31093 24041 31096
rect 24075 31124 24087 31127
rect 24121 31127 24179 31133
rect 24121 31124 24133 31127
rect 24075 31096 24133 31124
rect 24075 31093 24087 31096
rect 24029 31087 24087 31093
rect 24121 31093 24133 31096
rect 24167 31093 24179 31127
rect 24121 31087 24179 31093
rect 26329 31127 26387 31133
rect 26329 31093 26341 31127
rect 26375 31124 26387 31127
rect 26694 31124 26700 31136
rect 26375 31096 26700 31124
rect 26375 31093 26387 31096
rect 26329 31087 26387 31093
rect 26694 31084 26700 31096
rect 26752 31084 26758 31136
rect 31018 31124 31024 31136
rect 30979 31096 31024 31124
rect 31018 31084 31024 31096
rect 31076 31084 31082 31136
rect 31570 31084 31576 31136
rect 31628 31124 31634 31136
rect 31665 31127 31723 31133
rect 31665 31124 31677 31127
rect 31628 31096 31677 31124
rect 31628 31084 31634 31096
rect 31665 31093 31677 31096
rect 31711 31124 31723 31127
rect 32048 31124 32076 31155
rect 39482 31152 39488 31164
rect 39540 31152 39546 31204
rect 41064 31136 41092 31232
rect 42150 31220 42156 31272
rect 42208 31260 42214 31272
rect 43318 31269 43346 31300
rect 43395 31297 43407 31331
rect 43441 31328 43453 31331
rect 43530 31328 43536 31340
rect 43441 31300 43536 31328
rect 43441 31297 43453 31300
rect 43395 31291 43453 31297
rect 43530 31288 43536 31300
rect 43588 31288 43594 31340
rect 42312 31263 42370 31269
rect 42312 31260 42324 31263
rect 42208 31232 42324 31260
rect 42208 31220 42214 31232
rect 42312 31229 42324 31232
rect 42358 31260 42370 31263
rect 43308 31263 43366 31269
rect 42358 31232 42748 31260
rect 42358 31229 42370 31232
rect 42312 31223 42370 31229
rect 42720 31136 42748 31232
rect 43308 31229 43320 31263
rect 43354 31260 43366 31263
rect 43622 31260 43628 31272
rect 43354 31232 43628 31260
rect 43354 31229 43366 31232
rect 43308 31223 43366 31229
rect 43622 31220 43628 31232
rect 43680 31220 43686 31272
rect 33502 31124 33508 31136
rect 31711 31096 32076 31124
rect 33463 31096 33508 31124
rect 31711 31093 31723 31096
rect 31665 31087 31723 31093
rect 33502 31084 33508 31096
rect 33560 31084 33566 31136
rect 37826 31084 37832 31136
rect 37884 31124 37890 31136
rect 38335 31127 38393 31133
rect 38335 31124 38347 31127
rect 37884 31096 38347 31124
rect 37884 31084 37890 31096
rect 38335 31093 38347 31096
rect 38381 31093 38393 31127
rect 41046 31124 41052 31136
rect 41007 31096 41052 31124
rect 38335 31087 38393 31093
rect 41046 31084 41052 31096
rect 41104 31084 41110 31136
rect 42702 31124 42708 31136
rect 42663 31096 42708 31124
rect 42702 31084 42708 31096
rect 42760 31084 42766 31136
rect 1104 31034 48852 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 48852 31034
rect 1104 30960 48852 30982
rect 4614 30920 4620 30932
rect 4575 30892 4620 30920
rect 4614 30880 4620 30892
rect 4672 30880 4678 30932
rect 5169 30923 5227 30929
rect 5169 30889 5181 30923
rect 5215 30920 5227 30923
rect 5721 30923 5779 30929
rect 5721 30920 5733 30923
rect 5215 30892 5733 30920
rect 5215 30889 5227 30892
rect 5169 30883 5227 30889
rect 5721 30889 5733 30892
rect 5767 30920 5779 30923
rect 5810 30920 5816 30932
rect 5767 30892 5816 30920
rect 5767 30889 5779 30892
rect 5721 30883 5779 30889
rect 5810 30880 5816 30892
rect 5868 30880 5874 30932
rect 6178 30880 6184 30932
rect 6236 30920 6242 30932
rect 6917 30923 6975 30929
rect 6917 30920 6929 30923
rect 6236 30892 6929 30920
rect 6236 30880 6242 30892
rect 6917 30889 6929 30892
rect 6963 30889 6975 30923
rect 6917 30883 6975 30889
rect 7006 30880 7012 30932
rect 7064 30920 7070 30932
rect 8846 30920 8852 30932
rect 7064 30892 7972 30920
rect 8807 30892 8852 30920
rect 7064 30880 7070 30892
rect 5902 30812 5908 30864
rect 5960 30852 5966 30864
rect 6318 30855 6376 30861
rect 6318 30852 6330 30855
rect 5960 30824 6330 30852
rect 5960 30812 5966 30824
rect 6318 30821 6330 30824
rect 6364 30821 6376 30855
rect 7834 30852 7840 30864
rect 7795 30824 7840 30852
rect 6318 30815 6376 30821
rect 7834 30812 7840 30824
rect 7892 30812 7898 30864
rect 7944 30861 7972 30892
rect 8846 30880 8852 30892
rect 8904 30880 8910 30932
rect 10091 30923 10149 30929
rect 10091 30889 10103 30923
rect 10137 30920 10149 30923
rect 12526 30920 12532 30932
rect 10137 30892 12532 30920
rect 10137 30889 10149 30892
rect 10091 30883 10149 30889
rect 12526 30880 12532 30892
rect 12584 30880 12590 30932
rect 19242 30920 19248 30932
rect 19203 30892 19248 30920
rect 19242 30880 19248 30892
rect 19300 30880 19306 30932
rect 24486 30880 24492 30932
rect 24544 30920 24550 30932
rect 25041 30923 25099 30929
rect 25041 30920 25053 30923
rect 24544 30892 25053 30920
rect 24544 30880 24550 30892
rect 25041 30889 25053 30892
rect 25087 30889 25099 30923
rect 29546 30920 29552 30932
rect 29507 30892 29552 30920
rect 25041 30883 25099 30889
rect 29546 30880 29552 30892
rect 29604 30880 29610 30932
rect 31938 30920 31944 30932
rect 31899 30892 31944 30920
rect 31938 30880 31944 30892
rect 31996 30880 32002 30932
rect 33413 30923 33471 30929
rect 33413 30889 33425 30923
rect 33459 30920 33471 30923
rect 33962 30920 33968 30932
rect 33459 30892 33968 30920
rect 33459 30889 33471 30892
rect 33413 30883 33471 30889
rect 33962 30880 33968 30892
rect 34020 30880 34026 30932
rect 34977 30923 35035 30929
rect 34977 30889 34989 30923
rect 35023 30920 35035 30923
rect 35434 30920 35440 30932
rect 35023 30892 35440 30920
rect 35023 30889 35035 30892
rect 34977 30883 35035 30889
rect 35434 30880 35440 30892
rect 35492 30880 35498 30932
rect 36446 30920 36452 30932
rect 36407 30892 36452 30920
rect 36446 30880 36452 30892
rect 36504 30880 36510 30932
rect 38286 30920 38292 30932
rect 38199 30892 38292 30920
rect 38286 30880 38292 30892
rect 38344 30920 38350 30932
rect 39206 30920 39212 30932
rect 38344 30892 39212 30920
rect 38344 30880 38350 30892
rect 39206 30880 39212 30892
rect 39264 30880 39270 30932
rect 7929 30855 7987 30861
rect 7929 30821 7941 30855
rect 7975 30852 7987 30855
rect 8478 30852 8484 30864
rect 7975 30824 8484 30852
rect 7975 30821 7987 30824
rect 7929 30815 7987 30821
rect 8478 30812 8484 30824
rect 8536 30812 8542 30864
rect 11238 30852 11244 30864
rect 11199 30824 11244 30852
rect 11238 30812 11244 30824
rect 11296 30812 11302 30864
rect 12250 30852 12256 30864
rect 12211 30824 12256 30852
rect 12250 30812 12256 30824
rect 12308 30812 12314 30864
rect 23842 30852 23848 30864
rect 23803 30824 23848 30852
rect 23842 30812 23848 30824
rect 23900 30812 23906 30864
rect 26694 30852 26700 30864
rect 26655 30824 26700 30852
rect 26694 30812 26700 30824
rect 26752 30812 26758 30864
rect 27246 30852 27252 30864
rect 27207 30824 27252 30852
rect 27246 30812 27252 30824
rect 27304 30812 27310 30864
rect 32398 30852 32404 30864
rect 32359 30824 32404 30852
rect 32398 30812 32404 30824
rect 32456 30812 32462 30864
rect 32766 30812 32772 30864
rect 32824 30852 32830 30864
rect 32953 30855 33011 30861
rect 32953 30852 32965 30855
rect 32824 30824 32965 30852
rect 32824 30812 32830 30824
rect 32953 30821 32965 30824
rect 32999 30821 33011 30855
rect 32953 30815 33011 30821
rect 33502 30812 33508 30864
rect 33560 30852 33566 30864
rect 34057 30855 34115 30861
rect 34057 30852 34069 30855
rect 33560 30824 34069 30852
rect 33560 30812 33566 30824
rect 34057 30821 34069 30824
rect 34103 30852 34115 30855
rect 35253 30855 35311 30861
rect 35253 30852 35265 30855
rect 34103 30824 35265 30852
rect 34103 30821 34115 30824
rect 34057 30815 34115 30821
rect 35253 30821 35265 30824
rect 35299 30852 35311 30855
rect 35621 30855 35679 30861
rect 35621 30852 35633 30855
rect 35299 30824 35633 30852
rect 35299 30821 35311 30824
rect 35253 30815 35311 30821
rect 35621 30821 35633 30824
rect 35667 30821 35679 30855
rect 35621 30815 35679 30821
rect 6086 30744 6092 30796
rect 6144 30784 6150 30796
rect 7466 30784 7472 30796
rect 6144 30756 7472 30784
rect 6144 30744 6150 30756
rect 7466 30744 7472 30756
rect 7524 30784 7530 30796
rect 10042 30793 10048 30796
rect 7561 30787 7619 30793
rect 7561 30784 7573 30787
rect 7524 30756 7573 30784
rect 7524 30744 7530 30756
rect 7561 30753 7573 30756
rect 7607 30753 7619 30787
rect 10020 30787 10048 30793
rect 10020 30784 10032 30787
rect 9955 30756 10032 30784
rect 7561 30747 7619 30753
rect 10020 30753 10032 30756
rect 10100 30784 10106 30796
rect 11885 30787 11943 30793
rect 11885 30784 11897 30787
rect 10100 30756 11897 30784
rect 10020 30747 10048 30753
rect 10042 30744 10048 30747
rect 10100 30744 10106 30756
rect 11885 30753 11897 30756
rect 11931 30753 11943 30787
rect 13262 30784 13268 30796
rect 13223 30756 13268 30784
rect 11885 30747 11943 30753
rect 13262 30744 13268 30756
rect 13320 30744 13326 30796
rect 13354 30744 13360 30796
rect 13412 30784 13418 30796
rect 13725 30787 13783 30793
rect 13725 30784 13737 30787
rect 13412 30756 13737 30784
rect 13412 30744 13418 30756
rect 13725 30753 13737 30756
rect 13771 30753 13783 30787
rect 15470 30784 15476 30796
rect 15431 30756 15476 30784
rect 13725 30747 13783 30753
rect 15470 30744 15476 30756
rect 15528 30744 15534 30796
rect 17126 30784 17132 30796
rect 17087 30756 17132 30784
rect 17126 30744 17132 30756
rect 17184 30744 17190 30796
rect 19797 30787 19855 30793
rect 19797 30753 19809 30787
rect 19843 30784 19855 30787
rect 19886 30784 19892 30796
rect 19843 30756 19892 30784
rect 19843 30753 19855 30756
rect 19797 30747 19855 30753
rect 19886 30744 19892 30756
rect 19944 30744 19950 30796
rect 20901 30787 20959 30793
rect 20901 30753 20913 30787
rect 20947 30784 20959 30787
rect 21726 30784 21732 30796
rect 20947 30756 21732 30784
rect 20947 30753 20959 30756
rect 20901 30747 20959 30753
rect 21726 30744 21732 30756
rect 21784 30744 21790 30796
rect 22624 30787 22682 30793
rect 22624 30753 22636 30787
rect 22670 30784 22682 30787
rect 22738 30784 22744 30796
rect 22670 30756 22744 30784
rect 22670 30753 22682 30756
rect 22624 30747 22682 30753
rect 22738 30744 22744 30756
rect 22796 30744 22802 30796
rect 24394 30744 24400 30796
rect 24452 30784 24458 30796
rect 25444 30787 25502 30793
rect 25444 30784 25456 30787
rect 24452 30756 25456 30784
rect 24452 30744 24458 30756
rect 25444 30753 25456 30756
rect 25490 30784 25502 30787
rect 26234 30784 26240 30796
rect 25490 30756 26240 30784
rect 25490 30753 25502 30756
rect 25444 30747 25502 30753
rect 26234 30744 26240 30756
rect 26292 30744 26298 30796
rect 28905 30787 28963 30793
rect 28905 30753 28917 30787
rect 28951 30784 28963 30787
rect 29086 30784 29092 30796
rect 28951 30756 29092 30784
rect 28951 30753 28963 30756
rect 28905 30747 28963 30753
rect 29086 30744 29092 30756
rect 29144 30744 29150 30796
rect 30190 30784 30196 30796
rect 30151 30756 30196 30784
rect 30190 30744 30196 30756
rect 30248 30744 30254 30796
rect 30466 30784 30472 30796
rect 30427 30756 30472 30784
rect 30466 30744 30472 30756
rect 30524 30744 30530 30796
rect 37734 30784 37740 30796
rect 37695 30756 37740 30784
rect 37734 30744 37740 30756
rect 37792 30744 37798 30796
rect 38749 30787 38807 30793
rect 38749 30753 38761 30787
rect 38795 30784 38807 30787
rect 38930 30784 38936 30796
rect 38795 30756 38936 30784
rect 38795 30753 38807 30756
rect 38749 30747 38807 30753
rect 38930 30744 38936 30756
rect 38988 30744 38994 30796
rect 39758 30784 39764 30796
rect 39719 30756 39764 30784
rect 39758 30744 39764 30756
rect 39816 30744 39822 30796
rect 41138 30784 41144 30796
rect 41099 30756 41144 30784
rect 41138 30744 41144 30756
rect 41196 30744 41202 30796
rect 4249 30719 4307 30725
rect 4249 30685 4261 30719
rect 4295 30716 4307 30719
rect 4890 30716 4896 30728
rect 4295 30688 4896 30716
rect 4295 30685 4307 30688
rect 4249 30679 4307 30685
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 5994 30716 6000 30728
rect 5955 30688 6000 30716
rect 5994 30676 6000 30688
rect 6052 30676 6058 30728
rect 8110 30716 8116 30728
rect 8071 30688 8116 30716
rect 8110 30676 8116 30688
rect 8168 30676 8174 30728
rect 10962 30716 10968 30728
rect 10923 30688 10968 30716
rect 10962 30676 10968 30688
rect 11020 30676 11026 30728
rect 13814 30676 13820 30728
rect 13872 30716 13878 30728
rect 13872 30688 13917 30716
rect 13872 30676 13878 30688
rect 14734 30676 14740 30728
rect 14792 30716 14798 30728
rect 15381 30719 15439 30725
rect 15381 30716 15393 30719
rect 14792 30688 15393 30716
rect 14792 30676 14798 30688
rect 15381 30685 15393 30688
rect 15427 30685 15439 30719
rect 16942 30716 16948 30728
rect 16903 30688 16948 30716
rect 15381 30679 15439 30685
rect 16942 30676 16948 30688
rect 17000 30676 17006 30728
rect 18874 30716 18880 30728
rect 18835 30688 18880 30716
rect 18874 30676 18880 30688
rect 18932 30676 18938 30728
rect 23753 30719 23811 30725
rect 23753 30685 23765 30719
rect 23799 30716 23811 30719
rect 23934 30716 23940 30728
rect 23799 30688 23940 30716
rect 23799 30685 23811 30688
rect 23753 30679 23811 30685
rect 23934 30676 23940 30688
rect 23992 30676 23998 30728
rect 24118 30716 24124 30728
rect 24079 30688 24124 30716
rect 24118 30676 24124 30688
rect 24176 30676 24182 30728
rect 26605 30719 26663 30725
rect 26605 30716 26617 30719
rect 26252 30688 26617 30716
rect 17770 30608 17776 30660
rect 17828 30648 17834 30660
rect 21910 30648 21916 30660
rect 17828 30620 21916 30648
rect 17828 30608 17834 30620
rect 21910 30608 21916 30620
rect 21968 30648 21974 30660
rect 26252 30657 26280 30688
rect 26605 30685 26617 30688
rect 26651 30685 26663 30719
rect 30650 30716 30656 30728
rect 30563 30688 30656 30716
rect 26605 30679 26663 30685
rect 30650 30676 30656 30688
rect 30708 30716 30714 30728
rect 30929 30719 30987 30725
rect 30929 30716 30941 30719
rect 30708 30688 30941 30716
rect 30708 30676 30714 30688
rect 30929 30685 30941 30688
rect 30975 30685 30987 30719
rect 30929 30679 30987 30685
rect 31938 30676 31944 30728
rect 31996 30716 32002 30728
rect 32309 30719 32367 30725
rect 32309 30716 32321 30719
rect 31996 30688 32321 30716
rect 31996 30676 32002 30688
rect 32309 30685 32321 30688
rect 32355 30716 32367 30719
rect 33781 30719 33839 30725
rect 32355 30688 32996 30716
rect 32355 30685 32367 30688
rect 32309 30679 32367 30685
rect 32968 30660 32996 30688
rect 33781 30685 33793 30719
rect 33827 30716 33839 30719
rect 33962 30716 33968 30728
rect 33827 30688 33968 30716
rect 33827 30685 33839 30688
rect 33781 30679 33839 30685
rect 33962 30676 33968 30688
rect 34020 30676 34026 30728
rect 34238 30716 34244 30728
rect 34199 30688 34244 30716
rect 34238 30676 34244 30688
rect 34296 30676 34302 30728
rect 34606 30676 34612 30728
rect 34664 30716 34670 30728
rect 35529 30719 35587 30725
rect 35529 30716 35541 30719
rect 34664 30688 35541 30716
rect 34664 30676 34670 30688
rect 35529 30685 35541 30688
rect 35575 30685 35587 30719
rect 35802 30716 35808 30728
rect 35715 30688 35808 30716
rect 35529 30679 35587 30685
rect 35802 30676 35808 30688
rect 35860 30676 35866 30728
rect 25547 30651 25605 30657
rect 21968 30620 25268 30648
rect 21968 30608 21974 30620
rect 6730 30540 6736 30592
rect 6788 30580 6794 30592
rect 7193 30583 7251 30589
rect 7193 30580 7205 30583
rect 6788 30552 7205 30580
rect 6788 30540 6794 30552
rect 7193 30549 7205 30552
rect 7239 30580 7251 30583
rect 7374 30580 7380 30592
rect 7239 30552 7380 30580
rect 7239 30549 7251 30552
rect 7193 30543 7251 30549
rect 7374 30540 7380 30552
rect 7432 30580 7438 30592
rect 10134 30580 10140 30592
rect 7432 30552 10140 30580
rect 7432 30540 7438 30552
rect 10134 30540 10140 30552
rect 10192 30540 10198 30592
rect 10318 30540 10324 30592
rect 10376 30580 10382 30592
rect 10781 30583 10839 30589
rect 10781 30580 10793 30583
rect 10376 30552 10793 30580
rect 10376 30540 10382 30552
rect 10781 30549 10793 30552
rect 10827 30580 10839 30583
rect 11146 30580 11152 30592
rect 10827 30552 11152 30580
rect 10827 30549 10839 30552
rect 10781 30543 10839 30549
rect 11146 30540 11152 30552
rect 11204 30540 11210 30592
rect 18322 30580 18328 30592
rect 18283 30552 18328 30580
rect 18322 30540 18328 30552
rect 18380 30540 18386 30592
rect 18782 30540 18788 30592
rect 18840 30580 18846 30592
rect 21085 30583 21143 30589
rect 21085 30580 21097 30583
rect 18840 30552 21097 30580
rect 18840 30540 18846 30552
rect 21085 30549 21097 30552
rect 21131 30549 21143 30583
rect 21085 30543 21143 30549
rect 22695 30583 22753 30589
rect 22695 30549 22707 30583
rect 22741 30580 22753 30583
rect 23014 30580 23020 30592
rect 22741 30552 23020 30580
rect 22741 30549 22753 30552
rect 22695 30543 22753 30549
rect 23014 30540 23020 30552
rect 23072 30540 23078 30592
rect 24578 30540 24584 30592
rect 24636 30580 24642 30592
rect 24673 30583 24731 30589
rect 24673 30580 24685 30583
rect 24636 30552 24685 30580
rect 24636 30540 24642 30552
rect 24673 30549 24685 30552
rect 24719 30549 24731 30583
rect 25240 30580 25268 30620
rect 25547 30617 25559 30651
rect 25593 30648 25605 30651
rect 26237 30651 26295 30657
rect 26237 30648 26249 30651
rect 25593 30620 26249 30648
rect 25593 30617 25605 30620
rect 25547 30611 25605 30617
rect 26237 30617 26249 30620
rect 26283 30617 26295 30651
rect 26237 30611 26295 30617
rect 29089 30651 29147 30657
rect 29089 30617 29101 30651
rect 29135 30648 29147 30651
rect 30466 30648 30472 30660
rect 29135 30620 30472 30648
rect 29135 30617 29147 30620
rect 29089 30611 29147 30617
rect 30466 30608 30472 30620
rect 30524 30608 30530 30660
rect 32950 30608 32956 30660
rect 33008 30648 33014 30660
rect 35820 30648 35848 30676
rect 33008 30620 35848 30648
rect 33008 30608 33014 30620
rect 36446 30608 36452 30660
rect 36504 30648 36510 30660
rect 39945 30651 40003 30657
rect 39945 30648 39957 30651
rect 36504 30620 39957 30648
rect 36504 30608 36510 30620
rect 39945 30617 39957 30620
rect 39991 30617 40003 30651
rect 39945 30611 40003 30617
rect 28166 30580 28172 30592
rect 25240 30552 28172 30580
rect 24673 30543 24731 30549
rect 28166 30540 28172 30552
rect 28224 30540 28230 30592
rect 35342 30540 35348 30592
rect 35400 30580 35406 30592
rect 37921 30583 37979 30589
rect 37921 30580 37933 30583
rect 35400 30552 37933 30580
rect 35400 30540 35406 30552
rect 37921 30549 37933 30552
rect 37967 30549 37979 30583
rect 37921 30543 37979 30549
rect 38838 30540 38844 30592
rect 38896 30580 38902 30592
rect 38933 30583 38991 30589
rect 38933 30580 38945 30583
rect 38896 30552 38945 30580
rect 38896 30540 38902 30552
rect 38933 30549 38945 30552
rect 38979 30549 38991 30583
rect 39206 30580 39212 30592
rect 39167 30552 39212 30580
rect 38933 30543 38991 30549
rect 39206 30540 39212 30552
rect 39264 30540 39270 30592
rect 40954 30580 40960 30592
rect 40915 30552 40960 30580
rect 40954 30540 40960 30552
rect 41012 30540 41018 30592
rect 41279 30583 41337 30589
rect 41279 30549 41291 30583
rect 41325 30580 41337 30583
rect 41782 30580 41788 30592
rect 41325 30552 41788 30580
rect 41325 30549 41337 30552
rect 41279 30543 41337 30549
rect 41782 30540 41788 30552
rect 41840 30540 41846 30592
rect 1104 30490 48852 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 48852 30490
rect 1104 30416 48852 30438
rect 5994 30336 6000 30388
rect 6052 30376 6058 30388
rect 6365 30379 6423 30385
rect 6365 30376 6377 30379
rect 6052 30348 6377 30376
rect 6052 30336 6058 30348
rect 6365 30345 6377 30348
rect 6411 30345 6423 30379
rect 10042 30376 10048 30388
rect 10003 30348 10048 30376
rect 6365 30339 6423 30345
rect 10042 30336 10048 30348
rect 10100 30336 10106 30388
rect 11514 30376 11520 30388
rect 11475 30348 11520 30376
rect 11514 30336 11520 30348
rect 11572 30336 11578 30388
rect 15470 30376 15476 30388
rect 15431 30348 15476 30376
rect 15470 30336 15476 30348
rect 15528 30336 15534 30388
rect 19242 30336 19248 30388
rect 19300 30376 19306 30388
rect 19337 30379 19395 30385
rect 19337 30376 19349 30379
rect 19300 30348 19349 30376
rect 19300 30336 19306 30348
rect 19337 30345 19349 30348
rect 19383 30376 19395 30379
rect 20257 30379 20315 30385
rect 20257 30376 20269 30379
rect 19383 30348 20269 30376
rect 19383 30345 19395 30348
rect 19337 30339 19395 30345
rect 20257 30345 20269 30348
rect 20303 30345 20315 30379
rect 21358 30376 21364 30388
rect 21319 30348 21364 30376
rect 20257 30339 20315 30345
rect 3050 30268 3056 30320
rect 3108 30308 3114 30320
rect 3694 30308 3700 30320
rect 3108 30280 3700 30308
rect 3108 30268 3114 30280
rect 3694 30268 3700 30280
rect 3752 30308 3758 30320
rect 3752 30280 5212 30308
rect 3752 30268 3758 30280
rect 3252 30212 4154 30240
rect 3252 30181 3280 30212
rect 3237 30175 3295 30181
rect 3237 30172 3249 30175
rect 3068 30144 3249 30172
rect 2958 29996 2964 30048
rect 3016 30036 3022 30048
rect 3068 30045 3096 30144
rect 3237 30141 3249 30144
rect 3283 30141 3295 30175
rect 3237 30135 3295 30141
rect 3697 30175 3755 30181
rect 3697 30141 3709 30175
rect 3743 30141 3755 30175
rect 4126 30172 4154 30212
rect 4709 30175 4767 30181
rect 4709 30172 4721 30175
rect 4126 30144 4721 30172
rect 3697 30135 3755 30141
rect 4709 30141 4721 30144
rect 4755 30172 4767 30175
rect 5074 30172 5080 30184
rect 4755 30144 5080 30172
rect 4755 30141 4767 30144
rect 4709 30135 4767 30141
rect 3142 30064 3148 30116
rect 3200 30104 3206 30116
rect 3510 30104 3516 30116
rect 3200 30076 3516 30104
rect 3200 30064 3206 30076
rect 3510 30064 3516 30076
rect 3568 30104 3574 30116
rect 3712 30104 3740 30135
rect 5074 30132 5080 30144
rect 5132 30132 5138 30184
rect 5184 30172 5212 30280
rect 10778 30268 10784 30320
rect 10836 30308 10842 30320
rect 12250 30308 12256 30320
rect 10836 30280 12256 30308
rect 10836 30268 10842 30280
rect 12250 30268 12256 30280
rect 12308 30308 12314 30320
rect 13081 30311 13139 30317
rect 13081 30308 13093 30311
rect 12308 30280 13093 30308
rect 12308 30268 12314 30280
rect 13081 30277 13093 30280
rect 13127 30308 13139 30311
rect 13262 30308 13268 30320
rect 13127 30280 13268 30308
rect 13127 30277 13139 30280
rect 13081 30271 13139 30277
rect 13262 30268 13268 30280
rect 13320 30268 13326 30320
rect 7466 30240 7472 30252
rect 7427 30212 7472 30240
rect 7466 30200 7472 30212
rect 7524 30200 7530 30252
rect 8110 30240 8116 30252
rect 8071 30212 8116 30240
rect 8110 30200 8116 30212
rect 8168 30240 8174 30252
rect 9030 30240 9036 30252
rect 8168 30212 9036 30240
rect 8168 30200 8174 30212
rect 9030 30200 9036 30212
rect 9088 30200 9094 30252
rect 10597 30243 10655 30249
rect 10597 30209 10609 30243
rect 10643 30240 10655 30243
rect 10870 30240 10876 30252
rect 10643 30212 10876 30240
rect 10643 30209 10655 30212
rect 10597 30203 10655 30209
rect 10870 30200 10876 30212
rect 10928 30200 10934 30252
rect 13633 30243 13691 30249
rect 13633 30209 13645 30243
rect 13679 30240 13691 30243
rect 13814 30240 13820 30252
rect 13679 30212 13820 30240
rect 13679 30209 13691 30212
rect 13633 30203 13691 30209
rect 13814 30200 13820 30212
rect 13872 30200 13878 30252
rect 17862 30240 17868 30252
rect 17775 30212 17868 30240
rect 17862 30200 17868 30212
rect 17920 30240 17926 30252
rect 17920 30212 18828 30240
rect 17920 30200 17926 30212
rect 18800 30184 18828 30212
rect 18874 30200 18880 30252
rect 18932 30240 18938 30252
rect 19061 30243 19119 30249
rect 19061 30240 19073 30243
rect 18932 30212 19073 30240
rect 18932 30200 18938 30212
rect 19061 30209 19073 30212
rect 19107 30240 19119 30243
rect 19705 30243 19763 30249
rect 19705 30240 19717 30243
rect 19107 30212 19717 30240
rect 19107 30209 19119 30212
rect 19061 30203 19119 30209
rect 19705 30209 19717 30212
rect 19751 30209 19763 30243
rect 19705 30203 19763 30209
rect 5258 30172 5264 30184
rect 5171 30144 5264 30172
rect 5258 30132 5264 30144
rect 5316 30132 5322 30184
rect 12253 30175 12311 30181
rect 12253 30141 12265 30175
rect 12299 30172 12311 30175
rect 12688 30175 12746 30181
rect 12688 30172 12700 30175
rect 12299 30144 12700 30172
rect 12299 30141 12311 30144
rect 12253 30135 12311 30141
rect 12688 30141 12700 30144
rect 12734 30172 12746 30175
rect 14553 30175 14611 30181
rect 14553 30172 14565 30175
rect 12734 30144 14565 30172
rect 12734 30141 12746 30144
rect 12688 30135 12746 30141
rect 14553 30141 14565 30144
rect 14599 30141 14611 30175
rect 14553 30135 14611 30141
rect 14642 30132 14648 30184
rect 14700 30172 14706 30184
rect 15105 30175 15163 30181
rect 15105 30172 15117 30175
rect 14700 30144 15117 30172
rect 14700 30132 14706 30144
rect 15105 30141 15117 30144
rect 15151 30172 15163 30175
rect 15749 30175 15807 30181
rect 15749 30172 15761 30175
rect 15151 30144 15761 30172
rect 15151 30141 15163 30144
rect 15105 30135 15163 30141
rect 15749 30141 15761 30144
rect 15795 30141 15807 30175
rect 15749 30135 15807 30141
rect 17678 30132 17684 30184
rect 17736 30172 17742 30184
rect 18322 30172 18328 30184
rect 17736 30144 18328 30172
rect 17736 30132 17742 30144
rect 18322 30132 18328 30144
rect 18380 30132 18386 30184
rect 18782 30172 18788 30184
rect 18743 30144 18788 30172
rect 18782 30132 18788 30144
rect 18840 30132 18846 30184
rect 3568 30076 3740 30104
rect 3568 30064 3574 30076
rect 3878 30064 3884 30116
rect 3936 30104 3942 30116
rect 3973 30107 4031 30113
rect 3973 30104 3985 30107
rect 3936 30076 3985 30104
rect 3936 30064 3942 30076
rect 3973 30073 3985 30076
rect 4019 30073 4031 30107
rect 5902 30104 5908 30116
rect 3973 30067 4031 30073
rect 4632 30076 5908 30104
rect 4632 30048 4660 30076
rect 5902 30064 5908 30076
rect 5960 30104 5966 30116
rect 5997 30107 6055 30113
rect 5997 30104 6009 30107
rect 5960 30076 6009 30104
rect 5960 30064 5966 30076
rect 5997 30073 6009 30076
rect 6043 30073 6055 30107
rect 5997 30067 6055 30073
rect 7285 30107 7343 30113
rect 7285 30073 7297 30107
rect 7331 30104 7343 30107
rect 7558 30104 7564 30116
rect 7331 30076 7564 30104
rect 7331 30073 7343 30076
rect 7285 30067 7343 30073
rect 7558 30064 7564 30076
rect 7616 30064 7622 30116
rect 8849 30107 8907 30113
rect 8849 30073 8861 30107
rect 8895 30104 8907 30107
rect 9125 30107 9183 30113
rect 9125 30104 9137 30107
rect 8895 30076 9137 30104
rect 8895 30073 8907 30076
rect 8849 30067 8907 30073
rect 9125 30073 9137 30076
rect 9171 30104 9183 30107
rect 9490 30104 9496 30116
rect 9171 30076 9496 30104
rect 9171 30073 9183 30076
rect 9125 30067 9183 30073
rect 9490 30064 9496 30076
rect 9548 30064 9554 30116
rect 9674 30104 9680 30116
rect 9635 30076 9680 30104
rect 9674 30064 9680 30076
rect 9732 30064 9738 30116
rect 10505 30107 10563 30113
rect 10505 30073 10517 30107
rect 10551 30104 10563 30107
rect 10959 30107 11017 30113
rect 10959 30104 10971 30107
rect 10551 30076 10971 30104
rect 10551 30073 10563 30076
rect 10505 30067 10563 30073
rect 10959 30073 10971 30076
rect 11005 30104 11017 30107
rect 11238 30104 11244 30116
rect 11005 30076 11244 30104
rect 11005 30073 11017 30076
rect 10959 30067 11017 30073
rect 11238 30064 11244 30076
rect 11296 30104 11302 30116
rect 11885 30107 11943 30113
rect 11885 30104 11897 30107
rect 11296 30076 11897 30104
rect 11296 30064 11302 30076
rect 11885 30073 11897 30076
rect 11931 30104 11943 30107
rect 13541 30107 13599 30113
rect 13541 30104 13553 30107
rect 11931 30076 13553 30104
rect 11931 30073 11943 30076
rect 11885 30067 11943 30073
rect 13541 30073 13553 30076
rect 13587 30104 13599 30107
rect 13722 30104 13728 30116
rect 13587 30076 13728 30104
rect 13587 30073 13599 30076
rect 13541 30067 13599 30073
rect 13722 30064 13728 30076
rect 13780 30104 13786 30116
rect 13954 30107 14012 30113
rect 13954 30104 13966 30107
rect 13780 30076 13966 30104
rect 13780 30064 13786 30076
rect 13954 30073 13966 30076
rect 14000 30104 14012 30107
rect 14090 30104 14096 30116
rect 14000 30076 14096 30104
rect 14000 30073 14012 30076
rect 13954 30067 14012 30073
rect 14090 30064 14096 30076
rect 14148 30064 14154 30116
rect 15654 30104 15660 30116
rect 15615 30076 15660 30104
rect 15654 30064 15660 30076
rect 15712 30064 15718 30116
rect 20272 30104 20300 30339
rect 21358 30336 21364 30348
rect 21416 30336 21422 30388
rect 22738 30336 22744 30388
rect 22796 30376 22802 30388
rect 23017 30379 23075 30385
rect 23017 30376 23029 30379
rect 22796 30348 23029 30376
rect 22796 30336 22802 30348
rect 23017 30345 23029 30348
rect 23063 30345 23075 30379
rect 23017 30339 23075 30345
rect 23474 30336 23480 30388
rect 23532 30376 23538 30388
rect 23842 30376 23848 30388
rect 23532 30348 23848 30376
rect 23532 30336 23538 30348
rect 23842 30336 23848 30348
rect 23900 30336 23906 30388
rect 23934 30336 23940 30388
rect 23992 30376 23998 30388
rect 24857 30379 24915 30385
rect 24857 30376 24869 30379
rect 23992 30348 24869 30376
rect 23992 30336 23998 30348
rect 24857 30345 24869 30348
rect 24903 30376 24915 30379
rect 27246 30376 27252 30388
rect 24903 30348 27252 30376
rect 24903 30345 24915 30348
rect 24857 30339 24915 30345
rect 27246 30336 27252 30348
rect 27304 30336 27310 30388
rect 28258 30336 28264 30388
rect 28316 30376 28322 30388
rect 28445 30379 28503 30385
rect 28445 30376 28457 30379
rect 28316 30348 28457 30376
rect 28316 30336 28322 30348
rect 28445 30345 28457 30348
rect 28491 30345 28503 30379
rect 28445 30339 28503 30345
rect 30282 30336 30288 30388
rect 30340 30376 30346 30388
rect 30469 30379 30527 30385
rect 30469 30376 30481 30379
rect 30340 30348 30481 30376
rect 30340 30336 30346 30348
rect 30469 30345 30481 30348
rect 30515 30345 30527 30379
rect 31570 30376 31576 30388
rect 31531 30348 31576 30376
rect 30469 30339 30527 30345
rect 31570 30336 31576 30348
rect 31628 30336 31634 30388
rect 32217 30379 32275 30385
rect 32217 30345 32229 30379
rect 32263 30376 32275 30379
rect 32398 30376 32404 30388
rect 32263 30348 32404 30376
rect 32263 30345 32275 30348
rect 32217 30339 32275 30345
rect 32398 30336 32404 30348
rect 32456 30336 32462 30388
rect 33502 30336 33508 30388
rect 33560 30376 33566 30388
rect 33965 30379 34023 30385
rect 33965 30376 33977 30379
rect 33560 30348 33977 30376
rect 33560 30336 33566 30348
rect 33965 30345 33977 30348
rect 34011 30376 34023 30379
rect 34146 30376 34152 30388
rect 34011 30348 34152 30376
rect 34011 30345 34023 30348
rect 33965 30339 34023 30345
rect 34146 30336 34152 30348
rect 34204 30336 34210 30388
rect 36446 30376 36452 30388
rect 36407 30348 36452 30376
rect 36446 30336 36452 30348
rect 36504 30336 36510 30388
rect 39666 30336 39672 30388
rect 39724 30376 39730 30388
rect 40773 30379 40831 30385
rect 40773 30376 40785 30379
rect 39724 30348 40785 30376
rect 39724 30336 39730 30348
rect 40773 30345 40785 30348
rect 40819 30345 40831 30379
rect 40773 30339 40831 30345
rect 26234 30308 26240 30320
rect 26195 30280 26240 30308
rect 26234 30268 26240 30280
rect 26292 30268 26298 30320
rect 27065 30311 27123 30317
rect 27065 30277 27077 30311
rect 27111 30308 27123 30311
rect 27154 30308 27160 30320
rect 27111 30280 27160 30308
rect 27111 30277 27123 30280
rect 27065 30271 27123 30277
rect 27154 30268 27160 30280
rect 27212 30268 27218 30320
rect 29457 30311 29515 30317
rect 29457 30277 29469 30311
rect 29503 30308 29515 30311
rect 30190 30308 30196 30320
rect 29503 30280 30196 30308
rect 29503 30277 29515 30280
rect 29457 30271 29515 30277
rect 30190 30268 30196 30280
rect 30248 30308 30254 30320
rect 36906 30308 36912 30320
rect 30248 30280 36912 30308
rect 30248 30268 30254 30280
rect 36906 30268 36912 30280
rect 36964 30268 36970 30320
rect 40788 30308 40816 30339
rect 40788 30280 41092 30308
rect 22465 30243 22523 30249
rect 22465 30209 22477 30243
rect 22511 30240 22523 30243
rect 24118 30240 24124 30252
rect 22511 30212 24124 30240
rect 22511 30209 22523 30212
rect 22465 30203 22523 30209
rect 20438 30172 20444 30184
rect 20399 30144 20444 30172
rect 20438 30132 20444 30144
rect 20496 30132 20502 30184
rect 22639 30181 22667 30212
rect 24118 30200 24124 30212
rect 24176 30200 24182 30252
rect 26326 30200 26332 30252
rect 26384 30240 26390 30252
rect 26513 30243 26571 30249
rect 26513 30240 26525 30243
rect 26384 30212 26525 30240
rect 26384 30200 26390 30212
rect 26513 30209 26525 30212
rect 26559 30240 26571 30243
rect 28123 30243 28181 30249
rect 28123 30240 28135 30243
rect 26559 30212 28135 30240
rect 26559 30209 26571 30212
rect 26513 30203 26571 30209
rect 28123 30209 28135 30212
rect 28169 30209 28181 30243
rect 30650 30240 30656 30252
rect 30611 30212 30656 30240
rect 28123 30203 28181 30209
rect 30650 30200 30656 30212
rect 30708 30200 30714 30252
rect 32769 30243 32827 30249
rect 32769 30209 32781 30243
rect 32815 30240 32827 30243
rect 33502 30240 33508 30252
rect 32815 30212 33508 30240
rect 32815 30209 32827 30212
rect 32769 30203 32827 30209
rect 33502 30200 33508 30212
rect 33560 30200 33566 30252
rect 35713 30243 35771 30249
rect 35713 30209 35725 30243
rect 35759 30240 35771 30243
rect 40954 30240 40960 30252
rect 35759 30212 40960 30240
rect 35759 30209 35771 30212
rect 35713 30203 35771 30209
rect 40954 30200 40960 30212
rect 41012 30200 41018 30252
rect 22624 30175 22682 30181
rect 22624 30172 22636 30175
rect 22602 30144 22636 30172
rect 22624 30141 22636 30144
rect 22670 30141 22682 30175
rect 22624 30135 22682 30141
rect 25476 30175 25534 30181
rect 25476 30141 25488 30175
rect 25522 30172 25534 30175
rect 25774 30172 25780 30184
rect 25522 30144 25780 30172
rect 25522 30141 25534 30144
rect 25476 30135 25534 30141
rect 25774 30132 25780 30144
rect 25832 30172 25838 30184
rect 28036 30175 28094 30181
rect 25832 30144 26004 30172
rect 25832 30132 25838 30144
rect 20763 30107 20821 30113
rect 20763 30104 20775 30107
rect 20272 30076 20775 30104
rect 20763 30073 20775 30076
rect 20809 30073 20821 30107
rect 20763 30067 20821 30073
rect 20990 30064 20996 30116
rect 21048 30104 21054 30116
rect 23842 30104 23848 30116
rect 21048 30076 21950 30104
rect 23803 30076 23848 30104
rect 21048 30064 21054 30076
rect 3053 30039 3111 30045
rect 3053 30036 3065 30039
rect 3016 30008 3065 30036
rect 3016 29996 3022 30008
rect 3053 30005 3065 30008
rect 3099 30005 3111 30039
rect 3053 29999 3111 30005
rect 4341 30039 4399 30045
rect 4341 30005 4353 30039
rect 4387 30036 4399 30039
rect 4614 30036 4620 30048
rect 4387 30008 4620 30036
rect 4387 30005 4399 30008
rect 4341 29999 4399 30005
rect 4614 29996 4620 30008
rect 4672 29996 4678 30048
rect 4890 30036 4896 30048
rect 4851 30008 4896 30036
rect 4890 29996 4896 30008
rect 4948 29996 4954 30048
rect 8478 30036 8484 30048
rect 8391 30008 8484 30036
rect 8478 29996 8484 30008
rect 8536 30036 8542 30048
rect 10686 30036 10692 30048
rect 8536 30008 10692 30036
rect 8536 29996 8542 30008
rect 10686 29996 10692 30008
rect 10744 29996 10750 30048
rect 12759 30039 12817 30045
rect 12759 30005 12771 30039
rect 12805 30036 12817 30039
rect 12986 30036 12992 30048
rect 12805 30008 12992 30036
rect 12805 30005 12817 30008
rect 12759 29999 12817 30005
rect 12986 29996 12992 30008
rect 13044 29996 13050 30048
rect 17037 30039 17095 30045
rect 17037 30005 17049 30039
rect 17083 30036 17095 30039
rect 17126 30036 17132 30048
rect 17083 30008 17132 30036
rect 17083 30005 17095 30008
rect 17037 29999 17095 30005
rect 17126 29996 17132 30008
rect 17184 29996 17190 30048
rect 21726 30036 21732 30048
rect 21687 30008 21732 30036
rect 21726 29996 21732 30008
rect 21784 29996 21790 30048
rect 21922 30036 21950 30076
rect 23842 30064 23848 30076
rect 23900 30064 23906 30116
rect 23937 30107 23995 30113
rect 23937 30073 23949 30107
rect 23983 30104 23995 30107
rect 24118 30104 24124 30116
rect 23983 30076 24124 30104
rect 23983 30073 23995 30076
rect 23937 30067 23995 30073
rect 24118 30064 24124 30076
rect 24176 30064 24182 30116
rect 22695 30039 22753 30045
rect 22695 30036 22707 30039
rect 21922 30008 22707 30036
rect 22695 30005 22707 30008
rect 22741 30005 22753 30039
rect 22695 29999 22753 30005
rect 25547 30039 25605 30045
rect 25547 30005 25559 30039
rect 25593 30036 25605 30039
rect 25774 30036 25780 30048
rect 25593 30008 25780 30036
rect 25593 30005 25605 30008
rect 25547 29999 25605 30005
rect 25774 29996 25780 30008
rect 25832 29996 25838 30048
rect 25976 30045 26004 30144
rect 28036 30141 28048 30175
rect 28082 30172 28094 30175
rect 28258 30172 28264 30184
rect 28082 30144 28264 30172
rect 28082 30141 28094 30144
rect 28036 30135 28094 30141
rect 28258 30132 28264 30144
rect 28316 30172 28322 30184
rect 28534 30172 28540 30184
rect 28316 30144 28540 30172
rect 28316 30132 28322 30144
rect 28534 30132 28540 30144
rect 28592 30132 28598 30184
rect 29273 30175 29331 30181
rect 29273 30141 29285 30175
rect 29319 30141 29331 30175
rect 29273 30135 29331 30141
rect 32585 30175 32643 30181
rect 32585 30141 32597 30175
rect 32631 30172 32643 30175
rect 32858 30172 32864 30184
rect 32631 30144 32864 30172
rect 32631 30141 32643 30144
rect 32585 30135 32643 30141
rect 26510 30064 26516 30116
rect 26568 30104 26574 30116
rect 26605 30107 26663 30113
rect 26605 30104 26617 30107
rect 26568 30076 26617 30104
rect 26568 30064 26574 30076
rect 26605 30073 26617 30076
rect 26651 30073 26663 30107
rect 26605 30067 26663 30073
rect 25961 30039 26019 30045
rect 25961 30005 25973 30039
rect 26007 30036 26019 30039
rect 26050 30036 26056 30048
rect 26007 30008 26056 30036
rect 26007 30005 26019 30008
rect 25961 29999 26019 30005
rect 26050 29996 26056 30008
rect 26108 29996 26114 30048
rect 26620 30036 26648 30067
rect 28166 30064 28172 30116
rect 28224 30104 28230 30116
rect 29288 30104 29316 30135
rect 32858 30132 32864 30144
rect 32916 30172 32922 30184
rect 33045 30175 33103 30181
rect 33045 30172 33057 30175
rect 32916 30144 33057 30172
rect 32916 30132 32922 30144
rect 33045 30141 33057 30144
rect 33091 30141 33103 30175
rect 34701 30175 34759 30181
rect 34701 30172 34713 30175
rect 33045 30135 33103 30141
rect 33244 30144 34713 30172
rect 29733 30107 29791 30113
rect 29733 30104 29745 30107
rect 28224 30076 29745 30104
rect 28224 30064 28230 30076
rect 29733 30073 29745 30076
rect 29779 30073 29791 30107
rect 29733 30067 29791 30073
rect 30282 30064 30288 30116
rect 30340 30104 30346 30116
rect 30974 30107 31032 30113
rect 30974 30104 30986 30107
rect 30340 30076 30986 30104
rect 30340 30064 30346 30076
rect 30974 30073 30986 30076
rect 31020 30104 31032 30107
rect 31020 30076 32076 30104
rect 31020 30073 31032 30076
rect 30974 30067 31032 30073
rect 27433 30039 27491 30045
rect 27433 30036 27445 30039
rect 26620 30008 27445 30036
rect 27433 30005 27445 30008
rect 27479 30005 27491 30039
rect 27433 29999 27491 30005
rect 27893 30039 27951 30045
rect 27893 30005 27905 30039
rect 27939 30036 27951 30039
rect 28074 30036 28080 30048
rect 27939 30008 28080 30036
rect 27939 30005 27951 30008
rect 27893 29999 27951 30005
rect 28074 29996 28080 30008
rect 28132 29996 28138 30048
rect 28997 30039 29055 30045
rect 28997 30005 29009 30039
rect 29043 30036 29055 30039
rect 29086 30036 29092 30048
rect 29043 30008 29092 30036
rect 29043 30005 29055 30008
rect 28997 29999 29055 30005
rect 29086 29996 29092 30008
rect 29144 29996 29150 30048
rect 32048 30036 32076 30076
rect 32490 30064 32496 30116
rect 32548 30104 32554 30116
rect 33244 30104 33272 30144
rect 34701 30141 34713 30144
rect 34747 30172 34759 30175
rect 35250 30172 35256 30184
rect 34747 30144 35256 30172
rect 34747 30141 34759 30144
rect 34701 30135 34759 30141
rect 35250 30132 35256 30144
rect 35308 30132 35314 30184
rect 35529 30175 35587 30181
rect 35529 30141 35541 30175
rect 35575 30172 35587 30175
rect 35575 30144 36032 30172
rect 35575 30141 35587 30144
rect 35529 30135 35587 30141
rect 32548 30076 33272 30104
rect 33407 30107 33465 30113
rect 32548 30064 32554 30076
rect 33407 30073 33419 30107
rect 33453 30104 33465 30107
rect 33502 30104 33508 30116
rect 33453 30076 33508 30104
rect 33453 30073 33465 30076
rect 33407 30067 33465 30073
rect 33502 30064 33508 30076
rect 33560 30064 33566 30116
rect 34333 30107 34391 30113
rect 34333 30073 34345 30107
rect 34379 30104 34391 30107
rect 35544 30104 35572 30135
rect 34379 30076 35572 30104
rect 34379 30073 34391 30076
rect 34333 30067 34391 30073
rect 36004 30048 36032 30144
rect 36446 30132 36452 30184
rect 36504 30172 36510 30184
rect 36541 30175 36599 30181
rect 36541 30172 36553 30175
rect 36504 30144 36553 30172
rect 36504 30132 36510 30144
rect 36541 30141 36553 30144
rect 36587 30141 36599 30175
rect 36541 30135 36599 30141
rect 37093 30175 37151 30181
rect 37093 30141 37105 30175
rect 37139 30172 37151 30175
rect 38172 30175 38230 30181
rect 37139 30144 37412 30172
rect 37139 30141 37151 30144
rect 37093 30135 37151 30141
rect 37274 30104 37280 30116
rect 37235 30076 37280 30104
rect 37274 30064 37280 30076
rect 37332 30064 37338 30116
rect 37384 30104 37412 30144
rect 38172 30141 38184 30175
rect 38218 30172 38230 30175
rect 38562 30172 38568 30184
rect 38218 30144 38568 30172
rect 38218 30141 38230 30144
rect 38172 30135 38230 30141
rect 38562 30132 38568 30144
rect 38620 30132 38626 30184
rect 39117 30175 39175 30181
rect 39117 30141 39129 30175
rect 39163 30172 39175 30175
rect 39206 30172 39212 30184
rect 39163 30144 39212 30172
rect 39163 30141 39175 30144
rect 39117 30135 39175 30141
rect 39206 30132 39212 30144
rect 39264 30132 39270 30184
rect 37550 30104 37556 30116
rect 37384 30076 37556 30104
rect 37550 30064 37556 30076
rect 37608 30104 37614 30116
rect 41064 30104 41092 30280
rect 41322 30200 41328 30252
rect 41380 30240 41386 30252
rect 43346 30240 43352 30252
rect 41380 30212 43352 30240
rect 41380 30200 41386 30212
rect 43346 30200 43352 30212
rect 43404 30200 43410 30252
rect 41966 30132 41972 30184
rect 42024 30172 42030 30184
rect 42740 30175 42798 30181
rect 42740 30172 42752 30175
rect 42024 30144 42752 30172
rect 42024 30132 42030 30144
rect 42740 30141 42752 30144
rect 42786 30172 42798 30175
rect 43165 30175 43223 30181
rect 43165 30172 43177 30175
rect 42786 30144 43177 30172
rect 42786 30141 42798 30144
rect 42740 30135 42798 30141
rect 43165 30141 43177 30144
rect 43211 30141 43223 30175
rect 43165 30135 43223 30141
rect 41278 30107 41336 30113
rect 41278 30104 41290 30107
rect 37608 30076 39252 30104
rect 41064 30076 41290 30104
rect 37608 30064 37614 30076
rect 32769 30039 32827 30045
rect 32769 30036 32781 30039
rect 32048 30008 32781 30036
rect 32769 30005 32781 30008
rect 32815 30036 32827 30039
rect 32861 30039 32919 30045
rect 32861 30036 32873 30039
rect 32815 30008 32873 30036
rect 32815 30005 32827 30008
rect 32769 29999 32827 30005
rect 32861 30005 32873 30008
rect 32907 30005 32919 30039
rect 35986 30036 35992 30048
rect 35947 30008 35992 30036
rect 32861 29999 32919 30005
rect 35986 29996 35992 30008
rect 36044 29996 36050 30048
rect 37734 30036 37740 30048
rect 37695 30008 37740 30036
rect 37734 29996 37740 30008
rect 37792 29996 37798 30048
rect 38243 30039 38301 30045
rect 38243 30005 38255 30039
rect 38289 30036 38301 30039
rect 38378 30036 38384 30048
rect 38289 30008 38384 30036
rect 38289 30005 38301 30008
rect 38243 29999 38301 30005
rect 38378 29996 38384 30008
rect 38436 29996 38442 30048
rect 38930 30036 38936 30048
rect 38891 30008 38936 30036
rect 38930 29996 38936 30008
rect 38988 29996 38994 30048
rect 39224 30036 39252 30076
rect 41278 30073 41290 30076
rect 41324 30073 41336 30107
rect 41278 30067 41336 30073
rect 39301 30039 39359 30045
rect 39301 30036 39313 30039
rect 39224 30008 39313 30036
rect 39301 30005 39313 30008
rect 39347 30005 39359 30039
rect 39758 30036 39764 30048
rect 39719 30008 39764 30036
rect 39301 29999 39359 30005
rect 39758 29996 39764 30008
rect 39816 29996 39822 30048
rect 41874 30036 41880 30048
rect 41835 30008 41880 30036
rect 41874 29996 41880 30008
rect 41932 29996 41938 30048
rect 42518 29996 42524 30048
rect 42576 30036 42582 30048
rect 42843 30039 42901 30045
rect 42843 30036 42855 30039
rect 42576 30008 42855 30036
rect 42576 29996 42582 30008
rect 42843 30005 42855 30008
rect 42889 30005 42901 30039
rect 42843 29999 42901 30005
rect 1104 29946 48852 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 48852 29946
rect 1104 29872 48852 29894
rect 3881 29835 3939 29841
rect 3881 29801 3893 29835
rect 3927 29832 3939 29835
rect 4890 29832 4896 29844
rect 3927 29804 4896 29832
rect 3927 29801 3939 29804
rect 3881 29795 3939 29801
rect 4890 29792 4896 29804
rect 4948 29792 4954 29844
rect 5258 29832 5264 29844
rect 5219 29804 5264 29832
rect 5258 29792 5264 29804
rect 5316 29792 5322 29844
rect 5994 29792 6000 29844
rect 6052 29832 6058 29844
rect 6089 29835 6147 29841
rect 6089 29832 6101 29835
rect 6052 29804 6101 29832
rect 6052 29792 6058 29804
rect 6089 29801 6101 29804
rect 6135 29801 6147 29835
rect 6089 29795 6147 29801
rect 7834 29792 7840 29844
rect 7892 29832 7898 29844
rect 8389 29835 8447 29841
rect 8389 29832 8401 29835
rect 7892 29804 8401 29832
rect 7892 29792 7898 29804
rect 8389 29801 8401 29804
rect 8435 29801 8447 29835
rect 9030 29832 9036 29844
rect 8991 29804 9036 29832
rect 8389 29795 8447 29801
rect 9030 29792 9036 29804
rect 9088 29792 9094 29844
rect 10689 29835 10747 29841
rect 10689 29801 10701 29835
rect 10735 29832 10747 29835
rect 10870 29832 10876 29844
rect 10735 29804 10876 29832
rect 10735 29801 10747 29804
rect 10689 29795 10747 29801
rect 10870 29792 10876 29804
rect 10928 29792 10934 29844
rect 10962 29792 10968 29844
rect 11020 29832 11026 29844
rect 11057 29835 11115 29841
rect 11057 29832 11069 29835
rect 11020 29804 11069 29832
rect 11020 29792 11026 29804
rect 11057 29801 11069 29804
rect 11103 29832 11115 29835
rect 11793 29835 11851 29841
rect 11793 29832 11805 29835
rect 11103 29804 11805 29832
rect 11103 29801 11115 29804
rect 11057 29795 11115 29801
rect 11793 29801 11805 29804
rect 11839 29801 11851 29835
rect 11793 29795 11851 29801
rect 13814 29792 13820 29844
rect 13872 29832 13878 29844
rect 18325 29835 18383 29841
rect 13872 29804 13917 29832
rect 13872 29792 13878 29804
rect 18325 29801 18337 29835
rect 18371 29832 18383 29835
rect 18874 29832 18880 29844
rect 18371 29804 18880 29832
rect 18371 29801 18383 29804
rect 18325 29795 18383 29801
rect 18874 29792 18880 29804
rect 18932 29832 18938 29844
rect 20898 29832 20904 29844
rect 18932 29804 20904 29832
rect 18932 29792 18938 29804
rect 20898 29792 20904 29804
rect 20956 29792 20962 29844
rect 23474 29792 23480 29844
rect 23532 29832 23538 29844
rect 26326 29832 26332 29844
rect 23532 29804 23577 29832
rect 26287 29804 26332 29832
rect 23532 29792 23538 29804
rect 26326 29792 26332 29804
rect 26384 29792 26390 29844
rect 31938 29832 31944 29844
rect 31899 29804 31944 29832
rect 31938 29792 31944 29804
rect 31996 29792 32002 29844
rect 34146 29832 34152 29844
rect 34107 29804 34152 29832
rect 34146 29792 34152 29804
rect 34204 29792 34210 29844
rect 34606 29832 34612 29844
rect 34567 29804 34612 29832
rect 34606 29792 34612 29804
rect 34664 29792 34670 29844
rect 34885 29835 34943 29841
rect 34885 29801 34897 29835
rect 34931 29832 34943 29835
rect 35250 29832 35256 29844
rect 34931 29804 35256 29832
rect 34931 29801 34943 29804
rect 34885 29795 34943 29801
rect 35250 29792 35256 29804
rect 35308 29832 35314 29844
rect 36078 29832 36084 29844
rect 35308 29804 36084 29832
rect 35308 29792 35314 29804
rect 36078 29792 36084 29804
rect 36136 29792 36142 29844
rect 37642 29792 37648 29844
rect 37700 29832 37706 29844
rect 38194 29832 38200 29844
rect 37700 29804 38200 29832
rect 37700 29792 37706 29804
rect 38194 29792 38200 29804
rect 38252 29832 38258 29844
rect 41138 29832 41144 29844
rect 38252 29804 41144 29832
rect 38252 29792 38258 29804
rect 41138 29792 41144 29804
rect 41196 29832 41202 29844
rect 41417 29835 41475 29841
rect 41417 29832 41429 29835
rect 41196 29804 41429 29832
rect 41196 29792 41202 29804
rect 41417 29801 41429 29804
rect 41463 29801 41475 29835
rect 42518 29832 42524 29844
rect 42479 29804 42524 29832
rect 41417 29795 41475 29801
rect 42518 29792 42524 29804
rect 42576 29792 42582 29844
rect 4427 29767 4485 29773
rect 4427 29733 4439 29767
rect 4473 29764 4485 29767
rect 4614 29764 4620 29776
rect 4473 29736 4620 29764
rect 4473 29733 4485 29736
rect 4427 29727 4485 29733
rect 4614 29724 4620 29736
rect 4672 29724 4678 29776
rect 7558 29764 7564 29776
rect 7471 29736 7564 29764
rect 7558 29724 7564 29736
rect 7616 29764 7622 29776
rect 7926 29764 7932 29776
rect 7616 29736 7932 29764
rect 7616 29724 7622 29736
rect 7926 29724 7932 29736
rect 7984 29724 7990 29776
rect 8113 29767 8171 29773
rect 8113 29733 8125 29767
rect 8159 29764 8171 29767
rect 8846 29764 8852 29776
rect 8159 29736 8852 29764
rect 8159 29733 8171 29736
rect 8113 29727 8171 29733
rect 8846 29724 8852 29736
rect 8904 29724 8910 29776
rect 12538 29767 12596 29773
rect 12538 29733 12550 29767
rect 12584 29764 12596 29767
rect 12710 29764 12716 29776
rect 12584 29736 12716 29764
rect 12584 29733 12596 29736
rect 12538 29727 12596 29733
rect 12710 29724 12716 29736
rect 12768 29724 12774 29776
rect 13081 29767 13139 29773
rect 13081 29733 13093 29767
rect 13127 29764 13139 29767
rect 13170 29764 13176 29776
rect 13127 29736 13176 29764
rect 13127 29733 13139 29736
rect 13081 29727 13139 29733
rect 5074 29656 5080 29708
rect 5132 29696 5138 29708
rect 5813 29699 5871 29705
rect 5813 29696 5825 29699
rect 5132 29668 5825 29696
rect 5132 29656 5138 29668
rect 5813 29665 5825 29668
rect 5859 29665 5871 29699
rect 5813 29659 5871 29665
rect 5902 29656 5908 29708
rect 5960 29696 5966 29708
rect 6270 29696 6276 29708
rect 5960 29668 6276 29696
rect 5960 29656 5966 29668
rect 6270 29656 6276 29668
rect 6328 29656 6334 29708
rect 9836 29699 9894 29705
rect 9836 29665 9848 29699
rect 9882 29696 9894 29699
rect 10134 29696 10140 29708
rect 9882 29668 10140 29696
rect 9882 29665 9894 29668
rect 9836 29659 9894 29665
rect 10134 29656 10140 29668
rect 10192 29656 10198 29708
rect 10778 29696 10784 29708
rect 10739 29668 10784 29696
rect 10778 29656 10784 29668
rect 10836 29656 10842 29708
rect 11333 29699 11391 29705
rect 11333 29665 11345 29699
rect 11379 29696 11391 29699
rect 11422 29696 11428 29708
rect 11379 29668 11428 29696
rect 11379 29665 11391 29668
rect 11333 29659 11391 29665
rect 11422 29656 11428 29668
rect 11480 29656 11486 29708
rect 3878 29588 3884 29640
rect 3936 29628 3942 29640
rect 4065 29631 4123 29637
rect 4065 29628 4077 29631
rect 3936 29600 4077 29628
rect 3936 29588 3942 29600
rect 4065 29597 4077 29600
rect 4111 29597 4123 29631
rect 4065 29591 4123 29597
rect 6454 29588 6460 29640
rect 6512 29628 6518 29640
rect 7469 29631 7527 29637
rect 7469 29628 7481 29631
rect 6512 29600 7481 29628
rect 6512 29588 6518 29600
rect 7469 29597 7481 29600
rect 7515 29628 7527 29631
rect 8202 29628 8208 29640
rect 7515 29600 8208 29628
rect 7515 29597 7527 29600
rect 7469 29591 7527 29597
rect 8202 29588 8208 29600
rect 8260 29588 8266 29640
rect 12434 29628 12440 29640
rect 12395 29600 12440 29628
rect 12434 29588 12440 29600
rect 12492 29588 12498 29640
rect 12526 29588 12532 29640
rect 12584 29628 12590 29640
rect 13096 29628 13124 29727
rect 13170 29724 13176 29736
rect 13228 29724 13234 29776
rect 15470 29764 15476 29776
rect 15383 29736 15476 29764
rect 15470 29724 15476 29736
rect 15528 29764 15534 29776
rect 16942 29764 16948 29776
rect 15528 29736 16948 29764
rect 15528 29724 15534 29736
rect 16942 29724 16948 29736
rect 17000 29724 17006 29776
rect 17037 29767 17095 29773
rect 17037 29733 17049 29767
rect 17083 29764 17095 29767
rect 17402 29764 17408 29776
rect 17083 29736 17408 29764
rect 17083 29733 17095 29736
rect 17037 29727 17095 29733
rect 17402 29724 17408 29736
rect 17460 29724 17466 29776
rect 22278 29724 22284 29776
rect 22336 29764 22342 29776
rect 22878 29767 22936 29773
rect 22878 29764 22890 29767
rect 22336 29736 22890 29764
rect 22336 29724 22342 29736
rect 22878 29733 22890 29736
rect 22924 29764 22936 29767
rect 23106 29764 23112 29776
rect 22924 29736 23112 29764
rect 22924 29733 22936 29736
rect 22878 29727 22936 29733
rect 23106 29724 23112 29736
rect 23164 29764 23170 29776
rect 24626 29767 24684 29773
rect 24626 29764 24638 29767
rect 23164 29736 24638 29764
rect 23164 29724 23170 29736
rect 24626 29733 24638 29736
rect 24672 29764 24684 29767
rect 24854 29764 24860 29776
rect 24672 29736 24860 29764
rect 24672 29733 24684 29736
rect 24626 29727 24684 29733
rect 24854 29724 24860 29736
rect 24912 29724 24918 29776
rect 25774 29724 25780 29776
rect 25832 29764 25838 29776
rect 26234 29764 26240 29776
rect 25832 29736 26240 29764
rect 25832 29724 25838 29736
rect 26234 29724 26240 29736
rect 26292 29764 26298 29776
rect 26605 29767 26663 29773
rect 26605 29764 26617 29767
rect 26292 29736 26617 29764
rect 26292 29724 26298 29736
rect 26605 29733 26617 29736
rect 26651 29733 26663 29767
rect 26605 29727 26663 29733
rect 26694 29724 26700 29776
rect 26752 29764 26758 29776
rect 28074 29764 28080 29776
rect 26752 29736 28080 29764
rect 26752 29724 26758 29736
rect 28074 29724 28080 29736
rect 28132 29724 28138 29776
rect 30009 29767 30067 29773
rect 30009 29733 30021 29767
rect 30055 29764 30067 29767
rect 30190 29764 30196 29776
rect 30055 29736 30196 29764
rect 30055 29733 30067 29736
rect 30009 29727 30067 29733
rect 30190 29724 30196 29736
rect 30248 29764 30254 29776
rect 30466 29764 30472 29776
rect 30248 29736 30472 29764
rect 30248 29724 30254 29736
rect 30466 29724 30472 29736
rect 30524 29764 30530 29776
rect 32858 29764 32864 29776
rect 30524 29736 32720 29764
rect 32819 29736 32864 29764
rect 30524 29724 30530 29736
rect 13630 29656 13636 29708
rect 13688 29696 13694 29708
rect 13976 29699 14034 29705
rect 13976 29696 13988 29699
rect 13688 29668 13988 29696
rect 13688 29656 13694 29668
rect 13976 29665 13988 29668
rect 14022 29696 14034 29699
rect 14369 29699 14427 29705
rect 14369 29696 14381 29699
rect 14022 29668 14381 29696
rect 14022 29665 14034 29668
rect 13976 29659 14034 29665
rect 14369 29665 14381 29668
rect 14415 29665 14427 29699
rect 18690 29696 18696 29708
rect 18651 29668 18696 29696
rect 14369 29659 14427 29665
rect 18690 29656 18696 29668
rect 18748 29656 18754 29708
rect 18782 29656 18788 29708
rect 18840 29696 18846 29708
rect 18877 29699 18935 29705
rect 18877 29696 18889 29699
rect 18840 29668 18889 29696
rect 18840 29656 18846 29668
rect 18877 29665 18889 29668
rect 18923 29665 18935 29699
rect 21082 29696 21088 29708
rect 21043 29668 21088 29696
rect 18877 29659 18935 29665
rect 21082 29656 21088 29668
rect 21140 29656 21146 29708
rect 21450 29656 21456 29708
rect 21508 29696 21514 29708
rect 21545 29699 21603 29705
rect 21545 29696 21557 29699
rect 21508 29668 21557 29696
rect 21508 29656 21514 29668
rect 21545 29665 21557 29668
rect 21591 29696 21603 29699
rect 22094 29696 22100 29708
rect 21591 29668 22100 29696
rect 21591 29665 21603 29668
rect 21545 29659 21603 29665
rect 22094 29656 22100 29668
rect 22152 29656 22158 29708
rect 23845 29699 23903 29705
rect 23845 29665 23857 29699
rect 23891 29696 23903 29699
rect 24118 29696 24124 29708
rect 23891 29668 24124 29696
rect 23891 29665 23903 29668
rect 23845 29659 23903 29665
rect 24118 29656 24124 29668
rect 24176 29696 24182 29708
rect 25225 29699 25283 29705
rect 25225 29696 25237 29699
rect 24176 29668 25237 29696
rect 24176 29656 24182 29668
rect 25225 29665 25237 29668
rect 25271 29665 25283 29699
rect 28166 29696 28172 29708
rect 28127 29668 28172 29696
rect 25225 29659 25283 29665
rect 28166 29656 28172 29668
rect 28224 29656 28230 29708
rect 28626 29696 28632 29708
rect 28587 29668 28632 29696
rect 28626 29656 28632 29668
rect 28684 29656 28690 29708
rect 30558 29696 30564 29708
rect 30519 29668 30564 29696
rect 30558 29656 30564 29668
rect 30616 29656 30622 29708
rect 30944 29705 30972 29736
rect 30929 29699 30987 29705
rect 30929 29665 30941 29699
rect 30975 29665 30987 29699
rect 30929 29659 30987 29665
rect 31018 29656 31024 29708
rect 31076 29696 31082 29708
rect 32125 29699 32183 29705
rect 32125 29696 32137 29699
rect 31076 29668 32137 29696
rect 31076 29656 31082 29668
rect 32125 29665 32137 29668
rect 32171 29696 32183 29699
rect 32490 29696 32496 29708
rect 32171 29668 32496 29696
rect 32171 29665 32183 29668
rect 32125 29659 32183 29665
rect 32490 29656 32496 29668
rect 32548 29656 32554 29708
rect 32692 29705 32720 29736
rect 32858 29724 32864 29736
rect 32916 29724 32922 29776
rect 33827 29767 33885 29773
rect 33827 29733 33839 29767
rect 33873 29764 33885 29767
rect 33962 29764 33968 29776
rect 33873 29736 33968 29764
rect 33873 29733 33885 29736
rect 33827 29727 33885 29733
rect 33962 29724 33968 29736
rect 34020 29724 34026 29776
rect 35621 29767 35679 29773
rect 35621 29733 35633 29767
rect 35667 29764 35679 29767
rect 35986 29764 35992 29776
rect 35667 29736 35992 29764
rect 35667 29733 35679 29736
rect 35621 29727 35679 29733
rect 35986 29724 35992 29736
rect 36044 29764 36050 29776
rect 36044 29736 36676 29764
rect 36044 29724 36050 29736
rect 32677 29699 32735 29705
rect 32677 29665 32689 29699
rect 32723 29696 32735 29699
rect 32766 29696 32772 29708
rect 32723 29668 32772 29696
rect 32723 29665 32735 29668
rect 32677 29659 32735 29665
rect 32766 29656 32772 29668
rect 32824 29656 32830 29708
rect 33502 29656 33508 29708
rect 33560 29696 33566 29708
rect 33724 29699 33782 29705
rect 33724 29696 33736 29699
rect 33560 29668 33736 29696
rect 33560 29656 33566 29668
rect 33724 29665 33736 29668
rect 33770 29665 33782 29699
rect 33724 29659 33782 29665
rect 34701 29699 34759 29705
rect 34701 29665 34713 29699
rect 34747 29696 34759 29699
rect 35161 29699 35219 29705
rect 35161 29696 35173 29699
rect 34747 29668 35173 29696
rect 34747 29665 34759 29668
rect 34701 29659 34759 29665
rect 35161 29665 35173 29668
rect 35207 29665 35219 29699
rect 36078 29696 36084 29708
rect 36039 29668 36084 29696
rect 35161 29659 35219 29665
rect 15378 29628 15384 29640
rect 12584 29600 13124 29628
rect 15339 29600 15384 29628
rect 12584 29588 12590 29600
rect 15378 29588 15384 29600
rect 15436 29588 15442 29640
rect 16025 29631 16083 29637
rect 16025 29597 16037 29631
rect 16071 29628 16083 29631
rect 16114 29628 16120 29640
rect 16071 29600 16120 29628
rect 16071 29597 16083 29600
rect 16025 29591 16083 29597
rect 16114 29588 16120 29600
rect 16172 29628 16178 29640
rect 16945 29631 17003 29637
rect 16945 29628 16957 29631
rect 16172 29600 16957 29628
rect 16172 29588 16178 29600
rect 16945 29597 16957 29600
rect 16991 29597 17003 29631
rect 17586 29628 17592 29640
rect 17547 29600 17592 29628
rect 16945 29591 17003 29597
rect 17586 29588 17592 29600
rect 17644 29588 17650 29640
rect 18966 29628 18972 29640
rect 18927 29600 18972 29628
rect 18966 29588 18972 29600
rect 19024 29588 19030 29640
rect 21729 29631 21787 29637
rect 21729 29597 21741 29631
rect 21775 29628 21787 29631
rect 22557 29631 22615 29637
rect 22557 29628 22569 29631
rect 21775 29600 22569 29628
rect 21775 29597 21787 29600
rect 21729 29591 21787 29597
rect 22557 29597 22569 29600
rect 22603 29628 22615 29631
rect 23382 29628 23388 29640
rect 22603 29600 23388 29628
rect 22603 29597 22615 29600
rect 22557 29591 22615 29597
rect 23382 29588 23388 29600
rect 23440 29588 23446 29640
rect 23934 29588 23940 29640
rect 23992 29628 23998 29640
rect 24305 29631 24363 29637
rect 24305 29628 24317 29631
rect 23992 29600 24317 29628
rect 23992 29588 23998 29600
rect 24305 29597 24317 29600
rect 24351 29597 24363 29631
rect 28902 29628 28908 29640
rect 28863 29600 28908 29628
rect 24305 29591 24363 29597
rect 28902 29588 28908 29600
rect 28960 29588 28966 29640
rect 31202 29628 31208 29640
rect 31163 29600 31208 29628
rect 31202 29588 31208 29600
rect 31260 29588 31266 29640
rect 33870 29588 33876 29640
rect 33928 29628 33934 29640
rect 34716 29628 34744 29659
rect 36078 29656 36084 29668
rect 36136 29656 36142 29708
rect 36648 29705 36676 29736
rect 38470 29724 38476 29776
rect 38528 29764 38534 29776
rect 38978 29767 39036 29773
rect 38978 29764 38990 29767
rect 38528 29736 38990 29764
rect 38528 29724 38534 29736
rect 38978 29733 38990 29736
rect 39024 29733 39036 29767
rect 40586 29764 40592 29776
rect 40547 29736 40592 29764
rect 38978 29727 39036 29733
rect 40586 29724 40592 29736
rect 40644 29724 40650 29776
rect 43530 29764 43536 29776
rect 43491 29736 43536 29764
rect 43530 29724 43536 29736
rect 43588 29724 43594 29776
rect 36633 29699 36691 29705
rect 36633 29665 36645 29699
rect 36679 29696 36691 29699
rect 37550 29696 37556 29708
rect 36679 29668 37556 29696
rect 36679 29665 36691 29668
rect 36633 29659 36691 29665
rect 37550 29656 37556 29668
rect 37608 29656 37614 29708
rect 41690 29656 41696 29708
rect 41748 29696 41754 29708
rect 42004 29699 42062 29705
rect 42004 29696 42016 29699
rect 41748 29668 42016 29696
rect 41748 29656 41754 29668
rect 42004 29665 42016 29668
rect 42050 29665 42062 29699
rect 42004 29659 42062 29665
rect 36814 29628 36820 29640
rect 33928 29600 34744 29628
rect 36775 29600 36820 29628
rect 33928 29588 33934 29600
rect 36814 29588 36820 29600
rect 36872 29588 36878 29640
rect 37182 29588 37188 29640
rect 37240 29628 37246 29640
rect 38657 29631 38715 29637
rect 38657 29628 38669 29631
rect 37240 29600 38669 29628
rect 37240 29588 37246 29600
rect 38657 29597 38669 29600
rect 38703 29628 38715 29631
rect 39666 29628 39672 29640
rect 38703 29600 39672 29628
rect 38703 29597 38715 29600
rect 38657 29591 38715 29597
rect 39666 29588 39672 29600
rect 39724 29588 39730 29640
rect 40497 29631 40555 29637
rect 40497 29628 40509 29631
rect 40328 29600 40509 29628
rect 14047 29563 14105 29569
rect 14047 29560 14059 29563
rect 13786 29532 14059 29560
rect 13786 29504 13814 29532
rect 14047 29529 14059 29532
rect 14093 29529 14105 29563
rect 14047 29523 14105 29529
rect 18230 29520 18236 29572
rect 18288 29560 18294 29572
rect 22462 29560 22468 29572
rect 18288 29532 22468 29560
rect 18288 29520 18294 29532
rect 22462 29520 22468 29532
rect 22520 29560 22526 29572
rect 23750 29560 23756 29572
rect 22520 29532 23756 29560
rect 22520 29520 22526 29532
rect 23750 29520 23756 29532
rect 23808 29520 23814 29572
rect 23842 29520 23848 29572
rect 23900 29560 23906 29572
rect 24213 29563 24271 29569
rect 24213 29560 24225 29563
rect 23900 29532 24225 29560
rect 23900 29520 23906 29532
rect 24213 29529 24225 29532
rect 24259 29560 24271 29563
rect 27154 29560 27160 29572
rect 24259 29532 27160 29560
rect 24259 29529 24271 29532
rect 24213 29523 24271 29529
rect 27154 29520 27160 29532
rect 27212 29520 27218 29572
rect 40328 29504 40356 29600
rect 40497 29597 40509 29600
rect 40543 29597 40555 29631
rect 41138 29628 41144 29640
rect 41099 29600 41144 29628
rect 40497 29591 40555 29597
rect 41138 29588 41144 29600
rect 41196 29588 41202 29640
rect 42107 29631 42165 29637
rect 42107 29597 42119 29631
rect 42153 29628 42165 29631
rect 43438 29628 43444 29640
rect 42153 29600 43444 29628
rect 42153 29597 42165 29600
rect 42107 29591 42165 29597
rect 43438 29588 43444 29600
rect 43496 29588 43502 29640
rect 43717 29631 43775 29637
rect 43717 29628 43729 29631
rect 43548 29600 43729 29628
rect 41230 29520 41236 29572
rect 41288 29560 41294 29572
rect 42334 29560 42340 29572
rect 41288 29532 42340 29560
rect 41288 29520 41294 29532
rect 42334 29520 42340 29532
rect 42392 29560 42398 29572
rect 43548 29560 43576 29600
rect 43717 29597 43729 29600
rect 43763 29597 43775 29631
rect 43717 29591 43775 29597
rect 42392 29532 43576 29560
rect 42392 29520 42398 29532
rect 3142 29452 3148 29504
rect 3200 29492 3206 29504
rect 3237 29495 3295 29501
rect 3237 29492 3249 29495
rect 3200 29464 3249 29492
rect 3200 29452 3206 29464
rect 3237 29461 3249 29464
rect 3283 29461 3295 29495
rect 3237 29455 3295 29461
rect 4062 29452 4068 29504
rect 4120 29492 4126 29504
rect 4985 29495 5043 29501
rect 4985 29492 4997 29495
rect 4120 29464 4997 29492
rect 4120 29452 4126 29464
rect 4985 29461 4997 29464
rect 5031 29461 5043 29495
rect 6914 29492 6920 29504
rect 6875 29464 6920 29492
rect 4985 29455 5043 29461
rect 6914 29452 6920 29464
rect 6972 29452 6978 29504
rect 9907 29495 9965 29501
rect 9907 29461 9919 29495
rect 9953 29492 9965 29495
rect 11514 29492 11520 29504
rect 9953 29464 11520 29492
rect 9953 29461 9965 29464
rect 9907 29455 9965 29461
rect 11514 29452 11520 29464
rect 11572 29452 11578 29504
rect 13170 29452 13176 29504
rect 13228 29492 13234 29504
rect 13354 29492 13360 29504
rect 13228 29464 13360 29492
rect 13228 29452 13234 29464
rect 13354 29452 13360 29464
rect 13412 29452 13418 29504
rect 13722 29452 13728 29504
rect 13780 29464 13814 29504
rect 19981 29495 20039 29501
rect 13780 29452 13786 29464
rect 19981 29461 19993 29495
rect 20027 29492 20039 29495
rect 20254 29492 20260 29504
rect 20027 29464 20260 29492
rect 20027 29461 20039 29464
rect 19981 29455 20039 29461
rect 20254 29452 20260 29464
rect 20312 29452 20318 29504
rect 20438 29492 20444 29504
rect 20399 29464 20444 29492
rect 20438 29452 20444 29464
rect 20496 29452 20502 29504
rect 25498 29492 25504 29504
rect 25459 29464 25504 29492
rect 25498 29452 25504 29464
rect 25556 29452 25562 29504
rect 39574 29492 39580 29504
rect 39535 29464 39580 29492
rect 39574 29452 39580 29464
rect 39632 29452 39638 29504
rect 40310 29492 40316 29504
rect 40271 29464 40316 29492
rect 40310 29452 40316 29464
rect 40368 29452 40374 29504
rect 1104 29402 48852 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 48852 29402
rect 1104 29328 48852 29350
rect 5166 29288 5172 29300
rect 5127 29260 5172 29288
rect 5166 29248 5172 29260
rect 5224 29248 5230 29300
rect 8202 29288 8208 29300
rect 8163 29260 8208 29288
rect 8202 29248 8208 29260
rect 8260 29248 8266 29300
rect 10778 29288 10784 29300
rect 10739 29260 10784 29288
rect 10778 29248 10784 29260
rect 10836 29248 10842 29300
rect 12986 29248 12992 29300
rect 13044 29288 13050 29300
rect 13725 29291 13783 29297
rect 13725 29288 13737 29291
rect 13044 29260 13737 29288
rect 13044 29248 13050 29260
rect 13725 29257 13737 29260
rect 13771 29288 13783 29291
rect 15381 29291 15439 29297
rect 13771 29260 14412 29288
rect 13771 29257 13783 29260
rect 13725 29251 13783 29257
rect 11606 29180 11612 29232
rect 11664 29220 11670 29232
rect 12253 29223 12311 29229
rect 12253 29220 12265 29223
rect 11664 29192 12265 29220
rect 11664 29180 11670 29192
rect 12253 29189 12265 29192
rect 12299 29220 12311 29223
rect 12710 29220 12716 29232
rect 12299 29192 12716 29220
rect 12299 29189 12311 29192
rect 12253 29183 12311 29189
rect 12710 29180 12716 29192
rect 12768 29220 12774 29232
rect 12768 29192 13814 29220
rect 12768 29180 12774 29192
rect 3421 29155 3479 29161
rect 3421 29121 3433 29155
rect 3467 29152 3479 29155
rect 7190 29152 7196 29164
rect 3467 29124 4154 29152
rect 7151 29124 7196 29152
rect 3467 29121 3479 29124
rect 3421 29115 3479 29121
rect 2593 29087 2651 29093
rect 2593 29053 2605 29087
rect 2639 29084 2651 29087
rect 2958 29084 2964 29096
rect 2639 29056 2964 29084
rect 2639 29053 2651 29056
rect 2593 29047 2651 29053
rect 2958 29044 2964 29056
rect 3016 29044 3022 29096
rect 3234 29084 3240 29096
rect 3195 29056 3240 29084
rect 3234 29044 3240 29056
rect 3292 29044 3298 29096
rect 4126 29084 4154 29124
rect 7190 29112 7196 29124
rect 7248 29112 7254 29164
rect 9769 29155 9827 29161
rect 9769 29121 9781 29155
rect 9815 29152 9827 29155
rect 12802 29152 12808 29164
rect 9815 29124 12808 29152
rect 9815 29121 9827 29124
rect 9769 29115 9827 29121
rect 12802 29112 12808 29124
rect 12860 29112 12866 29164
rect 4249 29087 4307 29093
rect 4249 29084 4261 29087
rect 4126 29056 4261 29084
rect 4249 29053 4261 29056
rect 4295 29084 4307 29087
rect 5445 29087 5503 29093
rect 5445 29084 5457 29087
rect 4295 29056 5457 29084
rect 4295 29053 4307 29056
rect 4249 29047 4307 29053
rect 5445 29053 5457 29056
rect 5491 29053 5503 29087
rect 5445 29047 5503 29053
rect 10778 29044 10784 29096
rect 10836 29084 10842 29096
rect 11000 29087 11058 29093
rect 11000 29084 11012 29087
rect 10836 29056 11012 29084
rect 10836 29044 10842 29056
rect 11000 29053 11012 29056
rect 11046 29084 11058 29087
rect 11793 29087 11851 29093
rect 11793 29084 11805 29087
rect 11046 29056 11805 29084
rect 11046 29053 11058 29056
rect 11000 29047 11058 29053
rect 11793 29053 11805 29056
rect 11839 29053 11851 29087
rect 13786 29084 13814 29192
rect 14384 29161 14412 29260
rect 15381 29257 15393 29291
rect 15427 29288 15439 29291
rect 15470 29288 15476 29300
rect 15427 29260 15476 29288
rect 15427 29257 15439 29260
rect 15381 29251 15439 29257
rect 15470 29248 15476 29260
rect 15528 29248 15534 29300
rect 17862 29288 17868 29300
rect 17823 29260 17868 29288
rect 17862 29248 17868 29260
rect 17920 29248 17926 29300
rect 21450 29288 21456 29300
rect 21411 29260 21456 29288
rect 21450 29248 21456 29260
rect 21508 29248 21514 29300
rect 23106 29288 23112 29300
rect 23067 29260 23112 29288
rect 23106 29248 23112 29260
rect 23164 29248 23170 29300
rect 23382 29288 23388 29300
rect 23343 29260 23388 29288
rect 23382 29248 23388 29260
rect 23440 29248 23446 29300
rect 23934 29288 23940 29300
rect 23895 29260 23940 29288
rect 23934 29248 23940 29260
rect 23992 29248 23998 29300
rect 24578 29288 24584 29300
rect 24539 29260 24584 29288
rect 24578 29248 24584 29260
rect 24636 29248 24642 29300
rect 24854 29288 24860 29300
rect 24815 29260 24860 29288
rect 24854 29248 24860 29260
rect 24912 29288 24918 29300
rect 25225 29291 25283 29297
rect 25225 29288 25237 29291
rect 24912 29260 25237 29288
rect 24912 29248 24918 29260
rect 25225 29257 25237 29260
rect 25271 29257 25283 29291
rect 25225 29251 25283 29257
rect 26329 29291 26387 29297
rect 26329 29257 26341 29291
rect 26375 29288 26387 29291
rect 26418 29288 26424 29300
rect 26375 29260 26424 29288
rect 26375 29257 26387 29260
rect 26329 29251 26387 29257
rect 14369 29155 14427 29161
rect 14369 29121 14381 29155
rect 14415 29121 14427 29155
rect 14642 29152 14648 29164
rect 14603 29124 14648 29152
rect 14369 29115 14427 29121
rect 14642 29112 14648 29124
rect 14700 29152 14706 29164
rect 15378 29152 15384 29164
rect 14700 29124 15384 29152
rect 14700 29112 14706 29124
rect 15378 29112 15384 29124
rect 15436 29152 15442 29164
rect 15657 29155 15715 29161
rect 15657 29152 15669 29155
rect 15436 29124 15669 29152
rect 15436 29112 15442 29124
rect 15657 29121 15669 29124
rect 15703 29121 15715 29155
rect 20438 29152 20444 29164
rect 20399 29124 20444 29152
rect 15657 29115 15715 29121
rect 20438 29112 20444 29124
rect 20496 29112 20502 29164
rect 22741 29155 22799 29161
rect 22741 29121 22753 29155
rect 22787 29152 22799 29155
rect 23952 29152 23980 29248
rect 22787 29124 23980 29152
rect 22787 29121 22799 29124
rect 22741 29115 22799 29121
rect 18874 29084 18880 29096
rect 13786 29056 14228 29084
rect 18835 29056 18880 29084
rect 11793 29047 11851 29053
rect 4522 28976 4528 29028
rect 4580 29016 4586 29028
rect 6914 29016 6920 29028
rect 4580 28988 4660 29016
rect 6875 28988 6920 29016
rect 4580 28976 4586 28988
rect 3789 28951 3847 28957
rect 3789 28917 3801 28951
rect 3835 28948 3847 28951
rect 3970 28948 3976 28960
rect 3835 28920 3976 28948
rect 3835 28917 3847 28920
rect 3789 28911 3847 28917
rect 3970 28908 3976 28920
rect 4028 28948 4034 28960
rect 4632 28957 4660 28988
rect 6914 28976 6920 28988
rect 6972 28976 6978 29028
rect 7009 29019 7067 29025
rect 7009 28985 7021 29019
rect 7055 29016 7067 29019
rect 8478 29016 8484 29028
rect 7055 28988 8484 29016
rect 7055 28985 7067 28988
rect 7009 28979 7067 28985
rect 4065 28951 4123 28957
rect 4065 28948 4077 28951
rect 4028 28920 4077 28948
rect 4028 28908 4034 28920
rect 4065 28917 4077 28920
rect 4111 28917 4123 28951
rect 4065 28911 4123 28917
rect 4617 28951 4675 28957
rect 4617 28917 4629 28951
rect 4663 28917 4675 28951
rect 5810 28948 5816 28960
rect 5771 28920 5816 28948
rect 4617 28911 4675 28917
rect 5810 28908 5816 28920
rect 5868 28908 5874 28960
rect 5902 28908 5908 28960
rect 5960 28948 5966 28960
rect 6181 28951 6239 28957
rect 6181 28948 6193 28951
rect 5960 28920 6193 28948
rect 5960 28908 5966 28920
rect 6181 28917 6193 28920
rect 6227 28917 6239 28951
rect 6181 28911 6239 28917
rect 6641 28951 6699 28957
rect 6641 28917 6653 28951
rect 6687 28948 6699 28951
rect 7024 28948 7052 28979
rect 8478 28976 8484 28988
rect 8536 28976 8542 29028
rect 9122 29016 9128 29028
rect 9083 28988 9128 29016
rect 9122 28976 9128 28988
rect 9180 28976 9186 29028
rect 9217 29019 9275 29025
rect 9217 28985 9229 29019
rect 9263 29016 9275 29019
rect 9858 29016 9864 29028
rect 9263 28988 9864 29016
rect 9263 28985 9275 28988
rect 9217 28979 9275 28985
rect 7926 28948 7932 28960
rect 6687 28920 7052 28948
rect 7887 28920 7932 28948
rect 6687 28917 6699 28920
rect 6641 28911 6699 28917
rect 7926 28908 7932 28920
rect 7984 28908 7990 28960
rect 8938 28948 8944 28960
rect 8851 28920 8944 28948
rect 8938 28908 8944 28920
rect 8996 28948 9002 28960
rect 9232 28948 9260 28979
rect 9858 28976 9864 28988
rect 9916 28976 9922 29028
rect 12526 29016 12532 29028
rect 12487 28988 12532 29016
rect 12526 28976 12532 28988
rect 12584 28976 12590 29028
rect 12621 29019 12679 29025
rect 12621 28985 12633 29019
rect 12667 29016 12679 29019
rect 13814 29016 13820 29028
rect 12667 28988 13032 29016
rect 12667 28985 12679 28988
rect 12621 28979 12679 28985
rect 10134 28948 10140 28960
rect 8996 28920 9260 28948
rect 10095 28920 10140 28948
rect 8996 28908 9002 28920
rect 10134 28908 10140 28920
rect 10192 28908 10198 28960
rect 10870 28908 10876 28960
rect 10928 28948 10934 28960
rect 11103 28951 11161 28957
rect 11103 28948 11115 28951
rect 10928 28920 11115 28948
rect 10928 28908 10934 28920
rect 11103 28917 11115 28920
rect 11149 28917 11161 28951
rect 11422 28948 11428 28960
rect 11383 28920 11428 28948
rect 11103 28911 11161 28917
rect 11422 28908 11428 28920
rect 11480 28908 11486 28960
rect 13004 28948 13032 28988
rect 13280 28988 13820 29016
rect 13280 28948 13308 28988
rect 13814 28976 13820 28988
rect 13872 28976 13878 29028
rect 14200 29025 14228 29056
rect 18874 29044 18880 29056
rect 18932 29044 18938 29096
rect 19797 29087 19855 29093
rect 19797 29053 19809 29087
rect 19843 29084 19855 29087
rect 20162 29084 20168 29096
rect 19843 29056 20168 29084
rect 19843 29053 19855 29056
rect 19797 29047 19855 29053
rect 20162 29044 20168 29056
rect 20220 29044 20226 29096
rect 20254 29044 20260 29096
rect 20312 29084 20318 29096
rect 20349 29087 20407 29093
rect 20349 29084 20361 29087
rect 20312 29056 20361 29084
rect 20312 29044 20318 29056
rect 20349 29053 20361 29056
rect 20395 29084 20407 29087
rect 21726 29084 21732 29096
rect 20395 29056 21732 29084
rect 20395 29053 20407 29056
rect 20349 29047 20407 29053
rect 21726 29044 21732 29056
rect 21784 29044 21790 29096
rect 22002 29084 22008 29096
rect 21836 29056 22008 29084
rect 14185 29019 14243 29025
rect 14185 28985 14197 29019
rect 14231 29016 14243 29019
rect 14461 29019 14519 29025
rect 14461 29016 14473 29019
rect 14231 28988 14473 29016
rect 14231 28985 14243 28988
rect 14185 28979 14243 28985
rect 14461 28985 14473 28988
rect 14507 29016 14519 29019
rect 14734 29016 14740 29028
rect 14507 28988 14740 29016
rect 14507 28985 14519 28988
rect 14461 28979 14519 28985
rect 14715 28976 14740 28988
rect 14792 28976 14798 29028
rect 16482 29016 16488 29028
rect 16443 28988 16488 29016
rect 16482 28976 16488 28988
rect 16540 28976 16546 29028
rect 16577 29019 16635 29025
rect 16577 28985 16589 29019
rect 16623 28985 16635 29019
rect 16577 28979 16635 28985
rect 17129 29019 17187 29025
rect 17129 28985 17141 29019
rect 17175 29016 17187 29019
rect 17218 29016 17224 29028
rect 17175 28988 17224 29016
rect 17175 28985 17187 28988
rect 17129 28979 17187 28985
rect 14715 28966 14780 28976
rect 13004 28920 13308 28948
rect 14752 28948 14780 28966
rect 15470 28948 15476 28960
rect 14752 28920 15476 28948
rect 15470 28908 15476 28920
rect 15528 28908 15534 28960
rect 16301 28951 16359 28957
rect 16301 28917 16313 28951
rect 16347 28948 16359 28951
rect 16592 28948 16620 28979
rect 17218 28976 17224 28988
rect 17276 28976 17282 29028
rect 17494 29016 17500 29028
rect 17407 28988 17500 29016
rect 17494 28976 17500 28988
rect 17552 29016 17558 29028
rect 18233 29019 18291 29025
rect 18233 29016 18245 29019
rect 17552 28988 18245 29016
rect 17552 28976 17558 28988
rect 18233 28985 18245 28988
rect 18279 28985 18291 29019
rect 18233 28979 18291 28985
rect 17034 28948 17040 28960
rect 16347 28920 17040 28948
rect 16347 28917 16359 28920
rect 16301 28911 16359 28917
rect 17034 28908 17040 28920
rect 17092 28908 17098 28960
rect 18690 28908 18696 28960
rect 18748 28948 18754 28960
rect 19337 28951 19395 28957
rect 19337 28948 19349 28951
rect 18748 28920 19349 28948
rect 18748 28908 18754 28920
rect 19337 28917 19349 28920
rect 19383 28948 19395 28951
rect 19426 28948 19432 28960
rect 19383 28920 19432 28948
rect 19383 28917 19395 28920
rect 19337 28911 19395 28917
rect 19426 28908 19432 28920
rect 19484 28948 19490 28960
rect 21082 28948 21088 28960
rect 19484 28920 21088 28948
rect 19484 28908 19490 28920
rect 21082 28908 21088 28920
rect 21140 28908 21146 28960
rect 21174 28908 21180 28960
rect 21232 28948 21238 28960
rect 21836 28957 21864 29056
rect 22002 29044 22008 29056
rect 22060 29044 22066 29096
rect 22094 29044 22100 29096
rect 22152 29084 22158 29096
rect 22465 29087 22523 29093
rect 22465 29084 22477 29087
rect 22152 29056 22477 29084
rect 22152 29044 22158 29056
rect 22465 29053 22477 29056
rect 22511 29053 22523 29087
rect 22465 29047 22523 29053
rect 24397 29087 24455 29093
rect 24397 29053 24409 29087
rect 24443 29053 24455 29087
rect 24397 29047 24455 29053
rect 21821 28951 21879 28957
rect 21821 28948 21833 28951
rect 21232 28920 21833 28948
rect 21232 28908 21238 28920
rect 21821 28917 21833 28920
rect 21867 28917 21879 28951
rect 21821 28911 21879 28917
rect 24305 28951 24363 28957
rect 24305 28917 24317 28951
rect 24351 28948 24363 28951
rect 24412 28948 24440 29047
rect 25240 29016 25268 29251
rect 26418 29248 26424 29260
rect 26476 29248 26482 29300
rect 26694 29288 26700 29300
rect 26655 29260 26700 29288
rect 26694 29248 26700 29260
rect 26752 29248 26758 29300
rect 28074 29288 28080 29300
rect 28035 29260 28080 29288
rect 28074 29248 28080 29260
rect 28132 29248 28138 29300
rect 30190 29288 30196 29300
rect 30151 29260 30196 29288
rect 30190 29248 30196 29260
rect 30248 29248 30254 29300
rect 32125 29291 32183 29297
rect 32125 29257 32137 29291
rect 32171 29288 32183 29291
rect 32398 29288 32404 29300
rect 32171 29260 32404 29288
rect 32171 29257 32183 29260
rect 32125 29251 32183 29257
rect 32398 29248 32404 29260
rect 32456 29248 32462 29300
rect 32490 29248 32496 29300
rect 32548 29288 32554 29300
rect 32766 29288 32772 29300
rect 32548 29260 32593 29288
rect 32727 29260 32772 29288
rect 32548 29248 32554 29260
rect 32766 29248 32772 29260
rect 32824 29248 32830 29300
rect 33735 29291 33793 29297
rect 33735 29257 33747 29291
rect 33781 29288 33793 29291
rect 34606 29288 34612 29300
rect 33781 29260 34612 29288
rect 33781 29257 33793 29260
rect 33735 29251 33793 29257
rect 34606 29248 34612 29260
rect 34664 29248 34670 29300
rect 37550 29288 37556 29300
rect 37511 29260 37556 29288
rect 37550 29248 37556 29260
rect 37608 29248 37614 29300
rect 39574 29248 39580 29300
rect 39632 29288 39638 29300
rect 40221 29291 40279 29297
rect 40221 29288 40233 29291
rect 39632 29260 40233 29288
rect 39632 29248 39638 29260
rect 40221 29257 40233 29260
rect 40267 29288 40279 29291
rect 40586 29288 40592 29300
rect 40267 29260 40592 29288
rect 40267 29257 40279 29260
rect 40221 29251 40279 29257
rect 40586 29248 40592 29260
rect 40644 29248 40650 29300
rect 41601 29291 41659 29297
rect 41601 29257 41613 29291
rect 41647 29288 41659 29291
rect 41874 29288 41880 29300
rect 41647 29260 41880 29288
rect 41647 29257 41659 29260
rect 41601 29251 41659 29257
rect 41874 29248 41880 29260
rect 41932 29288 41938 29300
rect 43441 29291 43499 29297
rect 43441 29288 43453 29291
rect 41932 29260 43453 29288
rect 41932 29248 41938 29260
rect 43441 29257 43453 29260
rect 43487 29288 43499 29291
rect 43530 29288 43536 29300
rect 43487 29260 43536 29288
rect 43487 29257 43499 29260
rect 43441 29251 43499 29257
rect 43530 29248 43536 29260
rect 43588 29248 43594 29300
rect 39666 29220 39672 29232
rect 39627 29192 39672 29220
rect 39666 29180 39672 29192
rect 39724 29180 39730 29232
rect 42518 29220 42524 29232
rect 42168 29192 42524 29220
rect 25409 29155 25467 29161
rect 25409 29121 25421 29155
rect 25455 29152 25467 29155
rect 25498 29152 25504 29164
rect 25455 29124 25504 29152
rect 25455 29121 25467 29124
rect 25409 29115 25467 29121
rect 25498 29112 25504 29124
rect 25556 29112 25562 29164
rect 25866 29112 25872 29164
rect 25924 29152 25930 29164
rect 31202 29152 31208 29164
rect 25924 29124 29316 29152
rect 31163 29124 31208 29152
rect 25924 29112 25930 29124
rect 27154 29084 27160 29096
rect 27115 29056 27160 29084
rect 27154 29044 27160 29056
rect 27212 29044 27218 29096
rect 29288 29093 29316 29124
rect 31202 29112 31208 29124
rect 31260 29112 31266 29164
rect 32950 29112 32956 29164
rect 33008 29152 33014 29164
rect 33410 29152 33416 29164
rect 33008 29124 33416 29152
rect 33008 29112 33014 29124
rect 33410 29112 33416 29124
rect 33468 29112 33474 29164
rect 37182 29152 37188 29164
rect 37143 29124 37188 29152
rect 37182 29112 37188 29124
rect 37240 29112 37246 29164
rect 37274 29112 37280 29164
rect 37332 29152 37338 29164
rect 38102 29152 38108 29164
rect 37332 29124 38108 29152
rect 37332 29112 37338 29124
rect 38102 29112 38108 29124
rect 38160 29112 38166 29164
rect 40034 29112 40040 29164
rect 40092 29152 40098 29164
rect 40589 29155 40647 29161
rect 40589 29152 40601 29155
rect 40092 29124 40601 29152
rect 40092 29112 40098 29124
rect 40589 29121 40601 29124
rect 40635 29152 40647 29155
rect 41230 29152 41236 29164
rect 40635 29124 41236 29152
rect 40635 29121 40647 29124
rect 40589 29115 40647 29121
rect 41230 29112 41236 29124
rect 41288 29112 41294 29164
rect 42168 29161 42196 29192
rect 42518 29180 42524 29192
rect 42576 29180 42582 29232
rect 42153 29155 42211 29161
rect 42153 29121 42165 29155
rect 42199 29121 42211 29155
rect 42426 29152 42432 29164
rect 42387 29124 42432 29152
rect 42153 29115 42211 29121
rect 42426 29112 42432 29124
rect 42484 29112 42490 29164
rect 43438 29112 43444 29164
rect 43496 29152 43502 29164
rect 43717 29155 43775 29161
rect 43717 29152 43729 29155
rect 43496 29124 43729 29152
rect 43496 29112 43502 29124
rect 43717 29121 43729 29124
rect 43763 29121 43775 29155
rect 43717 29115 43775 29121
rect 29273 29087 29331 29093
rect 29273 29053 29285 29087
rect 29319 29084 29331 29087
rect 29733 29087 29791 29093
rect 29733 29084 29745 29087
rect 29319 29056 29745 29084
rect 29319 29053 29331 29056
rect 29273 29047 29331 29053
rect 29733 29053 29745 29056
rect 29779 29053 29791 29087
rect 29733 29047 29791 29053
rect 33664 29087 33722 29093
rect 33664 29053 33676 29087
rect 33710 29084 33722 29087
rect 34146 29084 34152 29096
rect 33710 29056 34152 29084
rect 33710 29053 33722 29056
rect 33664 29047 33722 29053
rect 34146 29044 34152 29056
rect 34204 29044 34210 29096
rect 35250 29084 35256 29096
rect 35211 29056 35256 29084
rect 35250 29044 35256 29056
rect 35308 29044 35314 29096
rect 35529 29087 35587 29093
rect 35529 29053 35541 29087
rect 35575 29084 35587 29087
rect 35986 29084 35992 29096
rect 35575 29056 35992 29084
rect 35575 29053 35587 29056
rect 35529 29047 35587 29053
rect 35986 29044 35992 29056
rect 36044 29044 36050 29096
rect 36817 29087 36875 29093
rect 36817 29053 36829 29087
rect 36863 29084 36875 29087
rect 36906 29084 36912 29096
rect 36863 29056 36912 29084
rect 36863 29053 36875 29056
rect 36817 29047 36875 29053
rect 36906 29044 36912 29056
rect 36964 29044 36970 29096
rect 37093 29087 37151 29093
rect 37093 29053 37105 29087
rect 37139 29084 37151 29087
rect 37550 29084 37556 29096
rect 37139 29056 37556 29084
rect 37139 29053 37151 29056
rect 37093 29047 37151 29053
rect 37550 29044 37556 29056
rect 37608 29044 37614 29096
rect 39025 29087 39083 29093
rect 39025 29053 39037 29087
rect 39071 29084 39083 29087
rect 39071 29056 39849 29084
rect 39071 29053 39083 29056
rect 39025 29047 39083 29053
rect 25730 29019 25788 29025
rect 25730 29016 25742 29019
rect 25240 28988 25742 29016
rect 25730 28985 25742 28988
rect 25776 29016 25788 29019
rect 26973 29019 27031 29025
rect 26973 29016 26985 29019
rect 25776 28988 26985 29016
rect 25776 28985 25788 28988
rect 25730 28979 25788 28985
rect 26973 28985 26985 28988
rect 27019 29016 27031 29019
rect 27478 29019 27536 29025
rect 27478 29016 27490 29019
rect 27019 28988 27490 29016
rect 27019 28985 27031 28988
rect 26973 28979 27031 28985
rect 27478 28985 27490 28988
rect 27524 28985 27536 29019
rect 27478 28979 27536 28985
rect 28258 28976 28264 29028
rect 28316 29016 28322 29028
rect 28626 29016 28632 29028
rect 28316 28988 28632 29016
rect 28316 28976 28322 28988
rect 28626 28976 28632 28988
rect 28684 29016 28690 29028
rect 28721 29019 28779 29025
rect 28721 29016 28733 29019
rect 28684 28988 28733 29016
rect 28684 28976 28690 28988
rect 28721 28985 28733 28988
rect 28767 28985 28779 29019
rect 30558 29016 30564 29028
rect 30519 28988 30564 29016
rect 28721 28979 28779 28985
rect 30558 28976 30564 28988
rect 30616 28976 30622 29028
rect 31526 29019 31584 29025
rect 31526 29016 31538 29019
rect 31036 28988 31538 29016
rect 25406 28948 25412 28960
rect 24351 28920 25412 28948
rect 24351 28917 24363 28920
rect 24305 28911 24363 28917
rect 25406 28908 25412 28920
rect 25464 28908 25470 28960
rect 28074 28908 28080 28960
rect 28132 28948 28138 28960
rect 28353 28951 28411 28957
rect 28353 28948 28365 28951
rect 28132 28920 28365 28948
rect 28132 28908 28138 28920
rect 28353 28917 28365 28920
rect 28399 28917 28411 28951
rect 29454 28948 29460 28960
rect 29415 28920 29460 28948
rect 28353 28911 28411 28917
rect 29454 28908 29460 28920
rect 29512 28908 29518 28960
rect 30374 28908 30380 28960
rect 30432 28948 30438 28960
rect 31036 28948 31064 28988
rect 31526 28985 31538 28988
rect 31572 28985 31584 29019
rect 31526 28979 31584 28985
rect 33502 28976 33508 29028
rect 33560 29016 33566 29028
rect 34425 29019 34483 29025
rect 34425 29016 34437 29019
rect 33560 28988 34437 29016
rect 33560 28976 33566 28988
rect 34425 28985 34437 28988
rect 34471 28985 34483 29019
rect 35710 29016 35716 29028
rect 35671 28988 35716 29016
rect 34425 28979 34483 28985
rect 31110 28948 31116 28960
rect 30432 28920 31116 28948
rect 30432 28908 30438 28920
rect 31110 28908 31116 28920
rect 31168 28908 31174 28960
rect 34146 28948 34152 28960
rect 34107 28920 34152 28948
rect 34146 28908 34152 28920
rect 34204 28908 34210 28960
rect 34440 28948 34468 28979
rect 35710 28976 35716 28988
rect 35768 28976 35774 29028
rect 36078 29016 36084 29028
rect 36039 28988 36084 29016
rect 36078 28976 36084 28988
rect 36136 28976 36142 29028
rect 38467 28997 38525 29003
rect 38467 28994 38479 28997
rect 38396 28966 38479 28994
rect 37642 28948 37648 28960
rect 34440 28920 37648 28948
rect 37642 28908 37648 28920
rect 37700 28908 37706 28960
rect 38013 28951 38071 28957
rect 38013 28917 38025 28951
rect 38059 28948 38071 28951
rect 38194 28948 38200 28960
rect 38059 28920 38200 28948
rect 38059 28917 38071 28920
rect 38013 28911 38071 28917
rect 38194 28908 38200 28920
rect 38252 28948 38258 28960
rect 38396 28948 38424 28966
rect 38467 28963 38479 28966
rect 38513 28963 38525 28997
rect 38467 28957 38525 28963
rect 38252 28920 38424 28948
rect 38252 28908 38258 28920
rect 38562 28908 38568 28960
rect 38620 28948 38626 28960
rect 39301 28951 39359 28957
rect 39301 28948 39313 28951
rect 38620 28920 39313 28948
rect 38620 28908 38626 28920
rect 39301 28917 39313 28920
rect 39347 28917 39359 28951
rect 39821 28948 39849 29056
rect 40681 29019 40739 29025
rect 40681 28985 40693 29019
rect 40727 28985 40739 29019
rect 41230 29016 41236 29028
rect 41191 28988 41236 29016
rect 40681 28979 40739 28985
rect 40696 28948 40724 28979
rect 41230 28976 41236 28988
rect 41288 28976 41294 29028
rect 41966 28976 41972 29028
rect 42024 29016 42030 29028
rect 42245 29019 42303 29025
rect 42245 29016 42257 29019
rect 42024 28988 42257 29016
rect 42024 28976 42030 28988
rect 42245 28985 42257 28988
rect 42291 28985 42303 29019
rect 42245 28979 42303 28985
rect 41138 28948 41144 28960
rect 39821 28920 41144 28948
rect 39301 28911 39359 28917
rect 41138 28908 41144 28920
rect 41196 28908 41202 28960
rect 41690 28908 41696 28960
rect 41748 28948 41754 28960
rect 41877 28951 41935 28957
rect 41877 28948 41889 28951
rect 41748 28920 41889 28948
rect 41748 28908 41754 28920
rect 41877 28917 41889 28920
rect 41923 28917 41935 28951
rect 41877 28911 41935 28917
rect 1104 28858 48852 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 48852 28858
rect 1104 28784 48852 28806
rect 4479 28747 4537 28753
rect 4479 28713 4491 28747
rect 4525 28744 4537 28747
rect 6914 28744 6920 28756
rect 4525 28716 6920 28744
rect 4525 28713 4537 28716
rect 4479 28707 4537 28713
rect 6914 28704 6920 28716
rect 6972 28704 6978 28756
rect 7926 28744 7932 28756
rect 7024 28716 7932 28744
rect 4062 28636 4068 28688
rect 4120 28676 4126 28688
rect 5166 28676 5172 28688
rect 4120 28648 5172 28676
rect 4120 28636 4126 28648
rect 5166 28636 5172 28648
rect 5224 28676 5230 28688
rect 5491 28679 5549 28685
rect 5224 28648 5431 28676
rect 5224 28636 5230 28648
rect 4408 28611 4466 28617
rect 4408 28577 4420 28611
rect 4454 28608 4466 28611
rect 4614 28608 4620 28620
rect 4454 28580 4620 28608
rect 4454 28577 4466 28580
rect 4408 28571 4466 28577
rect 4614 28568 4620 28580
rect 4672 28568 4678 28620
rect 5403 28617 5431 28648
rect 5491 28645 5503 28679
rect 5537 28676 5549 28679
rect 6454 28676 6460 28688
rect 5537 28648 6460 28676
rect 5537 28645 5549 28648
rect 5491 28639 5549 28645
rect 6454 28636 6460 28648
rect 6512 28636 6518 28688
rect 6546 28636 6552 28688
rect 6604 28676 6610 28688
rect 7024 28676 7052 28716
rect 7926 28704 7932 28716
rect 7984 28704 7990 28756
rect 9490 28704 9496 28756
rect 9548 28744 9554 28756
rect 12158 28744 12164 28756
rect 9548 28716 12164 28744
rect 9548 28704 9554 28716
rect 12158 28704 12164 28716
rect 12216 28744 12222 28756
rect 12437 28747 12495 28753
rect 12437 28744 12449 28747
rect 12216 28716 12449 28744
rect 12216 28704 12222 28716
rect 12437 28713 12449 28716
rect 12483 28713 12495 28747
rect 12437 28707 12495 28713
rect 12802 28704 12808 28756
rect 12860 28744 12866 28756
rect 12860 28716 15608 28744
rect 12860 28704 12866 28716
rect 6604 28648 7052 28676
rect 7101 28679 7159 28685
rect 6604 28636 6610 28648
rect 7101 28645 7113 28679
rect 7147 28676 7159 28679
rect 7190 28676 7196 28688
rect 7147 28648 7196 28676
rect 7147 28645 7159 28648
rect 7101 28639 7159 28645
rect 7190 28636 7196 28648
rect 7248 28676 7254 28688
rect 9033 28679 9091 28685
rect 9033 28676 9045 28679
rect 7248 28648 9045 28676
rect 7248 28636 7254 28648
rect 9033 28645 9045 28648
rect 9079 28676 9091 28679
rect 9122 28676 9128 28688
rect 9079 28648 9128 28676
rect 9079 28645 9091 28648
rect 9033 28639 9091 28645
rect 9122 28636 9128 28648
rect 9180 28636 9186 28688
rect 9858 28676 9864 28688
rect 9819 28648 9864 28676
rect 9858 28636 9864 28648
rect 9916 28636 9922 28688
rect 11514 28676 11520 28688
rect 11475 28648 11520 28676
rect 11514 28636 11520 28648
rect 11572 28636 11578 28688
rect 11606 28636 11612 28688
rect 11664 28676 11670 28688
rect 11664 28648 11709 28676
rect 11664 28636 11670 28648
rect 12526 28636 12532 28688
rect 12584 28676 12590 28688
rect 13173 28679 13231 28685
rect 13173 28676 13185 28679
rect 12584 28648 13185 28676
rect 12584 28636 12590 28648
rect 13173 28645 13185 28648
rect 13219 28645 13231 28679
rect 13173 28639 13231 28645
rect 13817 28679 13875 28685
rect 13817 28645 13829 28679
rect 13863 28676 13875 28679
rect 13906 28676 13912 28688
rect 13863 28648 13912 28676
rect 13863 28645 13875 28648
rect 13817 28639 13875 28645
rect 13906 28636 13912 28648
rect 13964 28636 13970 28688
rect 14369 28679 14427 28685
rect 14369 28645 14381 28679
rect 14415 28676 14427 28679
rect 14642 28676 14648 28688
rect 14415 28648 14648 28676
rect 14415 28645 14427 28648
rect 14369 28639 14427 28645
rect 14642 28636 14648 28648
rect 14700 28636 14706 28688
rect 15580 28676 15608 28716
rect 16114 28704 16120 28756
rect 16172 28744 16178 28756
rect 17681 28747 17739 28753
rect 17681 28744 17693 28747
rect 16172 28716 17693 28744
rect 16172 28704 16178 28716
rect 17681 28713 17693 28716
rect 17727 28713 17739 28747
rect 22094 28744 22100 28756
rect 22055 28716 22100 28744
rect 17681 28707 17739 28713
rect 22094 28704 22100 28716
rect 22152 28704 22158 28756
rect 26234 28744 26240 28756
rect 26195 28716 26240 28744
rect 26234 28704 26240 28716
rect 26292 28704 26298 28756
rect 31202 28704 31208 28756
rect 31260 28744 31266 28756
rect 31481 28747 31539 28753
rect 31481 28744 31493 28747
rect 31260 28716 31493 28744
rect 31260 28704 31266 28716
rect 31481 28713 31493 28716
rect 31527 28713 31539 28747
rect 31481 28707 31539 28713
rect 34977 28747 35035 28753
rect 34977 28713 34989 28747
rect 35023 28744 35035 28747
rect 35434 28744 35440 28756
rect 35023 28716 35440 28744
rect 35023 28713 35035 28716
rect 34977 28707 35035 28713
rect 35434 28704 35440 28716
rect 35492 28704 35498 28756
rect 36906 28744 36912 28756
rect 36867 28716 36912 28744
rect 36906 28704 36912 28716
rect 36964 28704 36970 28756
rect 38102 28744 38108 28756
rect 38063 28716 38108 28744
rect 38102 28704 38108 28716
rect 38160 28704 38166 28756
rect 39301 28747 39359 28753
rect 39301 28713 39313 28747
rect 39347 28744 39359 28747
rect 40126 28744 40132 28756
rect 39347 28716 40132 28744
rect 39347 28713 39359 28716
rect 39301 28707 39359 28713
rect 40126 28704 40132 28716
rect 40184 28744 40190 28756
rect 41138 28744 41144 28756
rect 40184 28716 40356 28744
rect 41099 28716 41144 28744
rect 40184 28704 40190 28716
rect 16393 28679 16451 28685
rect 16393 28676 16405 28679
rect 15580 28648 16405 28676
rect 16393 28645 16405 28648
rect 16439 28676 16451 28679
rect 16482 28676 16488 28688
rect 16439 28648 16488 28676
rect 16439 28645 16451 28648
rect 16393 28639 16451 28645
rect 16482 28636 16488 28648
rect 16540 28636 16546 28688
rect 16758 28636 16764 28688
rect 16816 28676 16822 28688
rect 16853 28679 16911 28685
rect 16853 28676 16865 28679
rect 16816 28648 16865 28676
rect 16816 28636 16822 28648
rect 16853 28645 16865 28648
rect 16899 28676 16911 28679
rect 17494 28676 17500 28688
rect 16899 28648 17500 28676
rect 16899 28645 16911 28648
rect 16853 28639 16911 28645
rect 17494 28636 17500 28648
rect 17552 28636 17558 28688
rect 19981 28679 20039 28685
rect 19981 28645 19993 28679
rect 20027 28676 20039 28679
rect 20070 28676 20076 28688
rect 20027 28648 20076 28676
rect 20027 28645 20039 28648
rect 19981 28639 20039 28645
rect 20070 28636 20076 28648
rect 20128 28636 20134 28688
rect 25593 28679 25651 28685
rect 25593 28645 25605 28679
rect 25639 28676 25651 28679
rect 27154 28676 27160 28688
rect 25639 28648 27160 28676
rect 25639 28645 25651 28648
rect 25593 28639 25651 28645
rect 27154 28636 27160 28648
rect 27212 28636 27218 28688
rect 29635 28679 29693 28685
rect 29635 28645 29647 28679
rect 29681 28676 29693 28679
rect 30374 28676 30380 28688
rect 29681 28648 30380 28676
rect 29681 28645 29693 28648
rect 29635 28639 29693 28645
rect 30374 28636 30380 28648
rect 30432 28636 30438 28688
rect 33410 28676 33416 28688
rect 33371 28648 33416 28676
rect 33410 28636 33416 28648
rect 33468 28636 33474 28688
rect 35250 28676 35256 28688
rect 35211 28648 35256 28676
rect 35250 28636 35256 28648
rect 35308 28636 35314 28688
rect 38194 28636 38200 28688
rect 38252 28676 38258 28688
rect 38470 28676 38476 28688
rect 38252 28648 38476 28676
rect 38252 28636 38258 28648
rect 38470 28636 38476 28648
rect 38528 28676 38534 28688
rect 38702 28679 38760 28685
rect 38702 28676 38714 28679
rect 38528 28648 38714 28676
rect 38528 28636 38534 28648
rect 38702 28645 38714 28648
rect 38748 28645 38760 28679
rect 40034 28676 40040 28688
rect 39995 28648 40040 28676
rect 38702 28639 38760 28645
rect 40034 28636 40040 28648
rect 40092 28636 40098 28688
rect 40328 28685 40356 28716
rect 41138 28704 41144 28716
rect 41196 28704 41202 28756
rect 40313 28679 40371 28685
rect 40313 28645 40325 28679
rect 40359 28645 40371 28679
rect 41782 28676 41788 28688
rect 41743 28648 41788 28676
rect 40313 28639 40371 28645
rect 41782 28636 41788 28648
rect 41840 28636 41846 28688
rect 41874 28636 41880 28688
rect 41932 28676 41938 28688
rect 42794 28676 42800 28688
rect 41932 28648 42800 28676
rect 41932 28636 41938 28648
rect 42794 28636 42800 28648
rect 42852 28636 42858 28688
rect 5388 28611 5446 28617
rect 5388 28577 5400 28611
rect 5434 28577 5446 28611
rect 5388 28571 5446 28577
rect 7650 28568 7656 28620
rect 7708 28608 7714 28620
rect 7964 28611 8022 28617
rect 7964 28608 7976 28611
rect 7708 28580 7976 28608
rect 7708 28568 7714 28580
rect 7964 28577 7976 28580
rect 8010 28577 8022 28611
rect 7964 28571 8022 28577
rect 12434 28568 12440 28620
rect 12492 28608 12498 28620
rect 12805 28611 12863 28617
rect 12805 28608 12817 28611
rect 12492 28580 12817 28608
rect 12492 28568 12498 28580
rect 12805 28577 12817 28580
rect 12851 28577 12863 28611
rect 12805 28571 12863 28577
rect 14918 28568 14924 28620
rect 14976 28608 14982 28620
rect 15324 28611 15382 28617
rect 15324 28608 15336 28611
rect 14976 28580 15336 28608
rect 14976 28568 14982 28580
rect 15324 28577 15336 28580
rect 15370 28577 15382 28611
rect 15324 28571 15382 28577
rect 18138 28568 18144 28620
rect 18196 28608 18202 28620
rect 18233 28611 18291 28617
rect 18233 28608 18245 28611
rect 18196 28580 18245 28608
rect 18196 28568 18202 28580
rect 18233 28577 18245 28580
rect 18279 28577 18291 28611
rect 18233 28571 18291 28577
rect 18966 28568 18972 28620
rect 19024 28608 19030 28620
rect 19245 28611 19303 28617
rect 19245 28608 19257 28611
rect 19024 28580 19257 28608
rect 19024 28568 19030 28580
rect 19245 28577 19257 28580
rect 19291 28577 19303 28611
rect 19245 28571 19303 28577
rect 19334 28568 19340 28620
rect 19392 28608 19398 28620
rect 19797 28611 19855 28617
rect 19797 28608 19809 28611
rect 19392 28580 19809 28608
rect 19392 28568 19398 28580
rect 19797 28577 19809 28580
rect 19843 28608 19855 28611
rect 20254 28608 20260 28620
rect 19843 28580 20260 28608
rect 19843 28577 19855 28580
rect 19797 28571 19855 28577
rect 20254 28568 20260 28580
rect 20312 28568 20318 28620
rect 20901 28611 20959 28617
rect 20901 28577 20913 28611
rect 20947 28577 20959 28611
rect 21450 28608 21456 28620
rect 21411 28580 21456 28608
rect 20901 28571 20959 28577
rect 3878 28500 3884 28552
rect 3936 28540 3942 28552
rect 4801 28543 4859 28549
rect 4801 28540 4813 28543
rect 3936 28512 4813 28540
rect 3936 28500 3942 28512
rect 4801 28509 4813 28512
rect 4847 28509 4859 28543
rect 6454 28540 6460 28552
rect 6415 28512 6460 28540
rect 4801 28503 4859 28509
rect 6454 28500 6460 28512
rect 6512 28500 6518 28552
rect 9306 28500 9312 28552
rect 9364 28540 9370 28552
rect 9769 28543 9827 28549
rect 9769 28540 9781 28543
rect 9364 28512 9781 28540
rect 9364 28500 9370 28512
rect 9769 28509 9781 28512
rect 9815 28509 9827 28543
rect 9769 28503 9827 28509
rect 10413 28543 10471 28549
rect 10413 28509 10425 28543
rect 10459 28540 10471 28543
rect 11974 28540 11980 28552
rect 10459 28512 11980 28540
rect 10459 28509 10471 28512
rect 10413 28503 10471 28509
rect 11974 28500 11980 28512
rect 12032 28500 12038 28552
rect 12161 28543 12219 28549
rect 12161 28509 12173 28543
rect 12207 28540 12219 28543
rect 12526 28540 12532 28552
rect 12207 28512 12532 28540
rect 12207 28509 12219 28512
rect 12161 28503 12219 28509
rect 12526 28500 12532 28512
rect 12584 28500 12590 28552
rect 13722 28540 13728 28552
rect 13635 28512 13728 28540
rect 13722 28500 13728 28512
rect 13780 28540 13786 28552
rect 14366 28540 14372 28552
rect 13780 28512 14372 28540
rect 13780 28500 13786 28512
rect 14366 28500 14372 28512
rect 14424 28500 14430 28552
rect 16574 28500 16580 28552
rect 16632 28540 16638 28552
rect 16761 28543 16819 28549
rect 16761 28540 16773 28543
rect 16632 28512 16773 28540
rect 16632 28500 16638 28512
rect 16761 28509 16773 28512
rect 16807 28509 16819 28543
rect 17218 28540 17224 28552
rect 17179 28512 17224 28540
rect 16761 28503 16819 28509
rect 17218 28500 17224 28512
rect 17276 28500 17282 28552
rect 17678 28500 17684 28552
rect 17736 28540 17742 28552
rect 20916 28540 20944 28571
rect 21450 28568 21456 28580
rect 21508 28568 21514 28620
rect 22462 28608 22468 28620
rect 22423 28580 22468 28608
rect 22462 28568 22468 28580
rect 22520 28568 22526 28620
rect 23017 28611 23075 28617
rect 23017 28577 23029 28611
rect 23063 28608 23075 28611
rect 23106 28608 23112 28620
rect 23063 28580 23112 28608
rect 23063 28577 23075 28580
rect 23017 28571 23075 28577
rect 23106 28568 23112 28580
rect 23164 28568 23170 28620
rect 25133 28611 25191 28617
rect 25133 28577 25145 28611
rect 25179 28608 25191 28611
rect 25406 28608 25412 28620
rect 25179 28580 25268 28608
rect 25367 28580 25412 28608
rect 25179 28577 25191 28580
rect 25133 28571 25191 28577
rect 25240 28552 25268 28580
rect 25406 28568 25412 28580
rect 25464 28568 25470 28620
rect 26580 28611 26638 28617
rect 26580 28577 26592 28611
rect 26626 28577 26638 28611
rect 26580 28571 26638 28577
rect 21174 28540 21180 28552
rect 17736 28512 21180 28540
rect 17736 28500 17742 28512
rect 21174 28500 21180 28512
rect 21232 28500 21238 28552
rect 21542 28540 21548 28552
rect 21503 28512 21548 28540
rect 21542 28500 21548 28512
rect 21600 28500 21606 28552
rect 23198 28540 23204 28552
rect 23159 28512 23204 28540
rect 23198 28500 23204 28512
rect 23256 28500 23262 28552
rect 25222 28540 25228 28552
rect 23446 28512 25228 28540
rect 20162 28432 20168 28484
rect 20220 28472 20226 28484
rect 23446 28472 23474 28512
rect 25222 28500 25228 28512
rect 25280 28500 25286 28552
rect 26595 28540 26623 28571
rect 27522 28568 27528 28620
rect 27580 28608 27586 28620
rect 27982 28608 27988 28620
rect 27580 28580 27988 28608
rect 27580 28568 27586 28580
rect 27982 28568 27988 28580
rect 28040 28568 28046 28620
rect 28258 28608 28264 28620
rect 28219 28580 28264 28608
rect 28258 28568 28264 28580
rect 28316 28568 28322 28620
rect 31018 28608 31024 28620
rect 30979 28580 31024 28608
rect 31018 28568 31024 28580
rect 31076 28568 31082 28620
rect 32284 28611 32342 28617
rect 32284 28577 32296 28611
rect 32330 28608 32342 28611
rect 32950 28608 32956 28620
rect 32330 28580 32956 28608
rect 32330 28577 32342 28580
rect 32284 28571 32342 28577
rect 32950 28568 32956 28580
rect 33008 28568 33014 28620
rect 34606 28568 34612 28620
rect 34664 28608 34670 28620
rect 34793 28611 34851 28617
rect 34793 28608 34805 28611
rect 34664 28580 34805 28608
rect 34664 28568 34670 28580
rect 34793 28577 34805 28580
rect 34839 28577 34851 28611
rect 34793 28571 34851 28577
rect 35618 28568 35624 28620
rect 35676 28608 35682 28620
rect 35897 28611 35955 28617
rect 35897 28608 35909 28611
rect 35676 28580 35909 28608
rect 35676 28568 35682 28580
rect 35897 28577 35909 28580
rect 35943 28577 35955 28611
rect 35897 28571 35955 28577
rect 35986 28568 35992 28620
rect 36044 28608 36050 28620
rect 36357 28611 36415 28617
rect 36357 28608 36369 28611
rect 36044 28580 36369 28608
rect 36044 28568 36050 28580
rect 36357 28577 36369 28580
rect 36403 28577 36415 28611
rect 36357 28571 36415 28577
rect 36814 28568 36820 28620
rect 36872 28608 36878 28620
rect 38381 28611 38439 28617
rect 38381 28608 38393 28611
rect 36872 28580 38393 28608
rect 36872 28568 36878 28580
rect 38381 28577 38393 28580
rect 38427 28608 38439 28611
rect 38838 28608 38844 28620
rect 38427 28580 38844 28608
rect 38427 28577 38439 28580
rect 38381 28571 38439 28577
rect 38838 28568 38844 28580
rect 38896 28568 38902 28620
rect 27154 28540 27160 28552
rect 26595 28512 27160 28540
rect 27154 28500 27160 28512
rect 27212 28500 27218 28552
rect 28445 28543 28503 28549
rect 28445 28509 28457 28543
rect 28491 28540 28503 28543
rect 29178 28540 29184 28552
rect 28491 28512 29184 28540
rect 28491 28509 28503 28512
rect 28445 28503 28503 28509
rect 29178 28500 29184 28512
rect 29236 28540 29242 28552
rect 29273 28543 29331 28549
rect 29273 28540 29285 28543
rect 29236 28512 29285 28540
rect 29236 28500 29242 28512
rect 29273 28509 29285 28512
rect 29319 28509 29331 28543
rect 33318 28540 33324 28552
rect 33279 28512 33324 28540
rect 29273 28503 29331 28509
rect 33318 28500 33324 28512
rect 33376 28500 33382 28552
rect 33686 28540 33692 28552
rect 33647 28512 33692 28540
rect 33686 28500 33692 28512
rect 33744 28500 33750 28552
rect 36446 28540 36452 28552
rect 36407 28512 36452 28540
rect 36446 28500 36452 28512
rect 36504 28500 36510 28552
rect 40221 28543 40279 28549
rect 40221 28509 40233 28543
rect 40267 28540 40279 28543
rect 40678 28540 40684 28552
rect 40267 28512 40684 28540
rect 40267 28509 40279 28512
rect 40221 28503 40279 28509
rect 40678 28500 40684 28512
rect 40736 28500 40742 28552
rect 42429 28543 42487 28549
rect 42429 28509 42441 28543
rect 42475 28540 42487 28543
rect 42518 28540 42524 28552
rect 42475 28512 42524 28540
rect 42475 28509 42487 28512
rect 42429 28503 42487 28509
rect 42518 28500 42524 28512
rect 42576 28500 42582 28552
rect 20220 28444 23474 28472
rect 32355 28475 32413 28481
rect 20220 28432 20226 28444
rect 32355 28441 32367 28475
rect 32401 28472 32413 28475
rect 32401 28444 33134 28472
rect 32401 28441 32413 28444
rect 32355 28435 32413 28441
rect 33106 28416 33134 28444
rect 39942 28432 39948 28484
rect 40000 28472 40006 28484
rect 40773 28475 40831 28481
rect 40773 28472 40785 28475
rect 40000 28444 40785 28472
rect 40000 28432 40006 28444
rect 40773 28441 40785 28444
rect 40819 28472 40831 28475
rect 41230 28472 41236 28484
rect 40819 28444 41236 28472
rect 40819 28441 40831 28444
rect 40773 28435 40831 28441
rect 41230 28432 41236 28444
rect 41288 28432 41294 28484
rect 2777 28407 2835 28413
rect 2777 28373 2789 28407
rect 2823 28404 2835 28407
rect 3234 28404 3240 28416
rect 2823 28376 3240 28404
rect 2823 28373 2835 28376
rect 2777 28367 2835 28373
rect 3234 28364 3240 28376
rect 3292 28404 3298 28416
rect 5350 28404 5356 28416
rect 3292 28376 5356 28404
rect 3292 28364 3298 28376
rect 5350 28364 5356 28376
rect 5408 28364 5414 28416
rect 8067 28407 8125 28413
rect 8067 28373 8079 28407
rect 8113 28404 8125 28407
rect 8202 28404 8208 28416
rect 8113 28376 8208 28404
rect 8113 28373 8125 28376
rect 8067 28367 8125 28373
rect 8202 28364 8208 28376
rect 8260 28404 8266 28416
rect 8389 28407 8447 28413
rect 8389 28404 8401 28407
rect 8260 28376 8401 28404
rect 8260 28364 8266 28376
rect 8389 28373 8401 28376
rect 8435 28373 8447 28407
rect 8389 28367 8447 28373
rect 15286 28364 15292 28416
rect 15344 28404 15350 28416
rect 15427 28407 15485 28413
rect 15427 28404 15439 28407
rect 15344 28376 15439 28404
rect 15344 28364 15350 28376
rect 15427 28373 15439 28376
rect 15473 28373 15485 28407
rect 15427 28367 15485 28373
rect 15841 28407 15899 28413
rect 15841 28373 15853 28407
rect 15887 28404 15899 28407
rect 16022 28404 16028 28416
rect 15887 28376 16028 28404
rect 15887 28373 15899 28376
rect 15841 28367 15899 28373
rect 16022 28364 16028 28376
rect 16080 28364 16086 28416
rect 18230 28364 18236 28416
rect 18288 28404 18294 28416
rect 18371 28407 18429 28413
rect 18371 28404 18383 28407
rect 18288 28376 18383 28404
rect 18288 28364 18294 28376
rect 18371 28373 18383 28376
rect 18417 28373 18429 28407
rect 18371 28367 18429 28373
rect 24210 28364 24216 28416
rect 24268 28404 24274 28416
rect 26651 28407 26709 28413
rect 26651 28404 26663 28407
rect 24268 28376 26663 28404
rect 24268 28364 24274 28376
rect 26651 28373 26663 28376
rect 26697 28373 26709 28407
rect 26651 28367 26709 28373
rect 27617 28407 27675 28413
rect 27617 28373 27629 28407
rect 27663 28404 27675 28407
rect 28258 28404 28264 28416
rect 27663 28376 28264 28404
rect 27663 28373 27675 28376
rect 27617 28367 27675 28373
rect 28258 28364 28264 28376
rect 28316 28364 28322 28416
rect 30190 28404 30196 28416
rect 30151 28376 30196 28404
rect 30190 28364 30196 28376
rect 30248 28364 30254 28416
rect 30466 28404 30472 28416
rect 30427 28376 30472 28404
rect 30466 28364 30472 28376
rect 30524 28364 30530 28416
rect 31202 28404 31208 28416
rect 31163 28376 31208 28404
rect 31202 28364 31208 28376
rect 31260 28364 31266 28416
rect 32490 28364 32496 28416
rect 32548 28404 32554 28416
rect 32677 28407 32735 28413
rect 32677 28404 32689 28407
rect 32548 28376 32689 28404
rect 32548 28364 32554 28376
rect 32677 28373 32689 28376
rect 32723 28373 32735 28407
rect 33106 28376 33140 28416
rect 32677 28367 32735 28373
rect 33134 28364 33140 28376
rect 33192 28364 33198 28416
rect 1104 28314 48852 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 48852 28314
rect 1104 28240 48852 28262
rect 5166 28200 5172 28212
rect 5127 28172 5172 28200
rect 5166 28160 5172 28172
rect 5224 28160 5230 28212
rect 6365 28203 6423 28209
rect 6365 28169 6377 28203
rect 6411 28200 6423 28203
rect 6546 28200 6552 28212
rect 6411 28172 6552 28200
rect 6411 28169 6423 28172
rect 6365 28163 6423 28169
rect 6546 28160 6552 28172
rect 6604 28160 6610 28212
rect 7650 28200 7656 28212
rect 7611 28172 7656 28200
rect 7650 28160 7656 28172
rect 7708 28160 7714 28212
rect 9306 28200 9312 28212
rect 8772 28172 9312 28200
rect 8772 28144 8800 28172
rect 9306 28160 9312 28172
rect 9364 28160 9370 28212
rect 9858 28160 9864 28212
rect 9916 28200 9922 28212
rect 10229 28203 10287 28209
rect 10229 28200 10241 28203
rect 9916 28172 10241 28200
rect 9916 28160 9922 28172
rect 10229 28169 10241 28172
rect 10275 28169 10287 28203
rect 10229 28163 10287 28169
rect 11514 28160 11520 28212
rect 11572 28200 11578 28212
rect 12161 28203 12219 28209
rect 12161 28200 12173 28203
rect 11572 28172 12173 28200
rect 11572 28160 11578 28172
rect 12161 28169 12173 28172
rect 12207 28169 12219 28203
rect 12161 28163 12219 28169
rect 13630 28160 13636 28212
rect 13688 28200 13694 28212
rect 13725 28203 13783 28209
rect 13725 28200 13737 28203
rect 13688 28172 13737 28200
rect 13688 28160 13694 28172
rect 13725 28169 13737 28172
rect 13771 28169 13783 28203
rect 13725 28163 13783 28169
rect 13906 28160 13912 28212
rect 13964 28200 13970 28212
rect 14001 28203 14059 28209
rect 14001 28200 14013 28203
rect 13964 28172 14013 28200
rect 13964 28160 13970 28172
rect 14001 28169 14013 28172
rect 14047 28169 14059 28203
rect 14366 28200 14372 28212
rect 14327 28172 14372 28200
rect 14001 28163 14059 28169
rect 14366 28160 14372 28172
rect 14424 28160 14430 28212
rect 15289 28203 15347 28209
rect 15289 28169 15301 28203
rect 15335 28200 15347 28203
rect 15654 28200 15660 28212
rect 15335 28172 15660 28200
rect 15335 28169 15347 28172
rect 15289 28163 15347 28169
rect 5491 28135 5549 28141
rect 5491 28101 5503 28135
rect 5537 28132 5549 28135
rect 6454 28132 6460 28144
rect 5537 28104 6460 28132
rect 5537 28101 5549 28104
rect 5491 28095 5549 28101
rect 6454 28092 6460 28104
rect 6512 28092 6518 28144
rect 8754 28132 8760 28144
rect 8667 28104 8760 28132
rect 8754 28092 8760 28104
rect 8812 28092 8818 28144
rect 11606 28132 11612 28144
rect 9324 28104 11612 28132
rect 4062 28064 4068 28076
rect 4023 28036 4068 28064
rect 4062 28024 4068 28036
rect 4120 28024 4126 28076
rect 8202 28064 8208 28076
rect 8163 28036 8208 28064
rect 8202 28024 8208 28036
rect 8260 28024 8266 28076
rect 2958 27956 2964 28008
rect 3016 27996 3022 28008
rect 3421 27999 3479 28005
rect 3421 27996 3433 27999
rect 3016 27968 3433 27996
rect 3016 27956 3022 27968
rect 3421 27965 3433 27968
rect 3467 27996 3479 27999
rect 3786 27996 3792 28008
rect 3467 27968 3792 27996
rect 3467 27965 3479 27968
rect 3421 27959 3479 27965
rect 3786 27956 3792 27968
rect 3844 27956 3850 28008
rect 3878 27956 3884 28008
rect 3936 27996 3942 28008
rect 3973 27999 4031 28005
rect 3973 27996 3985 27999
rect 3936 27968 3985 27996
rect 3936 27956 3942 27968
rect 3973 27965 3985 27968
rect 4019 27965 4031 27999
rect 3973 27959 4031 27965
rect 5166 27956 5172 28008
rect 5224 27996 5230 28008
rect 5420 27999 5478 28005
rect 5420 27996 5432 27999
rect 5224 27968 5432 27996
rect 5224 27956 5230 27968
rect 5420 27965 5432 27968
rect 5466 27996 5478 27999
rect 5813 27999 5871 28005
rect 5813 27996 5825 27999
rect 5466 27968 5825 27996
rect 5466 27965 5478 27968
rect 5420 27959 5478 27965
rect 5813 27965 5825 27968
rect 5859 27965 5871 27999
rect 5813 27959 5871 27965
rect 7168 27999 7226 28005
rect 7168 27965 7180 27999
rect 7214 27996 7226 27999
rect 7558 27996 7564 28008
rect 7214 27968 7564 27996
rect 7214 27965 7226 27968
rect 7168 27959 7226 27965
rect 7558 27956 7564 27968
rect 7616 27956 7622 28008
rect 7926 27888 7932 27940
rect 7984 27928 7990 27940
rect 8021 27931 8079 27937
rect 8021 27928 8033 27931
rect 7984 27900 8033 27928
rect 7984 27888 7990 27900
rect 8021 27897 8033 27900
rect 8067 27928 8079 27931
rect 8297 27931 8355 27937
rect 8297 27928 8309 27931
rect 8067 27900 8309 27928
rect 8067 27897 8079 27900
rect 8021 27891 8079 27897
rect 8297 27897 8309 27900
rect 8343 27928 8355 27931
rect 9324 27928 9352 28104
rect 11606 28092 11612 28104
rect 11664 28132 11670 28144
rect 11793 28135 11851 28141
rect 11793 28132 11805 28135
rect 11664 28104 11805 28132
rect 11664 28092 11670 28104
rect 11793 28101 11805 28104
rect 11839 28101 11851 28135
rect 11793 28095 11851 28101
rect 10870 28064 10876 28076
rect 10831 28036 10876 28064
rect 10870 28024 10876 28036
rect 10928 28024 10934 28076
rect 12158 28024 12164 28076
rect 12216 28064 12222 28076
rect 13814 28064 13820 28076
rect 12216 28036 13820 28064
rect 12216 28024 12222 28036
rect 13814 28024 13820 28036
rect 13872 28064 13878 28076
rect 15304 28064 15332 28163
rect 15654 28160 15660 28172
rect 15712 28160 15718 28212
rect 16758 28200 16764 28212
rect 16719 28172 16764 28200
rect 16758 28160 16764 28172
rect 16816 28160 16822 28212
rect 17126 28200 17132 28212
rect 17087 28172 17132 28200
rect 17126 28160 17132 28172
rect 17184 28160 17190 28212
rect 17865 28203 17923 28209
rect 17865 28169 17877 28203
rect 17911 28200 17923 28203
rect 18138 28200 18144 28212
rect 17911 28172 18144 28200
rect 17911 28169 17923 28172
rect 17865 28163 17923 28169
rect 18138 28160 18144 28172
rect 18196 28200 18202 28212
rect 21634 28200 21640 28212
rect 18196 28172 21640 28200
rect 18196 28160 18202 28172
rect 21634 28160 21640 28172
rect 21692 28200 21698 28212
rect 26743 28203 26801 28209
rect 26743 28200 26755 28203
rect 21692 28172 26755 28200
rect 21692 28160 21698 28172
rect 26743 28169 26755 28172
rect 26789 28169 26801 28203
rect 27154 28200 27160 28212
rect 27115 28172 27160 28200
rect 26743 28163 26801 28169
rect 27154 28160 27160 28172
rect 27212 28160 27218 28212
rect 27246 28160 27252 28212
rect 27304 28200 27310 28212
rect 27522 28200 27528 28212
rect 27304 28172 27528 28200
rect 27304 28160 27310 28172
rect 27522 28160 27528 28172
rect 27580 28160 27586 28212
rect 31849 28203 31907 28209
rect 31849 28169 31861 28203
rect 31895 28200 31907 28203
rect 32950 28200 32956 28212
rect 31895 28172 32956 28200
rect 31895 28169 31907 28172
rect 31849 28163 31907 28169
rect 32950 28160 32956 28172
rect 33008 28160 33014 28212
rect 33318 28160 33324 28212
rect 33376 28200 33382 28212
rect 33873 28203 33931 28209
rect 33873 28200 33885 28203
rect 33376 28172 33885 28200
rect 33376 28160 33382 28172
rect 33873 28169 33885 28172
rect 33919 28200 33931 28203
rect 35023 28203 35081 28209
rect 35023 28200 35035 28203
rect 33919 28172 35035 28200
rect 33919 28169 33931 28172
rect 33873 28163 33931 28169
rect 35023 28169 35035 28172
rect 35069 28169 35081 28203
rect 35023 28163 35081 28169
rect 35618 28160 35624 28212
rect 35676 28200 35682 28212
rect 35713 28203 35771 28209
rect 35713 28200 35725 28203
rect 35676 28172 35725 28200
rect 35676 28160 35682 28172
rect 35713 28169 35725 28172
rect 35759 28169 35771 28203
rect 38838 28200 38844 28212
rect 38799 28172 38844 28200
rect 35713 28163 35771 28169
rect 38838 28160 38844 28172
rect 38896 28160 38902 28212
rect 40126 28200 40132 28212
rect 40087 28172 40132 28200
rect 40126 28160 40132 28172
rect 40184 28160 40190 28212
rect 42794 28160 42800 28212
rect 42852 28200 42858 28212
rect 42852 28172 42897 28200
rect 42852 28160 42858 28172
rect 16942 28132 16948 28144
rect 16855 28104 16948 28132
rect 16942 28092 16948 28104
rect 17000 28132 17006 28144
rect 17497 28135 17555 28141
rect 17497 28132 17509 28135
rect 17000 28104 17509 28132
rect 17000 28092 17006 28104
rect 17497 28101 17509 28104
rect 17543 28132 17555 28135
rect 20990 28132 20996 28144
rect 17543 28104 20996 28132
rect 17543 28101 17555 28104
rect 17497 28095 17555 28101
rect 20990 28092 20996 28104
rect 21048 28092 21054 28144
rect 21174 28132 21180 28144
rect 21135 28104 21180 28132
rect 21174 28092 21180 28104
rect 21232 28092 21238 28144
rect 21450 28092 21456 28144
rect 21508 28132 21514 28144
rect 21545 28135 21603 28141
rect 21545 28132 21557 28135
rect 21508 28104 21557 28132
rect 21508 28092 21514 28104
rect 21545 28101 21557 28104
rect 21591 28132 21603 28135
rect 23106 28132 23112 28144
rect 21591 28104 23112 28132
rect 21591 28101 21603 28104
rect 21545 28095 21603 28101
rect 23106 28092 23112 28104
rect 23164 28092 23170 28144
rect 24673 28135 24731 28141
rect 24673 28101 24685 28135
rect 24719 28132 24731 28135
rect 25130 28132 25136 28144
rect 24719 28104 25136 28132
rect 24719 28101 24731 28104
rect 24673 28095 24731 28101
rect 25130 28092 25136 28104
rect 25188 28092 25194 28144
rect 25406 28132 25412 28144
rect 25319 28104 25412 28132
rect 16114 28064 16120 28076
rect 13872 28036 15332 28064
rect 16075 28036 16120 28064
rect 13872 28024 13878 28036
rect 16114 28024 16120 28036
rect 16172 28024 16178 28076
rect 9769 27999 9827 28005
rect 9769 27996 9781 27999
rect 8343 27900 9352 27928
rect 9692 27968 9781 27996
rect 8343 27897 8355 27900
rect 8297 27891 8355 27897
rect 9692 27872 9720 27968
rect 9769 27965 9781 27968
rect 9815 27965 9827 27999
rect 12802 27996 12808 28008
rect 12763 27968 12808 27996
rect 9769 27959 9827 27965
rect 12802 27956 12808 27968
rect 12860 27956 12866 28008
rect 16960 28005 16988 28092
rect 17034 28024 17040 28076
rect 17092 28064 17098 28076
rect 18141 28067 18199 28073
rect 18141 28064 18153 28067
rect 17092 28036 18153 28064
rect 17092 28024 17098 28036
rect 18141 28033 18153 28036
rect 18187 28033 18199 28067
rect 18141 28027 18199 28033
rect 19058 28024 19064 28076
rect 19116 28064 19122 28076
rect 22097 28067 22155 28073
rect 22097 28064 22109 28067
rect 19116 28036 22109 28064
rect 19116 28024 19122 28036
rect 22097 28033 22109 28036
rect 22143 28064 22155 28067
rect 22278 28064 22284 28076
rect 22143 28036 22284 28064
rect 22143 28033 22155 28036
rect 22097 28027 22155 28033
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 22462 28024 22468 28076
rect 22520 28064 22526 28076
rect 22741 28067 22799 28073
rect 22741 28064 22753 28067
rect 22520 28036 22753 28064
rect 22520 28024 22526 28036
rect 22741 28033 22753 28036
rect 22787 28064 22799 28067
rect 25222 28064 25228 28076
rect 22787 28036 25228 28064
rect 22787 28033 22799 28036
rect 22741 28027 22799 28033
rect 25222 28024 25228 28036
rect 25280 28024 25286 28076
rect 16945 27999 17003 28005
rect 16945 27965 16957 27999
rect 16991 27965 17003 27999
rect 18230 27996 18236 28008
rect 18191 27968 18236 27996
rect 16945 27959 17003 27965
rect 18230 27956 18236 27968
rect 18288 27956 18294 28008
rect 20073 27999 20131 28005
rect 20073 27965 20085 27999
rect 20119 27965 20131 27999
rect 20073 27959 20131 27965
rect 20625 27999 20683 28005
rect 20625 27965 20637 27999
rect 20671 27965 20683 27999
rect 20625 27959 20683 27965
rect 20809 27999 20867 28005
rect 20809 27965 20821 27999
rect 20855 27996 20867 27999
rect 21082 27996 21088 28008
rect 20855 27968 21088 27996
rect 20855 27965 20867 27968
rect 20809 27959 20867 27965
rect 10686 27928 10692 27940
rect 10599 27900 10692 27928
rect 10686 27888 10692 27900
rect 10744 27928 10750 27940
rect 10965 27931 11023 27937
rect 10965 27928 10977 27931
rect 10744 27900 10977 27928
rect 10744 27888 10750 27900
rect 10965 27897 10977 27900
rect 11011 27897 11023 27931
rect 10965 27891 11023 27897
rect 11517 27931 11575 27937
rect 11517 27897 11529 27931
rect 11563 27928 11575 27931
rect 12526 27928 12532 27940
rect 11563 27900 12532 27928
rect 11563 27897 11575 27900
rect 11517 27891 11575 27897
rect 4614 27860 4620 27872
rect 4575 27832 4620 27860
rect 4614 27820 4620 27832
rect 4672 27820 4678 27872
rect 7239 27863 7297 27869
rect 7239 27829 7251 27863
rect 7285 27860 7297 27863
rect 7834 27860 7840 27872
rect 7285 27832 7840 27860
rect 7285 27829 7297 27832
rect 7239 27823 7297 27829
rect 7834 27820 7840 27832
rect 7892 27820 7898 27872
rect 9674 27860 9680 27872
rect 9635 27832 9680 27860
rect 9674 27820 9680 27832
rect 9732 27820 9738 27872
rect 9950 27860 9956 27872
rect 9911 27832 9956 27860
rect 9950 27820 9956 27832
rect 10008 27820 10014 27872
rect 10980 27860 11008 27891
rect 12526 27888 12532 27900
rect 12584 27888 12590 27940
rect 12713 27931 12771 27937
rect 12713 27897 12725 27931
rect 12759 27928 12771 27931
rect 13126 27931 13184 27937
rect 13126 27928 13138 27931
rect 12759 27900 13138 27928
rect 12759 27897 12771 27900
rect 12713 27891 12771 27897
rect 13126 27897 13138 27900
rect 13172 27928 13184 27931
rect 14090 27928 14096 27940
rect 13172 27900 14096 27928
rect 13172 27897 13184 27900
rect 13126 27891 13184 27897
rect 14090 27888 14096 27900
rect 14148 27888 14154 27940
rect 15473 27931 15531 27937
rect 15473 27897 15485 27931
rect 15519 27897 15531 27931
rect 15473 27891 15531 27897
rect 15565 27931 15623 27937
rect 15565 27897 15577 27931
rect 15611 27928 15623 27931
rect 15654 27928 15660 27940
rect 15611 27900 15660 27928
rect 15611 27897 15623 27900
rect 15565 27891 15623 27897
rect 12894 27860 12900 27872
rect 10980 27832 12900 27860
rect 12894 27820 12900 27832
rect 12952 27820 12958 27872
rect 14918 27860 14924 27872
rect 14879 27832 14924 27860
rect 14918 27820 14924 27832
rect 14976 27820 14982 27872
rect 15488 27860 15516 27891
rect 15654 27888 15660 27900
rect 15712 27888 15718 27940
rect 17862 27888 17868 27940
rect 17920 27928 17926 27940
rect 19889 27931 19947 27937
rect 19889 27928 19901 27931
rect 17920 27900 19901 27928
rect 17920 27888 17926 27900
rect 19889 27897 19901 27900
rect 19935 27928 19947 27931
rect 20088 27928 20116 27959
rect 19935 27900 20116 27928
rect 19935 27897 19947 27900
rect 19889 27891 19947 27897
rect 20346 27888 20352 27940
rect 20404 27928 20410 27940
rect 20640 27928 20668 27959
rect 21082 27956 21088 27968
rect 21140 27956 21146 28008
rect 23820 27999 23878 28005
rect 23820 27965 23832 27999
rect 23866 27996 23878 27999
rect 25038 27996 25044 28008
rect 23866 27968 24348 27996
rect 24999 27968 25044 27996
rect 23866 27965 23878 27968
rect 23820 27959 23878 27965
rect 21450 27928 21456 27940
rect 20404 27900 21456 27928
rect 20404 27888 20410 27900
rect 21450 27888 21456 27900
rect 21508 27888 21514 27940
rect 21818 27928 21824 27940
rect 21779 27900 21824 27928
rect 21818 27888 21824 27900
rect 21876 27888 21882 27940
rect 21910 27888 21916 27940
rect 21968 27928 21974 27940
rect 21968 27900 22013 27928
rect 21968 27888 21974 27900
rect 16022 27860 16028 27872
rect 15488 27832 16028 27860
rect 16022 27820 16028 27832
rect 16080 27820 16086 27872
rect 18966 27820 18972 27872
rect 19024 27860 19030 27872
rect 19245 27863 19303 27869
rect 19245 27860 19257 27863
rect 19024 27832 19257 27860
rect 19024 27820 19030 27832
rect 19245 27829 19257 27832
rect 19291 27829 19303 27863
rect 19245 27823 19303 27829
rect 23891 27863 23949 27869
rect 23891 27829 23903 27863
rect 23937 27860 23949 27863
rect 24118 27860 24124 27872
rect 23937 27832 24124 27860
rect 23937 27829 23949 27832
rect 23891 27823 23949 27829
rect 24118 27820 24124 27832
rect 24176 27820 24182 27872
rect 24320 27869 24348 27968
rect 25038 27956 25044 27968
rect 25096 27956 25102 28008
rect 25332 28005 25360 28104
rect 25406 28092 25412 28104
rect 25464 28132 25470 28144
rect 25869 28135 25927 28141
rect 25869 28132 25881 28135
rect 25464 28104 25881 28132
rect 25464 28092 25470 28104
rect 25869 28101 25881 28104
rect 25915 28132 25927 28135
rect 29454 28132 29460 28144
rect 25915 28104 29460 28132
rect 25915 28101 25927 28104
rect 25869 28095 25927 28101
rect 29454 28092 29460 28104
rect 29512 28092 29518 28144
rect 34606 28132 34612 28144
rect 34567 28104 34612 28132
rect 34606 28092 34612 28104
rect 34664 28092 34670 28144
rect 35437 28135 35495 28141
rect 35437 28101 35449 28135
rect 35483 28132 35495 28135
rect 35802 28132 35808 28144
rect 35483 28104 35808 28132
rect 35483 28101 35495 28104
rect 35437 28095 35495 28101
rect 25498 28064 25504 28076
rect 25459 28036 25504 28064
rect 25498 28024 25504 28036
rect 25556 28024 25562 28076
rect 28902 28024 28908 28076
rect 28960 28064 28966 28076
rect 29641 28067 29699 28073
rect 29641 28064 29653 28067
rect 28960 28036 29653 28064
rect 28960 28024 28966 28036
rect 29641 28033 29653 28036
rect 29687 28064 29699 28067
rect 30466 28064 30472 28076
rect 29687 28036 30472 28064
rect 29687 28033 29699 28036
rect 29641 28027 29699 28033
rect 30466 28024 30472 28036
rect 30524 28024 30530 28076
rect 25317 27999 25375 28005
rect 25317 27965 25329 27999
rect 25363 27965 25375 27999
rect 25317 27959 25375 27965
rect 26513 27999 26571 28005
rect 26513 27965 26525 27999
rect 26559 27996 26571 27999
rect 26640 27999 26698 28005
rect 26640 27996 26652 27999
rect 26559 27968 26652 27996
rect 26559 27965 26571 27968
rect 26513 27959 26571 27965
rect 26640 27965 26652 27968
rect 26686 27996 26698 27999
rect 27522 27996 27528 28008
rect 26686 27968 27528 27996
rect 26686 27965 26698 27968
rect 26640 27959 26698 27965
rect 27522 27956 27528 27968
rect 27580 27956 27586 28008
rect 27798 27996 27804 28008
rect 27759 27968 27804 27996
rect 27798 27956 27804 27968
rect 27856 27956 27862 28008
rect 28169 27999 28227 28005
rect 28169 27965 28181 27999
rect 28215 27996 28227 27999
rect 28258 27996 28264 28008
rect 28215 27968 28264 27996
rect 28215 27965 28227 27968
rect 28169 27959 28227 27965
rect 28258 27956 28264 27968
rect 28316 27956 28322 28008
rect 28353 27999 28411 28005
rect 28353 27965 28365 27999
rect 28399 27996 28411 27999
rect 32309 27999 32367 28005
rect 32309 27996 32321 27999
rect 28399 27968 32321 27996
rect 28399 27965 28411 27968
rect 28353 27959 28411 27965
rect 32309 27965 32321 27968
rect 32355 27996 32367 27999
rect 32490 27996 32496 28008
rect 32355 27968 32496 27996
rect 32355 27965 32367 27968
rect 32309 27959 32367 27965
rect 32490 27956 32496 27968
rect 32548 27956 32554 28008
rect 34146 27956 34152 28008
rect 34204 27996 34210 28008
rect 34952 27999 35010 28005
rect 34952 27996 34964 27999
rect 34204 27968 34964 27996
rect 34204 27956 34210 27968
rect 34952 27965 34964 27968
rect 34998 27996 35010 27999
rect 35452 27996 35480 28095
rect 35802 28092 35808 28104
rect 35860 28132 35866 28144
rect 38010 28132 38016 28144
rect 35860 28104 38016 28132
rect 35860 28092 35866 28104
rect 38010 28092 38016 28104
rect 38068 28092 38074 28144
rect 35710 28024 35716 28076
rect 35768 28064 35774 28076
rect 36265 28067 36323 28073
rect 36265 28064 36277 28067
rect 35768 28036 36277 28064
rect 35768 28024 35774 28036
rect 36265 28033 36277 28036
rect 36311 28064 36323 28067
rect 36630 28064 36636 28076
rect 36311 28036 36636 28064
rect 36311 28033 36323 28036
rect 36265 28027 36323 28033
rect 36630 28024 36636 28036
rect 36688 28024 36694 28076
rect 41877 28067 41935 28073
rect 41877 28033 41889 28067
rect 41923 28064 41935 28067
rect 41923 28036 42794 28064
rect 41923 28033 41935 28036
rect 41877 28027 41935 28033
rect 34998 27968 35480 27996
rect 37185 27999 37243 28005
rect 34998 27965 35010 27968
rect 34952 27959 35010 27965
rect 37185 27965 37197 27999
rect 37231 27996 37243 27999
rect 38286 27996 38292 28008
rect 37231 27968 38292 27996
rect 37231 27965 37243 27968
rect 37185 27959 37243 27965
rect 38286 27956 38292 27968
rect 38344 27956 38350 28008
rect 39276 27999 39334 28005
rect 39276 27965 39288 27999
rect 39322 27996 39334 27999
rect 39322 27968 39712 27996
rect 39322 27965 39334 27968
rect 39276 27959 39334 27965
rect 28276 27928 28304 27956
rect 28629 27931 28687 27937
rect 28629 27928 28641 27931
rect 28276 27900 28641 27928
rect 28629 27897 28641 27900
rect 28675 27897 28687 27931
rect 28629 27891 28687 27897
rect 29089 27931 29147 27937
rect 29089 27897 29101 27931
rect 29135 27928 29147 27931
rect 29549 27931 29607 27937
rect 29549 27928 29561 27931
rect 29135 27900 29561 27928
rect 29135 27897 29147 27900
rect 29089 27891 29147 27897
rect 29549 27897 29561 27900
rect 29595 27928 29607 27931
rect 29730 27928 29736 27940
rect 29595 27900 29736 27928
rect 29595 27897 29607 27900
rect 29549 27891 29607 27897
rect 29730 27888 29736 27900
rect 29788 27928 29794 27940
rect 30003 27931 30061 27937
rect 30003 27928 30015 27931
rect 29788 27900 30015 27928
rect 29788 27888 29794 27900
rect 30003 27897 30015 27900
rect 30049 27928 30061 27931
rect 31110 27928 31116 27940
rect 30049 27900 31116 27928
rect 30049 27897 30061 27900
rect 30003 27891 30061 27897
rect 31110 27888 31116 27900
rect 31168 27928 31174 27940
rect 32217 27931 32275 27937
rect 32217 27928 32229 27931
rect 31168 27900 32229 27928
rect 31168 27888 31174 27900
rect 32217 27897 32229 27900
rect 32263 27928 32275 27931
rect 32671 27931 32729 27937
rect 32671 27928 32683 27931
rect 32263 27900 32683 27928
rect 32263 27897 32275 27900
rect 32217 27891 32275 27897
rect 32671 27897 32683 27900
rect 32717 27928 32729 27931
rect 36586 27931 36644 27937
rect 36586 27928 36598 27931
rect 32717 27900 36598 27928
rect 32717 27897 32729 27900
rect 32671 27891 32729 27897
rect 36188 27872 36216 27900
rect 36586 27897 36598 27900
rect 36632 27928 36644 27931
rect 38470 27928 38476 27940
rect 36632 27900 38476 27928
rect 36632 27897 36644 27900
rect 36586 27891 36644 27897
rect 38470 27888 38476 27900
rect 38528 27888 38534 27940
rect 39684 27872 39712 27968
rect 40402 27956 40408 28008
rect 40460 27996 40466 28008
rect 40532 27999 40590 28005
rect 40532 27996 40544 27999
rect 40460 27968 40544 27996
rect 40460 27956 40466 27968
rect 40532 27965 40544 27968
rect 40578 27996 40590 27999
rect 40957 27999 41015 28005
rect 40957 27996 40969 27999
rect 40578 27968 40969 27996
rect 40578 27965 40590 27968
rect 40532 27959 40590 27965
rect 40957 27965 40969 27968
rect 41003 27996 41015 27999
rect 41046 27996 41052 28008
rect 41003 27968 41052 27996
rect 41003 27965 41015 27968
rect 40957 27959 41015 27965
rect 41046 27956 41052 27968
rect 41104 27956 41110 28008
rect 39758 27888 39764 27940
rect 39816 27928 39822 27940
rect 40635 27931 40693 27937
rect 40635 27928 40647 27931
rect 39816 27900 40647 27928
rect 39816 27888 39822 27900
rect 40635 27897 40647 27900
rect 40681 27897 40693 27931
rect 41969 27931 42027 27937
rect 41969 27928 41981 27931
rect 40635 27891 40693 27897
rect 41616 27900 41981 27928
rect 24305 27863 24363 27869
rect 24305 27829 24317 27863
rect 24351 27860 24363 27863
rect 25590 27860 25596 27872
rect 24351 27832 25596 27860
rect 24351 27829 24363 27832
rect 24305 27823 24363 27829
rect 25590 27820 25596 27832
rect 25648 27860 25654 27872
rect 28350 27860 28356 27872
rect 25648 27832 28356 27860
rect 25648 27820 25654 27832
rect 28350 27820 28356 27832
rect 28408 27820 28414 27872
rect 30561 27863 30619 27869
rect 30561 27829 30573 27863
rect 30607 27860 30619 27863
rect 30926 27860 30932 27872
rect 30607 27832 30932 27860
rect 30607 27829 30619 27832
rect 30561 27823 30619 27829
rect 30926 27820 30932 27832
rect 30984 27820 30990 27872
rect 31018 27820 31024 27872
rect 31076 27860 31082 27872
rect 33229 27863 33287 27869
rect 31076 27832 31121 27860
rect 31076 27820 31082 27832
rect 33229 27829 33241 27863
rect 33275 27860 33287 27863
rect 33410 27860 33416 27872
rect 33275 27832 33416 27860
rect 33275 27829 33287 27832
rect 33229 27823 33287 27829
rect 33410 27820 33416 27832
rect 33468 27860 33474 27872
rect 33597 27863 33655 27869
rect 33597 27860 33609 27863
rect 33468 27832 33609 27860
rect 33468 27820 33474 27832
rect 33597 27829 33609 27832
rect 33643 27860 33655 27863
rect 33778 27860 33784 27872
rect 33643 27832 33784 27860
rect 33643 27829 33655 27832
rect 33597 27823 33655 27829
rect 33778 27820 33784 27832
rect 33836 27820 33842 27872
rect 36170 27860 36176 27872
rect 36131 27832 36176 27860
rect 36170 27820 36176 27832
rect 36228 27820 36234 27872
rect 38010 27860 38016 27872
rect 37971 27832 38016 27860
rect 38010 27820 38016 27832
rect 38068 27820 38074 27872
rect 39347 27863 39405 27869
rect 39347 27829 39359 27863
rect 39393 27860 39405 27863
rect 39574 27860 39580 27872
rect 39393 27832 39580 27860
rect 39393 27829 39405 27832
rect 39347 27823 39405 27829
rect 39574 27820 39580 27832
rect 39632 27820 39638 27872
rect 39666 27820 39672 27872
rect 39724 27860 39730 27872
rect 39724 27832 39769 27860
rect 39724 27820 39730 27832
rect 41506 27820 41512 27872
rect 41564 27860 41570 27872
rect 41616 27869 41644 27900
rect 41969 27897 41981 27900
rect 42015 27897 42027 27931
rect 42518 27928 42524 27940
rect 42479 27900 42524 27928
rect 41969 27891 42027 27897
rect 42518 27888 42524 27900
rect 42576 27888 42582 27940
rect 42766 27928 42794 28036
rect 43400 27999 43458 28005
rect 43400 27965 43412 27999
rect 43446 27996 43458 27999
rect 43446 27968 43944 27996
rect 43446 27965 43458 27968
rect 43400 27959 43458 27965
rect 43257 27931 43315 27937
rect 43257 27928 43269 27931
rect 42766 27900 43269 27928
rect 43257 27897 43269 27900
rect 43303 27928 43315 27931
rect 43487 27931 43545 27937
rect 43487 27928 43499 27931
rect 43303 27900 43499 27928
rect 43303 27897 43315 27900
rect 43257 27891 43315 27897
rect 43487 27897 43499 27900
rect 43533 27897 43545 27931
rect 43487 27891 43545 27897
rect 43916 27869 43944 27968
rect 41601 27863 41659 27869
rect 41601 27860 41613 27863
rect 41564 27832 41613 27860
rect 41564 27820 41570 27832
rect 41601 27829 41613 27832
rect 41647 27829 41659 27863
rect 41601 27823 41659 27829
rect 43901 27863 43959 27869
rect 43901 27829 43913 27863
rect 43947 27860 43959 27863
rect 44818 27860 44824 27872
rect 43947 27832 44824 27860
rect 43947 27829 43959 27832
rect 43901 27823 43959 27829
rect 44818 27820 44824 27832
rect 44876 27820 44882 27872
rect 1104 27770 48852 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 48852 27770
rect 1104 27696 48852 27718
rect 4614 27616 4620 27668
rect 4672 27656 4678 27668
rect 4985 27659 5043 27665
rect 4985 27656 4997 27659
rect 4672 27628 4997 27656
rect 4672 27616 4678 27628
rect 4985 27625 4997 27628
rect 5031 27625 5043 27659
rect 4985 27619 5043 27625
rect 6454 27616 6460 27668
rect 6512 27656 6518 27668
rect 6917 27659 6975 27665
rect 6917 27656 6929 27659
rect 6512 27628 6929 27656
rect 6512 27616 6518 27628
rect 6917 27625 6929 27628
rect 6963 27625 6975 27659
rect 9766 27656 9772 27668
rect 9727 27628 9772 27656
rect 6917 27619 6975 27625
rect 9766 27616 9772 27628
rect 9824 27616 9830 27668
rect 10870 27656 10876 27668
rect 10831 27628 10876 27656
rect 10870 27616 10876 27628
rect 10928 27616 10934 27668
rect 15286 27616 15292 27668
rect 15344 27656 15350 27668
rect 15344 27628 15424 27656
rect 15344 27616 15350 27628
rect 3970 27548 3976 27600
rect 4028 27588 4034 27600
rect 4427 27591 4485 27597
rect 4427 27588 4439 27591
rect 4028 27560 4439 27588
rect 4028 27548 4034 27560
rect 4427 27557 4439 27560
rect 4473 27588 4485 27591
rect 4798 27588 4804 27600
rect 4473 27560 4804 27588
rect 4473 27557 4485 27560
rect 4427 27551 4485 27557
rect 4798 27548 4804 27560
rect 4856 27548 4862 27600
rect 7834 27548 7840 27600
rect 7892 27588 7898 27600
rect 8113 27591 8171 27597
rect 8113 27588 8125 27591
rect 7892 27560 8125 27588
rect 7892 27548 7898 27560
rect 8113 27557 8125 27560
rect 8159 27557 8171 27591
rect 8113 27551 8171 27557
rect 8205 27591 8263 27597
rect 8205 27557 8217 27591
rect 8251 27588 8263 27591
rect 8478 27588 8484 27600
rect 8251 27560 8484 27588
rect 8251 27557 8263 27560
rect 8205 27551 8263 27557
rect 8478 27548 8484 27560
rect 8536 27548 8542 27600
rect 8754 27588 8760 27600
rect 8715 27560 8760 27588
rect 8754 27548 8760 27560
rect 8812 27548 8818 27600
rect 12802 27548 12808 27600
rect 12860 27588 12866 27600
rect 15396 27597 15424 27628
rect 16574 27616 16580 27668
rect 16632 27656 16638 27668
rect 16669 27659 16727 27665
rect 16669 27656 16681 27659
rect 16632 27628 16681 27656
rect 16632 27616 16638 27628
rect 16669 27625 16681 27628
rect 16715 27625 16727 27659
rect 18230 27656 18236 27668
rect 18191 27628 18236 27656
rect 16669 27619 16727 27625
rect 18230 27616 18236 27628
rect 18288 27616 18294 27668
rect 19334 27656 19340 27668
rect 19295 27628 19340 27656
rect 19334 27616 19340 27628
rect 19392 27616 19398 27668
rect 20346 27656 20352 27668
rect 20307 27628 20352 27656
rect 20346 27616 20352 27628
rect 20404 27616 20410 27668
rect 21174 27616 21180 27668
rect 21232 27656 21238 27668
rect 21269 27659 21327 27665
rect 21269 27656 21281 27659
rect 21232 27628 21281 27656
rect 21232 27616 21238 27628
rect 21269 27625 21281 27628
rect 21315 27625 21327 27659
rect 21269 27619 21327 27625
rect 21821 27659 21879 27665
rect 21821 27625 21833 27659
rect 21867 27656 21879 27659
rect 21910 27656 21916 27668
rect 21867 27628 21916 27656
rect 21867 27625 21879 27628
rect 21821 27619 21879 27625
rect 21910 27616 21916 27628
rect 21968 27656 21974 27668
rect 22097 27659 22155 27665
rect 22097 27656 22109 27659
rect 21968 27628 22109 27656
rect 21968 27616 21974 27628
rect 22097 27625 22109 27628
rect 22143 27625 22155 27659
rect 22097 27619 22155 27625
rect 23198 27616 23204 27668
rect 23256 27656 23262 27668
rect 23658 27656 23664 27668
rect 23256 27628 23664 27656
rect 23256 27616 23262 27628
rect 23658 27616 23664 27628
rect 23716 27616 23722 27668
rect 25038 27656 25044 27668
rect 24999 27628 25044 27656
rect 25038 27616 25044 27628
rect 25096 27616 25102 27668
rect 25406 27656 25412 27668
rect 25367 27628 25412 27656
rect 25406 27616 25412 27628
rect 25464 27616 25470 27668
rect 27614 27616 27620 27668
rect 27672 27656 27678 27668
rect 27709 27659 27767 27665
rect 27709 27656 27721 27659
rect 27672 27628 27721 27656
rect 27672 27616 27678 27628
rect 27709 27625 27721 27628
rect 27755 27656 27767 27659
rect 27798 27656 27804 27668
rect 27755 27628 27804 27656
rect 27755 27625 27767 27628
rect 27709 27619 27767 27625
rect 27798 27616 27804 27628
rect 27856 27616 27862 27668
rect 29178 27656 29184 27668
rect 29139 27628 29184 27656
rect 29178 27616 29184 27628
rect 29236 27616 29242 27668
rect 29730 27656 29736 27668
rect 29691 27628 29736 27656
rect 29730 27616 29736 27628
rect 29788 27616 29794 27668
rect 35986 27616 35992 27668
rect 36044 27656 36050 27668
rect 36265 27659 36323 27665
rect 36265 27656 36277 27659
rect 36044 27628 36277 27656
rect 36044 27616 36050 27628
rect 36265 27625 36277 27628
rect 36311 27625 36323 27659
rect 36630 27656 36636 27668
rect 36591 27628 36636 27656
rect 36265 27619 36323 27625
rect 36630 27616 36636 27628
rect 36688 27616 36694 27668
rect 39206 27656 39212 27668
rect 37746 27628 39212 27656
rect 12897 27591 12955 27597
rect 12897 27588 12909 27591
rect 12860 27560 12909 27588
rect 12860 27548 12866 27560
rect 12897 27557 12909 27560
rect 12943 27588 12955 27591
rect 13173 27591 13231 27597
rect 13173 27588 13185 27591
rect 12943 27560 13185 27588
rect 12943 27557 12955 27560
rect 12897 27551 12955 27557
rect 13173 27557 13185 27560
rect 13219 27557 13231 27591
rect 13173 27551 13231 27557
rect 15381 27591 15439 27597
rect 15381 27557 15393 27591
rect 15427 27557 15439 27591
rect 15381 27551 15439 27557
rect 15470 27548 15476 27600
rect 15528 27588 15534 27600
rect 17034 27588 17040 27600
rect 15528 27560 15573 27588
rect 16995 27560 17040 27588
rect 15528 27548 15534 27560
rect 17034 27548 17040 27560
rect 17092 27548 17098 27600
rect 17586 27588 17592 27600
rect 17547 27560 17592 27588
rect 17586 27548 17592 27560
rect 17644 27548 17650 27600
rect 24121 27591 24179 27597
rect 24121 27557 24133 27591
rect 24167 27588 24179 27591
rect 24486 27588 24492 27600
rect 24167 27560 24492 27588
rect 24167 27557 24179 27560
rect 24121 27551 24179 27557
rect 24486 27548 24492 27560
rect 24544 27548 24550 27600
rect 32306 27588 32312 27600
rect 32267 27560 32312 27588
rect 32306 27548 32312 27560
rect 32364 27548 32370 27600
rect 33778 27548 33784 27600
rect 33836 27588 33842 27600
rect 33873 27591 33931 27597
rect 33873 27588 33885 27591
rect 33836 27560 33885 27588
rect 33836 27548 33842 27560
rect 33873 27557 33885 27560
rect 33919 27557 33931 27591
rect 33873 27551 33931 27557
rect 4062 27520 4068 27532
rect 4023 27492 4068 27520
rect 4062 27480 4068 27492
rect 4120 27480 4126 27532
rect 5626 27480 5632 27532
rect 5684 27520 5690 27532
rect 5905 27523 5963 27529
rect 5905 27520 5917 27523
rect 5684 27492 5917 27520
rect 5684 27480 5690 27492
rect 5905 27489 5917 27492
rect 5951 27489 5963 27523
rect 5905 27483 5963 27489
rect 6362 27480 6368 27532
rect 6420 27520 6426 27532
rect 6457 27523 6515 27529
rect 6457 27520 6469 27523
rect 6420 27492 6469 27520
rect 6420 27480 6426 27492
rect 6457 27489 6469 27492
rect 6503 27520 6515 27523
rect 7006 27520 7012 27532
rect 6503 27492 7012 27520
rect 6503 27489 6515 27492
rect 6457 27483 6515 27489
rect 7006 27480 7012 27492
rect 7064 27480 7070 27532
rect 9858 27520 9864 27532
rect 9819 27492 9864 27520
rect 9858 27480 9864 27492
rect 9916 27480 9922 27532
rect 10137 27523 10195 27529
rect 10137 27489 10149 27523
rect 10183 27489 10195 27523
rect 12250 27520 12256 27532
rect 12211 27492 12256 27520
rect 10137 27483 10195 27489
rect 6641 27455 6699 27461
rect 6641 27421 6653 27455
rect 6687 27452 6699 27455
rect 6822 27452 6828 27464
rect 6687 27424 6828 27452
rect 6687 27421 6699 27424
rect 6641 27415 6699 27421
rect 6822 27412 6828 27424
rect 6880 27452 6886 27464
rect 7653 27455 7711 27461
rect 7653 27452 7665 27455
rect 6880 27424 7665 27452
rect 6880 27412 6886 27424
rect 7653 27421 7665 27424
rect 7699 27421 7711 27455
rect 7653 27415 7711 27421
rect 9582 27412 9588 27464
rect 9640 27452 9646 27464
rect 10152 27452 10180 27483
rect 12250 27480 12256 27492
rect 12308 27480 12314 27532
rect 12710 27520 12716 27532
rect 12671 27492 12716 27520
rect 12710 27480 12716 27492
rect 12768 27480 12774 27532
rect 13722 27520 13728 27532
rect 13683 27492 13728 27520
rect 13722 27480 13728 27492
rect 13780 27480 13786 27532
rect 18576 27523 18634 27529
rect 18576 27489 18588 27523
rect 18622 27520 18634 27523
rect 19058 27520 19064 27532
rect 18622 27492 19064 27520
rect 18622 27489 18634 27492
rect 18576 27483 18634 27489
rect 19058 27480 19064 27492
rect 19116 27480 19122 27532
rect 19797 27523 19855 27529
rect 19797 27489 19809 27523
rect 19843 27520 19855 27523
rect 19886 27520 19892 27532
rect 19843 27492 19892 27520
rect 19843 27489 19855 27492
rect 19797 27483 19855 27489
rect 19886 27480 19892 27492
rect 19944 27480 19950 27532
rect 26142 27480 26148 27532
rect 26200 27520 26206 27532
rect 26548 27523 26606 27529
rect 26548 27520 26560 27523
rect 26200 27492 26560 27520
rect 26200 27480 26206 27492
rect 26548 27489 26560 27492
rect 26594 27520 26606 27523
rect 27338 27520 27344 27532
rect 26594 27492 27344 27520
rect 26594 27489 26606 27492
rect 26548 27483 26606 27489
rect 27338 27480 27344 27492
rect 27396 27480 27402 27532
rect 27982 27520 27988 27532
rect 27943 27492 27988 27520
rect 27982 27480 27988 27492
rect 28040 27480 28046 27532
rect 28258 27520 28264 27532
rect 28219 27492 28264 27520
rect 28258 27480 28264 27492
rect 28316 27480 28322 27532
rect 35342 27520 35348 27532
rect 35303 27492 35348 27520
rect 35342 27480 35348 27492
rect 35400 27480 35406 27532
rect 35710 27480 35716 27532
rect 35768 27520 35774 27532
rect 35805 27523 35863 27529
rect 35805 27520 35817 27523
rect 35768 27492 35817 27520
rect 35768 27480 35774 27492
rect 35805 27489 35817 27492
rect 35851 27520 35863 27523
rect 37746 27520 37774 27628
rect 39206 27616 39212 27628
rect 39264 27616 39270 27668
rect 41601 27659 41659 27665
rect 41601 27625 41613 27659
rect 41647 27656 41659 27659
rect 41782 27656 41788 27668
rect 41647 27628 41788 27656
rect 41647 27625 41659 27628
rect 41601 27619 41659 27625
rect 41782 27616 41788 27628
rect 41840 27616 41846 27668
rect 38010 27548 38016 27600
rect 38068 27588 38074 27600
rect 38197 27591 38255 27597
rect 38197 27588 38209 27591
rect 38068 27560 38209 27588
rect 38068 27548 38074 27560
rect 38197 27557 38209 27560
rect 38243 27557 38255 27591
rect 38197 27551 38255 27557
rect 38286 27548 38292 27600
rect 38344 27588 38350 27600
rect 39758 27588 39764 27600
rect 38344 27560 38389 27588
rect 39719 27560 39764 27588
rect 38344 27548 38350 27560
rect 39758 27548 39764 27560
rect 39816 27548 39822 27600
rect 39850 27548 39856 27600
rect 39908 27588 39914 27600
rect 39908 27560 39953 27588
rect 39908 27548 39914 27560
rect 41506 27548 41512 27600
rect 41564 27588 41570 27600
rect 41877 27591 41935 27597
rect 41877 27588 41889 27591
rect 41564 27560 41889 27588
rect 41564 27548 41570 27560
rect 41877 27557 41889 27560
rect 41923 27557 41935 27591
rect 42426 27588 42432 27600
rect 42387 27560 42432 27588
rect 41877 27551 41935 27557
rect 42426 27548 42432 27560
rect 42484 27548 42490 27600
rect 35851 27492 37774 27520
rect 43416 27523 43474 27529
rect 35851 27489 35863 27492
rect 35805 27483 35863 27489
rect 43416 27489 43428 27523
rect 43462 27520 43474 27523
rect 43898 27520 43904 27532
rect 43462 27492 43904 27520
rect 43462 27489 43474 27492
rect 43416 27483 43474 27489
rect 43898 27480 43904 27492
rect 43956 27480 43962 27532
rect 16022 27452 16028 27464
rect 9640 27424 10180 27452
rect 15983 27424 16028 27452
rect 9640 27412 9646 27424
rect 16022 27412 16028 27424
rect 16080 27412 16086 27464
rect 16945 27455 17003 27461
rect 16945 27421 16957 27455
rect 16991 27421 17003 27455
rect 16945 27415 17003 27421
rect 20901 27455 20959 27461
rect 20901 27421 20913 27455
rect 20947 27452 20959 27455
rect 21082 27452 21088 27464
rect 20947 27424 21088 27452
rect 20947 27421 20959 27424
rect 20901 27415 20959 27421
rect 12802 27344 12808 27396
rect 12860 27384 12866 27396
rect 16850 27384 16856 27396
rect 12860 27356 16856 27384
rect 12860 27344 12866 27356
rect 16850 27344 16856 27356
rect 16908 27384 16914 27396
rect 16960 27384 16988 27415
rect 21082 27412 21088 27424
rect 21140 27412 21146 27464
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27452 22983 27455
rect 24026 27452 24032 27464
rect 22971 27424 24032 27452
rect 22971 27421 22983 27424
rect 22925 27415 22983 27421
rect 24026 27412 24032 27424
rect 24084 27412 24090 27464
rect 24302 27452 24308 27464
rect 24263 27424 24308 27452
rect 24302 27412 24308 27424
rect 24360 27412 24366 27464
rect 28537 27455 28595 27461
rect 28537 27421 28549 27455
rect 28583 27452 28595 27455
rect 28994 27452 29000 27464
rect 28583 27424 29000 27452
rect 28583 27421 28595 27424
rect 28537 27415 28595 27421
rect 28994 27412 29000 27424
rect 29052 27452 29058 27464
rect 29365 27455 29423 27461
rect 29365 27452 29377 27455
rect 29052 27424 29377 27452
rect 29052 27412 29058 27424
rect 29365 27421 29377 27424
rect 29411 27421 29423 27455
rect 32214 27452 32220 27464
rect 32175 27424 32220 27452
rect 29365 27415 29423 27421
rect 32214 27412 32220 27424
rect 32272 27412 32278 27464
rect 32493 27455 32551 27461
rect 32493 27421 32505 27455
rect 32539 27421 32551 27455
rect 32493 27415 32551 27421
rect 16908 27356 16988 27384
rect 19935 27387 19993 27393
rect 16908 27344 16914 27356
rect 19935 27353 19947 27387
rect 19981 27384 19993 27387
rect 24394 27384 24400 27396
rect 19981 27356 24400 27384
rect 19981 27353 19993 27356
rect 19935 27347 19993 27353
rect 24394 27344 24400 27356
rect 24452 27344 24458 27396
rect 25958 27344 25964 27396
rect 26016 27384 26022 27396
rect 31018 27384 31024 27396
rect 26016 27356 31024 27384
rect 26016 27344 26022 27356
rect 31018 27344 31024 27356
rect 31076 27344 31082 27396
rect 31110 27344 31116 27396
rect 31168 27384 31174 27396
rect 32508 27384 32536 27415
rect 33410 27412 33416 27464
rect 33468 27452 33474 27464
rect 33781 27455 33839 27461
rect 33781 27452 33793 27455
rect 33468 27424 33793 27452
rect 33468 27412 33474 27424
rect 33781 27421 33793 27424
rect 33827 27421 33839 27455
rect 34422 27452 34428 27464
rect 34383 27424 34428 27452
rect 33781 27415 33839 27421
rect 34422 27412 34428 27424
rect 34480 27412 34486 27464
rect 35894 27452 35900 27464
rect 35855 27424 35900 27452
rect 35894 27412 35900 27424
rect 35952 27412 35958 27464
rect 38562 27452 38568 27464
rect 38523 27424 38568 27452
rect 38562 27412 38568 27424
rect 38620 27412 38626 27464
rect 40034 27452 40040 27464
rect 39995 27424 40040 27452
rect 40034 27412 40040 27424
rect 40092 27412 40098 27464
rect 41785 27455 41843 27461
rect 41785 27421 41797 27455
rect 41831 27452 41843 27455
rect 41831 27424 42794 27452
rect 41831 27421 41843 27424
rect 41785 27415 41843 27421
rect 32766 27384 32772 27396
rect 31168 27356 32772 27384
rect 31168 27344 31174 27356
rect 32766 27344 32772 27356
rect 32824 27344 32830 27396
rect 40770 27384 40776 27396
rect 40683 27356 40776 27384
rect 40770 27344 40776 27356
rect 40828 27384 40834 27396
rect 42426 27384 42432 27396
rect 40828 27356 42432 27384
rect 40828 27344 40834 27356
rect 42426 27344 42432 27356
rect 42484 27344 42490 27396
rect 3605 27319 3663 27325
rect 3605 27285 3617 27319
rect 3651 27316 3663 27319
rect 3970 27316 3976 27328
rect 3651 27288 3976 27316
rect 3651 27285 3663 27288
rect 3605 27279 3663 27285
rect 3970 27276 3976 27288
rect 4028 27276 4034 27328
rect 7377 27319 7435 27325
rect 7377 27285 7389 27319
rect 7423 27316 7435 27319
rect 7558 27316 7564 27328
rect 7423 27288 7564 27316
rect 7423 27285 7435 27288
rect 7377 27279 7435 27285
rect 7558 27276 7564 27288
rect 7616 27276 7622 27328
rect 12710 27276 12716 27328
rect 12768 27316 12774 27328
rect 13446 27316 13452 27328
rect 12768 27288 13452 27316
rect 12768 27276 12774 27288
rect 13446 27276 13452 27288
rect 13504 27316 13510 27328
rect 13909 27319 13967 27325
rect 13909 27316 13921 27319
rect 13504 27288 13921 27316
rect 13504 27276 13510 27288
rect 13909 27285 13921 27288
rect 13955 27285 13967 27319
rect 14182 27316 14188 27328
rect 14143 27288 14188 27316
rect 13909 27279 13967 27285
rect 14182 27276 14188 27288
rect 14240 27276 14246 27328
rect 17954 27276 17960 27328
rect 18012 27316 18018 27328
rect 18647 27319 18705 27325
rect 18647 27316 18659 27319
rect 18012 27288 18659 27316
rect 18012 27276 18018 27288
rect 18647 27285 18659 27288
rect 18693 27285 18705 27319
rect 18647 27279 18705 27285
rect 21910 27276 21916 27328
rect 21968 27316 21974 27328
rect 22465 27319 22523 27325
rect 22465 27316 22477 27319
rect 21968 27288 22477 27316
rect 21968 27276 21974 27288
rect 22465 27285 22477 27288
rect 22511 27285 22523 27319
rect 22465 27279 22523 27285
rect 25590 27276 25596 27328
rect 25648 27316 25654 27328
rect 26651 27319 26709 27325
rect 26651 27316 26663 27319
rect 25648 27288 26663 27316
rect 25648 27276 25654 27288
rect 26651 27285 26663 27288
rect 26697 27285 26709 27319
rect 26651 27279 26709 27285
rect 30285 27319 30343 27325
rect 30285 27285 30297 27319
rect 30331 27316 30343 27319
rect 30558 27316 30564 27328
rect 30331 27288 30564 27316
rect 30331 27285 30343 27288
rect 30285 27279 30343 27285
rect 30558 27276 30564 27288
rect 30616 27276 30622 27328
rect 30834 27316 30840 27328
rect 30795 27288 30840 27316
rect 30834 27276 30840 27288
rect 30892 27276 30898 27328
rect 32674 27276 32680 27328
rect 32732 27316 32738 27328
rect 34422 27316 34428 27328
rect 32732 27288 34428 27316
rect 32732 27276 32738 27288
rect 34422 27276 34428 27288
rect 34480 27276 34486 27328
rect 35986 27276 35992 27328
rect 36044 27316 36050 27328
rect 37826 27316 37832 27328
rect 36044 27288 37832 27316
rect 36044 27276 36050 27288
rect 37826 27276 37832 27288
rect 37884 27276 37890 27328
rect 38654 27276 38660 27328
rect 38712 27316 38718 27328
rect 39117 27319 39175 27325
rect 39117 27316 39129 27319
rect 38712 27288 39129 27316
rect 38712 27276 38718 27288
rect 39117 27285 39129 27288
rect 39163 27285 39175 27319
rect 42766 27316 42794 27424
rect 43162 27316 43168 27328
rect 42766 27288 43168 27316
rect 39117 27279 39175 27285
rect 43162 27276 43168 27288
rect 43220 27316 43226 27328
rect 43487 27319 43545 27325
rect 43487 27316 43499 27319
rect 43220 27288 43499 27316
rect 43220 27276 43226 27288
rect 43487 27285 43499 27288
rect 43533 27285 43545 27319
rect 43487 27279 43545 27285
rect 1104 27226 48852 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 48852 27226
rect 1104 27152 48852 27174
rect 5166 27112 5172 27124
rect 5127 27084 5172 27112
rect 5166 27072 5172 27084
rect 5224 27072 5230 27124
rect 5629 27115 5687 27121
rect 5629 27081 5641 27115
rect 5675 27112 5687 27115
rect 7006 27112 7012 27124
rect 5675 27084 7012 27112
rect 5675 27081 5687 27084
rect 5629 27075 5687 27081
rect 7006 27072 7012 27084
rect 7064 27072 7070 27124
rect 7650 27072 7656 27124
rect 7708 27112 7714 27124
rect 7745 27115 7803 27121
rect 7745 27112 7757 27115
rect 7708 27084 7757 27112
rect 7708 27072 7714 27084
rect 7745 27081 7757 27084
rect 7791 27081 7803 27115
rect 7745 27075 7803 27081
rect 7834 27072 7840 27124
rect 7892 27112 7898 27124
rect 8389 27115 8447 27121
rect 8389 27112 8401 27115
rect 7892 27084 8401 27112
rect 7892 27072 7898 27084
rect 8389 27081 8401 27084
rect 8435 27081 8447 27115
rect 10778 27112 10784 27124
rect 10739 27084 10784 27112
rect 8389 27075 8447 27081
rect 10778 27072 10784 27084
rect 10836 27072 10842 27124
rect 12158 27112 12164 27124
rect 12119 27084 12164 27112
rect 12158 27072 12164 27084
rect 12216 27112 12222 27124
rect 12618 27112 12624 27124
rect 12216 27084 12624 27112
rect 12216 27072 12222 27084
rect 12618 27072 12624 27084
rect 12676 27072 12682 27124
rect 14090 27112 14096 27124
rect 14051 27084 14096 27112
rect 14090 27072 14096 27084
rect 14148 27072 14154 27124
rect 15286 27072 15292 27124
rect 15344 27112 15350 27124
rect 15749 27115 15807 27121
rect 15749 27112 15761 27115
rect 15344 27084 15761 27112
rect 15344 27072 15350 27084
rect 15749 27081 15761 27084
rect 15795 27081 15807 27115
rect 15749 27075 15807 27081
rect 17034 27072 17040 27124
rect 17092 27112 17098 27124
rect 17405 27115 17463 27121
rect 17405 27112 17417 27115
rect 17092 27084 17417 27112
rect 17092 27072 17098 27084
rect 17405 27081 17417 27084
rect 17451 27081 17463 27115
rect 19058 27112 19064 27124
rect 19019 27084 19064 27112
rect 17405 27075 17463 27081
rect 19058 27072 19064 27084
rect 19116 27072 19122 27124
rect 24486 27072 24492 27124
rect 24544 27112 24550 27124
rect 24581 27115 24639 27121
rect 24581 27112 24593 27115
rect 24544 27084 24593 27112
rect 24544 27072 24550 27084
rect 24581 27081 24593 27084
rect 24627 27081 24639 27115
rect 24581 27075 24639 27081
rect 26970 27072 26976 27124
rect 27028 27112 27034 27124
rect 27801 27115 27859 27121
rect 27801 27112 27813 27115
rect 27028 27084 27813 27112
rect 27028 27072 27034 27084
rect 27801 27081 27813 27084
rect 27847 27112 27859 27115
rect 27982 27112 27988 27124
rect 27847 27084 27988 27112
rect 27847 27081 27859 27084
rect 27801 27075 27859 27081
rect 27982 27072 27988 27084
rect 28040 27072 28046 27124
rect 28994 27112 29000 27124
rect 28955 27084 29000 27112
rect 28994 27072 29000 27084
rect 29052 27072 29058 27124
rect 29730 27112 29736 27124
rect 29691 27084 29736 27112
rect 29730 27072 29736 27084
rect 29788 27072 29794 27124
rect 30558 27112 30564 27124
rect 30519 27084 30564 27112
rect 30558 27072 30564 27084
rect 30616 27072 30622 27124
rect 30926 27072 30932 27124
rect 30984 27112 30990 27124
rect 32125 27115 32183 27121
rect 32125 27112 32137 27115
rect 30984 27084 32137 27112
rect 30984 27072 30990 27084
rect 32125 27081 32137 27084
rect 32171 27112 32183 27115
rect 32490 27112 32496 27124
rect 32171 27084 32496 27112
rect 32171 27081 32183 27084
rect 32125 27075 32183 27081
rect 32490 27072 32496 27084
rect 32548 27072 32554 27124
rect 33410 27112 33416 27124
rect 33371 27084 33416 27112
rect 33410 27072 33416 27084
rect 33468 27072 33474 27124
rect 36265 27115 36323 27121
rect 36265 27081 36277 27115
rect 36311 27112 36323 27115
rect 36446 27112 36452 27124
rect 36311 27084 36452 27112
rect 36311 27081 36323 27084
rect 36265 27075 36323 27081
rect 36446 27072 36452 27084
rect 36504 27112 36510 27124
rect 36504 27084 36768 27112
rect 36504 27072 36510 27084
rect 8113 27047 8171 27053
rect 8113 27013 8125 27047
rect 8159 27044 8171 27047
rect 8478 27044 8484 27056
rect 8159 27016 8484 27044
rect 8159 27013 8171 27016
rect 8113 27007 8171 27013
rect 8478 27004 8484 27016
rect 8536 27004 8542 27056
rect 9674 27004 9680 27056
rect 9732 27044 9738 27056
rect 16761 27047 16819 27053
rect 16761 27044 16773 27047
rect 9732 27016 16773 27044
rect 9732 27004 9738 27016
rect 16761 27013 16773 27016
rect 16807 27013 16819 27047
rect 16761 27007 16819 27013
rect 20441 27047 20499 27053
rect 20441 27013 20453 27047
rect 20487 27044 20499 27047
rect 23934 27044 23940 27056
rect 20487 27016 23940 27044
rect 20487 27013 20499 27016
rect 20441 27007 20499 27013
rect 3789 26979 3847 26985
rect 3789 26945 3801 26979
rect 3835 26976 3847 26979
rect 6822 26976 6828 26988
rect 3835 26948 4384 26976
rect 6783 26948 6828 26976
rect 3835 26945 3847 26948
rect 3789 26939 3847 26945
rect 3421 26911 3479 26917
rect 3421 26877 3433 26911
rect 3467 26908 3479 26911
rect 4246 26908 4252 26920
rect 3467 26880 4252 26908
rect 3467 26877 3479 26880
rect 3421 26871 3479 26877
rect 4246 26868 4252 26880
rect 4304 26868 4310 26920
rect 4157 26843 4215 26849
rect 4157 26809 4169 26843
rect 4203 26840 4215 26843
rect 4356 26840 4384 26948
rect 6822 26936 6828 26948
rect 6880 26936 6886 26988
rect 9766 26936 9772 26988
rect 9824 26976 9830 26988
rect 9861 26979 9919 26985
rect 9861 26976 9873 26979
rect 9824 26948 9873 26976
rect 9824 26936 9830 26948
rect 9861 26945 9873 26948
rect 9907 26976 9919 26979
rect 11425 26979 11483 26985
rect 11425 26976 11437 26979
rect 9907 26948 11437 26976
rect 9907 26945 9919 26948
rect 9861 26939 9919 26945
rect 11425 26945 11437 26948
rect 11471 26945 11483 26979
rect 11425 26939 11483 26945
rect 11974 26936 11980 26988
rect 12032 26976 12038 26988
rect 12802 26976 12808 26988
rect 12032 26948 12808 26976
rect 12032 26936 12038 26948
rect 12802 26936 12808 26948
rect 12860 26936 12866 26988
rect 14182 26976 14188 26988
rect 14143 26948 14188 26976
rect 14182 26936 14188 26948
rect 14240 26936 14246 26988
rect 15470 26976 15476 26988
rect 15431 26948 15476 26976
rect 15470 26936 15476 26948
rect 15528 26936 15534 26988
rect 7742 26868 7748 26920
rect 7800 26908 7806 26920
rect 8573 26911 8631 26917
rect 8573 26908 8585 26911
rect 7800 26880 8585 26908
rect 7800 26868 7806 26880
rect 8573 26877 8585 26880
rect 8619 26908 8631 26911
rect 9033 26911 9091 26917
rect 9033 26908 9045 26911
rect 8619 26880 9045 26908
rect 8619 26877 8631 26880
rect 8573 26871 8631 26877
rect 9033 26877 9045 26880
rect 9079 26877 9091 26911
rect 9033 26871 9091 26877
rect 9582 26868 9588 26920
rect 9640 26908 9646 26920
rect 11057 26911 11115 26917
rect 11057 26908 11069 26911
rect 9640 26880 11069 26908
rect 9640 26868 9646 26880
rect 11057 26877 11069 26880
rect 11103 26877 11115 26911
rect 11057 26871 11115 26877
rect 11885 26911 11943 26917
rect 11885 26877 11897 26911
rect 11931 26908 11943 26911
rect 12250 26908 12256 26920
rect 11931 26880 12256 26908
rect 11931 26877 11943 26880
rect 11885 26871 11943 26877
rect 12250 26868 12256 26880
rect 12308 26868 12314 26920
rect 15105 26911 15163 26917
rect 15105 26877 15117 26911
rect 15151 26908 15163 26911
rect 15968 26911 16026 26917
rect 15968 26908 15980 26911
rect 15151 26880 15980 26908
rect 15151 26877 15163 26880
rect 15105 26871 15163 26877
rect 15968 26877 15980 26880
rect 16014 26908 16026 26911
rect 16393 26911 16451 26917
rect 16393 26908 16405 26911
rect 16014 26880 16405 26908
rect 16014 26877 16026 26880
rect 15968 26871 16026 26877
rect 16393 26877 16405 26880
rect 16439 26877 16451 26911
rect 16776 26908 16804 27007
rect 17586 26936 17592 26988
rect 17644 26976 17650 26988
rect 18138 26976 18144 26988
rect 17644 26948 18144 26976
rect 17644 26936 17650 26948
rect 18138 26936 18144 26948
rect 18196 26936 18202 26988
rect 18414 26976 18420 26988
rect 18375 26948 18420 26976
rect 18414 26936 18420 26948
rect 18472 26936 18478 26988
rect 16980 26911 17038 26917
rect 16980 26908 16992 26911
rect 16776 26880 16992 26908
rect 16393 26871 16451 26877
rect 16980 26877 16992 26880
rect 17026 26908 17038 26911
rect 17954 26908 17960 26920
rect 17026 26880 17960 26908
rect 17026 26877 17038 26880
rect 16980 26871 17038 26877
rect 17954 26868 17960 26880
rect 18012 26868 18018 26920
rect 20615 26917 20643 27016
rect 23934 27004 23940 27016
rect 23992 27004 23998 27056
rect 24854 27004 24860 27056
rect 24912 27044 24918 27056
rect 29411 27047 29469 27053
rect 29411 27044 29423 27047
rect 24912 27016 29423 27044
rect 24912 27004 24918 27016
rect 29411 27013 29423 27016
rect 29457 27013 29469 27047
rect 29411 27007 29469 27013
rect 30190 27004 30196 27056
rect 30248 27044 30254 27056
rect 31757 27047 31815 27053
rect 31757 27044 31769 27047
rect 30248 27016 31769 27044
rect 30248 27004 30254 27016
rect 31757 27013 31769 27016
rect 31803 27044 31815 27047
rect 32306 27044 32312 27056
rect 31803 27016 32312 27044
rect 31803 27013 31815 27016
rect 31757 27007 31815 27013
rect 32306 27004 32312 27016
rect 32364 27004 32370 27056
rect 21542 26976 21548 26988
rect 21503 26948 21548 26976
rect 21542 26936 21548 26948
rect 21600 26936 21606 26988
rect 23658 26976 23664 26988
rect 23619 26948 23664 26976
rect 23658 26936 23664 26948
rect 23716 26936 23722 26988
rect 26878 26976 26884 26988
rect 26839 26948 26884 26976
rect 26878 26936 26884 26948
rect 26936 26936 26942 26988
rect 27338 26976 27344 26988
rect 27299 26948 27344 26976
rect 27338 26936 27344 26948
rect 27396 26936 27402 26988
rect 30834 26976 30840 26988
rect 30795 26948 30840 26976
rect 30834 26936 30840 26948
rect 30892 26936 30898 26988
rect 31110 26976 31116 26988
rect 31071 26948 31116 26976
rect 31110 26936 31116 26948
rect 31168 26936 31174 26988
rect 32401 26979 32459 26985
rect 32401 26945 32413 26979
rect 32447 26976 32459 26979
rect 32674 26976 32680 26988
rect 32447 26948 32680 26976
rect 32447 26945 32459 26948
rect 32401 26939 32459 26945
rect 32674 26936 32680 26948
rect 32732 26936 32738 26988
rect 32766 26936 32772 26988
rect 32824 26976 32830 26988
rect 36740 26985 36768 27084
rect 38010 27072 38016 27124
rect 38068 27112 38074 27124
rect 38105 27115 38163 27121
rect 38105 27112 38117 27115
rect 38068 27084 38117 27112
rect 38068 27072 38074 27084
rect 38105 27081 38117 27084
rect 38151 27081 38163 27115
rect 38105 27075 38163 27081
rect 39758 27072 39764 27124
rect 39816 27112 39822 27124
rect 40037 27115 40095 27121
rect 40037 27112 40049 27115
rect 39816 27084 40049 27112
rect 39816 27072 39822 27084
rect 40037 27081 40049 27084
rect 40083 27081 40095 27115
rect 43162 27112 43168 27124
rect 43123 27084 43168 27112
rect 40037 27075 40095 27081
rect 43162 27072 43168 27084
rect 43220 27072 43226 27124
rect 43809 27115 43867 27121
rect 43809 27081 43821 27115
rect 43855 27112 43867 27115
rect 43898 27112 43904 27124
rect 43855 27084 43904 27112
rect 43855 27081 43867 27084
rect 43809 27075 43867 27081
rect 43898 27072 43904 27084
rect 43956 27072 43962 27124
rect 38286 27004 38292 27056
rect 38344 27044 38350 27056
rect 41506 27044 41512 27056
rect 38344 27016 41512 27044
rect 38344 27004 38350 27016
rect 41506 27004 41512 27016
rect 41564 27004 41570 27056
rect 42334 27044 42340 27056
rect 42295 27016 42340 27044
rect 42334 27004 42340 27016
rect 42392 27004 42398 27056
rect 34333 26979 34391 26985
rect 32824 26948 32869 26976
rect 32824 26936 32830 26948
rect 34333 26945 34345 26979
rect 34379 26976 34391 26979
rect 36725 26979 36783 26985
rect 34379 26948 35756 26976
rect 34379 26945 34391 26948
rect 34333 26939 34391 26945
rect 35728 26920 35756 26948
rect 36725 26945 36737 26979
rect 36771 26945 36783 26979
rect 38562 26976 38568 26988
rect 38523 26948 38568 26976
rect 36725 26939 36783 26945
rect 38562 26936 38568 26948
rect 38620 26936 38626 26988
rect 40589 26979 40647 26985
rect 40589 26945 40601 26979
rect 40635 26976 40647 26979
rect 40635 26948 40908 26976
rect 40635 26945 40647 26948
rect 40589 26939 40647 26945
rect 40880 26920 40908 26948
rect 41598 26936 41604 26988
rect 41656 26976 41662 26988
rect 41785 26979 41843 26985
rect 41785 26976 41797 26979
rect 41656 26948 41797 26976
rect 41656 26936 41662 26948
rect 41785 26945 41797 26948
rect 41831 26976 41843 26979
rect 43395 26979 43453 26985
rect 43395 26976 43407 26979
rect 41831 26948 43407 26976
rect 41831 26945 41843 26948
rect 41785 26939 41843 26945
rect 43395 26945 43407 26948
rect 43441 26945 43453 26979
rect 43395 26939 43453 26945
rect 20600 26911 20658 26917
rect 20600 26877 20612 26911
rect 20646 26877 20658 26911
rect 26050 26908 26056 26920
rect 20600 26871 20658 26877
rect 21054 26880 26056 26908
rect 4611 26843 4669 26849
rect 4611 26840 4623 26843
rect 4203 26812 4623 26840
rect 4203 26809 4215 26812
rect 4157 26803 4215 26809
rect 4611 26809 4623 26812
rect 4657 26840 4669 26843
rect 4798 26840 4804 26852
rect 4657 26812 4804 26840
rect 4657 26809 4669 26812
rect 4611 26803 4669 26809
rect 4798 26800 4804 26812
rect 4856 26840 4862 26852
rect 5442 26840 5448 26852
rect 4856 26812 5448 26840
rect 4856 26800 4862 26812
rect 5442 26800 5448 26812
rect 5500 26840 5506 26852
rect 6641 26843 6699 26849
rect 6641 26840 6653 26843
rect 5500 26812 6653 26840
rect 5500 26800 5506 26812
rect 6641 26809 6653 26812
rect 6687 26840 6699 26843
rect 6914 26840 6920 26852
rect 6687 26812 6920 26840
rect 6687 26809 6699 26812
rect 6641 26803 6699 26809
rect 6914 26800 6920 26812
rect 6972 26840 6978 26852
rect 7187 26843 7245 26849
rect 7187 26840 7199 26843
rect 6972 26812 7199 26840
rect 6972 26800 6978 26812
rect 7187 26809 7199 26812
rect 7233 26840 7245 26843
rect 9769 26843 9827 26849
rect 9769 26840 9781 26843
rect 7233 26812 9781 26840
rect 7233 26809 7245 26812
rect 7187 26803 7245 26809
rect 9769 26809 9781 26812
rect 9815 26840 9827 26843
rect 10223 26843 10281 26849
rect 10223 26840 10235 26843
rect 9815 26812 10235 26840
rect 9815 26809 9827 26812
rect 9769 26803 9827 26809
rect 10223 26809 10235 26812
rect 10269 26840 10281 26843
rect 10594 26840 10600 26852
rect 10269 26812 10600 26840
rect 10269 26809 10281 26812
rect 10223 26803 10281 26809
rect 10594 26800 10600 26812
rect 10652 26800 10658 26852
rect 12526 26840 12532 26852
rect 12487 26812 12532 26840
rect 12526 26800 12532 26812
rect 12584 26800 12590 26852
rect 12618 26800 12624 26852
rect 12676 26840 12682 26852
rect 12676 26812 12721 26840
rect 12676 26800 12682 26812
rect 14090 26800 14096 26852
rect 14148 26840 14154 26852
rect 14506 26843 14564 26849
rect 14506 26840 14518 26843
rect 14148 26812 14518 26840
rect 14148 26800 14154 26812
rect 14506 26809 14518 26812
rect 14552 26809 14564 26843
rect 14506 26803 14564 26809
rect 18230 26800 18236 26852
rect 18288 26840 18294 26852
rect 19886 26840 19892 26852
rect 18288 26812 18333 26840
rect 19799 26812 19892 26840
rect 18288 26800 18294 26812
rect 19886 26800 19892 26812
rect 19944 26840 19950 26852
rect 21054 26840 21082 26880
rect 26050 26868 26056 26880
rect 26108 26868 26114 26920
rect 26234 26908 26240 26920
rect 26147 26880 26240 26908
rect 26234 26868 26240 26880
rect 26292 26908 26298 26920
rect 26602 26908 26608 26920
rect 26292 26880 26608 26908
rect 26292 26868 26298 26880
rect 26602 26868 26608 26880
rect 26660 26868 26666 26920
rect 26786 26908 26792 26920
rect 26747 26880 26792 26908
rect 26786 26868 26792 26880
rect 26844 26868 26850 26920
rect 27706 26868 27712 26920
rect 27764 26908 27770 26920
rect 27928 26911 27986 26917
rect 27928 26908 27940 26911
rect 27764 26880 27940 26908
rect 27764 26868 27770 26880
rect 27928 26877 27940 26880
rect 27974 26908 27986 26911
rect 28353 26911 28411 26917
rect 28353 26908 28365 26911
rect 27974 26880 28365 26908
rect 27974 26877 27986 26880
rect 27928 26871 27986 26877
rect 28353 26877 28365 26880
rect 28399 26908 28411 26911
rect 28810 26908 28816 26920
rect 28399 26880 28816 26908
rect 28399 26877 28411 26880
rect 28353 26871 28411 26877
rect 28810 26868 28816 26880
rect 28868 26868 28874 26920
rect 29340 26911 29398 26917
rect 29340 26877 29352 26911
rect 29386 26908 29398 26911
rect 34701 26911 34759 26917
rect 29386 26880 30236 26908
rect 29386 26877 29398 26880
rect 29340 26871 29398 26877
rect 19944 26812 21082 26840
rect 21453 26843 21511 26849
rect 19944 26800 19950 26812
rect 21453 26809 21465 26843
rect 21499 26840 21511 26843
rect 21907 26843 21965 26849
rect 21907 26840 21919 26843
rect 21499 26812 21919 26840
rect 21499 26809 21511 26812
rect 21453 26803 21511 26809
rect 21907 26809 21919 26812
rect 21953 26840 21965 26843
rect 23477 26843 23535 26849
rect 23477 26840 23489 26843
rect 21953 26812 23489 26840
rect 21953 26809 21965 26812
rect 21907 26803 21965 26809
rect 23477 26809 23489 26812
rect 23523 26840 23535 26843
rect 23658 26840 23664 26852
rect 23523 26812 23664 26840
rect 23523 26809 23535 26812
rect 23477 26803 23535 26809
rect 5626 26732 5632 26784
rect 5684 26772 5690 26784
rect 5905 26775 5963 26781
rect 5905 26772 5917 26775
rect 5684 26744 5917 26772
rect 5684 26732 5690 26744
rect 5905 26741 5917 26744
rect 5951 26741 5963 26775
rect 8754 26772 8760 26784
rect 8715 26744 8760 26772
rect 5905 26735 5963 26741
rect 8754 26732 8760 26744
rect 8812 26732 8818 26784
rect 12342 26732 12348 26784
rect 12400 26772 12406 26784
rect 13633 26775 13691 26781
rect 13633 26772 13645 26775
rect 12400 26744 13645 26772
rect 12400 26732 12406 26744
rect 13633 26741 13645 26744
rect 13679 26772 13691 26775
rect 13722 26772 13728 26784
rect 13679 26744 13728 26772
rect 13679 26741 13691 26744
rect 13633 26735 13691 26741
rect 13722 26732 13728 26744
rect 13780 26732 13786 26784
rect 15930 26732 15936 26784
rect 15988 26772 15994 26784
rect 16071 26775 16129 26781
rect 16071 26772 16083 26775
rect 15988 26744 16083 26772
rect 15988 26732 15994 26744
rect 16071 26741 16083 26744
rect 16117 26741 16129 26775
rect 16071 26735 16129 26741
rect 17083 26775 17141 26781
rect 17083 26741 17095 26775
rect 17129 26772 17141 26775
rect 17310 26772 17316 26784
rect 17129 26744 17316 26772
rect 17129 26741 17141 26744
rect 17083 26735 17141 26741
rect 17310 26732 17316 26744
rect 17368 26732 17374 26784
rect 17865 26775 17923 26781
rect 17865 26741 17877 26775
rect 17911 26772 17923 26775
rect 18248 26772 18276 26800
rect 17911 26744 18276 26772
rect 20671 26775 20729 26781
rect 17911 26741 17923 26744
rect 17865 26735 17923 26741
rect 20671 26741 20683 26775
rect 20717 26772 20729 26775
rect 20898 26772 20904 26784
rect 20717 26744 20904 26772
rect 20717 26741 20729 26744
rect 20671 26735 20729 26741
rect 20898 26732 20904 26744
rect 20956 26732 20962 26784
rect 21085 26775 21143 26781
rect 21085 26741 21097 26775
rect 21131 26772 21143 26775
rect 21174 26772 21180 26784
rect 21131 26744 21180 26772
rect 21131 26741 21143 26744
rect 21085 26735 21143 26741
rect 21174 26732 21180 26744
rect 21232 26772 21238 26784
rect 21468 26772 21496 26803
rect 23658 26800 23664 26812
rect 23716 26840 23722 26852
rect 23982 26843 24040 26849
rect 23982 26840 23994 26843
rect 23716 26812 23994 26840
rect 23716 26800 23722 26812
rect 23982 26809 23994 26812
rect 24028 26840 24040 26843
rect 25774 26840 25780 26852
rect 24028 26812 25780 26840
rect 24028 26809 24040 26812
rect 23982 26803 24040 26809
rect 25774 26800 25780 26812
rect 25832 26800 25838 26852
rect 25869 26843 25927 26849
rect 25869 26809 25881 26843
rect 25915 26840 25927 26843
rect 26804 26840 26832 26868
rect 25915 26812 26832 26840
rect 25915 26809 25927 26812
rect 25869 26803 25927 26809
rect 27338 26800 27344 26852
rect 27396 26840 27402 26852
rect 29730 26840 29736 26852
rect 27396 26812 29736 26840
rect 27396 26800 27402 26812
rect 29730 26800 29736 26812
rect 29788 26800 29794 26852
rect 22462 26772 22468 26784
rect 21232 26744 21496 26772
rect 22423 26744 22468 26772
rect 21232 26732 21238 26744
rect 22462 26732 22468 26744
rect 22520 26732 22526 26784
rect 27798 26732 27804 26784
rect 27856 26772 27862 26784
rect 30208 26781 30236 26880
rect 34701 26877 34713 26911
rect 34747 26908 34759 26911
rect 35434 26908 35440 26920
rect 34747 26880 35440 26908
rect 34747 26877 34759 26880
rect 34701 26871 34759 26877
rect 35434 26868 35440 26880
rect 35492 26868 35498 26920
rect 35710 26908 35716 26920
rect 35671 26880 35716 26908
rect 35710 26868 35716 26880
rect 35768 26868 35774 26920
rect 40862 26868 40868 26920
rect 40920 26908 40926 26920
rect 41141 26911 41199 26917
rect 41141 26908 41153 26911
rect 40920 26880 41153 26908
rect 40920 26868 40926 26880
rect 41141 26877 41153 26880
rect 41187 26908 41199 26911
rect 41322 26908 41328 26920
rect 41187 26880 41328 26908
rect 41187 26877 41199 26880
rect 41141 26871 41199 26877
rect 41322 26868 41328 26880
rect 41380 26868 41386 26920
rect 42978 26868 42984 26920
rect 43036 26908 43042 26920
rect 43308 26911 43366 26917
rect 43308 26908 43320 26911
rect 43036 26880 43320 26908
rect 43036 26868 43042 26880
rect 43308 26877 43320 26880
rect 43354 26908 43366 26911
rect 44085 26911 44143 26917
rect 44085 26908 44097 26911
rect 43354 26880 44097 26908
rect 43354 26877 43366 26880
rect 43308 26871 43366 26877
rect 44085 26877 44097 26880
rect 44131 26877 44143 26911
rect 44085 26871 44143 26877
rect 30929 26843 30987 26849
rect 30929 26809 30941 26843
rect 30975 26809 30987 26843
rect 30929 26803 30987 26809
rect 28031 26775 28089 26781
rect 28031 26772 28043 26775
rect 27856 26744 28043 26772
rect 27856 26732 27862 26744
rect 28031 26741 28043 26744
rect 28077 26741 28089 26775
rect 28031 26735 28089 26741
rect 30193 26775 30251 26781
rect 30193 26741 30205 26775
rect 30239 26772 30251 26775
rect 30282 26772 30288 26784
rect 30239 26744 30288 26772
rect 30239 26741 30251 26744
rect 30193 26735 30251 26741
rect 30282 26732 30288 26744
rect 30340 26732 30346 26784
rect 30558 26732 30564 26784
rect 30616 26772 30622 26784
rect 30944 26772 30972 26803
rect 32490 26800 32496 26852
rect 32548 26840 32554 26852
rect 35897 26843 35955 26849
rect 32548 26812 32593 26840
rect 32548 26800 32554 26812
rect 35897 26809 35909 26843
rect 35943 26840 35955 26843
rect 36078 26840 36084 26852
rect 35943 26812 36084 26840
rect 35943 26809 35955 26812
rect 35897 26803 35955 26809
rect 36078 26800 36084 26812
rect 36136 26800 36142 26852
rect 37046 26843 37104 26849
rect 37046 26809 37058 26843
rect 37092 26809 37104 26843
rect 37046 26803 37104 26809
rect 33778 26772 33784 26784
rect 30616 26744 30972 26772
rect 33739 26744 33784 26772
rect 30616 26732 30622 26744
rect 33778 26732 33784 26744
rect 33836 26732 33842 26784
rect 36170 26732 36176 26784
rect 36228 26772 36234 26784
rect 36541 26775 36599 26781
rect 36541 26772 36553 26775
rect 36228 26744 36553 26772
rect 36228 26732 36234 26744
rect 36541 26741 36553 26744
rect 36587 26772 36599 26775
rect 37061 26772 37089 26803
rect 38654 26800 38660 26852
rect 38712 26840 38718 26852
rect 39209 26843 39267 26849
rect 38712 26812 38757 26840
rect 38712 26800 38718 26812
rect 39209 26809 39221 26843
rect 39255 26840 39267 26843
rect 39942 26840 39948 26852
rect 39255 26812 39948 26840
rect 39255 26809 39267 26812
rect 39209 26803 39267 26809
rect 39942 26800 39948 26812
rect 40000 26800 40006 26852
rect 41506 26800 41512 26852
rect 41564 26840 41570 26852
rect 41877 26843 41935 26849
rect 41877 26840 41889 26843
rect 41564 26812 41889 26840
rect 41564 26800 41570 26812
rect 41877 26809 41889 26812
rect 41923 26809 41935 26843
rect 41877 26803 41935 26809
rect 36587 26744 37089 26772
rect 37645 26775 37703 26781
rect 36587 26741 36599 26744
rect 36541 26735 36599 26741
rect 37645 26741 37657 26775
rect 37691 26772 37703 26775
rect 38672 26772 38700 26800
rect 39758 26772 39764 26784
rect 37691 26744 38700 26772
rect 39719 26744 39764 26772
rect 37691 26741 37703 26744
rect 37645 26735 37703 26741
rect 39758 26732 39764 26744
rect 39816 26732 39822 26784
rect 40819 26775 40877 26781
rect 40819 26741 40831 26775
rect 40865 26772 40877 26775
rect 41046 26772 41052 26784
rect 40865 26744 41052 26772
rect 40865 26741 40877 26744
rect 40819 26735 40877 26741
rect 41046 26732 41052 26744
rect 41104 26732 41110 26784
rect 41892 26772 41920 26803
rect 42705 26775 42763 26781
rect 42705 26772 42717 26775
rect 41892 26744 42717 26772
rect 42705 26741 42717 26744
rect 42751 26741 42763 26775
rect 42705 26735 42763 26741
rect 1104 26682 48852 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 48852 26682
rect 1104 26608 48852 26630
rect 3881 26571 3939 26577
rect 3881 26537 3893 26571
rect 3927 26568 3939 26571
rect 4062 26568 4068 26580
rect 3927 26540 4068 26568
rect 3927 26537 3939 26540
rect 3881 26531 3939 26537
rect 4062 26528 4068 26540
rect 4120 26528 4126 26580
rect 4246 26528 4252 26580
rect 4304 26568 4310 26580
rect 4341 26571 4399 26577
rect 4341 26568 4353 26571
rect 4304 26540 4353 26568
rect 4304 26528 4310 26540
rect 4341 26537 4353 26540
rect 4387 26537 4399 26571
rect 5810 26568 5816 26580
rect 5771 26540 5816 26568
rect 4341 26531 4399 26537
rect 5810 26528 5816 26540
rect 5868 26528 5874 26580
rect 6914 26528 6920 26580
rect 6972 26568 6978 26580
rect 7009 26571 7067 26577
rect 7009 26568 7021 26571
rect 6972 26540 7021 26568
rect 6972 26528 6978 26540
rect 7009 26537 7021 26540
rect 7055 26537 7067 26571
rect 7558 26568 7564 26580
rect 7519 26540 7564 26568
rect 7009 26531 7067 26537
rect 7558 26528 7564 26540
rect 7616 26528 7622 26580
rect 8757 26571 8815 26577
rect 8757 26537 8769 26571
rect 8803 26537 8815 26571
rect 8757 26531 8815 26537
rect 4706 26500 4712 26512
rect 4356 26472 4712 26500
rect 3786 26392 3792 26444
rect 3844 26432 3850 26444
rect 4356 26441 4384 26472
rect 4706 26460 4712 26472
rect 4764 26500 4770 26512
rect 5828 26500 5856 26528
rect 4764 26472 5856 26500
rect 8772 26500 8800 26531
rect 10134 26528 10140 26580
rect 10192 26568 10198 26580
rect 11149 26571 11207 26577
rect 11149 26568 11161 26571
rect 10192 26540 11161 26568
rect 10192 26528 10198 26540
rect 11149 26537 11161 26540
rect 11195 26537 11207 26571
rect 11149 26531 11207 26537
rect 12250 26528 12256 26580
rect 12308 26568 12314 26580
rect 12308 26540 12480 26568
rect 12308 26528 12314 26540
rect 10318 26500 10324 26512
rect 8772 26472 10324 26500
rect 4764 26460 4770 26472
rect 10318 26460 10324 26472
rect 10376 26460 10382 26512
rect 10594 26509 10600 26512
rect 10591 26500 10600 26509
rect 10555 26472 10600 26500
rect 10591 26463 10600 26472
rect 10594 26460 10600 26463
rect 10652 26460 10658 26512
rect 12452 26500 12480 26540
rect 12526 26528 12532 26580
rect 12584 26568 12590 26580
rect 12989 26571 13047 26577
rect 12989 26568 13001 26571
rect 12584 26540 13001 26568
rect 12584 26528 12590 26540
rect 12989 26537 13001 26540
rect 13035 26537 13047 26571
rect 12989 26531 13047 26537
rect 13906 26528 13912 26580
rect 13964 26568 13970 26580
rect 16850 26568 16856 26580
rect 13964 26540 15516 26568
rect 16811 26540 16856 26568
rect 13964 26528 13970 26540
rect 15488 26512 15516 26540
rect 16850 26528 16856 26540
rect 16908 26528 16914 26580
rect 18138 26528 18144 26580
rect 18196 26568 18202 26580
rect 18417 26571 18475 26577
rect 18417 26568 18429 26571
rect 18196 26540 18429 26568
rect 18196 26528 18202 26540
rect 18417 26537 18429 26540
rect 18463 26537 18475 26571
rect 21082 26568 21088 26580
rect 21043 26540 21088 26568
rect 18417 26531 18475 26537
rect 21082 26528 21088 26540
rect 21140 26528 21146 26580
rect 21542 26528 21548 26580
rect 21600 26568 21606 26580
rect 22189 26571 22247 26577
rect 22189 26568 22201 26571
rect 21600 26540 22201 26568
rect 21600 26528 21606 26540
rect 22189 26537 22201 26540
rect 22235 26537 22247 26571
rect 24026 26568 24032 26580
rect 23987 26540 24032 26568
rect 22189 26531 22247 26537
rect 24026 26528 24032 26540
rect 24084 26528 24090 26580
rect 24397 26571 24455 26577
rect 24397 26537 24409 26571
rect 24443 26568 24455 26571
rect 24486 26568 24492 26580
rect 24443 26540 24492 26568
rect 24443 26537 24455 26540
rect 24397 26531 24455 26537
rect 24486 26528 24492 26540
rect 24544 26528 24550 26580
rect 27801 26571 27859 26577
rect 27801 26537 27813 26571
rect 27847 26568 27859 26571
rect 28626 26568 28632 26580
rect 27847 26540 28632 26568
rect 27847 26537 27859 26540
rect 27801 26531 27859 26537
rect 28626 26528 28632 26540
rect 28684 26568 28690 26580
rect 32355 26571 32413 26577
rect 28684 26540 28856 26568
rect 28684 26528 28690 26540
rect 12452 26472 13584 26500
rect 13556 26444 13584 26472
rect 14182 26460 14188 26512
rect 14240 26500 14246 26512
rect 14277 26503 14335 26509
rect 14277 26500 14289 26503
rect 14240 26472 14289 26500
rect 14240 26460 14246 26472
rect 14277 26469 14289 26472
rect 14323 26469 14335 26503
rect 15470 26500 15476 26512
rect 15383 26472 15476 26500
rect 14277 26463 14335 26469
rect 15470 26460 15476 26472
rect 15528 26460 15534 26512
rect 16022 26500 16028 26512
rect 15983 26472 16028 26500
rect 16022 26460 16028 26472
rect 16080 26460 16086 26512
rect 17494 26460 17500 26512
rect 17552 26500 17558 26512
rect 17589 26503 17647 26509
rect 17589 26500 17601 26503
rect 17552 26472 17601 26500
rect 17552 26460 17558 26472
rect 17589 26469 17601 26472
rect 17635 26500 17647 26503
rect 18969 26503 19027 26509
rect 18969 26500 18981 26503
rect 17635 26472 18981 26500
rect 17635 26469 17647 26472
rect 17589 26463 17647 26469
rect 18969 26469 18981 26472
rect 19015 26469 19027 26503
rect 18969 26463 19027 26469
rect 22462 26460 22468 26512
rect 22520 26500 22526 26512
rect 22557 26503 22615 26509
rect 22557 26500 22569 26503
rect 22520 26472 22569 26500
rect 22520 26460 22526 26472
rect 22557 26469 22569 26472
rect 22603 26469 22615 26503
rect 24504 26500 24532 26528
rect 24673 26503 24731 26509
rect 24673 26500 24685 26503
rect 24504 26472 24685 26500
rect 22557 26463 22615 26469
rect 24673 26469 24685 26472
rect 24719 26469 24731 26503
rect 24673 26463 24731 26469
rect 25774 26460 25780 26512
rect 25832 26500 25838 26512
rect 27202 26503 27260 26509
rect 27202 26500 27214 26503
rect 25832 26472 27214 26500
rect 25832 26460 25838 26472
rect 27202 26469 27214 26472
rect 27248 26500 27260 26503
rect 27338 26500 27344 26512
rect 27248 26472 27344 26500
rect 27248 26469 27260 26472
rect 27202 26463 27260 26469
rect 27338 26460 27344 26472
rect 27396 26460 27402 26512
rect 28828 26509 28856 26540
rect 32355 26537 32367 26571
rect 32401 26568 32413 26571
rect 33318 26568 33324 26580
rect 32401 26540 33324 26568
rect 32401 26537 32413 26540
rect 32355 26531 32413 26537
rect 33318 26528 33324 26540
rect 33376 26528 33382 26580
rect 35342 26568 35348 26580
rect 35303 26540 35348 26568
rect 35342 26528 35348 26540
rect 35400 26528 35406 26580
rect 35710 26568 35716 26580
rect 35671 26540 35716 26568
rect 35710 26528 35716 26540
rect 35768 26528 35774 26580
rect 36170 26528 36176 26580
rect 36228 26568 36234 26580
rect 36265 26571 36323 26577
rect 36265 26568 36277 26571
rect 36228 26540 36277 26568
rect 36228 26528 36234 26540
rect 36265 26537 36277 26540
rect 36311 26537 36323 26571
rect 36265 26531 36323 26537
rect 38120 26540 39712 26568
rect 28813 26503 28871 26509
rect 28813 26469 28825 26503
rect 28859 26469 28871 26503
rect 28813 26463 28871 26469
rect 32030 26460 32036 26512
rect 32088 26500 32094 26512
rect 33413 26503 33471 26509
rect 32088 26472 32295 26500
rect 32088 26460 32094 26472
rect 4341 26435 4399 26441
rect 4341 26432 4353 26435
rect 3844 26404 4353 26432
rect 3844 26392 3850 26404
rect 4341 26401 4353 26404
rect 4387 26401 4399 26435
rect 4614 26432 4620 26444
rect 4575 26404 4620 26432
rect 4341 26395 4399 26401
rect 4614 26392 4620 26404
rect 4672 26392 4678 26444
rect 5626 26432 5632 26444
rect 5587 26404 5632 26432
rect 5626 26392 5632 26404
rect 5684 26392 5690 26444
rect 8570 26432 8576 26444
rect 8531 26404 8576 26432
rect 8570 26392 8576 26404
rect 8628 26392 8634 26444
rect 12250 26392 12256 26444
rect 12308 26432 12314 26444
rect 12529 26435 12587 26441
rect 12529 26432 12541 26435
rect 12308 26404 12541 26432
rect 12308 26392 12314 26404
rect 12529 26401 12541 26404
rect 12575 26401 12587 26435
rect 13538 26432 13544 26444
rect 13451 26404 13544 26432
rect 12529 26395 12587 26401
rect 13538 26392 13544 26404
rect 13596 26392 13602 26444
rect 13998 26432 14004 26444
rect 13786 26404 14004 26432
rect 13786 26376 13814 26404
rect 13998 26392 14004 26404
rect 14056 26392 14062 26444
rect 19058 26432 19064 26444
rect 18524 26404 19064 26432
rect 6641 26367 6699 26373
rect 6641 26333 6653 26367
rect 6687 26364 6699 26367
rect 6914 26364 6920 26376
rect 6687 26336 6920 26364
rect 6687 26333 6699 26336
rect 6641 26327 6699 26333
rect 6914 26324 6920 26336
rect 6972 26324 6978 26376
rect 10226 26364 10232 26376
rect 10187 26336 10232 26364
rect 10226 26324 10232 26336
rect 10284 26324 10290 26376
rect 13449 26367 13507 26373
rect 13449 26333 13461 26367
rect 13495 26364 13507 26367
rect 13722 26364 13728 26376
rect 13495 26336 13728 26364
rect 13495 26333 13507 26336
rect 13449 26327 13507 26333
rect 13722 26324 13728 26336
rect 13780 26336 13814 26376
rect 15381 26367 15439 26373
rect 13780 26324 13786 26336
rect 15381 26333 15393 26367
rect 15427 26364 15439 26367
rect 15838 26364 15844 26376
rect 15427 26336 15844 26364
rect 15427 26333 15439 26336
rect 15381 26327 15439 26333
rect 15838 26324 15844 26336
rect 15896 26324 15902 26376
rect 17218 26324 17224 26376
rect 17276 26364 17282 26376
rect 17497 26367 17555 26373
rect 17497 26364 17509 26367
rect 17276 26336 17509 26364
rect 17276 26324 17282 26336
rect 17497 26333 17509 26336
rect 17543 26333 17555 26367
rect 17497 26327 17555 26333
rect 18141 26367 18199 26373
rect 18141 26333 18153 26367
rect 18187 26364 18199 26367
rect 18414 26364 18420 26376
rect 18187 26336 18420 26364
rect 18187 26333 18199 26336
rect 18141 26327 18199 26333
rect 18414 26324 18420 26336
rect 18472 26324 18478 26376
rect 9950 26256 9956 26308
rect 10008 26296 10014 26308
rect 18524 26296 18552 26404
rect 19058 26392 19064 26404
rect 19116 26392 19122 26444
rect 21266 26392 21272 26444
rect 21324 26432 21330 26444
rect 21396 26435 21454 26441
rect 21396 26432 21408 26435
rect 21324 26404 21408 26432
rect 21324 26392 21330 26404
rect 21396 26401 21408 26404
rect 21442 26401 21454 26435
rect 21396 26395 21454 26401
rect 30742 26392 30748 26444
rect 30800 26432 30806 26444
rect 30872 26435 30930 26441
rect 30872 26432 30884 26435
rect 30800 26404 30884 26432
rect 30800 26392 30806 26404
rect 30872 26401 30884 26404
rect 30918 26432 30930 26435
rect 32122 26432 32128 26444
rect 30918 26404 32128 26432
rect 30918 26401 30930 26404
rect 30872 26395 30930 26401
rect 32122 26392 32128 26404
rect 32180 26392 32186 26444
rect 32267 26441 32295 26472
rect 33413 26469 33425 26503
rect 33459 26500 33471 26503
rect 33778 26500 33784 26512
rect 33459 26472 33784 26500
rect 33459 26469 33471 26472
rect 33413 26463 33471 26469
rect 33778 26460 33784 26472
rect 33836 26460 33842 26512
rect 38120 26509 38148 26540
rect 38105 26503 38163 26509
rect 38105 26469 38117 26503
rect 38151 26469 38163 26503
rect 38105 26463 38163 26469
rect 38286 26460 38292 26512
rect 38344 26500 38350 26512
rect 38933 26503 38991 26509
rect 38933 26500 38945 26503
rect 38344 26472 38945 26500
rect 38344 26460 38350 26472
rect 38933 26469 38945 26472
rect 38979 26469 38991 26503
rect 39574 26500 39580 26512
rect 39535 26472 39580 26500
rect 38933 26463 38991 26469
rect 39574 26460 39580 26472
rect 39632 26460 39638 26512
rect 39684 26509 39712 26540
rect 41046 26528 41052 26580
rect 41104 26568 41110 26580
rect 43070 26568 43076 26580
rect 41104 26540 43076 26568
rect 41104 26528 41110 26540
rect 43070 26528 43076 26540
rect 43128 26568 43134 26580
rect 43128 26540 43484 26568
rect 43128 26528 43134 26540
rect 39669 26503 39727 26509
rect 39669 26469 39681 26503
rect 39715 26500 39727 26503
rect 39758 26500 39764 26512
rect 39715 26472 39764 26500
rect 39715 26469 39727 26472
rect 39669 26463 39727 26469
rect 39758 26460 39764 26472
rect 39816 26460 39822 26512
rect 40221 26503 40279 26509
rect 40221 26469 40233 26503
rect 40267 26500 40279 26503
rect 40770 26500 40776 26512
rect 40267 26472 40776 26500
rect 40267 26469 40279 26472
rect 40221 26463 40279 26469
rect 40770 26460 40776 26472
rect 40828 26460 40834 26512
rect 41598 26500 41604 26512
rect 41559 26472 41604 26500
rect 41598 26460 41604 26472
rect 41656 26460 41662 26512
rect 41874 26500 41880 26512
rect 41835 26472 41880 26500
rect 41874 26460 41880 26472
rect 41932 26460 41938 26512
rect 42426 26500 42432 26512
rect 42387 26472 42432 26500
rect 42426 26460 42432 26472
rect 42484 26460 42490 26512
rect 43456 26509 43484 26540
rect 43441 26503 43499 26509
rect 43441 26469 43453 26503
rect 43487 26469 43499 26503
rect 43441 26463 43499 26469
rect 43530 26460 43536 26512
rect 43588 26500 43594 26512
rect 43588 26472 43633 26500
rect 43588 26460 43594 26472
rect 32252 26435 32310 26441
rect 32252 26401 32264 26435
rect 32298 26401 32310 26435
rect 34790 26432 34796 26444
rect 34751 26404 34796 26432
rect 32252 26395 32310 26401
rect 34790 26392 34796 26404
rect 34848 26392 34854 26444
rect 35894 26432 35900 26444
rect 35855 26404 35900 26432
rect 35894 26392 35900 26404
rect 35952 26392 35958 26444
rect 22465 26367 22523 26373
rect 22465 26333 22477 26367
rect 22511 26364 22523 26367
rect 22922 26364 22928 26376
rect 22511 26336 22928 26364
rect 22511 26333 22523 26336
rect 22465 26327 22523 26333
rect 22922 26324 22928 26336
rect 22980 26324 22986 26376
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26364 24639 26367
rect 25590 26364 25596 26376
rect 24627 26336 25596 26364
rect 24627 26333 24639 26336
rect 24581 26327 24639 26333
rect 25590 26324 25596 26336
rect 25648 26324 25654 26376
rect 26878 26364 26884 26376
rect 26839 26336 26884 26364
rect 26878 26324 26884 26336
rect 26936 26324 26942 26376
rect 28721 26367 28779 26373
rect 28721 26333 28733 26367
rect 28767 26364 28779 26367
rect 29086 26364 29092 26376
rect 28767 26336 29092 26364
rect 28767 26333 28779 26336
rect 28721 26327 28779 26333
rect 29086 26324 29092 26336
rect 29144 26324 29150 26376
rect 33134 26324 33140 26376
rect 33192 26364 33198 26376
rect 33321 26367 33379 26373
rect 33321 26364 33333 26367
rect 33192 26336 33333 26364
rect 33192 26324 33198 26336
rect 33321 26333 33333 26336
rect 33367 26333 33379 26367
rect 33321 26327 33379 26333
rect 38013 26367 38071 26373
rect 38013 26333 38025 26367
rect 38059 26364 38071 26367
rect 38470 26364 38476 26376
rect 38059 26336 38476 26364
rect 38059 26333 38071 26336
rect 38013 26327 38071 26333
rect 38470 26324 38476 26336
rect 38528 26324 38534 26376
rect 41782 26364 41788 26376
rect 41743 26336 41788 26364
rect 41782 26324 41788 26336
rect 41840 26324 41846 26376
rect 43717 26367 43775 26373
rect 43717 26364 43729 26367
rect 43548 26336 43729 26364
rect 10008 26268 18552 26296
rect 21499 26299 21557 26305
rect 10008 26256 10014 26268
rect 21499 26265 21511 26299
rect 21545 26296 21557 26299
rect 22830 26296 22836 26308
rect 21545 26268 22836 26296
rect 21545 26265 21557 26268
rect 21499 26259 21557 26265
rect 22830 26256 22836 26268
rect 22888 26256 22894 26308
rect 23017 26299 23075 26305
rect 23017 26265 23029 26299
rect 23063 26265 23075 26299
rect 25130 26296 25136 26308
rect 25091 26268 25136 26296
rect 23017 26259 23075 26265
rect 9858 26228 9864 26240
rect 9819 26200 9864 26228
rect 9858 26188 9864 26200
rect 9916 26188 9922 26240
rect 12253 26231 12311 26237
rect 12253 26197 12265 26231
rect 12299 26228 12311 26231
rect 12526 26228 12532 26240
rect 12299 26200 12532 26228
rect 12299 26197 12311 26200
rect 12253 26191 12311 26197
rect 12526 26188 12532 26200
rect 12584 26188 12590 26240
rect 12710 26228 12716 26240
rect 12671 26200 12716 26228
rect 12710 26188 12716 26200
rect 12768 26188 12774 26240
rect 14550 26228 14556 26240
rect 14511 26200 14556 26228
rect 14550 26188 14556 26200
rect 14608 26188 14614 26240
rect 19978 26228 19984 26240
rect 19939 26200 19984 26228
rect 19978 26188 19984 26200
rect 20036 26188 20042 26240
rect 21818 26228 21824 26240
rect 21779 26200 21824 26228
rect 21818 26188 21824 26200
rect 21876 26188 21882 26240
rect 22278 26188 22284 26240
rect 22336 26228 22342 26240
rect 23032 26228 23060 26259
rect 25130 26256 25136 26268
rect 25188 26256 25194 26308
rect 27522 26256 27528 26308
rect 27580 26296 27586 26308
rect 29273 26299 29331 26305
rect 29273 26296 29285 26299
rect 27580 26268 29285 26296
rect 27580 26256 27586 26268
rect 29273 26265 29285 26268
rect 29319 26296 29331 26299
rect 31110 26296 31116 26308
rect 29319 26268 31116 26296
rect 29319 26265 29331 26268
rect 29273 26259 29331 26265
rect 31110 26256 31116 26268
rect 31168 26256 31174 26308
rect 31941 26299 31999 26305
rect 31941 26265 31953 26299
rect 31987 26296 31999 26299
rect 32214 26296 32220 26308
rect 31987 26268 32220 26296
rect 31987 26265 31999 26268
rect 31941 26259 31999 26265
rect 32214 26256 32220 26268
rect 32272 26296 32278 26308
rect 33870 26296 33876 26308
rect 32272 26268 33876 26296
rect 32272 26256 32278 26268
rect 33870 26256 33876 26268
rect 33928 26256 33934 26308
rect 38562 26296 38568 26308
rect 38523 26268 38568 26296
rect 38562 26256 38568 26268
rect 38620 26296 38626 26308
rect 39301 26299 39359 26305
rect 39301 26296 39313 26299
rect 38620 26268 39313 26296
rect 38620 26256 38626 26268
rect 39301 26265 39313 26268
rect 39347 26265 39359 26299
rect 39301 26259 39359 26265
rect 40310 26256 40316 26308
rect 40368 26296 40374 26308
rect 42518 26296 42524 26308
rect 40368 26268 42524 26296
rect 40368 26256 40374 26268
rect 42518 26256 42524 26268
rect 42576 26296 42582 26308
rect 43548 26296 43576 26336
rect 43717 26333 43729 26336
rect 43763 26333 43775 26367
rect 43717 26327 43775 26333
rect 42576 26268 43576 26296
rect 42576 26256 42582 26268
rect 22336 26200 23060 26228
rect 28169 26231 28227 26237
rect 22336 26188 22342 26200
rect 28169 26197 28181 26231
rect 28215 26228 28227 26231
rect 28258 26228 28264 26240
rect 28215 26200 28264 26228
rect 28215 26197 28227 26200
rect 28169 26191 28227 26197
rect 28258 26188 28264 26200
rect 28316 26188 28322 26240
rect 30975 26231 31033 26237
rect 30975 26197 30987 26231
rect 31021 26228 31033 26231
rect 31294 26228 31300 26240
rect 31021 26200 31300 26228
rect 31021 26197 31033 26200
rect 30975 26191 31033 26197
rect 31294 26188 31300 26200
rect 31352 26188 31358 26240
rect 32674 26228 32680 26240
rect 32635 26200 32680 26228
rect 32674 26188 32680 26200
rect 32732 26188 32738 26240
rect 33410 26188 33416 26240
rect 33468 26228 33474 26240
rect 34931 26231 34989 26237
rect 34931 26228 34943 26231
rect 33468 26200 34943 26228
rect 33468 26188 33474 26200
rect 34931 26197 34943 26200
rect 34977 26197 34989 26231
rect 34931 26191 34989 26197
rect 36817 26231 36875 26237
rect 36817 26197 36829 26231
rect 36863 26228 36875 26231
rect 37734 26228 37740 26240
rect 36863 26200 37740 26228
rect 36863 26197 36875 26200
rect 36817 26191 36875 26197
rect 37734 26188 37740 26200
rect 37792 26188 37798 26240
rect 1104 26138 48852 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 48852 26138
rect 1104 26064 48852 26086
rect 4706 26024 4712 26036
rect 4667 25996 4712 26024
rect 4706 25984 4712 25996
rect 4764 25984 4770 26036
rect 4798 25984 4804 26036
rect 4856 26024 4862 26036
rect 5350 26024 5356 26036
rect 4856 25996 5356 26024
rect 4856 25984 4862 25996
rect 5350 25984 5356 25996
rect 5408 25984 5414 26036
rect 6641 26027 6699 26033
rect 6641 25993 6653 26027
rect 6687 26024 6699 26027
rect 6822 26024 6828 26036
rect 6687 25996 6828 26024
rect 6687 25993 6699 25996
rect 6641 25987 6699 25993
rect 6822 25984 6828 25996
rect 6880 25984 6886 26036
rect 8573 26027 8631 26033
rect 8573 26024 8585 26027
rect 7852 25996 8585 26024
rect 3970 25916 3976 25968
rect 4028 25956 4034 25968
rect 4341 25959 4399 25965
rect 4341 25956 4353 25959
rect 4028 25928 4353 25956
rect 4028 25916 4034 25928
rect 4341 25925 4353 25928
rect 4387 25925 4399 25959
rect 4341 25919 4399 25925
rect 5626 25848 5632 25900
rect 5684 25888 5690 25900
rect 5721 25891 5779 25897
rect 5721 25888 5733 25891
rect 5684 25860 5733 25888
rect 5684 25848 5690 25860
rect 5721 25857 5733 25860
rect 5767 25888 5779 25891
rect 5767 25860 7052 25888
rect 5767 25857 5779 25860
rect 5721 25851 5779 25857
rect 3145 25823 3203 25829
rect 3145 25789 3157 25823
rect 3191 25820 3203 25823
rect 4157 25823 4215 25829
rect 3191 25792 3740 25820
rect 3191 25789 3203 25792
rect 3145 25783 3203 25789
rect 3712 25696 3740 25792
rect 4157 25789 4169 25823
rect 4203 25820 4215 25823
rect 4338 25820 4344 25832
rect 4203 25792 4344 25820
rect 4203 25789 4215 25792
rect 4157 25783 4215 25789
rect 4338 25780 4344 25792
rect 4396 25820 4402 25832
rect 7024 25829 7052 25860
rect 4985 25823 5043 25829
rect 4985 25820 4997 25823
rect 4396 25792 4997 25820
rect 4396 25780 4402 25792
rect 4985 25789 4997 25792
rect 5031 25789 5043 25823
rect 4985 25783 5043 25789
rect 5169 25823 5227 25829
rect 5169 25789 5181 25823
rect 5215 25820 5227 25823
rect 7009 25823 7067 25829
rect 5215 25792 6040 25820
rect 5215 25789 5227 25792
rect 5169 25783 5227 25789
rect 6012 25696 6040 25792
rect 7009 25789 7021 25823
rect 7055 25789 7067 25823
rect 7009 25783 7067 25789
rect 7377 25823 7435 25829
rect 7377 25789 7389 25823
rect 7423 25820 7435 25823
rect 7650 25820 7656 25832
rect 7423 25792 7656 25820
rect 7423 25789 7435 25792
rect 7377 25783 7435 25789
rect 6822 25712 6828 25764
rect 6880 25752 6886 25764
rect 7024 25752 7052 25783
rect 7650 25780 7656 25792
rect 7708 25820 7714 25832
rect 7852 25829 7880 25996
rect 8573 25993 8585 25996
rect 8619 25993 8631 26027
rect 8573 25987 8631 25993
rect 11517 26027 11575 26033
rect 11517 25993 11529 26027
rect 11563 26024 11575 26027
rect 12158 26024 12164 26036
rect 11563 25996 12164 26024
rect 11563 25993 11575 25996
rect 11517 25987 11575 25993
rect 12158 25984 12164 25996
rect 12216 25984 12222 26036
rect 13538 26024 13544 26036
rect 13499 25996 13544 26024
rect 13538 25984 13544 25996
rect 13596 25984 13602 26036
rect 14090 26024 14096 26036
rect 14051 25996 14096 26024
rect 14090 25984 14096 25996
rect 14148 25984 14154 26036
rect 14918 25984 14924 26036
rect 14976 26024 14982 26036
rect 15197 26027 15255 26033
rect 15197 26024 15209 26027
rect 14976 25996 15209 26024
rect 14976 25984 14982 25996
rect 15197 25993 15209 25996
rect 15243 25993 15255 26027
rect 15470 26024 15476 26036
rect 15431 25996 15476 26024
rect 15197 25987 15255 25993
rect 15470 25984 15476 25996
rect 15528 25984 15534 26036
rect 15930 26024 15936 26036
rect 15891 25996 15936 26024
rect 15930 25984 15936 25996
rect 15988 25984 15994 26036
rect 16853 26027 16911 26033
rect 16853 25993 16865 26027
rect 16899 26024 16911 26027
rect 17218 26024 17224 26036
rect 16899 25996 17224 26024
rect 16899 25993 16911 25996
rect 16853 25987 16911 25993
rect 17218 25984 17224 25996
rect 17276 25984 17282 26036
rect 17494 26024 17500 26036
rect 17455 25996 17500 26024
rect 17494 25984 17500 25996
rect 17552 25984 17558 26036
rect 18230 25984 18236 26036
rect 18288 26024 18294 26036
rect 18325 26027 18383 26033
rect 18325 26024 18337 26027
rect 18288 25996 18337 26024
rect 18288 25984 18294 25996
rect 18325 25993 18337 25996
rect 18371 25993 18383 26027
rect 19058 26024 19064 26036
rect 19019 25996 19064 26024
rect 18325 25987 18383 25993
rect 19058 25984 19064 25996
rect 19116 25984 19122 26036
rect 21266 25984 21272 26036
rect 21324 26024 21330 26036
rect 21361 26027 21419 26033
rect 21361 26024 21373 26027
rect 21324 25996 21373 26024
rect 21324 25984 21330 25996
rect 21361 25993 21373 25996
rect 21407 25993 21419 26027
rect 21361 25987 21419 25993
rect 22462 25984 22468 26036
rect 22520 26024 22526 26036
rect 22649 26027 22707 26033
rect 22649 26024 22661 26027
rect 22520 25996 22661 26024
rect 22520 25984 22526 25996
rect 22649 25993 22661 25996
rect 22695 25993 22707 26027
rect 22649 25987 22707 25993
rect 22922 25984 22928 26036
rect 22980 26024 22986 26036
rect 23017 26027 23075 26033
rect 23017 26024 23029 26027
rect 22980 25996 23029 26024
rect 22980 25984 22986 25996
rect 23017 25993 23029 25996
rect 23063 25993 23075 26027
rect 23017 25987 23075 25993
rect 24029 26027 24087 26033
rect 24029 25993 24041 26027
rect 24075 26024 24087 26027
rect 24486 26024 24492 26036
rect 24075 25996 24492 26024
rect 24075 25993 24087 25996
rect 24029 25987 24087 25993
rect 24486 25984 24492 25996
rect 24544 26024 24550 26036
rect 25133 26027 25191 26033
rect 25133 26024 25145 26027
rect 24544 25996 25145 26024
rect 24544 25984 24550 25996
rect 25133 25993 25145 25996
rect 25179 25993 25191 26027
rect 25590 26024 25596 26036
rect 25551 25996 25596 26024
rect 25133 25987 25191 25993
rect 25590 25984 25596 25996
rect 25648 25984 25654 26036
rect 26878 25984 26884 26036
rect 26936 26024 26942 26036
rect 27801 26027 27859 26033
rect 27801 26024 27813 26027
rect 26936 25996 27813 26024
rect 26936 25984 26942 25996
rect 27801 25993 27813 25996
rect 27847 25993 27859 26027
rect 28626 26024 28632 26036
rect 28587 25996 28632 26024
rect 27801 25987 27859 25993
rect 28626 25984 28632 25996
rect 28684 25984 28690 26036
rect 33778 26024 33784 26036
rect 33739 25996 33784 26024
rect 33778 25984 33784 25996
rect 33836 25984 33842 26036
rect 34790 25984 34796 26036
rect 34848 26024 34854 26036
rect 35342 26024 35348 26036
rect 34848 25996 35348 26024
rect 34848 25984 34854 25996
rect 35342 25984 35348 25996
rect 35400 25984 35406 26036
rect 37734 26024 37740 26036
rect 37695 25996 37740 26024
rect 37734 25984 37740 25996
rect 37792 25984 37798 26036
rect 39574 25984 39580 26036
rect 39632 26024 39638 26036
rect 39853 26027 39911 26033
rect 39853 26024 39865 26027
rect 39632 25996 39865 26024
rect 39632 25984 39638 25996
rect 39853 25993 39865 25996
rect 39899 25993 39911 26027
rect 39853 25987 39911 25993
rect 41782 25984 41788 26036
rect 41840 26024 41846 26036
rect 42334 26024 42340 26036
rect 41840 25996 42340 26024
rect 41840 25984 41846 25996
rect 42334 25984 42340 25996
rect 42392 26024 42398 26036
rect 42613 26027 42671 26033
rect 42613 26024 42625 26027
rect 42392 25996 42625 26024
rect 42392 25984 42398 25996
rect 42613 25993 42625 25996
rect 42659 25993 42671 26027
rect 43070 26024 43076 26036
rect 43031 25996 43076 26024
rect 42613 25987 42671 25993
rect 43070 25984 43076 25996
rect 43128 25984 43134 26036
rect 10594 25956 10600 25968
rect 10507 25928 10600 25956
rect 10594 25916 10600 25928
rect 10652 25956 10658 25968
rect 14108 25956 14136 25984
rect 10652 25928 14136 25956
rect 10652 25916 10658 25928
rect 7944 25860 8524 25888
rect 7837 25823 7895 25829
rect 7837 25820 7849 25823
rect 7708 25792 7849 25820
rect 7708 25780 7714 25792
rect 7837 25789 7849 25792
rect 7883 25789 7895 25823
rect 7837 25783 7895 25789
rect 6880 25724 7052 25752
rect 6880 25712 6886 25724
rect 3050 25644 3056 25696
rect 3108 25684 3114 25696
rect 3329 25687 3387 25693
rect 3329 25684 3341 25687
rect 3108 25656 3341 25684
rect 3108 25644 3114 25656
rect 3329 25653 3341 25656
rect 3375 25653 3387 25687
rect 3694 25684 3700 25696
rect 3655 25656 3700 25684
rect 3329 25647 3387 25653
rect 3694 25644 3700 25656
rect 3752 25644 3758 25696
rect 4065 25687 4123 25693
rect 4065 25653 4077 25687
rect 4111 25684 4123 25687
rect 4614 25684 4620 25696
rect 4111 25656 4620 25684
rect 4111 25653 4123 25656
rect 4065 25647 4123 25653
rect 4614 25644 4620 25656
rect 4672 25644 4678 25696
rect 5994 25684 6000 25696
rect 5955 25656 6000 25684
rect 5994 25644 6000 25656
rect 6052 25644 6058 25696
rect 6914 25684 6920 25696
rect 6875 25656 6920 25684
rect 6914 25644 6920 25656
rect 6972 25644 6978 25696
rect 7024 25684 7052 25724
rect 7944 25684 7972 25860
rect 8389 25823 8447 25829
rect 8389 25820 8401 25823
rect 8220 25792 8401 25820
rect 8220 25696 8248 25792
rect 8389 25789 8401 25792
rect 8435 25789 8447 25823
rect 8496 25820 8524 25860
rect 8570 25848 8576 25900
rect 8628 25888 8634 25900
rect 8941 25891 8999 25897
rect 8941 25888 8953 25891
rect 8628 25860 8953 25888
rect 8628 25848 8634 25860
rect 8941 25857 8953 25860
rect 8987 25888 8999 25891
rect 11146 25888 11152 25900
rect 8987 25860 11152 25888
rect 8987 25857 8999 25860
rect 8941 25851 8999 25857
rect 11146 25848 11152 25860
rect 11204 25848 11210 25900
rect 9401 25823 9459 25829
rect 9401 25820 9413 25823
rect 8496 25792 9413 25820
rect 8389 25783 8447 25789
rect 9401 25789 9413 25792
rect 9447 25820 9459 25823
rect 9677 25823 9735 25829
rect 9677 25820 9689 25823
rect 9447 25792 9689 25820
rect 9447 25789 9459 25792
rect 9401 25783 9459 25789
rect 9677 25789 9689 25792
rect 9723 25789 9735 25823
rect 9677 25783 9735 25789
rect 8202 25684 8208 25696
rect 7024 25656 7972 25684
rect 8163 25656 8208 25684
rect 8202 25644 8208 25656
rect 8260 25644 8266 25696
rect 9692 25684 9720 25783
rect 9950 25780 9956 25832
rect 10008 25820 10014 25832
rect 10045 25823 10103 25829
rect 10045 25820 10057 25823
rect 10008 25792 10057 25820
rect 10008 25780 10014 25792
rect 10045 25789 10057 25792
rect 10091 25820 10103 25823
rect 10873 25823 10931 25829
rect 10873 25820 10885 25823
rect 10091 25792 10885 25820
rect 10091 25789 10103 25792
rect 10045 25783 10103 25789
rect 10873 25789 10885 25792
rect 10919 25789 10931 25823
rect 10873 25783 10931 25789
rect 11333 25823 11391 25829
rect 11333 25789 11345 25823
rect 11379 25820 11391 25823
rect 11379 25792 11928 25820
rect 11379 25789 11391 25792
rect 11333 25783 11391 25789
rect 10226 25752 10232 25764
rect 10187 25724 10232 25752
rect 10226 25712 10232 25724
rect 10284 25712 10290 25764
rect 9858 25684 9864 25696
rect 9692 25656 9864 25684
rect 9858 25644 9864 25656
rect 9916 25684 9922 25696
rect 11348 25684 11376 25783
rect 11900 25696 11928 25792
rect 12526 25780 12532 25832
rect 12584 25820 12590 25832
rect 12621 25823 12679 25829
rect 12621 25820 12633 25823
rect 12584 25792 12633 25820
rect 12584 25780 12590 25792
rect 12621 25789 12633 25792
rect 12667 25820 12679 25823
rect 13081 25823 13139 25829
rect 13081 25820 13093 25823
rect 12667 25792 13093 25820
rect 12667 25789 12679 25792
rect 12621 25783 12679 25789
rect 13081 25789 13093 25792
rect 13127 25789 13139 25823
rect 13081 25783 13139 25789
rect 14108 25752 14136 25928
rect 20809 25959 20867 25965
rect 20809 25925 20821 25959
rect 20855 25956 20867 25959
rect 21818 25956 21824 25968
rect 20855 25928 21824 25956
rect 20855 25925 20867 25928
rect 20809 25919 20867 25925
rect 21818 25916 21824 25928
rect 21876 25916 21882 25968
rect 22278 25956 22284 25968
rect 22239 25928 22284 25956
rect 22278 25916 22284 25928
rect 22336 25916 22342 25968
rect 24670 25916 24676 25968
rect 24728 25956 24734 25968
rect 25222 25956 25228 25968
rect 24728 25928 25228 25956
rect 24728 25916 24734 25928
rect 25222 25916 25228 25928
rect 25280 25956 25286 25968
rect 26329 25959 26387 25965
rect 26329 25956 26341 25959
rect 25280 25928 26341 25956
rect 25280 25916 25286 25928
rect 26329 25925 26341 25928
rect 26375 25956 26387 25959
rect 26602 25956 26608 25968
rect 26375 25928 26608 25956
rect 26375 25925 26387 25928
rect 26329 25919 26387 25925
rect 26602 25916 26608 25928
rect 26660 25916 26666 25968
rect 30834 25916 30840 25968
rect 30892 25956 30898 25968
rect 30892 25928 31616 25956
rect 30892 25916 30898 25928
rect 31588 25900 31616 25928
rect 32030 25916 32036 25968
rect 32088 25956 32094 25968
rect 32217 25959 32275 25965
rect 32217 25956 32229 25959
rect 32088 25928 32229 25956
rect 32088 25916 32094 25928
rect 32217 25925 32229 25928
rect 32263 25956 32275 25959
rect 32306 25956 32312 25968
rect 32263 25928 32312 25956
rect 32263 25925 32275 25928
rect 32217 25919 32275 25925
rect 32306 25916 32312 25928
rect 32364 25916 32370 25968
rect 33134 25916 33140 25968
rect 33192 25956 33198 25968
rect 34149 25959 34207 25965
rect 34149 25956 34161 25959
rect 33192 25928 34161 25956
rect 33192 25916 33198 25928
rect 34149 25925 34161 25928
rect 34195 25925 34207 25959
rect 38562 25956 38568 25968
rect 38523 25928 38568 25956
rect 34149 25919 34207 25925
rect 38562 25916 38568 25928
rect 38620 25916 38626 25968
rect 42242 25956 42248 25968
rect 42203 25928 42248 25956
rect 42242 25916 42248 25928
rect 42300 25916 42306 25968
rect 14277 25891 14335 25897
rect 14277 25857 14289 25891
rect 14323 25888 14335 25891
rect 14550 25888 14556 25900
rect 14323 25860 14556 25888
rect 14323 25857 14335 25860
rect 14277 25851 14335 25857
rect 14550 25848 14556 25860
rect 14608 25848 14614 25900
rect 19889 25891 19947 25897
rect 19889 25857 19901 25891
rect 19935 25888 19947 25891
rect 19978 25888 19984 25900
rect 19935 25860 19984 25888
rect 19935 25857 19947 25860
rect 19889 25851 19947 25857
rect 19978 25848 19984 25860
rect 20036 25848 20042 25900
rect 21726 25848 21732 25900
rect 21784 25888 21790 25900
rect 24489 25891 24547 25897
rect 24489 25888 24501 25891
rect 21784 25860 24501 25888
rect 21784 25848 21790 25860
rect 24489 25857 24501 25860
rect 24535 25857 24547 25891
rect 24489 25851 24547 25857
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25888 26019 25891
rect 26007 25860 26832 25888
rect 26007 25857 26019 25860
rect 25961 25851 26019 25857
rect 26804 25832 26832 25860
rect 27338 25848 27344 25900
rect 27396 25888 27402 25900
rect 27433 25891 27491 25897
rect 27433 25888 27445 25891
rect 27396 25860 27445 25888
rect 27396 25848 27402 25860
rect 27433 25857 27445 25860
rect 27479 25857 27491 25891
rect 31294 25888 31300 25900
rect 31255 25860 31300 25888
rect 27433 25851 27491 25857
rect 31294 25848 31300 25860
rect 31352 25848 31358 25900
rect 31570 25888 31576 25900
rect 31483 25860 31576 25888
rect 31570 25848 31576 25860
rect 31628 25888 31634 25900
rect 33686 25888 33692 25900
rect 31628 25860 33692 25888
rect 31628 25848 31634 25860
rect 33686 25848 33692 25860
rect 33744 25848 33750 25900
rect 35805 25891 35863 25897
rect 35805 25857 35817 25891
rect 35851 25888 35863 25891
rect 37826 25888 37832 25900
rect 35851 25860 37832 25888
rect 35851 25857 35863 25860
rect 35805 25851 35863 25857
rect 16945 25823 17003 25829
rect 16945 25789 16957 25823
rect 16991 25789 17003 25823
rect 16945 25783 17003 25789
rect 14598 25755 14656 25761
rect 14598 25752 14610 25755
rect 14108 25724 14610 25752
rect 14598 25721 14610 25724
rect 14644 25752 14656 25755
rect 14734 25752 14740 25764
rect 14644 25724 14740 25752
rect 14644 25721 14656 25724
rect 14598 25715 14656 25721
rect 14734 25712 14740 25724
rect 14792 25712 14798 25764
rect 16960 25752 16988 25783
rect 17310 25780 17316 25832
rect 17368 25820 17374 25832
rect 18046 25820 18052 25832
rect 17368 25792 18052 25820
rect 17368 25780 17374 25792
rect 18046 25780 18052 25792
rect 18104 25820 18110 25832
rect 18141 25823 18199 25829
rect 18141 25820 18153 25823
rect 18104 25792 18153 25820
rect 18104 25780 18110 25792
rect 18141 25789 18153 25792
rect 18187 25789 18199 25823
rect 26602 25820 26608 25832
rect 26563 25792 26608 25820
rect 18141 25783 18199 25789
rect 26602 25780 26608 25792
rect 26660 25780 26666 25832
rect 26786 25780 26792 25832
rect 26844 25820 26850 25832
rect 26973 25823 27031 25829
rect 26973 25820 26985 25823
rect 26844 25792 26985 25820
rect 26844 25780 26850 25792
rect 26973 25789 26985 25792
rect 27019 25820 27031 25823
rect 28258 25820 28264 25832
rect 27019 25792 28264 25820
rect 27019 25789 27031 25792
rect 26973 25783 27031 25789
rect 28258 25780 28264 25792
rect 28316 25780 28322 25832
rect 28350 25780 28356 25832
rect 28408 25820 28414 25832
rect 30260 25823 30318 25829
rect 30260 25820 30272 25823
rect 28408 25792 30272 25820
rect 28408 25780 28414 25792
rect 30260 25789 30272 25792
rect 30306 25820 30318 25823
rect 30745 25823 30803 25829
rect 30745 25820 30757 25823
rect 30306 25792 30757 25820
rect 30306 25789 30318 25792
rect 30260 25783 30318 25789
rect 30745 25789 30757 25792
rect 30791 25820 30803 25823
rect 31018 25820 31024 25832
rect 30791 25792 31024 25820
rect 30791 25789 30803 25792
rect 30745 25783 30803 25789
rect 31018 25780 31024 25792
rect 31076 25780 31082 25832
rect 34054 25780 34060 25832
rect 34112 25820 34118 25832
rect 34952 25823 35010 25829
rect 34952 25820 34964 25823
rect 34112 25792 34964 25820
rect 34112 25780 34118 25792
rect 34952 25789 34964 25792
rect 34998 25820 35010 25823
rect 35820 25820 35848 25851
rect 37826 25848 37832 25860
rect 37884 25848 37890 25900
rect 38013 25891 38071 25897
rect 38013 25857 38025 25891
rect 38059 25888 38071 25891
rect 38378 25888 38384 25900
rect 38059 25860 38384 25888
rect 38059 25857 38071 25860
rect 38013 25851 38071 25857
rect 38378 25848 38384 25860
rect 38436 25848 38442 25900
rect 38470 25848 38476 25900
rect 38528 25888 38534 25900
rect 39025 25891 39083 25897
rect 39025 25888 39037 25891
rect 38528 25860 39037 25888
rect 38528 25848 38534 25860
rect 39025 25857 39037 25860
rect 39071 25888 39083 25891
rect 44315 25891 44373 25897
rect 44315 25888 44327 25891
rect 39071 25860 44327 25888
rect 39071 25857 39083 25860
rect 39025 25851 39083 25857
rect 44315 25857 44327 25860
rect 44361 25857 44373 25891
rect 44315 25851 44373 25857
rect 36078 25820 36084 25832
rect 34998 25792 35848 25820
rect 36039 25792 36084 25820
rect 34998 25789 35010 25792
rect 34952 25783 35010 25789
rect 36078 25780 36084 25792
rect 36136 25780 36142 25832
rect 40564 25823 40622 25829
rect 40564 25789 40576 25823
rect 40610 25820 40622 25823
rect 40954 25820 40960 25832
rect 40610 25792 40960 25820
rect 40610 25789 40622 25792
rect 40564 25783 40622 25789
rect 40954 25780 40960 25792
rect 41012 25780 41018 25832
rect 42702 25780 42708 25832
rect 42760 25820 42766 25832
rect 43232 25823 43290 25829
rect 43232 25820 43244 25823
rect 42760 25792 43244 25820
rect 42760 25780 42766 25792
rect 43232 25789 43244 25792
rect 43278 25820 43290 25823
rect 43625 25823 43683 25829
rect 43625 25820 43637 25823
rect 43278 25792 43637 25820
rect 43278 25789 43290 25792
rect 43232 25783 43290 25789
rect 43625 25789 43637 25792
rect 43671 25789 43683 25823
rect 43625 25783 43683 25789
rect 44228 25823 44286 25829
rect 44228 25789 44240 25823
rect 44274 25820 44286 25823
rect 44634 25820 44640 25832
rect 44274 25792 44640 25820
rect 44274 25789 44286 25792
rect 44228 25783 44286 25789
rect 44634 25780 44640 25792
rect 44692 25780 44698 25832
rect 19797 25755 19855 25761
rect 16960 25724 17908 25752
rect 11882 25684 11888 25696
rect 9916 25656 11376 25684
rect 11843 25656 11888 25684
rect 9916 25644 9922 25656
rect 11882 25644 11888 25656
rect 11940 25644 11946 25696
rect 12250 25684 12256 25696
rect 12211 25656 12256 25684
rect 12250 25644 12256 25656
rect 12308 25644 12314 25696
rect 12805 25687 12863 25693
rect 12805 25653 12817 25687
rect 12851 25684 12863 25687
rect 13170 25684 13176 25696
rect 12851 25656 13176 25684
rect 12851 25653 12863 25656
rect 12805 25647 12863 25653
rect 13170 25644 13176 25656
rect 13228 25644 13234 25696
rect 17126 25684 17132 25696
rect 17087 25656 17132 25684
rect 17126 25644 17132 25656
rect 17184 25644 17190 25696
rect 17880 25693 17908 25724
rect 19797 25721 19809 25755
rect 19843 25752 19855 25755
rect 20251 25755 20309 25761
rect 20251 25752 20263 25755
rect 19843 25724 20263 25752
rect 19843 25721 19855 25724
rect 19797 25715 19855 25721
rect 20251 25721 20263 25724
rect 20297 25752 20309 25755
rect 21174 25752 21180 25764
rect 20297 25724 21180 25752
rect 20297 25721 20309 25724
rect 20251 25715 20309 25721
rect 21174 25712 21180 25724
rect 21232 25712 21238 25764
rect 21726 25752 21732 25764
rect 21687 25724 21732 25752
rect 21726 25712 21732 25724
rect 21784 25712 21790 25764
rect 21818 25712 21824 25764
rect 21876 25752 21882 25764
rect 24210 25752 24216 25764
rect 21876 25724 21921 25752
rect 24171 25724 24216 25752
rect 21876 25712 21882 25724
rect 24210 25712 24216 25724
rect 24268 25712 24274 25764
rect 24305 25755 24363 25761
rect 24305 25721 24317 25755
rect 24351 25752 24363 25755
rect 24486 25752 24492 25764
rect 24351 25724 24492 25752
rect 24351 25721 24363 25724
rect 24305 25715 24363 25721
rect 24486 25712 24492 25724
rect 24544 25712 24550 25764
rect 27154 25752 27160 25764
rect 27115 25724 27160 25752
rect 27154 25712 27160 25724
rect 27212 25712 27218 25764
rect 31389 25755 31447 25761
rect 31389 25721 31401 25755
rect 31435 25752 31447 25755
rect 32585 25755 32643 25761
rect 32585 25752 32597 25755
rect 31435 25724 32597 25752
rect 31435 25721 31447 25724
rect 31389 25715 31447 25721
rect 32585 25721 32597 25724
rect 32631 25721 32643 25755
rect 32858 25752 32864 25764
rect 32819 25724 32864 25752
rect 32585 25715 32643 25721
rect 17865 25687 17923 25693
rect 17865 25653 17877 25687
rect 17911 25684 17923 25687
rect 18874 25684 18880 25696
rect 17911 25656 18880 25684
rect 17911 25653 17923 25656
rect 17865 25647 17923 25653
rect 18874 25644 18880 25656
rect 18932 25644 18938 25696
rect 22922 25644 22928 25696
rect 22980 25684 22986 25696
rect 24026 25684 24032 25696
rect 22980 25656 24032 25684
rect 22980 25644 22986 25656
rect 24026 25644 24032 25656
rect 24084 25644 24090 25696
rect 27982 25684 27988 25696
rect 27943 25656 27988 25684
rect 27982 25644 27988 25656
rect 28040 25644 28046 25696
rect 29086 25684 29092 25696
rect 28999 25656 29092 25684
rect 29086 25644 29092 25656
rect 29144 25684 29150 25696
rect 29638 25684 29644 25696
rect 29144 25656 29644 25684
rect 29144 25644 29150 25656
rect 29638 25644 29644 25656
rect 29696 25644 29702 25696
rect 30331 25687 30389 25693
rect 30331 25653 30343 25687
rect 30377 25684 30389 25687
rect 30650 25684 30656 25696
rect 30377 25656 30656 25684
rect 30377 25653 30389 25656
rect 30331 25647 30389 25653
rect 30650 25644 30656 25656
rect 30708 25644 30714 25696
rect 30742 25644 30748 25696
rect 30800 25684 30806 25696
rect 31021 25687 31079 25693
rect 31021 25684 31033 25687
rect 30800 25656 31033 25684
rect 30800 25644 30806 25656
rect 31021 25653 31033 25656
rect 31067 25653 31079 25687
rect 31021 25647 31079 25653
rect 31202 25644 31208 25696
rect 31260 25684 31266 25696
rect 31404 25684 31432 25715
rect 31260 25656 31432 25684
rect 32600 25684 32628 25715
rect 32858 25712 32864 25724
rect 32916 25712 32922 25764
rect 32953 25755 33011 25761
rect 32953 25721 32965 25755
rect 32999 25721 33011 25755
rect 32953 25715 33011 25721
rect 32968 25684 32996 25715
rect 33134 25712 33140 25764
rect 33192 25752 33198 25764
rect 33505 25755 33563 25761
rect 33505 25752 33517 25755
rect 33192 25724 33517 25752
rect 33192 25712 33198 25724
rect 33505 25721 33517 25724
rect 33551 25752 33563 25755
rect 33870 25752 33876 25764
rect 33551 25724 33876 25752
rect 33551 25721 33563 25724
rect 33505 25715 33563 25721
rect 33870 25712 33876 25724
rect 33928 25752 33934 25764
rect 35158 25752 35164 25764
rect 33928 25724 35164 25752
rect 33928 25712 33934 25724
rect 35158 25712 35164 25724
rect 35216 25712 35222 25764
rect 36170 25712 36176 25764
rect 36228 25752 36234 25764
rect 36443 25755 36501 25761
rect 36443 25752 36455 25755
rect 36228 25724 36455 25752
rect 36228 25712 36234 25724
rect 36443 25721 36455 25724
rect 36489 25752 36501 25755
rect 36489 25724 37412 25752
rect 36489 25721 36501 25724
rect 36443 25715 36501 25721
rect 37384 25696 37412 25724
rect 37734 25712 37740 25764
rect 37792 25752 37798 25764
rect 38105 25755 38163 25761
rect 38105 25752 38117 25755
rect 37792 25724 38117 25752
rect 37792 25712 37798 25724
rect 38105 25721 38117 25724
rect 38151 25752 38163 25755
rect 41417 25755 41475 25761
rect 41417 25752 41429 25755
rect 38151 25724 41429 25752
rect 38151 25721 38163 25724
rect 38105 25715 38163 25721
rect 41417 25721 41429 25724
rect 41463 25721 41475 25755
rect 41690 25752 41696 25764
rect 41651 25724 41696 25752
rect 41417 25715 41475 25721
rect 32600 25656 32996 25684
rect 31260 25644 31266 25656
rect 34698 25644 34704 25696
rect 34756 25684 34762 25696
rect 35023 25687 35081 25693
rect 35023 25684 35035 25687
rect 34756 25656 35035 25684
rect 34756 25644 34762 25656
rect 35023 25653 35035 25656
rect 35069 25653 35081 25687
rect 36998 25684 37004 25696
rect 36959 25656 37004 25684
rect 35023 25647 35081 25653
rect 36998 25644 37004 25656
rect 37056 25644 37062 25696
rect 37366 25684 37372 25696
rect 37327 25656 37372 25684
rect 37366 25644 37372 25656
rect 37424 25644 37430 25696
rect 39577 25687 39635 25693
rect 39577 25653 39589 25687
rect 39623 25684 39635 25687
rect 39758 25684 39764 25696
rect 39623 25656 39764 25684
rect 39623 25653 39635 25656
rect 39577 25647 39635 25653
rect 39758 25644 39764 25656
rect 39816 25644 39822 25696
rect 40635 25687 40693 25693
rect 40635 25653 40647 25687
rect 40681 25684 40693 25687
rect 40770 25684 40776 25696
rect 40681 25656 40776 25684
rect 40681 25653 40693 25656
rect 40635 25647 40693 25653
rect 40770 25644 40776 25656
rect 40828 25644 40834 25696
rect 41432 25684 41460 25715
rect 41690 25712 41696 25724
rect 41748 25712 41754 25764
rect 41785 25755 41843 25761
rect 41785 25721 41797 25755
rect 41831 25752 41843 25755
rect 41874 25752 41880 25764
rect 41831 25724 41880 25752
rect 41831 25721 41843 25724
rect 41785 25715 41843 25721
rect 41598 25684 41604 25696
rect 41432 25656 41604 25684
rect 41598 25644 41604 25656
rect 41656 25684 41662 25696
rect 41800 25684 41828 25715
rect 41874 25712 41880 25724
rect 41932 25712 41938 25764
rect 43530 25752 43536 25764
rect 42766 25724 43536 25752
rect 42766 25684 42794 25724
rect 43530 25712 43536 25724
rect 43588 25752 43594 25764
rect 43993 25755 44051 25761
rect 43993 25752 44005 25755
rect 43588 25724 44005 25752
rect 43588 25712 43594 25724
rect 43993 25721 44005 25724
rect 44039 25721 44051 25755
rect 43993 25715 44051 25721
rect 41656 25656 42794 25684
rect 41656 25644 41662 25656
rect 43070 25644 43076 25696
rect 43128 25684 43134 25696
rect 43303 25687 43361 25693
rect 43303 25684 43315 25687
rect 43128 25656 43315 25684
rect 43128 25644 43134 25656
rect 43303 25653 43315 25656
rect 43349 25653 43361 25687
rect 43303 25647 43361 25653
rect 1104 25594 48852 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 48852 25594
rect 1104 25520 48852 25542
rect 4338 25480 4344 25492
rect 4299 25452 4344 25480
rect 4338 25440 4344 25452
rect 4396 25440 4402 25492
rect 6549 25483 6607 25489
rect 6549 25449 6561 25483
rect 6595 25480 6607 25483
rect 6914 25480 6920 25492
rect 6595 25452 6920 25480
rect 6595 25449 6607 25452
rect 6549 25443 6607 25449
rect 6914 25440 6920 25452
rect 6972 25440 6978 25492
rect 7377 25483 7435 25489
rect 7377 25449 7389 25483
rect 7423 25480 7435 25483
rect 7466 25480 7472 25492
rect 7423 25452 7472 25480
rect 7423 25449 7435 25452
rect 7377 25443 7435 25449
rect 7466 25440 7472 25452
rect 7524 25480 7530 25492
rect 8754 25480 8760 25492
rect 7524 25452 8760 25480
rect 7524 25440 7530 25452
rect 8754 25440 8760 25452
rect 8812 25440 8818 25492
rect 10226 25440 10232 25492
rect 10284 25480 10290 25492
rect 10689 25483 10747 25489
rect 10689 25480 10701 25483
rect 10284 25452 10701 25480
rect 10284 25440 10290 25452
rect 10689 25449 10701 25452
rect 10735 25449 10747 25483
rect 10689 25443 10747 25449
rect 11882 25440 11888 25492
rect 11940 25480 11946 25492
rect 16669 25483 16727 25489
rect 16669 25480 16681 25483
rect 11940 25452 16681 25480
rect 11940 25440 11946 25452
rect 16669 25449 16681 25452
rect 16715 25449 16727 25483
rect 17678 25480 17684 25492
rect 17639 25452 17684 25480
rect 16669 25443 16727 25449
rect 17678 25440 17684 25452
rect 17736 25440 17742 25492
rect 18046 25480 18052 25492
rect 18007 25452 18052 25480
rect 18046 25440 18052 25452
rect 18104 25440 18110 25492
rect 21174 25440 21180 25492
rect 21232 25480 21238 25492
rect 21269 25483 21327 25489
rect 21269 25480 21281 25483
rect 21232 25452 21281 25480
rect 21232 25440 21238 25452
rect 21269 25449 21281 25452
rect 21315 25449 21327 25483
rect 24210 25480 24216 25492
rect 24171 25452 24216 25480
rect 21269 25443 21327 25449
rect 24210 25440 24216 25452
rect 24268 25440 24274 25492
rect 27154 25480 27160 25492
rect 27115 25452 27160 25480
rect 27154 25440 27160 25452
rect 27212 25440 27218 25492
rect 28169 25483 28227 25489
rect 28169 25449 28181 25483
rect 28215 25480 28227 25483
rect 28215 25452 29224 25480
rect 28215 25449 28227 25452
rect 28169 25443 28227 25449
rect 3878 25372 3884 25424
rect 3936 25412 3942 25424
rect 5445 25415 5503 25421
rect 3936 25384 4292 25412
rect 3936 25372 3942 25384
rect 1949 25347 2007 25353
rect 1949 25313 1961 25347
rect 1995 25344 2007 25347
rect 2222 25344 2228 25356
rect 1995 25316 2228 25344
rect 1995 25313 2007 25316
rect 1949 25307 2007 25313
rect 2222 25304 2228 25316
rect 2280 25304 2286 25356
rect 2958 25344 2964 25356
rect 2919 25316 2964 25344
rect 2958 25304 2964 25316
rect 3016 25304 3022 25356
rect 4264 25353 4292 25384
rect 5445 25381 5457 25415
rect 5491 25412 5503 25415
rect 5994 25412 6000 25424
rect 5491 25384 5764 25412
rect 5955 25384 6000 25412
rect 5491 25381 5503 25384
rect 5445 25375 5503 25381
rect 4065 25347 4123 25353
rect 4065 25313 4077 25347
rect 4111 25313 4123 25347
rect 4065 25307 4123 25313
rect 4249 25347 4307 25353
rect 4249 25313 4261 25347
rect 4295 25313 4307 25347
rect 4249 25307 4307 25313
rect 4080 25276 4108 25307
rect 4264 25276 4292 25307
rect 5534 25304 5540 25356
rect 5592 25344 5598 25356
rect 5629 25347 5687 25353
rect 5629 25344 5641 25347
rect 5592 25316 5641 25344
rect 5592 25304 5598 25316
rect 5629 25313 5641 25316
rect 5675 25313 5687 25347
rect 5736 25344 5764 25384
rect 5994 25372 6000 25384
rect 6052 25372 6058 25424
rect 6822 25412 6828 25424
rect 6783 25384 6828 25412
rect 6822 25372 6828 25384
rect 6880 25372 6886 25424
rect 8205 25415 8263 25421
rect 8205 25381 8217 25415
rect 8251 25412 8263 25415
rect 8294 25412 8300 25424
rect 8251 25384 8300 25412
rect 8251 25381 8263 25384
rect 8205 25375 8263 25381
rect 8294 25372 8300 25384
rect 8352 25372 8358 25424
rect 10410 25412 10416 25424
rect 10371 25384 10416 25412
rect 10410 25372 10416 25384
rect 10468 25372 10474 25424
rect 12342 25412 12348 25424
rect 12303 25384 12348 25412
rect 12342 25372 12348 25384
rect 12400 25372 12406 25424
rect 12710 25372 12716 25424
rect 12768 25412 12774 25424
rect 14185 25415 14243 25421
rect 12768 25384 13814 25412
rect 12768 25372 12774 25384
rect 6362 25344 6368 25356
rect 5736 25316 6368 25344
rect 5629 25307 5687 25313
rect 6362 25304 6368 25316
rect 6420 25304 6426 25356
rect 7650 25344 7656 25356
rect 7611 25316 7656 25344
rect 7650 25304 7656 25316
rect 7708 25304 7714 25356
rect 8021 25347 8079 25353
rect 8021 25313 8033 25347
rect 8067 25313 8079 25347
rect 9950 25344 9956 25356
rect 9911 25316 9956 25344
rect 8021 25307 8079 25313
rect 5552 25276 5580 25304
rect 4080 25248 4154 25276
rect 4264 25248 5580 25276
rect 2130 25140 2136 25152
rect 2091 25112 2136 25140
rect 2130 25100 2136 25112
rect 2188 25100 2194 25152
rect 3145 25143 3203 25149
rect 3145 25109 3157 25143
rect 3191 25140 3203 25143
rect 3234 25140 3240 25152
rect 3191 25112 3240 25140
rect 3191 25109 3203 25112
rect 3145 25103 3203 25109
rect 3234 25100 3240 25112
rect 3292 25100 3298 25152
rect 4126 25140 4154 25248
rect 6730 25236 6736 25288
rect 6788 25276 6794 25288
rect 8036 25276 8064 25307
rect 9950 25304 9956 25316
rect 10008 25304 10014 25356
rect 10229 25347 10287 25353
rect 10229 25313 10241 25347
rect 10275 25313 10287 25347
rect 11790 25344 11796 25356
rect 11751 25316 11796 25344
rect 10229 25307 10287 25313
rect 9493 25279 9551 25285
rect 9493 25276 9505 25279
rect 6788 25248 9505 25276
rect 6788 25236 6794 25248
rect 9493 25245 9505 25248
rect 9539 25276 9551 25279
rect 10244 25276 10272 25307
rect 11790 25304 11796 25316
rect 11848 25304 11854 25356
rect 11974 25344 11980 25356
rect 11935 25316 11980 25344
rect 11974 25304 11980 25316
rect 12032 25304 12038 25356
rect 13538 25344 13544 25356
rect 13499 25316 13544 25344
rect 13538 25304 13544 25316
rect 13596 25304 13602 25356
rect 13786 25344 13814 25384
rect 14185 25381 14197 25415
rect 14231 25412 14243 25415
rect 14550 25412 14556 25424
rect 14231 25384 14556 25412
rect 14231 25381 14243 25384
rect 14185 25375 14243 25381
rect 14550 25372 14556 25384
rect 14608 25372 14614 25424
rect 19978 25412 19984 25424
rect 19939 25384 19984 25412
rect 19978 25372 19984 25384
rect 20036 25372 20042 25424
rect 24026 25372 24032 25424
rect 24084 25412 24090 25424
rect 24302 25412 24308 25424
rect 24084 25384 24308 25412
rect 24084 25372 24090 25384
rect 24302 25372 24308 25384
rect 24360 25372 24366 25424
rect 24486 25372 24492 25424
rect 24544 25412 24550 25424
rect 24765 25415 24823 25421
rect 24765 25412 24777 25415
rect 24544 25384 24777 25412
rect 24544 25372 24550 25384
rect 24765 25381 24777 25384
rect 24811 25381 24823 25415
rect 24765 25375 24823 25381
rect 14001 25347 14059 25353
rect 14001 25344 14013 25347
rect 13786 25316 14013 25344
rect 14001 25313 14013 25316
rect 14047 25344 14059 25347
rect 14458 25344 14464 25356
rect 14047 25316 14464 25344
rect 14047 25313 14059 25316
rect 14001 25307 14059 25313
rect 14458 25304 14464 25316
rect 14516 25344 14522 25356
rect 14826 25344 14832 25356
rect 14516 25316 14832 25344
rect 14516 25304 14522 25316
rect 14826 25304 14832 25316
rect 14884 25304 14890 25356
rect 15286 25344 15292 25356
rect 15247 25316 15292 25344
rect 15286 25304 15292 25316
rect 15344 25304 15350 25356
rect 16482 25344 16488 25356
rect 16443 25316 16488 25344
rect 16482 25304 16488 25316
rect 16540 25304 16546 25356
rect 17494 25344 17500 25356
rect 17455 25316 17500 25344
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 19426 25344 19432 25356
rect 19387 25316 19432 25344
rect 19426 25304 19432 25316
rect 19484 25304 19490 25356
rect 19797 25347 19855 25353
rect 19797 25313 19809 25347
rect 19843 25344 19855 25347
rect 20346 25344 20352 25356
rect 19843 25316 20352 25344
rect 19843 25313 19855 25316
rect 19797 25307 19855 25313
rect 20346 25304 20352 25316
rect 20404 25304 20410 25356
rect 23477 25347 23535 25353
rect 23477 25313 23489 25347
rect 23523 25344 23535 25347
rect 23566 25344 23572 25356
rect 23523 25316 23572 25344
rect 23523 25313 23535 25316
rect 23477 25307 23535 25313
rect 23566 25304 23572 25316
rect 23624 25304 23630 25356
rect 27172 25344 27200 25440
rect 29196 25424 29224 25452
rect 30650 25440 30656 25492
rect 30708 25480 30714 25492
rect 32490 25480 32496 25492
rect 30708 25452 32496 25480
rect 30708 25440 30714 25452
rect 32490 25440 32496 25452
rect 32548 25480 32554 25492
rect 33137 25483 33195 25489
rect 33137 25480 33149 25483
rect 32548 25452 33149 25480
rect 32548 25440 32554 25452
rect 33137 25449 33149 25452
rect 33183 25449 33195 25483
rect 33137 25443 33195 25449
rect 36078 25440 36084 25492
rect 36136 25480 36142 25492
rect 36909 25483 36967 25489
rect 36909 25480 36921 25483
rect 36136 25452 36921 25480
rect 36136 25440 36142 25452
rect 36909 25449 36921 25452
rect 36955 25449 36967 25483
rect 38378 25480 38384 25492
rect 38339 25452 38384 25480
rect 36909 25443 36967 25449
rect 38378 25440 38384 25452
rect 38436 25440 38442 25492
rect 41598 25480 41604 25492
rect 41559 25452 41604 25480
rect 41598 25440 41604 25452
rect 41656 25440 41662 25492
rect 41690 25440 41696 25492
rect 41748 25480 41754 25492
rect 41969 25483 42027 25489
rect 41969 25480 41981 25483
rect 41748 25452 41981 25480
rect 41748 25440 41754 25452
rect 41969 25449 41981 25452
rect 42015 25480 42027 25483
rect 43070 25480 43076 25492
rect 42015 25452 43076 25480
rect 42015 25449 42027 25452
rect 41969 25443 42027 25449
rect 43070 25440 43076 25452
rect 43128 25440 43134 25492
rect 44542 25480 44548 25492
rect 44503 25452 44548 25480
rect 44542 25440 44548 25452
rect 44600 25440 44606 25492
rect 27338 25372 27344 25424
rect 27396 25412 27402 25424
rect 27570 25415 27628 25421
rect 27570 25412 27582 25415
rect 27396 25384 27582 25412
rect 27396 25372 27402 25384
rect 27570 25381 27582 25384
rect 27616 25381 27628 25415
rect 27570 25375 27628 25381
rect 27982 25372 27988 25424
rect 28040 25412 28046 25424
rect 29086 25412 29092 25424
rect 28040 25384 29092 25412
rect 28040 25372 28046 25384
rect 29086 25372 29092 25384
rect 29144 25372 29150 25424
rect 29178 25372 29184 25424
rect 29236 25412 29242 25424
rect 33410 25412 33416 25424
rect 29236 25384 29281 25412
rect 33371 25384 33416 25412
rect 29236 25372 29242 25384
rect 33410 25372 33416 25384
rect 33468 25372 33474 25424
rect 33505 25415 33563 25421
rect 33505 25381 33517 25415
rect 33551 25412 33563 25415
rect 35069 25415 35127 25421
rect 35069 25412 35081 25415
rect 33551 25384 35081 25412
rect 33551 25381 33563 25384
rect 33505 25375 33563 25381
rect 35069 25381 35081 25384
rect 35115 25412 35127 25415
rect 35250 25412 35256 25424
rect 35115 25384 35256 25412
rect 35115 25381 35127 25384
rect 35069 25375 35127 25381
rect 35250 25372 35256 25384
rect 35308 25372 35314 25424
rect 36170 25412 36176 25424
rect 36131 25384 36176 25412
rect 36170 25372 36176 25384
rect 36228 25372 36234 25424
rect 36998 25372 37004 25424
rect 37056 25412 37062 25424
rect 38013 25415 38071 25421
rect 38013 25412 38025 25415
rect 37056 25384 38025 25412
rect 37056 25372 37062 25384
rect 38013 25381 38025 25384
rect 38059 25412 38071 25415
rect 39758 25412 39764 25424
rect 38059 25384 39764 25412
rect 38059 25381 38071 25384
rect 38013 25375 38071 25381
rect 39758 25372 39764 25384
rect 39816 25372 39822 25424
rect 40310 25412 40316 25424
rect 40271 25384 40316 25412
rect 40310 25372 40316 25384
rect 40368 25372 40374 25424
rect 43487 25415 43545 25421
rect 43487 25412 43499 25415
rect 40563 25384 43499 25412
rect 27249 25347 27307 25353
rect 27249 25344 27261 25347
rect 27172 25316 27261 25344
rect 27249 25313 27261 25316
rect 27295 25313 27307 25347
rect 30650 25344 30656 25356
rect 30611 25316 30656 25344
rect 27249 25307 27307 25313
rect 30650 25304 30656 25316
rect 30708 25304 30714 25356
rect 31754 25304 31760 25356
rect 31812 25344 31818 25356
rect 32122 25344 32128 25356
rect 32180 25353 32186 25356
rect 32180 25347 32218 25353
rect 31812 25316 32128 25344
rect 31812 25304 31818 25316
rect 32122 25304 32128 25316
rect 32206 25313 32218 25347
rect 32180 25307 32218 25313
rect 38565 25347 38623 25353
rect 38565 25313 38577 25347
rect 38611 25344 38623 25347
rect 38838 25344 38844 25356
rect 38611 25316 38844 25344
rect 38611 25313 38623 25316
rect 38565 25307 38623 25313
rect 32180 25304 32186 25307
rect 38838 25304 38844 25316
rect 38896 25304 38902 25356
rect 17126 25276 17132 25288
rect 9539 25248 17132 25276
rect 9539 25245 9551 25248
rect 9493 25239 9551 25245
rect 17126 25236 17132 25248
rect 17184 25236 17190 25288
rect 20254 25236 20260 25288
rect 20312 25276 20318 25288
rect 20901 25279 20959 25285
rect 20901 25276 20913 25279
rect 20312 25248 20913 25276
rect 20312 25236 20318 25248
rect 20901 25245 20913 25248
rect 20947 25276 20959 25279
rect 22094 25276 22100 25288
rect 20947 25248 22100 25276
rect 20947 25245 20959 25248
rect 20901 25239 20959 25245
rect 22094 25236 22100 25248
rect 22152 25236 22158 25288
rect 23707 25279 23765 25285
rect 23707 25245 23719 25279
rect 23753 25276 23765 25279
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 23753 25248 24685 25276
rect 23753 25245 23765 25248
rect 23707 25239 23765 25245
rect 24673 25245 24685 25248
rect 24719 25276 24731 25279
rect 25038 25276 25044 25288
rect 24719 25248 25044 25276
rect 24719 25245 24731 25248
rect 24673 25239 24731 25245
rect 25038 25236 25044 25248
rect 25096 25236 25102 25288
rect 30883 25279 30941 25285
rect 30883 25245 30895 25279
rect 30929 25276 30941 25279
rect 32769 25279 32827 25285
rect 32769 25276 32781 25279
rect 30929 25248 32781 25276
rect 30929 25245 30941 25248
rect 30883 25239 30941 25245
rect 32769 25245 32781 25248
rect 32815 25276 32827 25279
rect 32858 25276 32864 25288
rect 32815 25248 32864 25276
rect 32815 25245 32827 25248
rect 32769 25239 32827 25245
rect 32858 25236 32864 25248
rect 32916 25236 32922 25288
rect 33686 25276 33692 25288
rect 33647 25248 33692 25276
rect 33686 25236 33692 25248
rect 33744 25236 33750 25288
rect 34698 25236 34704 25288
rect 34756 25276 34762 25288
rect 34977 25279 35035 25285
rect 34977 25276 34989 25279
rect 34756 25248 34989 25276
rect 34756 25236 34762 25248
rect 34977 25245 34989 25248
rect 35023 25245 35035 25279
rect 34977 25239 35035 25245
rect 35158 25236 35164 25288
rect 35216 25276 35222 25288
rect 35253 25279 35311 25285
rect 35253 25276 35265 25279
rect 35216 25248 35265 25276
rect 35216 25236 35222 25248
rect 35253 25245 35265 25248
rect 35299 25245 35311 25279
rect 35253 25239 35311 25245
rect 39298 25236 39304 25288
rect 39356 25276 39362 25288
rect 39669 25279 39727 25285
rect 39669 25276 39681 25279
rect 39356 25248 39681 25276
rect 39356 25236 39362 25248
rect 39669 25245 39681 25248
rect 39715 25276 39727 25279
rect 40563 25276 40591 25384
rect 43487 25381 43499 25384
rect 43533 25381 43545 25415
rect 43487 25375 43545 25381
rect 41176 25347 41234 25353
rect 41176 25344 41188 25347
rect 39715 25248 40591 25276
rect 40650 25316 41188 25344
rect 39715 25245 39727 25248
rect 39669 25239 39727 25245
rect 13722 25168 13728 25220
rect 13780 25208 13786 25220
rect 13780 25180 14596 25208
rect 13780 25168 13786 25180
rect 14568 25152 14596 25180
rect 21726 25168 21732 25220
rect 21784 25208 21790 25220
rect 22189 25211 22247 25217
rect 22189 25208 22201 25211
rect 21784 25180 22201 25208
rect 21784 25168 21790 25180
rect 22189 25177 22201 25180
rect 22235 25177 22247 25211
rect 22189 25171 22247 25177
rect 23198 25168 23204 25220
rect 23256 25208 23262 25220
rect 24854 25208 24860 25220
rect 23256 25180 24860 25208
rect 23256 25168 23262 25180
rect 24854 25168 24860 25180
rect 24912 25168 24918 25220
rect 24946 25168 24952 25220
rect 25004 25208 25010 25220
rect 25225 25211 25283 25217
rect 25225 25208 25237 25211
rect 25004 25180 25237 25208
rect 25004 25168 25010 25180
rect 25225 25177 25237 25180
rect 25271 25177 25283 25211
rect 29638 25208 29644 25220
rect 29599 25180 29644 25208
rect 25225 25171 25283 25177
rect 29638 25168 29644 25180
rect 29696 25168 29702 25220
rect 31018 25168 31024 25220
rect 31076 25208 31082 25220
rect 35802 25208 35808 25220
rect 31076 25180 32812 25208
rect 31076 25168 31082 25180
rect 32784 25152 32812 25180
rect 33106 25180 35808 25208
rect 4982 25140 4988 25152
rect 4126 25112 4988 25140
rect 4982 25100 4988 25112
rect 5040 25100 5046 25152
rect 8757 25143 8815 25149
rect 8757 25109 8769 25143
rect 8803 25140 8815 25143
rect 8938 25140 8944 25152
rect 8803 25112 8944 25140
rect 8803 25109 8815 25112
rect 8757 25103 8815 25109
rect 8938 25100 8944 25112
rect 8996 25100 9002 25152
rect 14550 25100 14556 25152
rect 14608 25140 14614 25152
rect 15473 25143 15531 25149
rect 15473 25140 15485 25143
rect 14608 25112 15485 25140
rect 14608 25100 14614 25112
rect 15473 25109 15485 25112
rect 15519 25109 15531 25143
rect 15473 25103 15531 25109
rect 21266 25100 21272 25152
rect 21324 25140 21330 25152
rect 21821 25143 21879 25149
rect 21821 25140 21833 25143
rect 21324 25112 21833 25140
rect 21324 25100 21330 25112
rect 21821 25109 21833 25112
rect 21867 25109 21879 25143
rect 28442 25140 28448 25152
rect 28403 25112 28448 25140
rect 21821 25103 21879 25109
rect 28442 25100 28448 25112
rect 28500 25100 28506 25152
rect 31202 25140 31208 25152
rect 31163 25112 31208 25140
rect 31202 25100 31208 25112
rect 31260 25100 31266 25152
rect 31662 25140 31668 25152
rect 31575 25112 31668 25140
rect 31662 25100 31668 25112
rect 31720 25140 31726 25152
rect 32263 25143 32321 25149
rect 32263 25140 32275 25143
rect 31720 25112 32275 25140
rect 31720 25100 31726 25112
rect 32263 25109 32275 25112
rect 32309 25109 32321 25143
rect 32263 25103 32321 25109
rect 32766 25100 32772 25152
rect 32824 25140 32830 25152
rect 33106 25140 33134 25180
rect 35802 25168 35808 25180
rect 35860 25168 35866 25220
rect 36354 25208 36360 25220
rect 36315 25180 36360 25208
rect 36354 25168 36360 25180
rect 36412 25208 36418 25220
rect 40650 25208 40678 25316
rect 41176 25313 41188 25316
rect 41222 25344 41234 25347
rect 41966 25344 41972 25356
rect 41222 25316 41972 25344
rect 41222 25313 41234 25316
rect 41176 25307 41234 25313
rect 41966 25304 41972 25316
rect 42024 25304 42030 25356
rect 42058 25304 42064 25356
rect 42116 25344 42122 25356
rect 42188 25347 42246 25353
rect 42188 25344 42200 25347
rect 42116 25316 42200 25344
rect 42116 25304 42122 25316
rect 42188 25313 42200 25316
rect 42234 25313 42246 25347
rect 43254 25344 43260 25356
rect 43215 25316 43260 25344
rect 42188 25307 42246 25313
rect 43254 25304 43260 25316
rect 43312 25304 43318 25356
rect 44361 25347 44419 25353
rect 44361 25313 44373 25347
rect 44407 25344 44419 25347
rect 44634 25344 44640 25356
rect 44407 25316 44640 25344
rect 44407 25313 44419 25316
rect 44361 25307 44419 25313
rect 44634 25304 44640 25316
rect 44692 25304 44698 25356
rect 42334 25276 42340 25288
rect 36412 25180 40678 25208
rect 42306 25236 42340 25276
rect 42392 25236 42398 25288
rect 36412 25168 36418 25180
rect 32824 25112 33134 25140
rect 32824 25100 32830 25112
rect 34514 25100 34520 25152
rect 34572 25140 34578 25152
rect 34701 25143 34759 25149
rect 34701 25140 34713 25143
rect 34572 25112 34713 25140
rect 34572 25100 34578 25112
rect 34701 25109 34713 25112
rect 34747 25109 34759 25143
rect 34701 25103 34759 25109
rect 36170 25100 36176 25152
rect 36228 25140 36234 25152
rect 36587 25143 36645 25149
rect 36587 25140 36599 25143
rect 36228 25112 36599 25140
rect 36228 25100 36234 25112
rect 36587 25109 36599 25112
rect 36633 25109 36645 25143
rect 36587 25103 36645 25109
rect 38749 25143 38807 25149
rect 38749 25109 38761 25143
rect 38795 25140 38807 25143
rect 39206 25140 39212 25152
rect 38795 25112 39212 25140
rect 38795 25109 38807 25112
rect 38749 25103 38807 25109
rect 39206 25100 39212 25112
rect 39264 25100 39270 25152
rect 41046 25140 41052 25152
rect 41007 25112 41052 25140
rect 41046 25100 41052 25112
rect 41104 25100 41110 25152
rect 41138 25100 41144 25152
rect 41196 25140 41202 25152
rect 42306 25149 42334 25236
rect 41279 25143 41337 25149
rect 41279 25140 41291 25143
rect 41196 25112 41291 25140
rect 41196 25100 41202 25112
rect 41279 25109 41291 25112
rect 41325 25109 41337 25143
rect 41279 25103 41337 25109
rect 42291 25143 42349 25149
rect 42291 25109 42303 25143
rect 42337 25109 42349 25143
rect 42291 25103 42349 25109
rect 1104 25050 48852 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 48852 25050
rect 1104 24976 48852 24998
rect 3878 24936 3884 24948
rect 3839 24908 3884 24936
rect 3878 24896 3884 24908
rect 3936 24896 3942 24948
rect 9769 24939 9827 24945
rect 9769 24905 9781 24939
rect 9815 24936 9827 24939
rect 9950 24936 9956 24948
rect 9815 24908 9956 24936
rect 9815 24905 9827 24908
rect 9769 24899 9827 24905
rect 9950 24896 9956 24908
rect 10008 24896 10014 24948
rect 12250 24896 12256 24948
rect 12308 24936 12314 24948
rect 13081 24939 13139 24945
rect 13081 24936 13093 24939
rect 12308 24908 13093 24936
rect 12308 24896 12314 24908
rect 13081 24905 13093 24908
rect 13127 24905 13139 24939
rect 13081 24899 13139 24905
rect 13538 24896 13544 24948
rect 13596 24936 13602 24948
rect 14001 24939 14059 24945
rect 14001 24936 14013 24939
rect 13596 24908 14013 24936
rect 13596 24896 13602 24908
rect 14001 24905 14013 24908
rect 14047 24905 14059 24939
rect 14001 24899 14059 24905
rect 15933 24939 15991 24945
rect 15933 24905 15945 24939
rect 15979 24936 15991 24939
rect 17862 24936 17868 24948
rect 15979 24908 17868 24936
rect 15979 24905 15991 24908
rect 15933 24899 15991 24905
rect 17862 24896 17868 24908
rect 17920 24896 17926 24948
rect 18233 24939 18291 24945
rect 18233 24905 18245 24939
rect 18279 24936 18291 24939
rect 19337 24939 19395 24945
rect 19337 24936 19349 24939
rect 18279 24908 19349 24936
rect 18279 24905 18291 24908
rect 18233 24899 18291 24905
rect 19337 24905 19349 24908
rect 19383 24936 19395 24939
rect 19426 24936 19432 24948
rect 19383 24908 19432 24936
rect 19383 24905 19395 24908
rect 19337 24899 19395 24905
rect 19426 24896 19432 24908
rect 19484 24896 19490 24948
rect 20993 24939 21051 24945
rect 20993 24905 21005 24939
rect 21039 24936 21051 24939
rect 21174 24936 21180 24948
rect 21039 24908 21180 24936
rect 21039 24905 21051 24908
rect 20993 24899 21051 24905
rect 21174 24896 21180 24908
rect 21232 24896 21238 24948
rect 22094 24936 22100 24948
rect 22055 24908 22100 24936
rect 22094 24896 22100 24908
rect 22152 24896 22158 24948
rect 23014 24936 23020 24948
rect 22975 24908 23020 24936
rect 23014 24896 23020 24908
rect 23072 24896 23078 24948
rect 23477 24939 23535 24945
rect 23477 24905 23489 24939
rect 23523 24936 23535 24939
rect 23566 24936 23572 24948
rect 23523 24908 23572 24936
rect 23523 24905 23535 24908
rect 23477 24899 23535 24905
rect 23566 24896 23572 24908
rect 23624 24896 23630 24948
rect 24486 24896 24492 24948
rect 24544 24936 24550 24948
rect 24673 24939 24731 24945
rect 24673 24936 24685 24939
rect 24544 24908 24685 24936
rect 24544 24896 24550 24908
rect 24673 24905 24685 24908
rect 24719 24905 24731 24939
rect 25038 24936 25044 24948
rect 24999 24908 25044 24936
rect 24673 24899 24731 24905
rect 25038 24896 25044 24908
rect 25096 24896 25102 24948
rect 26145 24939 26203 24945
rect 26145 24936 26157 24939
rect 25643 24908 26157 24936
rect 106 24828 112 24880
rect 164 24868 170 24880
rect 2133 24871 2191 24877
rect 2133 24868 2145 24871
rect 164 24840 2145 24868
rect 164 24828 170 24840
rect 2133 24837 2145 24840
rect 2179 24868 2191 24871
rect 2317 24871 2375 24877
rect 2317 24868 2329 24871
rect 2179 24840 2329 24868
rect 2179 24837 2191 24840
rect 2133 24831 2191 24837
rect 2317 24837 2329 24840
rect 2363 24837 2375 24871
rect 2317 24831 2375 24837
rect 6273 24871 6331 24877
rect 6273 24837 6285 24871
rect 6319 24868 6331 24871
rect 6362 24868 6368 24880
rect 6319 24840 6368 24868
rect 6319 24837 6331 24840
rect 6273 24831 6331 24837
rect 6362 24828 6368 24840
rect 6420 24868 6426 24880
rect 11790 24868 11796 24880
rect 6420 24840 11796 24868
rect 6420 24828 6426 24840
rect 11790 24828 11796 24840
rect 11848 24868 11854 24880
rect 11885 24871 11943 24877
rect 11885 24868 11897 24871
rect 11848 24840 11897 24868
rect 11848 24828 11854 24840
rect 11885 24837 11897 24840
rect 11931 24868 11943 24871
rect 17494 24868 17500 24880
rect 11931 24840 17500 24868
rect 11931 24837 11943 24840
rect 11885 24831 11943 24837
rect 17494 24828 17500 24840
rect 17552 24828 17558 24880
rect 1949 24803 2007 24809
rect 1949 24769 1961 24803
rect 1995 24800 2007 24803
rect 2222 24800 2228 24812
rect 1995 24772 2228 24800
rect 1995 24769 2007 24772
rect 1949 24763 2007 24769
rect 2222 24760 2228 24772
rect 2280 24800 2286 24812
rect 3513 24803 3571 24809
rect 3513 24800 3525 24803
rect 2280 24772 3525 24800
rect 2280 24760 2286 24772
rect 3513 24769 3525 24772
rect 3559 24800 3571 24803
rect 4065 24803 4123 24809
rect 4065 24800 4077 24803
rect 3559 24772 4077 24800
rect 3559 24769 3571 24772
rect 3513 24763 3571 24769
rect 4065 24769 4077 24772
rect 4111 24769 4123 24803
rect 4065 24763 4123 24769
rect 4709 24803 4767 24809
rect 4709 24769 4721 24803
rect 4755 24800 4767 24803
rect 4982 24800 4988 24812
rect 4755 24772 4988 24800
rect 4755 24769 4767 24772
rect 4709 24763 4767 24769
rect 4982 24760 4988 24772
rect 5040 24800 5046 24812
rect 7837 24803 7895 24809
rect 5040 24772 7236 24800
rect 5040 24760 5046 24772
rect 2133 24735 2191 24741
rect 2133 24701 2145 24735
rect 2179 24732 2191 24735
rect 2501 24735 2559 24741
rect 2501 24732 2513 24735
rect 2179 24704 2513 24732
rect 2179 24701 2191 24704
rect 2133 24695 2191 24701
rect 2501 24701 2513 24704
rect 2547 24732 2559 24735
rect 3602 24732 3608 24744
rect 2547 24704 3608 24732
rect 2547 24701 2559 24704
rect 2501 24695 2559 24701
rect 3602 24692 3608 24704
rect 3660 24692 3666 24744
rect 3786 24692 3792 24744
rect 3844 24732 3850 24744
rect 3973 24735 4031 24741
rect 3973 24732 3985 24735
rect 3844 24704 3985 24732
rect 3844 24692 3850 24704
rect 3973 24701 3985 24704
rect 4019 24701 4031 24735
rect 3973 24695 4031 24701
rect 2406 24664 2412 24676
rect 2367 24636 2412 24664
rect 2406 24624 2412 24636
rect 2464 24624 2470 24676
rect 3988 24664 4016 24695
rect 4154 24692 4160 24744
rect 4212 24732 4218 24744
rect 4249 24735 4307 24741
rect 4249 24732 4261 24735
rect 4212 24704 4261 24732
rect 4212 24692 4218 24704
rect 4249 24701 4261 24704
rect 4295 24732 4307 24735
rect 5258 24732 5264 24744
rect 4295 24704 5264 24732
rect 4295 24701 4307 24704
rect 4249 24695 4307 24701
rect 5258 24692 5264 24704
rect 5316 24692 5322 24744
rect 5721 24735 5779 24741
rect 5721 24701 5733 24735
rect 5767 24732 5779 24735
rect 5767 24704 6684 24732
rect 5767 24701 5779 24704
rect 5721 24695 5779 24701
rect 4522 24664 4528 24676
rect 3988 24636 4528 24664
rect 4522 24624 4528 24636
rect 4580 24664 4586 24676
rect 4985 24667 5043 24673
rect 4985 24664 4997 24667
rect 4580 24636 4997 24664
rect 4580 24624 4586 24636
rect 4985 24633 4997 24636
rect 5031 24633 5043 24667
rect 4985 24627 5043 24633
rect 6656 24608 6684 24704
rect 7208 24673 7236 24772
rect 7837 24769 7849 24803
rect 7883 24800 7895 24803
rect 8202 24800 8208 24812
rect 7883 24772 8208 24800
rect 7883 24769 7895 24772
rect 7837 24763 7895 24769
rect 8202 24760 8208 24772
rect 8260 24760 8266 24812
rect 8757 24803 8815 24809
rect 8757 24800 8769 24803
rect 8312 24772 8769 24800
rect 7466 24732 7472 24744
rect 7427 24704 7472 24732
rect 7466 24692 7472 24704
rect 7524 24692 7530 24744
rect 7926 24692 7932 24744
rect 7984 24732 7990 24744
rect 8113 24735 8171 24741
rect 8113 24732 8125 24735
rect 7984 24704 8125 24732
rect 7984 24692 7990 24704
rect 8113 24701 8125 24704
rect 8159 24732 8171 24735
rect 8312 24732 8340 24772
rect 8757 24769 8769 24772
rect 8803 24769 8815 24803
rect 8757 24763 8815 24769
rect 9401 24803 9459 24809
rect 9401 24769 9413 24803
rect 9447 24800 9459 24803
rect 13630 24800 13636 24812
rect 9447 24772 13636 24800
rect 9447 24769 9459 24772
rect 9401 24763 9459 24769
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 18969 24803 19027 24809
rect 18969 24769 18981 24803
rect 19015 24800 19027 24803
rect 20254 24800 20260 24812
rect 19015 24772 20116 24800
rect 20215 24772 20260 24800
rect 19015 24769 19027 24772
rect 18969 24763 19027 24769
rect 8159 24704 8340 24732
rect 8665 24735 8723 24741
rect 8159 24701 8171 24704
rect 8113 24695 8171 24701
rect 8665 24701 8677 24735
rect 8711 24701 8723 24735
rect 8938 24732 8944 24744
rect 8899 24704 8944 24732
rect 8665 24695 8723 24701
rect 7193 24667 7251 24673
rect 7193 24633 7205 24667
rect 7239 24664 7251 24667
rect 7285 24667 7343 24673
rect 7285 24664 7297 24667
rect 7239 24636 7297 24664
rect 7239 24633 7251 24636
rect 7193 24627 7251 24633
rect 7285 24633 7297 24636
rect 7331 24664 7343 24667
rect 8570 24664 8576 24676
rect 7331 24636 8576 24664
rect 7331 24633 7343 24636
rect 7285 24627 7343 24633
rect 8570 24624 8576 24636
rect 8628 24624 8634 24676
rect 5534 24596 5540 24608
rect 5495 24568 5540 24596
rect 5534 24556 5540 24568
rect 5592 24556 5598 24608
rect 5902 24596 5908 24608
rect 5863 24568 5908 24596
rect 5902 24556 5908 24568
rect 5960 24556 5966 24608
rect 6638 24596 6644 24608
rect 6599 24568 6644 24596
rect 6638 24556 6644 24568
rect 6696 24556 6702 24608
rect 8110 24556 8116 24608
rect 8168 24596 8174 24608
rect 8481 24599 8539 24605
rect 8481 24596 8493 24599
rect 8168 24568 8493 24596
rect 8168 24556 8174 24568
rect 8481 24565 8493 24568
rect 8527 24596 8539 24599
rect 8680 24596 8708 24695
rect 8938 24692 8944 24704
rect 8996 24692 9002 24744
rect 10597 24735 10655 24741
rect 10597 24732 10609 24735
rect 10244 24704 10609 24732
rect 8754 24624 8760 24676
rect 8812 24664 8818 24676
rect 10244 24673 10272 24704
rect 10597 24701 10609 24704
rect 10643 24732 10655 24735
rect 11974 24732 11980 24744
rect 10643 24704 11980 24732
rect 10643 24701 10655 24704
rect 10597 24695 10655 24701
rect 11974 24692 11980 24704
rect 12032 24732 12038 24744
rect 12161 24735 12219 24741
rect 12161 24732 12173 24735
rect 12032 24704 12173 24732
rect 12032 24692 12038 24704
rect 12161 24701 12173 24704
rect 12207 24732 12219 24735
rect 12434 24732 12440 24744
rect 12207 24704 12440 24732
rect 12207 24701 12219 24704
rect 12161 24695 12219 24701
rect 12434 24692 12440 24704
rect 12492 24732 12498 24744
rect 12621 24735 12679 24741
rect 12621 24732 12633 24735
rect 12492 24704 12633 24732
rect 12492 24692 12498 24704
rect 12621 24701 12633 24704
rect 12667 24732 12679 24735
rect 12989 24735 13047 24741
rect 12989 24732 13001 24735
rect 12667 24704 13001 24732
rect 12667 24701 12679 24704
rect 12621 24695 12679 24701
rect 12989 24701 13001 24704
rect 13035 24701 13047 24735
rect 14458 24732 14464 24744
rect 14419 24704 14464 24732
rect 12989 24695 13047 24701
rect 14458 24692 14464 24704
rect 14516 24692 14522 24744
rect 14642 24732 14648 24744
rect 14603 24704 14648 24732
rect 14642 24692 14648 24704
rect 14700 24692 14706 24744
rect 14918 24732 14924 24744
rect 14879 24704 14924 24732
rect 14918 24692 14924 24704
rect 14976 24692 14982 24744
rect 15749 24735 15807 24741
rect 15749 24701 15761 24735
rect 15795 24701 15807 24735
rect 15749 24695 15807 24701
rect 17012 24735 17070 24741
rect 17012 24701 17024 24735
rect 17058 24732 17070 24735
rect 17126 24732 17132 24744
rect 17058 24704 17132 24732
rect 17058 24701 17070 24704
rect 17012 24695 17070 24701
rect 10229 24667 10287 24673
rect 10229 24664 10241 24667
rect 8812 24636 10241 24664
rect 8812 24624 8818 24636
rect 10229 24633 10241 24636
rect 10275 24633 10287 24667
rect 10229 24627 10287 24633
rect 10413 24667 10471 24673
rect 10413 24633 10425 24667
rect 10459 24664 10471 24667
rect 10459 24636 11284 24664
rect 10459 24633 10471 24636
rect 10413 24627 10471 24633
rect 11256 24608 11284 24636
rect 12066 24624 12072 24676
rect 12124 24664 12130 24676
rect 12805 24667 12863 24673
rect 12805 24664 12817 24667
rect 12124 24636 12817 24664
rect 12124 24624 12130 24636
rect 12805 24633 12817 24636
rect 12851 24664 12863 24667
rect 13633 24667 13691 24673
rect 13633 24664 13645 24667
rect 12851 24636 13645 24664
rect 12851 24633 12863 24636
rect 12805 24627 12863 24633
rect 13633 24633 13645 24636
rect 13679 24664 13691 24667
rect 15565 24667 15623 24673
rect 15565 24664 15577 24667
rect 13679 24636 15577 24664
rect 13679 24633 13691 24636
rect 13633 24627 13691 24633
rect 15565 24633 15577 24636
rect 15611 24664 15623 24667
rect 15764 24664 15792 24695
rect 17126 24692 17132 24704
rect 17184 24692 17190 24744
rect 17770 24692 17776 24744
rect 17828 24732 17834 24744
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 17828 24704 18061 24732
rect 17828 24692 17834 24704
rect 18049 24701 18061 24704
rect 18095 24732 18107 24735
rect 18509 24735 18567 24741
rect 18509 24732 18521 24735
rect 18095 24704 18521 24732
rect 18095 24701 18107 24704
rect 18049 24695 18107 24701
rect 18509 24701 18521 24704
rect 18555 24701 18567 24735
rect 19794 24732 19800 24744
rect 19755 24704 19800 24732
rect 18509 24695 18567 24701
rect 19794 24692 19800 24704
rect 19852 24692 19858 24744
rect 20088 24741 20116 24772
rect 20254 24760 20260 24772
rect 20312 24760 20318 24812
rect 20625 24803 20683 24809
rect 20625 24769 20637 24803
rect 20671 24800 20683 24803
rect 21266 24800 21272 24812
rect 20671 24772 21272 24800
rect 20671 24769 20683 24772
rect 20625 24763 20683 24769
rect 21266 24760 21272 24772
rect 21324 24760 21330 24812
rect 21821 24803 21879 24809
rect 21821 24769 21833 24803
rect 21867 24800 21879 24803
rect 22278 24800 22284 24812
rect 21867 24772 22284 24800
rect 21867 24769 21879 24772
rect 21821 24763 21879 24769
rect 22278 24760 22284 24772
rect 22336 24760 22342 24812
rect 23032 24800 23060 24896
rect 24302 24868 24308 24880
rect 24263 24840 24308 24868
rect 24302 24828 24308 24840
rect 24360 24868 24366 24880
rect 24854 24868 24860 24880
rect 24360 24840 24860 24868
rect 24360 24828 24366 24840
rect 24854 24828 24860 24840
rect 24912 24828 24918 24880
rect 23753 24803 23811 24809
rect 23753 24800 23765 24803
rect 23032 24772 23765 24800
rect 23753 24769 23765 24772
rect 23799 24769 23811 24803
rect 23753 24763 23811 24769
rect 20073 24735 20131 24741
rect 20073 24701 20085 24735
rect 20119 24732 20131 24735
rect 20346 24732 20352 24744
rect 20119 24704 20352 24732
rect 20119 24701 20131 24704
rect 20073 24695 20131 24701
rect 20346 24692 20352 24704
rect 20404 24692 20410 24744
rect 25643 24741 25671 24908
rect 26145 24905 26157 24908
rect 26191 24936 26203 24939
rect 28534 24936 28540 24948
rect 26191 24908 28540 24936
rect 26191 24905 26203 24908
rect 26145 24899 26203 24905
rect 28534 24896 28540 24908
rect 28592 24896 28598 24948
rect 29086 24936 29092 24948
rect 29047 24908 29092 24936
rect 29086 24896 29092 24908
rect 29144 24896 29150 24948
rect 33321 24939 33379 24945
rect 33321 24936 33333 24939
rect 29748 24908 33333 24936
rect 27338 24868 27344 24880
rect 27299 24840 27344 24868
rect 27338 24828 27344 24840
rect 27396 24828 27402 24880
rect 28721 24871 28779 24877
rect 28721 24837 28733 24871
rect 28767 24868 28779 24871
rect 29178 24868 29184 24880
rect 28767 24840 29184 24868
rect 28767 24837 28779 24840
rect 28721 24831 28779 24837
rect 29178 24828 29184 24840
rect 29236 24868 29242 24880
rect 29748 24868 29776 24908
rect 33321 24905 33333 24908
rect 33367 24905 33379 24939
rect 33321 24899 33379 24905
rect 33410 24896 33416 24948
rect 33468 24936 33474 24948
rect 33781 24939 33839 24945
rect 33781 24936 33793 24939
rect 33468 24908 33793 24936
rect 33468 24896 33474 24908
rect 33781 24905 33793 24908
rect 33827 24905 33839 24939
rect 35894 24936 35900 24948
rect 35855 24908 35900 24936
rect 33781 24899 33839 24905
rect 35894 24896 35900 24908
rect 35952 24896 35958 24948
rect 39298 24936 39304 24948
rect 39259 24908 39304 24936
rect 39298 24896 39304 24908
rect 39356 24896 39362 24948
rect 39758 24896 39764 24948
rect 39816 24936 39822 24948
rect 40221 24939 40279 24945
rect 40221 24936 40233 24939
rect 39816 24908 40233 24936
rect 39816 24896 39822 24908
rect 40221 24905 40233 24908
rect 40267 24905 40279 24939
rect 41966 24936 41972 24948
rect 41927 24908 41972 24936
rect 40221 24899 40279 24905
rect 41966 24896 41972 24908
rect 42024 24936 42030 24948
rect 43254 24936 43260 24948
rect 42024 24908 43260 24936
rect 42024 24896 42030 24908
rect 43254 24896 43260 24908
rect 43312 24936 43318 24948
rect 43349 24939 43407 24945
rect 43349 24936 43361 24939
rect 43312 24908 43361 24936
rect 43312 24896 43318 24908
rect 43349 24905 43361 24908
rect 43395 24905 43407 24939
rect 43349 24899 43407 24905
rect 29236 24840 29776 24868
rect 29236 24828 29242 24840
rect 34330 24828 34336 24880
rect 34388 24868 34394 24880
rect 36265 24871 36323 24877
rect 36265 24868 36277 24871
rect 34388 24840 36277 24868
rect 34388 24828 34394 24840
rect 36265 24837 36277 24840
rect 36311 24868 36323 24871
rect 36354 24868 36360 24880
rect 36311 24840 36360 24868
rect 36311 24837 36323 24840
rect 36265 24831 36323 24837
rect 36354 24828 36360 24840
rect 36412 24828 36418 24880
rect 38746 24828 38752 24880
rect 38804 24868 38810 24880
rect 43990 24868 43996 24880
rect 38804 24840 43996 24868
rect 38804 24828 38810 24840
rect 43990 24828 43996 24840
rect 44048 24828 44054 24880
rect 25731 24803 25789 24809
rect 25731 24769 25743 24803
rect 25777 24800 25789 24803
rect 27709 24803 27767 24809
rect 27709 24800 27721 24803
rect 25777 24772 27721 24800
rect 25777 24769 25789 24772
rect 25731 24763 25789 24769
rect 27709 24769 27721 24772
rect 27755 24800 27767 24803
rect 28442 24800 28448 24812
rect 27755 24772 28448 24800
rect 27755 24769 27767 24772
rect 27709 24763 27767 24769
rect 28442 24760 28448 24772
rect 28500 24760 28506 24812
rect 29638 24800 29644 24812
rect 29196 24772 29644 24800
rect 25628 24735 25686 24741
rect 25628 24701 25640 24735
rect 25674 24701 25686 24735
rect 25628 24695 25686 24701
rect 26050 24692 26056 24744
rect 26108 24732 26114 24744
rect 26640 24735 26698 24741
rect 26640 24732 26652 24735
rect 26108 24704 26652 24732
rect 26108 24692 26114 24704
rect 26640 24701 26652 24704
rect 26686 24701 26698 24735
rect 26640 24695 26698 24701
rect 28353 24735 28411 24741
rect 28353 24701 28365 24735
rect 28399 24732 28411 24735
rect 29196 24732 29224 24772
rect 29638 24760 29644 24772
rect 29696 24760 29702 24812
rect 30929 24803 30987 24809
rect 30929 24769 30941 24803
rect 30975 24800 30987 24803
rect 31662 24800 31668 24812
rect 30975 24772 31668 24800
rect 30975 24769 30987 24772
rect 30929 24763 30987 24769
rect 31662 24760 31668 24772
rect 31720 24760 31726 24812
rect 32122 24800 32128 24812
rect 32083 24772 32128 24800
rect 32122 24760 32128 24772
rect 32180 24760 32186 24812
rect 32490 24800 32496 24812
rect 32451 24772 32496 24800
rect 32490 24760 32496 24772
rect 32548 24760 32554 24812
rect 33134 24760 33140 24812
rect 33192 24800 33198 24812
rect 33192 24772 33237 24800
rect 33192 24760 33198 24772
rect 34422 24760 34428 24812
rect 34480 24800 34486 24812
rect 35253 24803 35311 24809
rect 35253 24800 35265 24803
rect 34480 24772 35265 24800
rect 34480 24760 34486 24772
rect 35253 24769 35265 24772
rect 35299 24769 35311 24803
rect 36814 24800 36820 24812
rect 36775 24772 36820 24800
rect 35253 24763 35311 24769
rect 36814 24760 36820 24772
rect 36872 24760 36878 24812
rect 39942 24760 39948 24812
rect 40000 24800 40006 24812
rect 40000 24772 44358 24800
rect 40000 24760 40006 24772
rect 28399 24704 29224 24732
rect 28399 24701 28411 24704
rect 28353 24695 28411 24701
rect 15611 24636 15792 24664
rect 15611 24633 15623 24636
rect 15565 24627 15623 24633
rect 16482 24624 16488 24676
rect 16540 24664 16546 24676
rect 16577 24667 16635 24673
rect 16577 24664 16589 24667
rect 16540 24636 16589 24664
rect 16540 24624 16546 24636
rect 16577 24633 16589 24636
rect 16623 24664 16635 24667
rect 17678 24664 17684 24676
rect 16623 24636 17684 24664
rect 16623 24633 16635 24636
rect 16577 24627 16635 24633
rect 17678 24624 17684 24636
rect 17736 24624 17742 24676
rect 21174 24664 21180 24676
rect 21135 24636 21180 24664
rect 21174 24624 21180 24636
rect 21232 24624 21238 24676
rect 21266 24624 21272 24676
rect 21324 24664 21330 24676
rect 23842 24664 23848 24676
rect 21324 24636 21369 24664
rect 23803 24636 23848 24664
rect 21324 24624 21330 24636
rect 23842 24624 23848 24636
rect 23900 24624 23906 24676
rect 26655 24664 26683 24695
rect 31570 24692 31576 24744
rect 31628 24732 31634 24744
rect 38010 24732 38016 24744
rect 31628 24704 31673 24732
rect 37971 24704 38016 24732
rect 31628 24692 31634 24704
rect 38010 24692 38016 24704
rect 38068 24732 38074 24744
rect 38473 24735 38531 24741
rect 38473 24732 38485 24735
rect 38068 24704 38485 24732
rect 38068 24692 38074 24704
rect 38473 24701 38485 24704
rect 38519 24701 38531 24735
rect 38473 24695 38531 24701
rect 39428 24735 39486 24741
rect 39428 24701 39440 24735
rect 39474 24732 39486 24735
rect 39853 24735 39911 24741
rect 39853 24732 39865 24735
rect 39474 24704 39865 24732
rect 39474 24701 39486 24704
rect 39428 24695 39486 24701
rect 39853 24701 39865 24704
rect 39899 24732 39911 24735
rect 40402 24732 40408 24744
rect 39899 24704 40408 24732
rect 39899 24701 39911 24704
rect 39853 24695 39911 24701
rect 26620 24636 26683 24664
rect 26743 24667 26801 24673
rect 10686 24596 10692 24608
rect 8527 24568 8708 24596
rect 10647 24568 10692 24596
rect 8527 24565 8539 24568
rect 8481 24559 8539 24565
rect 10686 24556 10692 24568
rect 10744 24556 10750 24608
rect 11238 24596 11244 24608
rect 11199 24568 11244 24596
rect 11238 24556 11244 24568
rect 11296 24556 11302 24608
rect 14182 24556 14188 24608
rect 14240 24596 14246 24608
rect 15197 24599 15255 24605
rect 15197 24596 15209 24599
rect 14240 24568 15209 24596
rect 14240 24556 14246 24568
rect 15197 24565 15209 24568
rect 15243 24596 15255 24599
rect 15286 24596 15292 24608
rect 15243 24568 15292 24596
rect 15243 24565 15255 24568
rect 15197 24559 15255 24565
rect 15286 24556 15292 24568
rect 15344 24556 15350 24608
rect 17083 24599 17141 24605
rect 17083 24565 17095 24599
rect 17129 24596 17141 24599
rect 17402 24596 17408 24608
rect 17129 24568 17408 24596
rect 17129 24565 17141 24568
rect 17083 24559 17141 24565
rect 17402 24556 17408 24568
rect 17460 24556 17466 24608
rect 21192 24596 21220 24624
rect 26620 24608 26648 24636
rect 26743 24633 26755 24667
rect 26789 24664 26801 24667
rect 26789 24636 27521 24664
rect 26789 24633 26801 24636
rect 26743 24627 26801 24633
rect 22465 24599 22523 24605
rect 22465 24596 22477 24599
rect 21192 24568 22477 24596
rect 22465 24565 22477 24568
rect 22511 24596 22523 24599
rect 22922 24596 22928 24608
rect 22511 24568 22928 24596
rect 22511 24565 22523 24568
rect 22465 24559 22523 24565
rect 22922 24556 22928 24568
rect 22980 24556 22986 24608
rect 26513 24599 26571 24605
rect 26513 24565 26525 24599
rect 26559 24596 26571 24599
rect 26602 24596 26608 24608
rect 26559 24568 26608 24596
rect 26559 24565 26571 24568
rect 26513 24559 26571 24565
rect 26602 24556 26608 24568
rect 26660 24556 26666 24608
rect 27493 24596 27521 24636
rect 27706 24624 27712 24676
rect 27764 24664 27770 24676
rect 27801 24667 27859 24673
rect 27801 24664 27813 24667
rect 27764 24636 27813 24664
rect 27764 24624 27770 24636
rect 27801 24633 27813 24636
rect 27847 24633 27859 24667
rect 29362 24664 29368 24676
rect 27801 24627 27859 24633
rect 28552 24636 29368 24664
rect 28552 24596 28580 24636
rect 29362 24624 29368 24636
rect 29420 24624 29426 24676
rect 29457 24667 29515 24673
rect 29457 24633 29469 24667
rect 29503 24633 29515 24667
rect 31021 24667 31079 24673
rect 31021 24664 31033 24667
rect 29457 24627 29515 24633
rect 30576 24636 31033 24664
rect 27493 24568 28580 24596
rect 29086 24556 29092 24608
rect 29144 24596 29150 24608
rect 29472 24596 29500 24627
rect 30576 24608 30604 24636
rect 31021 24633 31033 24636
rect 31067 24664 31079 24667
rect 31294 24664 31300 24676
rect 31067 24636 31300 24664
rect 31067 24633 31079 24636
rect 31021 24627 31079 24633
rect 31294 24624 31300 24636
rect 31352 24624 31358 24676
rect 32582 24664 32588 24676
rect 32543 24636 32588 24664
rect 32582 24624 32588 24636
rect 32640 24624 32646 24676
rect 34146 24664 34152 24676
rect 33244 24636 34152 24664
rect 30285 24599 30343 24605
rect 30285 24596 30297 24599
rect 29144 24568 30297 24596
rect 29144 24556 29150 24568
rect 30285 24565 30297 24568
rect 30331 24596 30343 24599
rect 30558 24596 30564 24608
rect 30331 24568 30564 24596
rect 30331 24565 30343 24568
rect 30285 24559 30343 24565
rect 30558 24556 30564 24568
rect 30616 24556 30622 24608
rect 30650 24556 30656 24608
rect 30708 24596 30714 24608
rect 30745 24599 30803 24605
rect 30745 24596 30757 24599
rect 30708 24568 30757 24596
rect 30708 24556 30714 24568
rect 30745 24565 30757 24568
rect 30791 24596 30803 24599
rect 31386 24596 31392 24608
rect 30791 24568 31392 24596
rect 30791 24565 30803 24568
rect 30745 24559 30803 24565
rect 31386 24556 31392 24568
rect 31444 24556 31450 24608
rect 32122 24556 32128 24608
rect 32180 24596 32186 24608
rect 33244 24596 33272 24636
rect 34146 24624 34152 24636
rect 34204 24624 34210 24676
rect 34514 24624 34520 24676
rect 34572 24664 34578 24676
rect 34977 24667 35035 24673
rect 34977 24664 34989 24667
rect 34572 24636 34989 24664
rect 34572 24624 34578 24636
rect 34977 24633 34989 24636
rect 35023 24633 35035 24667
rect 34977 24627 35035 24633
rect 35069 24667 35127 24673
rect 35069 24633 35081 24667
rect 35115 24664 35127 24667
rect 35250 24664 35256 24676
rect 35115 24636 35256 24664
rect 35115 24633 35127 24636
rect 35069 24627 35127 24633
rect 32180 24568 33272 24596
rect 33321 24599 33379 24605
rect 32180 24556 32186 24568
rect 33321 24565 33333 24599
rect 33367 24596 33379 24599
rect 33505 24599 33563 24605
rect 33505 24596 33517 24599
rect 33367 24568 33517 24596
rect 33367 24565 33379 24568
rect 33321 24559 33379 24565
rect 33505 24565 33517 24568
rect 33551 24596 33563 24599
rect 34333 24599 34391 24605
rect 34333 24596 34345 24599
rect 33551 24568 34345 24596
rect 33551 24565 33563 24568
rect 33505 24559 33563 24565
rect 34333 24565 34345 24568
rect 34379 24596 34391 24599
rect 34701 24599 34759 24605
rect 34701 24596 34713 24599
rect 34379 24568 34713 24596
rect 34379 24565 34391 24568
rect 34333 24559 34391 24565
rect 34701 24565 34713 24568
rect 34747 24596 34759 24599
rect 35084 24596 35112 24627
rect 35250 24624 35256 24636
rect 35308 24624 35314 24676
rect 36541 24667 36599 24673
rect 36541 24633 36553 24667
rect 36587 24633 36599 24667
rect 36541 24627 36599 24633
rect 36633 24667 36691 24673
rect 36633 24633 36645 24667
rect 36679 24664 36691 24667
rect 36906 24664 36912 24676
rect 36679 24636 36912 24664
rect 36679 24633 36691 24636
rect 36633 24627 36691 24633
rect 34747 24568 35112 24596
rect 36556 24596 36584 24627
rect 36906 24624 36912 24636
rect 36964 24624 36970 24676
rect 37642 24624 37648 24676
rect 37700 24664 37706 24676
rect 39443 24664 39471 24695
rect 40402 24692 40408 24704
rect 40460 24692 40466 24744
rect 42702 24692 42708 24744
rect 42760 24732 42766 24744
rect 42832 24735 42890 24741
rect 42832 24732 42844 24735
rect 42760 24704 42844 24732
rect 42760 24692 42794 24704
rect 42832 24701 42844 24704
rect 42878 24701 42890 24735
rect 42832 24695 42890 24701
rect 43876 24735 43934 24741
rect 43876 24701 43888 24735
rect 43922 24701 43934 24735
rect 44330 24732 44358 24772
rect 44856 24735 44914 24741
rect 44856 24732 44868 24735
rect 44330 24704 44868 24732
rect 43876 24695 43934 24701
rect 44856 24701 44868 24704
rect 44902 24732 44914 24735
rect 45281 24735 45339 24741
rect 45281 24732 45293 24735
rect 44902 24704 45293 24732
rect 44902 24701 44914 24704
rect 44856 24695 44914 24701
rect 45281 24701 45293 24704
rect 45327 24701 45339 24735
rect 45281 24695 45339 24701
rect 41046 24664 41052 24676
rect 37700 24636 39471 24664
rect 41007 24636 41052 24664
rect 37700 24624 37706 24636
rect 41046 24624 41052 24636
rect 41104 24624 41110 24676
rect 41141 24667 41199 24673
rect 41141 24633 41153 24667
rect 41187 24633 41199 24667
rect 41141 24627 41199 24633
rect 41693 24667 41751 24673
rect 41693 24633 41705 24667
rect 41739 24664 41751 24667
rect 41782 24664 41788 24676
rect 41739 24636 41788 24664
rect 41739 24633 41751 24636
rect 41693 24627 41751 24633
rect 37550 24596 37556 24608
rect 36556 24568 37556 24596
rect 34747 24565 34759 24568
rect 34701 24559 34759 24565
rect 37550 24556 37556 24568
rect 37608 24556 37614 24608
rect 38197 24599 38255 24605
rect 38197 24565 38209 24599
rect 38243 24596 38255 24599
rect 38838 24596 38844 24608
rect 38243 24568 38844 24596
rect 38243 24565 38255 24568
rect 38197 24559 38255 24565
rect 38838 24556 38844 24568
rect 38896 24556 38902 24608
rect 39531 24599 39589 24605
rect 39531 24565 39543 24599
rect 39577 24596 39589 24599
rect 39758 24596 39764 24608
rect 39577 24568 39764 24596
rect 39577 24565 39589 24568
rect 39531 24559 39589 24565
rect 39758 24556 39764 24568
rect 39816 24556 39822 24608
rect 40865 24599 40923 24605
rect 40865 24565 40877 24599
rect 40911 24596 40923 24599
rect 41156 24596 41184 24627
rect 41782 24624 41788 24636
rect 41840 24624 41846 24676
rect 41322 24596 41328 24608
rect 40911 24568 41328 24596
rect 40911 24565 40923 24568
rect 40865 24559 40923 24565
rect 41322 24556 41328 24568
rect 41380 24556 41386 24608
rect 41414 24556 41420 24608
rect 41472 24596 41478 24608
rect 42613 24599 42671 24605
rect 42613 24596 42625 24599
rect 41472 24568 42625 24596
rect 41472 24556 41478 24568
rect 42613 24565 42625 24568
rect 42659 24596 42671 24599
rect 42766 24596 42794 24692
rect 43891 24664 43919 24695
rect 44266 24664 44272 24676
rect 43891 24636 44272 24664
rect 44266 24624 44272 24636
rect 44324 24624 44330 24676
rect 42659 24568 42794 24596
rect 42935 24599 42993 24605
rect 42659 24565 42671 24568
rect 42613 24559 42671 24565
rect 42935 24565 42947 24599
rect 42981 24596 42993 24599
rect 43162 24596 43168 24608
rect 42981 24568 43168 24596
rect 42981 24565 42993 24568
rect 42935 24559 42993 24565
rect 43162 24556 43168 24568
rect 43220 24556 43226 24608
rect 43530 24556 43536 24608
rect 43588 24596 43594 24608
rect 43947 24599 44005 24605
rect 43947 24596 43959 24599
rect 43588 24568 43959 24596
rect 43588 24556 43594 24568
rect 43947 24565 43959 24568
rect 43993 24565 44005 24599
rect 44634 24596 44640 24608
rect 44595 24568 44640 24596
rect 43947 24559 44005 24565
rect 44634 24556 44640 24568
rect 44692 24556 44698 24608
rect 44726 24556 44732 24608
rect 44784 24596 44790 24608
rect 44959 24599 45017 24605
rect 44959 24596 44971 24599
rect 44784 24568 44971 24596
rect 44784 24556 44790 24568
rect 44959 24565 44971 24568
rect 45005 24565 45017 24599
rect 44959 24559 45017 24565
rect 1104 24506 48852 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 48852 24506
rect 1104 24432 48852 24454
rect 2222 24392 2228 24404
rect 2183 24364 2228 24392
rect 2222 24352 2228 24364
rect 2280 24352 2286 24404
rect 2958 24352 2964 24404
rect 3016 24392 3022 24404
rect 3329 24395 3387 24401
rect 3329 24392 3341 24395
rect 3016 24364 3341 24392
rect 3016 24352 3022 24364
rect 3329 24361 3341 24364
rect 3375 24392 3387 24395
rect 3418 24392 3424 24404
rect 3375 24364 3424 24392
rect 3375 24361 3387 24364
rect 3329 24355 3387 24361
rect 3418 24352 3424 24364
rect 3476 24352 3482 24404
rect 3694 24352 3700 24404
rect 3752 24392 3758 24404
rect 4709 24395 4767 24401
rect 4709 24392 4721 24395
rect 3752 24364 4721 24392
rect 3752 24352 3758 24364
rect 4709 24361 4721 24364
rect 4755 24361 4767 24395
rect 4709 24355 4767 24361
rect 6638 24352 6644 24404
rect 6696 24392 6702 24404
rect 7469 24395 7527 24401
rect 7469 24392 7481 24395
rect 6696 24364 7481 24392
rect 6696 24352 6702 24364
rect 7469 24361 7481 24364
rect 7515 24361 7527 24395
rect 7469 24355 7527 24361
rect 9950 24352 9956 24404
rect 10008 24392 10014 24404
rect 10045 24395 10103 24401
rect 10045 24392 10057 24395
rect 10008 24364 10057 24392
rect 10008 24352 10014 24364
rect 10045 24361 10057 24364
rect 10091 24361 10103 24395
rect 10045 24355 10103 24361
rect 10413 24395 10471 24401
rect 10413 24361 10425 24395
rect 10459 24392 10471 24395
rect 10686 24392 10692 24404
rect 10459 24364 10692 24392
rect 10459 24361 10471 24364
rect 10413 24355 10471 24361
rect 3970 24324 3976 24336
rect 1872 24296 3976 24324
rect 1486 24216 1492 24268
rect 1544 24256 1550 24268
rect 1872 24265 1900 24296
rect 3970 24284 3976 24296
rect 4028 24324 4034 24336
rect 4065 24327 4123 24333
rect 4065 24324 4077 24327
rect 4028 24296 4077 24324
rect 4028 24284 4034 24296
rect 4065 24293 4077 24296
rect 4111 24293 4123 24327
rect 6362 24324 6368 24336
rect 6323 24296 6368 24324
rect 4065 24287 4123 24293
rect 6362 24284 6368 24296
rect 6420 24284 6426 24336
rect 6730 24324 6736 24336
rect 6691 24296 6736 24324
rect 6730 24284 6736 24296
rect 6788 24284 6794 24336
rect 1857 24259 1915 24265
rect 1857 24256 1869 24259
rect 1544 24228 1869 24256
rect 1544 24216 1550 24228
rect 1857 24225 1869 24228
rect 1903 24225 1915 24259
rect 1857 24219 1915 24225
rect 2130 24216 2136 24268
rect 2188 24256 2194 24268
rect 2958 24256 2964 24268
rect 2188 24228 2964 24256
rect 2188 24216 2194 24228
rect 2958 24216 2964 24228
rect 3016 24216 3022 24268
rect 5629 24259 5687 24265
rect 5629 24256 5641 24259
rect 5460 24228 5641 24256
rect 3881 24191 3939 24197
rect 3881 24157 3893 24191
rect 3927 24188 3939 24191
rect 4154 24188 4160 24200
rect 3927 24160 4160 24188
rect 3927 24157 3939 24160
rect 3881 24151 3939 24157
rect 2498 24080 2504 24132
rect 2556 24120 2562 24132
rect 3896 24120 3924 24151
rect 4154 24148 4160 24160
rect 4212 24148 4218 24200
rect 4433 24191 4491 24197
rect 4433 24157 4445 24191
rect 4479 24188 4491 24191
rect 4614 24188 4620 24200
rect 4479 24160 4620 24188
rect 4479 24157 4491 24160
rect 4433 24151 4491 24157
rect 4614 24148 4620 24160
rect 4672 24148 4678 24200
rect 4341 24123 4399 24129
rect 4341 24120 4353 24123
rect 2556 24092 3924 24120
rect 4126 24092 4353 24120
rect 2556 24080 2562 24092
rect 4126 24064 4154 24092
rect 4341 24089 4353 24092
rect 4387 24089 4399 24123
rect 4522 24120 4528 24132
rect 4341 24083 4399 24089
rect 4448 24092 4528 24120
rect 4062 24012 4068 24064
rect 4120 24024 4154 24064
rect 4230 24055 4288 24061
rect 4120 24012 4126 24024
rect 4230 24021 4242 24055
rect 4276 24052 4288 24055
rect 4448 24052 4476 24092
rect 4522 24080 4528 24092
rect 4580 24120 4586 24132
rect 5460 24129 5488 24228
rect 5629 24225 5641 24228
rect 5675 24256 5687 24259
rect 5810 24256 5816 24268
rect 5675 24228 5816 24256
rect 5675 24225 5687 24228
rect 5629 24219 5687 24225
rect 5810 24216 5816 24228
rect 5868 24216 5874 24268
rect 5905 24259 5963 24265
rect 5905 24225 5917 24259
rect 5951 24256 5963 24259
rect 5994 24256 6000 24268
rect 5951 24228 6000 24256
rect 5951 24225 5963 24228
rect 5905 24219 5963 24225
rect 5994 24216 6000 24228
rect 6052 24216 6058 24268
rect 7190 24256 7196 24268
rect 7151 24228 7196 24256
rect 7190 24216 7196 24228
rect 7248 24216 7254 24268
rect 7374 24256 7380 24268
rect 7335 24228 7380 24256
rect 7374 24216 7380 24228
rect 7432 24216 7438 24268
rect 8570 24256 8576 24268
rect 8531 24228 8576 24256
rect 8570 24216 8576 24228
rect 8628 24216 8634 24268
rect 9861 24259 9919 24265
rect 9861 24225 9873 24259
rect 9907 24256 9919 24259
rect 10428 24256 10456 24355
rect 10686 24352 10692 24364
rect 10744 24352 10750 24404
rect 11146 24392 11152 24404
rect 11107 24364 11152 24392
rect 11146 24352 11152 24364
rect 11204 24352 11210 24404
rect 12526 24392 12532 24404
rect 12487 24364 12532 24392
rect 12526 24352 12532 24364
rect 12584 24352 12590 24404
rect 14550 24392 14556 24404
rect 13786 24364 14412 24392
rect 14511 24364 14556 24392
rect 10873 24327 10931 24333
rect 10873 24293 10885 24327
rect 10919 24324 10931 24327
rect 11238 24324 11244 24336
rect 10919 24296 11244 24324
rect 10919 24293 10931 24296
rect 10873 24287 10931 24293
rect 11238 24284 11244 24296
rect 11296 24284 11302 24336
rect 13630 24324 13636 24336
rect 13591 24296 13636 24324
rect 13630 24284 13636 24296
rect 13688 24324 13694 24336
rect 13786 24324 13814 24364
rect 14182 24324 14188 24336
rect 13688 24296 13814 24324
rect 14143 24296 14188 24324
rect 13688 24284 13694 24296
rect 14182 24284 14188 24296
rect 14240 24284 14246 24336
rect 14384 24324 14412 24364
rect 14550 24352 14556 24364
rect 14608 24352 14614 24404
rect 19061 24395 19119 24401
rect 15533 24364 18920 24392
rect 15533 24324 15561 24364
rect 15654 24333 15660 24336
rect 15651 24324 15660 24333
rect 14384 24296 15561 24324
rect 15615 24296 15660 24324
rect 15651 24287 15660 24296
rect 15654 24284 15660 24287
rect 15712 24284 15718 24336
rect 17037 24327 17095 24333
rect 17037 24293 17049 24327
rect 17083 24324 17095 24327
rect 17126 24324 17132 24336
rect 17083 24296 17132 24324
rect 17083 24293 17095 24296
rect 17037 24287 17095 24293
rect 17126 24284 17132 24296
rect 17184 24324 17190 24336
rect 18782 24324 18788 24336
rect 17184 24296 18788 24324
rect 17184 24284 17190 24296
rect 18782 24284 18788 24296
rect 18840 24284 18846 24336
rect 11054 24256 11060 24268
rect 9907 24228 10456 24256
rect 11015 24228 11060 24256
rect 9907 24225 9919 24228
rect 9861 24219 9919 24225
rect 11054 24216 11060 24228
rect 11112 24216 11118 24268
rect 12253 24259 12311 24265
rect 12253 24225 12265 24259
rect 12299 24225 12311 24259
rect 12434 24256 12440 24268
rect 12395 24228 12440 24256
rect 12253 24219 12311 24225
rect 10134 24148 10140 24200
rect 10192 24188 10198 24200
rect 12268 24188 12296 24219
rect 12434 24216 12440 24228
rect 12492 24216 12498 24268
rect 13814 24216 13820 24268
rect 13872 24256 13878 24268
rect 17770 24256 17776 24268
rect 13872 24228 13917 24256
rect 15120 24228 17776 24256
rect 13872 24216 13878 24228
rect 12342 24188 12348 24200
rect 10192 24160 12348 24188
rect 10192 24148 10198 24160
rect 12342 24148 12348 24160
rect 12400 24188 12406 24200
rect 15120 24188 15148 24228
rect 17770 24216 17776 24228
rect 17828 24216 17834 24268
rect 17954 24256 17960 24268
rect 17915 24228 17960 24256
rect 17954 24216 17960 24228
rect 18012 24216 18018 24268
rect 18892 24265 18920 24364
rect 19061 24361 19073 24395
rect 19107 24361 19119 24395
rect 19061 24355 19119 24361
rect 19981 24395 20039 24401
rect 19981 24361 19993 24395
rect 20027 24392 20039 24395
rect 20070 24392 20076 24404
rect 20027 24364 20076 24392
rect 20027 24361 20039 24364
rect 19981 24355 20039 24361
rect 19076 24324 19104 24355
rect 20070 24352 20076 24364
rect 20128 24392 20134 24404
rect 20346 24392 20352 24404
rect 20128 24364 20352 24392
rect 20128 24352 20134 24364
rect 20346 24352 20352 24364
rect 20404 24352 20410 24404
rect 24118 24352 24124 24404
rect 24176 24392 24182 24404
rect 24397 24395 24455 24401
rect 24397 24392 24409 24395
rect 24176 24364 24409 24392
rect 24176 24352 24182 24364
rect 24397 24361 24409 24364
rect 24443 24361 24455 24395
rect 27706 24392 27712 24404
rect 27667 24364 27712 24392
rect 24397 24355 24455 24361
rect 19613 24327 19671 24333
rect 19613 24324 19625 24327
rect 19076 24296 19625 24324
rect 19613 24293 19625 24296
rect 19659 24324 19671 24327
rect 19886 24324 19892 24336
rect 19659 24296 19892 24324
rect 19659 24293 19671 24296
rect 19613 24287 19671 24293
rect 19886 24284 19892 24296
rect 19944 24284 19950 24336
rect 21082 24284 21088 24336
rect 21140 24324 21146 24336
rect 21177 24327 21235 24333
rect 21177 24324 21189 24327
rect 21140 24296 21189 24324
rect 21140 24284 21146 24296
rect 21177 24293 21189 24296
rect 21223 24293 21235 24327
rect 22830 24324 22836 24336
rect 22791 24296 22836 24324
rect 21177 24287 21235 24293
rect 22830 24284 22836 24296
rect 22888 24284 22894 24336
rect 22925 24327 22983 24333
rect 22925 24293 22937 24327
rect 22971 24324 22983 24327
rect 23842 24324 23848 24336
rect 22971 24296 23848 24324
rect 22971 24293 22983 24296
rect 22925 24287 22983 24293
rect 23842 24284 23848 24296
rect 23900 24284 23906 24336
rect 18877 24259 18935 24265
rect 18877 24225 18889 24259
rect 18923 24256 18935 24259
rect 19058 24256 19064 24268
rect 18923 24228 19064 24256
rect 18923 24225 18935 24228
rect 18877 24219 18935 24225
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 15286 24188 15292 24200
rect 12400 24160 15148 24188
rect 15247 24160 15292 24188
rect 12400 24148 12406 24160
rect 15286 24148 15292 24160
rect 15344 24148 15350 24200
rect 17310 24188 17316 24200
rect 17271 24160 17316 24188
rect 17310 24148 17316 24160
rect 17368 24148 17374 24200
rect 20898 24148 20904 24200
rect 20956 24188 20962 24200
rect 21085 24191 21143 24197
rect 21085 24188 21097 24191
rect 20956 24160 21097 24188
rect 20956 24148 20962 24160
rect 21085 24157 21097 24160
rect 21131 24157 21143 24191
rect 21085 24151 21143 24157
rect 21729 24191 21787 24197
rect 21729 24157 21741 24191
rect 21775 24188 21787 24191
rect 21910 24188 21916 24200
rect 21775 24160 21916 24188
rect 21775 24157 21787 24160
rect 21729 24151 21787 24157
rect 21910 24148 21916 24160
rect 21968 24148 21974 24200
rect 22922 24148 22928 24200
rect 22980 24188 22986 24200
rect 23109 24191 23167 24197
rect 23109 24188 23121 24191
rect 22980 24160 23121 24188
rect 22980 24148 22986 24160
rect 23109 24157 23121 24160
rect 23155 24188 23167 24191
rect 24412 24188 24440 24355
rect 27706 24352 27712 24364
rect 27764 24392 27770 24404
rect 28902 24392 28908 24404
rect 27764 24364 28908 24392
rect 27764 24352 27770 24364
rect 28902 24352 28908 24364
rect 28960 24352 28966 24404
rect 29362 24352 29368 24404
rect 29420 24392 29426 24404
rect 29641 24395 29699 24401
rect 29641 24392 29653 24395
rect 29420 24364 29653 24392
rect 29420 24352 29426 24364
rect 29641 24361 29653 24364
rect 29687 24361 29699 24395
rect 29641 24355 29699 24361
rect 32907 24395 32965 24401
rect 32907 24361 32919 24395
rect 32953 24392 32965 24395
rect 34514 24392 34520 24404
rect 32953 24364 34520 24392
rect 32953 24361 32965 24364
rect 32907 24355 32965 24361
rect 34514 24352 34520 24364
rect 34572 24352 34578 24404
rect 34698 24392 34704 24404
rect 34659 24364 34704 24392
rect 34698 24352 34704 24364
rect 34756 24352 34762 24404
rect 42058 24352 42064 24404
rect 42116 24392 42122 24404
rect 42153 24395 42211 24401
rect 42153 24392 42165 24395
rect 42116 24364 42165 24392
rect 42116 24352 42122 24364
rect 42153 24361 42165 24364
rect 42199 24361 42211 24395
rect 42153 24355 42211 24361
rect 43990 24352 43996 24404
rect 44048 24392 44054 24404
rect 45097 24395 45155 24401
rect 45097 24392 45109 24395
rect 44048 24364 45109 24392
rect 44048 24352 44054 24364
rect 45097 24361 45109 24364
rect 45143 24361 45155 24395
rect 45097 24355 45155 24361
rect 24762 24324 24768 24336
rect 24723 24296 24768 24324
rect 24762 24284 24768 24296
rect 24820 24284 24826 24336
rect 27338 24284 27344 24336
rect 27396 24324 27402 24336
rect 28306 24327 28364 24333
rect 28306 24324 28318 24327
rect 27396 24296 28318 24324
rect 27396 24284 27402 24296
rect 28306 24293 28318 24296
rect 28352 24293 28364 24327
rect 28306 24287 28364 24293
rect 30558 24284 30564 24336
rect 30616 24324 30622 24336
rect 30653 24327 30711 24333
rect 30653 24324 30665 24327
rect 30616 24296 30665 24324
rect 30616 24284 30622 24296
rect 30653 24293 30665 24296
rect 30699 24293 30711 24327
rect 30653 24287 30711 24293
rect 32398 24284 32404 24336
rect 32456 24324 32462 24336
rect 32677 24327 32735 24333
rect 32677 24324 32689 24327
rect 32456 24296 32689 24324
rect 32456 24284 32462 24296
rect 32677 24293 32689 24296
rect 32723 24293 32735 24327
rect 32677 24287 32735 24293
rect 33321 24327 33379 24333
rect 33321 24293 33333 24327
rect 33367 24324 33379 24327
rect 33410 24324 33416 24336
rect 33367 24296 33416 24324
rect 33367 24293 33379 24296
rect 33321 24287 33379 24293
rect 33410 24284 33416 24296
rect 33468 24324 33474 24336
rect 34606 24324 34612 24336
rect 33468 24296 34612 24324
rect 33468 24284 33474 24296
rect 34606 24284 34612 24296
rect 34664 24324 34670 24336
rect 34977 24327 35035 24333
rect 34977 24324 34989 24327
rect 34664 24296 34989 24324
rect 34664 24284 34670 24296
rect 34977 24293 34989 24296
rect 35023 24324 35035 24327
rect 36906 24324 36912 24336
rect 35023 24296 36912 24324
rect 35023 24293 35035 24296
rect 34977 24287 35035 24293
rect 36906 24284 36912 24296
rect 36964 24284 36970 24336
rect 37366 24284 37372 24336
rect 37424 24324 37430 24336
rect 39298 24324 39304 24336
rect 37424 24296 39304 24324
rect 37424 24284 37430 24296
rect 39298 24284 39304 24296
rect 39356 24324 39362 24336
rect 39530 24327 39588 24333
rect 39530 24324 39542 24327
rect 39356 24296 39542 24324
rect 39356 24284 39362 24296
rect 39530 24293 39542 24296
rect 39576 24293 39588 24327
rect 41141 24327 41199 24333
rect 41141 24324 41153 24327
rect 39530 24287 39588 24293
rect 40144 24296 41153 24324
rect 26510 24256 26516 24268
rect 26471 24228 26516 24256
rect 26510 24216 26516 24228
rect 26568 24216 26574 24268
rect 33848 24259 33906 24265
rect 33848 24256 33860 24259
rect 31220 24228 32714 24256
rect 24673 24191 24731 24197
rect 24673 24188 24685 24191
rect 23155 24160 23474 24188
rect 24412 24160 24685 24188
rect 23155 24157 23167 24160
rect 23109 24151 23167 24157
rect 5445 24123 5503 24129
rect 5445 24120 5457 24123
rect 4580 24092 5457 24120
rect 4580 24080 4586 24092
rect 5445 24089 5457 24092
rect 5491 24089 5503 24123
rect 5718 24120 5724 24132
rect 5679 24092 5724 24120
rect 5445 24083 5503 24089
rect 5718 24080 5724 24092
rect 5776 24080 5782 24132
rect 7558 24080 7564 24132
rect 7616 24120 7622 24132
rect 8113 24123 8171 24129
rect 8113 24120 8125 24123
rect 7616 24092 8125 24120
rect 7616 24080 7622 24092
rect 8113 24089 8125 24092
rect 8159 24120 8171 24123
rect 10686 24120 10692 24132
rect 8159 24092 10692 24120
rect 8159 24089 8171 24092
rect 8113 24083 8171 24089
rect 10686 24080 10692 24092
rect 10744 24080 10750 24132
rect 13173 24123 13231 24129
rect 13173 24089 13185 24123
rect 13219 24120 13231 24123
rect 13722 24120 13728 24132
rect 13219 24092 13728 24120
rect 13219 24089 13231 24092
rect 13173 24083 13231 24089
rect 13722 24080 13728 24092
rect 13780 24120 13786 24132
rect 14642 24120 14648 24132
rect 13780 24092 14648 24120
rect 13780 24080 13786 24092
rect 14642 24080 14648 24092
rect 14700 24120 14706 24132
rect 14829 24123 14887 24129
rect 14829 24120 14841 24123
rect 14700 24092 14841 24120
rect 14700 24080 14706 24092
rect 14829 24089 14841 24092
rect 14875 24089 14887 24123
rect 23446 24120 23474 24160
rect 24673 24157 24685 24160
rect 24719 24157 24731 24191
rect 24946 24188 24952 24200
rect 24859 24160 24952 24188
rect 24673 24151 24731 24157
rect 24946 24148 24952 24160
rect 25004 24148 25010 24200
rect 27982 24188 27988 24200
rect 27943 24160 27988 24188
rect 27982 24148 27988 24160
rect 28040 24148 28046 24200
rect 30558 24188 30564 24200
rect 30519 24160 30564 24188
rect 30558 24148 30564 24160
rect 30616 24148 30622 24200
rect 30742 24148 30748 24200
rect 30800 24188 30806 24200
rect 31220 24188 31248 24228
rect 30800 24160 31248 24188
rect 30800 24148 30806 24160
rect 31294 24148 31300 24200
rect 31352 24188 31358 24200
rect 32401 24191 32459 24197
rect 32401 24188 32413 24191
rect 31352 24160 32413 24188
rect 31352 24148 31358 24160
rect 32401 24157 32413 24160
rect 32447 24188 32459 24191
rect 32582 24188 32588 24200
rect 32447 24160 32588 24188
rect 32447 24157 32459 24160
rect 32401 24151 32459 24157
rect 32582 24148 32588 24160
rect 32640 24148 32646 24200
rect 32686 24188 32714 24228
rect 33106 24228 33860 24256
rect 33106 24188 33134 24228
rect 33848 24225 33860 24228
rect 33894 24256 33906 24259
rect 34238 24256 34244 24268
rect 33894 24228 34244 24256
rect 33894 24225 33906 24228
rect 33848 24219 33906 24225
rect 34238 24216 34244 24228
rect 34296 24216 34302 24268
rect 35802 24216 35808 24268
rect 35860 24256 35866 24268
rect 36354 24256 36360 24268
rect 36412 24265 36418 24268
rect 36412 24259 36450 24265
rect 35860 24228 36360 24256
rect 35860 24216 35866 24228
rect 36354 24216 36360 24228
rect 36438 24256 36450 24259
rect 37642 24256 37648 24268
rect 36438 24228 37648 24256
rect 36438 24225 36450 24228
rect 36412 24219 36450 24225
rect 36412 24216 36418 24219
rect 37642 24216 37648 24228
rect 37700 24216 37706 24268
rect 40144 24265 40172 24296
rect 41141 24293 41153 24296
rect 41187 24324 41199 24327
rect 41322 24324 41328 24336
rect 41187 24296 41328 24324
rect 41187 24293 41199 24296
rect 41141 24287 41199 24293
rect 41322 24284 41328 24296
rect 41380 24284 41386 24336
rect 43533 24327 43591 24333
rect 43533 24293 43545 24327
rect 43579 24324 43591 24327
rect 43622 24324 43628 24336
rect 43579 24296 43628 24324
rect 43579 24293 43591 24296
rect 43533 24287 43591 24293
rect 43622 24284 43628 24296
rect 43680 24284 43686 24336
rect 40129 24259 40187 24265
rect 40129 24225 40141 24259
rect 40175 24225 40187 24259
rect 44910 24256 44916 24268
rect 44871 24228 44916 24256
rect 40129 24219 40187 24225
rect 44910 24216 44916 24228
rect 44968 24216 44974 24268
rect 32686 24160 33134 24188
rect 34885 24191 34943 24197
rect 34885 24157 34897 24191
rect 34931 24157 34943 24191
rect 34885 24151 34943 24157
rect 24964 24120 24992 24148
rect 23446 24092 24992 24120
rect 31113 24123 31171 24129
rect 14829 24083 14887 24089
rect 31113 24089 31125 24123
rect 31159 24120 31171 24123
rect 31570 24120 31576 24132
rect 31159 24092 31576 24120
rect 31159 24089 31171 24092
rect 31113 24083 31171 24089
rect 31570 24080 31576 24092
rect 31628 24120 31634 24132
rect 32674 24120 32680 24132
rect 31628 24092 32680 24120
rect 31628 24080 31634 24092
rect 32674 24080 32680 24092
rect 32732 24080 32738 24132
rect 33919 24123 33977 24129
rect 33919 24089 33931 24123
rect 33965 24120 33977 24123
rect 34900 24120 34928 24151
rect 39114 24148 39120 24200
rect 39172 24188 39178 24200
rect 39209 24191 39267 24197
rect 39209 24188 39221 24191
rect 39172 24160 39221 24188
rect 39172 24148 39178 24160
rect 39209 24157 39221 24160
rect 39255 24157 39267 24191
rect 39209 24151 39267 24157
rect 39758 24148 39764 24200
rect 39816 24188 39822 24200
rect 41049 24191 41107 24197
rect 41049 24188 41061 24191
rect 39816 24160 41061 24188
rect 39816 24148 39822 24160
rect 41049 24157 41061 24160
rect 41095 24188 41107 24191
rect 41506 24188 41512 24200
rect 41095 24160 41512 24188
rect 41095 24157 41107 24160
rect 41049 24151 41107 24157
rect 41506 24148 41512 24160
rect 41564 24148 41570 24200
rect 41693 24191 41751 24197
rect 41693 24157 41705 24191
rect 41739 24188 41751 24191
rect 43254 24188 43260 24200
rect 41739 24160 43260 24188
rect 41739 24157 41751 24160
rect 41693 24151 41751 24157
rect 43254 24148 43260 24160
rect 43312 24148 43318 24200
rect 43438 24188 43444 24200
rect 43399 24160 43444 24188
rect 43438 24148 43444 24160
rect 43496 24148 43502 24200
rect 43717 24191 43775 24197
rect 43717 24188 43729 24191
rect 43548 24160 43729 24188
rect 35250 24120 35256 24132
rect 33965 24092 35256 24120
rect 33965 24089 33977 24092
rect 33919 24083 33977 24089
rect 35250 24080 35256 24092
rect 35308 24080 35314 24132
rect 35434 24120 35440 24132
rect 35395 24092 35440 24120
rect 35434 24080 35440 24092
rect 35492 24080 35498 24132
rect 37553 24123 37611 24129
rect 37553 24089 37565 24123
rect 37599 24120 37611 24123
rect 37642 24120 37648 24132
rect 37599 24092 37648 24120
rect 37599 24089 37611 24092
rect 37553 24083 37611 24089
rect 37642 24080 37648 24092
rect 37700 24080 37706 24132
rect 37875 24123 37933 24129
rect 37875 24089 37887 24123
rect 37921 24120 37933 24123
rect 38102 24120 38108 24132
rect 37921 24092 38108 24120
rect 37921 24089 37933 24092
rect 37875 24083 37933 24089
rect 38102 24080 38108 24092
rect 38160 24120 38166 24132
rect 38565 24123 38623 24129
rect 38565 24120 38577 24123
rect 38160 24092 38577 24120
rect 38160 24080 38166 24092
rect 38565 24089 38577 24092
rect 38611 24089 38623 24123
rect 38565 24083 38623 24089
rect 41874 24080 41880 24132
rect 41932 24120 41938 24132
rect 43548 24120 43576 24160
rect 43717 24157 43729 24160
rect 43763 24188 43775 24191
rect 43806 24188 43812 24200
rect 43763 24160 43812 24188
rect 43763 24157 43775 24160
rect 43717 24151 43775 24157
rect 43806 24148 43812 24160
rect 43864 24148 43870 24200
rect 41932 24092 43576 24120
rect 41932 24080 41938 24092
rect 5074 24052 5080 24064
rect 4276 24024 4476 24052
rect 5035 24024 5080 24052
rect 4276 24021 4288 24024
rect 4230 24015 4288 24021
rect 5074 24012 5080 24024
rect 5132 24012 5138 24064
rect 7101 24055 7159 24061
rect 7101 24021 7113 24055
rect 7147 24052 7159 24055
rect 7650 24052 7656 24064
rect 7147 24024 7656 24052
rect 7147 24021 7159 24024
rect 7101 24015 7159 24021
rect 7650 24012 7656 24024
rect 7708 24012 7714 24064
rect 8754 24052 8760 24064
rect 8715 24024 8760 24052
rect 8754 24012 8760 24024
rect 8812 24012 8818 24064
rect 9122 24052 9128 24064
rect 9083 24024 9128 24052
rect 9122 24012 9128 24024
rect 9180 24012 9186 24064
rect 13541 24055 13599 24061
rect 13541 24021 13553 24055
rect 13587 24052 13599 24055
rect 14458 24052 14464 24064
rect 13587 24024 14464 24052
rect 13587 24021 13599 24024
rect 13541 24015 13599 24021
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 16206 24052 16212 24064
rect 16167 24024 16212 24052
rect 16206 24012 16212 24024
rect 16264 24012 16270 24064
rect 23842 24052 23848 24064
rect 23803 24024 23848 24052
rect 23842 24012 23848 24024
rect 23900 24012 23906 24064
rect 26694 24052 26700 24064
rect 26655 24024 26700 24052
rect 26694 24012 26700 24024
rect 26752 24012 26758 24064
rect 27062 24052 27068 24064
rect 27023 24024 27068 24052
rect 27062 24012 27068 24024
rect 27120 24012 27126 24064
rect 29086 24012 29092 24064
rect 29144 24052 29150 24064
rect 29273 24055 29331 24061
rect 29273 24052 29285 24055
rect 29144 24024 29285 24052
rect 29144 24012 29150 24024
rect 29273 24021 29285 24024
rect 29319 24021 29331 24055
rect 31478 24052 31484 24064
rect 31439 24024 31484 24052
rect 29273 24015 29331 24021
rect 31478 24012 31484 24024
rect 31536 24012 31542 24064
rect 36495 24055 36553 24061
rect 36495 24021 36507 24055
rect 36541 24052 36553 24055
rect 36630 24052 36636 24064
rect 36541 24024 36636 24052
rect 36541 24021 36553 24024
rect 36495 24015 36553 24021
rect 36630 24012 36636 24024
rect 36688 24012 36694 24064
rect 36906 24052 36912 24064
rect 36819 24024 36912 24052
rect 36906 24012 36912 24024
rect 36964 24052 36970 24064
rect 38194 24052 38200 24064
rect 36964 24024 38200 24052
rect 36964 24012 36970 24024
rect 38194 24012 38200 24024
rect 38252 24012 38258 24064
rect 1104 23962 48852 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 48852 23962
rect 1104 23888 48852 23910
rect 2406 23848 2412 23860
rect 2367 23820 2412 23848
rect 2406 23808 2412 23820
rect 2464 23848 2470 23860
rect 2777 23851 2835 23857
rect 2777 23848 2789 23851
rect 2464 23820 2789 23848
rect 2464 23808 2470 23820
rect 2777 23817 2789 23820
rect 2823 23817 2835 23851
rect 3418 23848 3424 23860
rect 3379 23820 3424 23848
rect 2777 23811 2835 23817
rect 2792 23712 2820 23811
rect 3418 23808 3424 23820
rect 3476 23808 3482 23860
rect 3970 23808 3976 23860
rect 4028 23848 4034 23860
rect 4157 23851 4215 23857
rect 4157 23848 4169 23851
rect 4028 23820 4169 23848
rect 4028 23808 4034 23820
rect 4157 23817 4169 23820
rect 4203 23848 4215 23851
rect 7377 23851 7435 23857
rect 7377 23848 7389 23851
rect 4203 23820 7389 23848
rect 4203 23817 4215 23820
rect 4157 23811 4215 23817
rect 7377 23817 7389 23820
rect 7423 23848 7435 23851
rect 7837 23851 7895 23857
rect 7837 23848 7849 23851
rect 7423 23820 7849 23848
rect 7423 23817 7435 23820
rect 7377 23811 7435 23817
rect 7837 23817 7849 23820
rect 7883 23848 7895 23851
rect 8110 23848 8116 23860
rect 7883 23820 8116 23848
rect 7883 23817 7895 23820
rect 7837 23811 7895 23817
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 8570 23848 8576 23860
rect 8531 23820 8576 23848
rect 8570 23808 8576 23820
rect 8628 23808 8634 23860
rect 11054 23808 11060 23860
rect 11112 23848 11118 23860
rect 11517 23851 11575 23857
rect 11517 23848 11529 23851
rect 11112 23820 11529 23848
rect 11112 23808 11118 23820
rect 11517 23817 11529 23820
rect 11563 23817 11575 23851
rect 11517 23811 11575 23817
rect 12253 23851 12311 23857
rect 12253 23817 12265 23851
rect 12299 23848 12311 23851
rect 12434 23848 12440 23860
rect 12299 23820 12440 23848
rect 12299 23817 12311 23820
rect 12253 23811 12311 23817
rect 12434 23808 12440 23820
rect 12492 23848 12498 23860
rect 13449 23851 13507 23857
rect 13449 23848 13461 23851
rect 12492 23820 13461 23848
rect 12492 23808 12498 23820
rect 13449 23817 13461 23820
rect 13495 23848 13507 23851
rect 13814 23848 13820 23860
rect 13495 23820 13820 23848
rect 13495 23817 13507 23820
rect 13449 23811 13507 23817
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 14734 23848 14740 23860
rect 14695 23820 14740 23848
rect 14734 23808 14740 23820
rect 14792 23848 14798 23860
rect 15013 23851 15071 23857
rect 15013 23848 15025 23851
rect 14792 23820 15025 23848
rect 14792 23808 14798 23820
rect 15013 23817 15025 23820
rect 15059 23817 15071 23851
rect 15013 23811 15071 23817
rect 15286 23808 15292 23860
rect 15344 23848 15350 23860
rect 16393 23851 16451 23857
rect 16393 23848 16405 23851
rect 15344 23820 16405 23848
rect 15344 23808 15350 23820
rect 16393 23817 16405 23820
rect 16439 23817 16451 23851
rect 16393 23811 16451 23817
rect 17402 23808 17408 23860
rect 17460 23848 17466 23860
rect 17773 23851 17831 23857
rect 17773 23848 17785 23851
rect 17460 23820 17785 23848
rect 17460 23808 17466 23820
rect 17773 23817 17785 23820
rect 17819 23817 17831 23851
rect 17773 23811 17831 23817
rect 3142 23740 3148 23792
rect 3200 23780 3206 23792
rect 3237 23783 3295 23789
rect 3237 23780 3249 23783
rect 3200 23752 3249 23780
rect 3200 23740 3206 23752
rect 3237 23749 3249 23752
rect 3283 23780 3295 23783
rect 4062 23780 4068 23792
rect 3283 23752 4068 23780
rect 3283 23749 3295 23752
rect 3237 23743 3295 23749
rect 4062 23740 4068 23752
rect 4120 23780 4126 23792
rect 4341 23783 4399 23789
rect 4341 23780 4353 23783
rect 4120 23752 4353 23780
rect 4120 23740 4126 23752
rect 4341 23749 4353 23752
rect 4387 23749 4399 23783
rect 4341 23743 4399 23749
rect 5077 23783 5135 23789
rect 5077 23749 5089 23783
rect 5123 23780 5135 23783
rect 5166 23780 5172 23792
rect 5123 23752 5172 23780
rect 5123 23749 5135 23752
rect 5077 23743 5135 23749
rect 5166 23740 5172 23752
rect 5224 23780 5230 23792
rect 5718 23780 5724 23792
rect 5224 23752 5724 23780
rect 5224 23740 5230 23752
rect 5718 23740 5724 23752
rect 5776 23740 5782 23792
rect 15304 23780 15332 23808
rect 14384 23752 15332 23780
rect 3329 23715 3387 23721
rect 3329 23712 3341 23715
rect 1964 23684 3341 23712
rect 1964 23653 1992 23684
rect 3329 23681 3341 23684
rect 3375 23712 3387 23715
rect 4433 23715 4491 23721
rect 4433 23712 4445 23715
rect 3375 23684 4445 23712
rect 3375 23681 3387 23684
rect 3329 23675 3387 23681
rect 4433 23681 4445 23684
rect 4479 23712 4491 23715
rect 4614 23712 4620 23724
rect 4479 23684 4620 23712
rect 4479 23681 4491 23684
rect 4433 23675 4491 23681
rect 4614 23672 4620 23684
rect 4672 23672 4678 23724
rect 5626 23672 5632 23724
rect 5684 23712 5690 23724
rect 7742 23721 7748 23724
rect 7009 23715 7067 23721
rect 7009 23712 7021 23715
rect 5684 23684 7021 23712
rect 5684 23672 5690 23684
rect 7009 23681 7021 23684
rect 7055 23712 7067 23715
rect 7708 23715 7748 23721
rect 7708 23712 7720 23715
rect 7055 23684 7720 23712
rect 7055 23681 7067 23684
rect 7009 23675 7067 23681
rect 7708 23681 7720 23684
rect 7708 23675 7748 23681
rect 7742 23672 7748 23675
rect 7800 23672 7806 23724
rect 7834 23672 7840 23724
rect 7892 23712 7898 23724
rect 7929 23715 7987 23721
rect 7929 23712 7941 23715
rect 7892 23684 7941 23712
rect 7892 23672 7898 23684
rect 7929 23681 7941 23684
rect 7975 23681 7987 23715
rect 8938 23712 8944 23724
rect 8899 23684 8944 23712
rect 7929 23675 7987 23681
rect 8938 23672 8944 23684
rect 8996 23712 9002 23724
rect 9861 23715 9919 23721
rect 8996 23684 9444 23712
rect 8996 23672 9002 23684
rect 1949 23647 2007 23653
rect 1949 23613 1961 23647
rect 1995 23613 2007 23647
rect 2958 23644 2964 23656
rect 2919 23616 2964 23644
rect 1949 23607 2007 23613
rect 2958 23604 2964 23616
rect 3016 23604 3022 23656
rect 3108 23647 3166 23653
rect 3108 23613 3120 23647
rect 3154 23644 3166 23647
rect 4985 23647 5043 23653
rect 4985 23644 4997 23647
rect 3154 23616 4997 23644
rect 3154 23613 3166 23616
rect 3108 23607 3166 23613
rect 3344 23588 3372 23616
rect 4985 23613 4997 23616
rect 5031 23644 5043 23647
rect 5074 23644 5080 23656
rect 5031 23616 5080 23644
rect 5031 23613 5043 23616
rect 4985 23607 5043 23613
rect 5074 23604 5080 23616
rect 5132 23604 5138 23656
rect 5258 23644 5264 23656
rect 5219 23616 5264 23644
rect 5258 23604 5264 23616
rect 5316 23604 5322 23656
rect 5534 23604 5540 23656
rect 5592 23644 5598 23656
rect 6638 23644 6644 23656
rect 5592 23616 6644 23644
rect 5592 23604 5598 23616
rect 6638 23604 6644 23616
rect 6696 23604 6702 23656
rect 6730 23604 6736 23656
rect 6788 23644 6794 23656
rect 7558 23644 7564 23656
rect 6788 23616 7564 23644
rect 6788 23604 6794 23616
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 8386 23604 8392 23656
rect 8444 23644 8450 23656
rect 9122 23644 9128 23656
rect 8444 23616 9128 23644
rect 8444 23604 8450 23616
rect 9122 23604 9128 23616
rect 9180 23604 9186 23656
rect 9214 23604 9220 23656
rect 9272 23644 9278 23656
rect 9416 23653 9444 23684
rect 9861 23681 9873 23715
rect 9907 23712 9919 23715
rect 10134 23712 10140 23724
rect 9907 23684 10140 23712
rect 9907 23681 9919 23684
rect 9861 23675 9919 23681
rect 10134 23672 10140 23684
rect 10192 23672 10198 23724
rect 14384 23721 14412 23752
rect 10229 23715 10287 23721
rect 10229 23681 10241 23715
rect 10275 23712 10287 23715
rect 14369 23715 14427 23721
rect 10275 23684 11284 23712
rect 10275 23681 10287 23684
rect 10229 23675 10287 23681
rect 11256 23656 11284 23684
rect 14369 23681 14381 23715
rect 14415 23681 14427 23715
rect 14369 23675 14427 23681
rect 14918 23672 14924 23724
rect 14976 23712 14982 23724
rect 15197 23715 15255 23721
rect 15197 23712 15209 23715
rect 14976 23684 15209 23712
rect 14976 23672 14982 23684
rect 15197 23681 15209 23684
rect 15243 23681 15255 23715
rect 15197 23675 15255 23681
rect 9401 23647 9459 23653
rect 9272 23616 9317 23644
rect 9272 23604 9278 23616
rect 9401 23613 9413 23647
rect 9447 23644 9459 23647
rect 9490 23644 9496 23656
rect 9447 23616 9496 23644
rect 9447 23613 9459 23616
rect 9401 23607 9459 23613
rect 9490 23604 9496 23616
rect 9548 23604 9554 23656
rect 10778 23604 10784 23656
rect 10836 23644 10842 23656
rect 10873 23647 10931 23653
rect 10873 23644 10885 23647
rect 10836 23616 10885 23644
rect 10836 23604 10842 23616
rect 10873 23613 10885 23616
rect 10919 23613 10931 23647
rect 11238 23644 11244 23656
rect 11151 23616 11244 23644
rect 10873 23607 10931 23613
rect 11238 23604 11244 23616
rect 11296 23644 11302 23656
rect 12437 23647 12495 23653
rect 12437 23644 12449 23647
rect 11296 23616 12449 23644
rect 11296 23604 11302 23616
rect 12437 23613 12449 23616
rect 12483 23644 12495 23647
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12483 23616 12909 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 12897 23613 12909 23616
rect 12943 23613 12955 23647
rect 12897 23607 12955 23613
rect 13633 23647 13691 23653
rect 13633 23613 13645 23647
rect 13679 23613 13691 23647
rect 13633 23607 13691 23613
rect 3326 23536 3332 23588
rect 3384 23536 3390 23588
rect 4246 23536 4252 23588
rect 4304 23576 4310 23588
rect 5721 23579 5779 23585
rect 5721 23576 5733 23579
rect 4304 23548 5733 23576
rect 4304 23536 4310 23548
rect 5721 23545 5733 23548
rect 5767 23576 5779 23579
rect 7098 23576 7104 23588
rect 5767 23548 7104 23576
rect 5767 23545 5779 23548
rect 5721 23539 5779 23545
rect 7098 23536 7104 23548
rect 7156 23536 7162 23588
rect 8294 23576 8300 23588
rect 8255 23548 8300 23576
rect 8294 23536 8300 23548
rect 8352 23536 8358 23588
rect 10689 23579 10747 23585
rect 10689 23545 10701 23579
rect 10735 23545 10747 23579
rect 13648 23576 13676 23607
rect 13722 23604 13728 23656
rect 13780 23644 13786 23656
rect 14093 23647 14151 23653
rect 14093 23644 14105 23647
rect 13780 23616 14105 23644
rect 13780 23604 13786 23616
rect 14093 23613 14105 23616
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 16117 23647 16175 23653
rect 16117 23613 16129 23647
rect 16163 23644 16175 23647
rect 16761 23647 16819 23653
rect 16761 23644 16773 23647
rect 16163 23616 16773 23644
rect 16163 23613 16175 23616
rect 16117 23607 16175 23613
rect 16761 23613 16773 23616
rect 16807 23644 16819 23647
rect 16980 23647 17038 23653
rect 16980 23644 16992 23647
rect 16807 23616 16992 23644
rect 16807 23613 16819 23616
rect 16761 23607 16819 23613
rect 16980 23613 16992 23616
rect 17026 23613 17038 23647
rect 17788 23644 17816 23811
rect 17954 23808 17960 23860
rect 18012 23848 18018 23860
rect 19797 23851 19855 23857
rect 19797 23848 19809 23851
rect 18012 23820 19809 23848
rect 18012 23808 18018 23820
rect 19797 23817 19809 23820
rect 19843 23817 19855 23851
rect 19797 23811 19855 23817
rect 22465 23851 22523 23857
rect 22465 23817 22477 23851
rect 22511 23848 22523 23851
rect 22830 23848 22836 23860
rect 22511 23820 22836 23848
rect 22511 23817 22523 23820
rect 22465 23811 22523 23817
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 25593 23851 25651 23857
rect 25593 23817 25605 23851
rect 25639 23848 25651 23851
rect 27798 23848 27804 23860
rect 25639 23820 27804 23848
rect 25639 23817 25651 23820
rect 25593 23811 25651 23817
rect 19058 23780 19064 23792
rect 19019 23752 19064 23780
rect 19058 23740 19064 23752
rect 19116 23740 19122 23792
rect 25130 23780 25136 23792
rect 25091 23752 25136 23780
rect 25130 23740 25136 23752
rect 25188 23740 25194 23792
rect 21174 23712 21180 23724
rect 21135 23684 21180 23712
rect 21174 23672 21180 23684
rect 21232 23672 21238 23724
rect 24581 23715 24639 23721
rect 24581 23681 24593 23715
rect 24627 23712 24639 23715
rect 25608 23712 25636 23811
rect 27798 23808 27804 23820
rect 27856 23808 27862 23860
rect 27982 23808 27988 23860
rect 28040 23848 28046 23860
rect 28350 23848 28356 23860
rect 28040 23820 28356 23848
rect 28040 23808 28046 23820
rect 28350 23808 28356 23820
rect 28408 23808 28414 23860
rect 28902 23808 28908 23860
rect 28960 23848 28966 23860
rect 30929 23851 30987 23857
rect 30929 23848 30941 23851
rect 28960 23820 30941 23848
rect 28960 23808 28966 23820
rect 30929 23817 30941 23820
rect 30975 23848 30987 23851
rect 31021 23851 31079 23857
rect 31021 23848 31033 23851
rect 30975 23820 31033 23848
rect 30975 23817 30987 23820
rect 30929 23811 30987 23817
rect 31021 23817 31033 23820
rect 31067 23848 31079 23851
rect 31202 23848 31208 23860
rect 31067 23820 31208 23848
rect 31067 23817 31079 23820
rect 31021 23811 31079 23817
rect 31202 23808 31208 23820
rect 31260 23808 31266 23860
rect 31386 23808 31392 23860
rect 31444 23848 31450 23860
rect 34238 23848 34244 23860
rect 31444 23820 33134 23848
rect 34199 23820 34244 23848
rect 31444 23808 31450 23820
rect 26237 23783 26295 23789
rect 26237 23749 26249 23783
rect 26283 23780 26295 23783
rect 26510 23780 26516 23792
rect 26283 23752 26516 23780
rect 26283 23749 26295 23752
rect 26237 23743 26295 23749
rect 26510 23740 26516 23752
rect 26568 23740 26574 23792
rect 27338 23740 27344 23792
rect 27396 23780 27402 23792
rect 30331 23783 30389 23789
rect 27396 23752 28028 23780
rect 27396 23740 27402 23752
rect 24627 23684 25636 23712
rect 24627 23681 24639 23684
rect 24581 23675 24639 23681
rect 18141 23647 18199 23653
rect 18141 23644 18153 23647
rect 17788 23616 18153 23644
rect 16980 23607 17038 23613
rect 18141 23613 18153 23616
rect 18187 23613 18199 23647
rect 18141 23607 18199 23613
rect 18782 23604 18788 23656
rect 18840 23644 18846 23656
rect 19613 23647 19671 23653
rect 19613 23644 19625 23647
rect 18840 23616 19625 23644
rect 18840 23604 18846 23616
rect 19613 23613 19625 23616
rect 19659 23644 19671 23647
rect 20073 23647 20131 23653
rect 20073 23644 20085 23647
rect 19659 23616 20085 23644
rect 19659 23613 19671 23616
rect 19613 23607 19671 23613
rect 20073 23613 20085 23616
rect 20119 23644 20131 23647
rect 20162 23644 20168 23656
rect 20119 23616 20168 23644
rect 20119 23613 20131 23616
rect 20073 23607 20131 23613
rect 20162 23604 20168 23616
rect 20220 23604 20226 23656
rect 22624 23647 22682 23653
rect 22624 23613 22636 23647
rect 22670 23644 22682 23647
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22670 23616 23029 23644
rect 22670 23613 22682 23616
rect 22624 23607 22682 23613
rect 23017 23613 23029 23616
rect 23063 23644 23075 23647
rect 23106 23644 23112 23656
rect 23063 23616 23112 23644
rect 23063 23613 23075 23616
rect 23017 23607 23075 23613
rect 23106 23604 23112 23616
rect 23164 23604 23170 23656
rect 26528 23644 26556 23740
rect 28000 23724 28028 23752
rect 30331 23749 30343 23783
rect 30377 23780 30389 23783
rect 30558 23780 30564 23792
rect 30377 23752 30564 23780
rect 30377 23749 30389 23752
rect 30331 23743 30389 23749
rect 30558 23740 30564 23752
rect 30616 23780 30622 23792
rect 32217 23783 32275 23789
rect 32217 23780 32229 23783
rect 30616 23752 32229 23780
rect 30616 23740 30622 23752
rect 32217 23749 32229 23752
rect 32263 23749 32275 23783
rect 32217 23743 32275 23749
rect 32398 23740 32404 23792
rect 32456 23780 32462 23792
rect 32769 23783 32827 23789
rect 32769 23780 32781 23783
rect 32456 23752 32781 23780
rect 32456 23740 32462 23752
rect 32769 23749 32781 23752
rect 32815 23749 32827 23783
rect 33106 23780 33134 23820
rect 34238 23808 34244 23820
rect 34296 23808 34302 23860
rect 34606 23848 34612 23860
rect 34567 23820 34612 23848
rect 34606 23808 34612 23820
rect 34664 23808 34670 23860
rect 36354 23848 36360 23860
rect 36315 23820 36360 23848
rect 36354 23808 36360 23820
rect 36412 23808 36418 23860
rect 37642 23848 37648 23860
rect 37384 23820 37648 23848
rect 37384 23780 37412 23820
rect 37642 23808 37648 23820
rect 37700 23848 37706 23860
rect 37737 23851 37795 23857
rect 37737 23848 37749 23851
rect 37700 23820 37749 23848
rect 37700 23808 37706 23820
rect 37737 23817 37749 23820
rect 37783 23848 37795 23851
rect 41414 23848 41420 23860
rect 37783 23820 41420 23848
rect 37783 23817 37795 23820
rect 37737 23811 37795 23817
rect 41414 23808 41420 23820
rect 41472 23808 41478 23860
rect 41506 23808 41512 23860
rect 41564 23848 41570 23860
rect 41969 23851 42027 23857
rect 41969 23848 41981 23851
rect 41564 23820 41981 23848
rect 41564 23808 41570 23820
rect 41969 23817 41981 23820
rect 42015 23817 42027 23851
rect 41969 23811 42027 23817
rect 42058 23808 42064 23860
rect 42116 23848 42122 23860
rect 42518 23848 42524 23860
rect 42116 23820 42524 23848
rect 42116 23808 42122 23820
rect 42518 23808 42524 23820
rect 42576 23848 42582 23860
rect 42576 23820 44220 23848
rect 42576 23808 42582 23820
rect 33106 23752 37412 23780
rect 32769 23743 32827 23749
rect 27982 23712 27988 23724
rect 27895 23684 27988 23712
rect 27982 23672 27988 23684
rect 28040 23672 28046 23724
rect 31297 23715 31355 23721
rect 31297 23681 31309 23715
rect 31343 23712 31355 23715
rect 31478 23712 31484 23724
rect 31343 23684 31484 23712
rect 31343 23681 31355 23684
rect 31297 23675 31355 23681
rect 31478 23672 31484 23684
rect 31536 23672 31542 23724
rect 31570 23672 31576 23724
rect 31628 23712 31634 23724
rect 32784 23712 32812 23743
rect 37458 23740 37464 23792
rect 37516 23780 37522 23792
rect 42613 23783 42671 23789
rect 37516 23752 38424 23780
rect 37516 23740 37522 23752
rect 34606 23712 34612 23724
rect 31628 23684 31673 23712
rect 32784 23684 34612 23712
rect 31628 23672 31634 23684
rect 34606 23672 34612 23684
rect 34664 23672 34670 23724
rect 35434 23712 35440 23724
rect 35395 23684 35440 23712
rect 35434 23672 35440 23684
rect 35492 23672 35498 23724
rect 36541 23715 36599 23721
rect 36541 23681 36553 23715
rect 36587 23712 36599 23715
rect 36630 23712 36636 23724
rect 36587 23684 36636 23712
rect 36587 23681 36599 23684
rect 36541 23675 36599 23681
rect 36630 23672 36636 23684
rect 36688 23672 36694 23724
rect 38102 23712 38108 23724
rect 38063 23684 38108 23712
rect 38102 23672 38108 23684
rect 38160 23672 38166 23724
rect 38396 23721 38424 23752
rect 42613 23749 42625 23783
rect 42659 23780 42671 23783
rect 43438 23780 43444 23792
rect 42659 23752 43444 23780
rect 42659 23749 42671 23752
rect 42613 23743 42671 23749
rect 43438 23740 43444 23752
rect 43496 23740 43502 23792
rect 38381 23715 38439 23721
rect 38381 23681 38393 23715
rect 38427 23681 38439 23715
rect 38381 23675 38439 23681
rect 38562 23672 38568 23724
rect 38620 23712 38626 23724
rect 39114 23712 39120 23724
rect 38620 23684 39120 23712
rect 38620 23672 38626 23684
rect 39114 23672 39120 23684
rect 39172 23712 39178 23724
rect 39577 23715 39635 23721
rect 39577 23712 39589 23715
rect 39172 23684 39589 23712
rect 39172 23672 39178 23684
rect 39577 23681 39589 23684
rect 39623 23681 39635 23715
rect 39577 23675 39635 23681
rect 40313 23715 40371 23721
rect 40313 23681 40325 23715
rect 40359 23712 40371 23715
rect 41049 23715 41107 23721
rect 41049 23712 41061 23715
rect 40359 23684 41061 23712
rect 40359 23681 40371 23684
rect 40313 23675 40371 23681
rect 41049 23681 41061 23684
rect 41095 23712 41107 23715
rect 41138 23712 41144 23724
rect 41095 23684 41144 23712
rect 41095 23681 41107 23684
rect 41049 23675 41107 23681
rect 41138 23672 41144 23684
rect 41196 23672 41202 23724
rect 43162 23712 43168 23724
rect 43123 23684 43168 23712
rect 43162 23672 43168 23684
rect 43220 23672 43226 23724
rect 43254 23672 43260 23724
rect 43312 23712 43318 23724
rect 43533 23715 43591 23721
rect 43533 23712 43545 23715
rect 43312 23684 43545 23712
rect 43312 23672 43318 23684
rect 43533 23681 43545 23684
rect 43579 23681 43591 23715
rect 43533 23675 43591 23681
rect 26697 23647 26755 23653
rect 26697 23644 26709 23647
rect 26528 23616 26709 23644
rect 26697 23613 26709 23616
rect 26743 23613 26755 23647
rect 26697 23607 26755 23613
rect 27062 23604 27068 23656
rect 27120 23644 27126 23656
rect 27157 23647 27215 23653
rect 27157 23644 27169 23647
rect 27120 23616 27169 23644
rect 27120 23604 27126 23616
rect 27157 23613 27169 23616
rect 27203 23644 27215 23647
rect 27338 23644 27344 23656
rect 27203 23616 27344 23644
rect 27203 23613 27215 23616
rect 27157 23607 27215 23613
rect 27338 23604 27344 23616
rect 27396 23604 27402 23656
rect 28810 23604 28816 23656
rect 28868 23644 28874 23656
rect 30228 23647 30286 23653
rect 30228 23644 30240 23647
rect 28868 23616 30240 23644
rect 28868 23604 28874 23616
rect 30228 23613 30240 23616
rect 30274 23644 30286 23647
rect 30653 23647 30711 23653
rect 30653 23644 30665 23647
rect 30274 23616 30665 23644
rect 30274 23613 30286 23616
rect 30228 23607 30286 23613
rect 30653 23613 30665 23616
rect 30699 23644 30711 23647
rect 30834 23644 30840 23656
rect 30699 23616 30840 23644
rect 30699 23613 30711 23616
rect 30653 23607 30711 23613
rect 30834 23604 30840 23616
rect 30892 23604 30898 23656
rect 44192 23644 44220 23820
rect 44910 23808 44916 23860
rect 44968 23848 44974 23860
rect 45462 23848 45468 23860
rect 44968 23820 45468 23848
rect 44968 23808 44974 23820
rect 45462 23808 45468 23820
rect 45520 23808 45526 23860
rect 44672 23647 44730 23653
rect 44672 23644 44684 23647
rect 44192 23616 44684 23644
rect 44672 23613 44684 23616
rect 44718 23644 44730 23647
rect 45097 23647 45155 23653
rect 45097 23644 45109 23647
rect 44718 23616 45109 23644
rect 44718 23613 44730 23616
rect 44672 23607 44730 23613
rect 45097 23613 45109 23616
rect 45143 23613 45155 23647
rect 45097 23607 45155 23613
rect 13814 23576 13820 23588
rect 10689 23539 10747 23545
rect 12820 23548 13584 23576
rect 13648 23548 13820 23576
rect 1486 23468 1492 23520
rect 1544 23508 1550 23520
rect 1765 23511 1823 23517
rect 1765 23508 1777 23511
rect 1544 23480 1777 23508
rect 1544 23468 1550 23480
rect 1765 23477 1777 23480
rect 1811 23477 1823 23511
rect 1765 23471 1823 23477
rect 2133 23511 2191 23517
rect 2133 23477 2145 23511
rect 2179 23508 2191 23511
rect 2314 23508 2320 23520
rect 2179 23480 2320 23508
rect 2179 23477 2191 23480
rect 2133 23471 2191 23477
rect 2314 23468 2320 23480
rect 2372 23468 2378 23520
rect 4341 23511 4399 23517
rect 4341 23477 4353 23511
rect 4387 23508 4399 23511
rect 4801 23511 4859 23517
rect 4801 23508 4813 23511
rect 4387 23480 4813 23508
rect 4387 23477 4399 23480
rect 4341 23471 4399 23477
rect 4801 23477 4813 23480
rect 4847 23508 4859 23511
rect 4890 23508 4896 23520
rect 4847 23480 4896 23508
rect 4847 23477 4859 23480
rect 4801 23471 4859 23477
rect 4890 23468 4896 23480
rect 4948 23468 4954 23520
rect 5074 23468 5080 23520
rect 5132 23508 5138 23520
rect 5902 23508 5908 23520
rect 5132 23480 5908 23508
rect 5132 23468 5138 23480
rect 5902 23468 5908 23480
rect 5960 23468 5966 23520
rect 5994 23468 6000 23520
rect 6052 23508 6058 23520
rect 6638 23508 6644 23520
rect 6052 23480 6097 23508
rect 6599 23480 6644 23508
rect 6052 23468 6058 23480
rect 6638 23468 6644 23480
rect 6696 23468 6702 23520
rect 10226 23468 10232 23520
rect 10284 23508 10290 23520
rect 10505 23511 10563 23517
rect 10505 23508 10517 23511
rect 10284 23480 10517 23508
rect 10284 23468 10290 23480
rect 10505 23477 10517 23480
rect 10551 23508 10563 23511
rect 10704 23508 10732 23539
rect 10551 23480 10732 23508
rect 12621 23511 12679 23517
rect 10551 23477 10563 23480
rect 10505 23471 10563 23477
rect 12621 23477 12633 23511
rect 12667 23508 12679 23511
rect 12820 23508 12848 23548
rect 12667 23480 12848 23508
rect 13556 23508 13584 23548
rect 13814 23536 13820 23548
rect 13872 23576 13878 23588
rect 14550 23576 14556 23588
rect 13872 23548 14556 23576
rect 13872 23536 13878 23548
rect 14550 23536 14556 23548
rect 14608 23536 14614 23588
rect 14734 23536 14740 23588
rect 14792 23576 14798 23588
rect 15518 23579 15576 23585
rect 15518 23576 15530 23579
rect 14792 23548 15530 23576
rect 14792 23536 14798 23548
rect 15518 23545 15530 23548
rect 15564 23576 15576 23579
rect 15654 23576 15660 23588
rect 15564 23548 15660 23576
rect 15564 23545 15576 23548
rect 15518 23539 15576 23545
rect 15654 23536 15660 23548
rect 15712 23536 15718 23588
rect 17083 23579 17141 23585
rect 17083 23545 17095 23579
rect 17129 23576 17141 23579
rect 18230 23576 18236 23588
rect 17129 23548 18236 23576
rect 17129 23545 17141 23548
rect 17083 23539 17141 23545
rect 18230 23536 18236 23548
rect 18288 23536 18294 23588
rect 20714 23576 20720 23588
rect 20675 23548 20720 23576
rect 20714 23536 20720 23548
rect 20772 23536 20778 23588
rect 20809 23579 20867 23585
rect 20809 23545 20821 23579
rect 20855 23545 20867 23579
rect 20809 23539 20867 23545
rect 24673 23579 24731 23585
rect 24673 23545 24685 23579
rect 24719 23576 24731 23579
rect 24762 23576 24768 23588
rect 24719 23548 24768 23576
rect 24719 23545 24731 23548
rect 24673 23539 24731 23545
rect 17402 23508 17408 23520
rect 13556 23480 17408 23508
rect 12667 23477 12679 23480
rect 12621 23471 12679 23477
rect 17402 23468 17408 23480
rect 17460 23468 17466 23520
rect 17497 23511 17555 23517
rect 17497 23477 17509 23511
rect 17543 23508 17555 23511
rect 17954 23508 17960 23520
rect 17543 23480 17960 23508
rect 17543 23477 17555 23480
rect 17497 23471 17555 23477
rect 17954 23468 17960 23480
rect 18012 23468 18018 23520
rect 18509 23511 18567 23517
rect 18509 23477 18521 23511
rect 18555 23508 18567 23511
rect 18598 23508 18604 23520
rect 18555 23480 18604 23508
rect 18555 23477 18567 23480
rect 18509 23471 18567 23477
rect 18598 23468 18604 23480
rect 18656 23468 18662 23520
rect 20533 23511 20591 23517
rect 20533 23477 20545 23511
rect 20579 23508 20591 23511
rect 20824 23508 20852 23539
rect 21082 23508 21088 23520
rect 20579 23480 21088 23508
rect 20579 23477 20591 23480
rect 20533 23471 20591 23477
rect 21082 23468 21088 23480
rect 21140 23508 21146 23520
rect 21637 23511 21695 23517
rect 21637 23508 21649 23511
rect 21140 23480 21649 23508
rect 21140 23468 21146 23480
rect 21637 23477 21649 23480
rect 21683 23477 21695 23511
rect 21637 23471 21695 23477
rect 22695 23511 22753 23517
rect 22695 23477 22707 23511
rect 22741 23508 22753 23511
rect 22830 23508 22836 23520
rect 22741 23480 22836 23508
rect 22741 23477 22753 23480
rect 22695 23471 22753 23477
rect 22830 23468 22836 23480
rect 22888 23468 22894 23520
rect 23477 23511 23535 23517
rect 23477 23477 23489 23511
rect 23523 23508 23535 23511
rect 23842 23508 23848 23520
rect 23523 23480 23848 23508
rect 23523 23477 23535 23480
rect 23477 23471 23535 23477
rect 23842 23468 23848 23480
rect 23900 23468 23906 23520
rect 24029 23511 24087 23517
rect 24029 23477 24041 23511
rect 24075 23508 24087 23511
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 24075 23480 24409 23508
rect 24075 23477 24087 23480
rect 24029 23471 24087 23477
rect 24397 23477 24409 23480
rect 24443 23508 24455 23511
rect 24688 23508 24716 23539
rect 24762 23536 24768 23548
rect 24820 23536 24826 23588
rect 27430 23576 27436 23588
rect 27391 23548 27436 23576
rect 27430 23536 27436 23548
rect 27488 23536 27494 23588
rect 30929 23579 30987 23585
rect 30929 23545 30941 23579
rect 30975 23576 30987 23579
rect 31389 23579 31447 23585
rect 31389 23576 31401 23579
rect 30975 23548 31401 23576
rect 30975 23545 30987 23548
rect 30929 23539 30987 23545
rect 31389 23545 31401 23548
rect 31435 23545 31447 23579
rect 33318 23576 33324 23588
rect 33279 23548 33324 23576
rect 31389 23539 31447 23545
rect 33318 23536 33324 23548
rect 33376 23536 33382 23588
rect 33410 23536 33416 23588
rect 33468 23576 33474 23588
rect 33965 23579 34023 23585
rect 33468 23548 33513 23576
rect 33468 23536 33474 23548
rect 33965 23545 33977 23579
rect 34011 23576 34023 23579
rect 34146 23576 34152 23588
rect 34011 23548 34152 23576
rect 34011 23545 34023 23548
rect 33965 23539 34023 23545
rect 34146 23536 34152 23548
rect 34204 23536 34210 23588
rect 34790 23536 34796 23588
rect 34848 23576 34854 23588
rect 34977 23579 35035 23585
rect 34977 23576 34989 23579
rect 34848 23548 34989 23576
rect 34848 23536 34854 23548
rect 34977 23545 34989 23548
rect 35023 23545 35035 23579
rect 34977 23539 35035 23545
rect 35069 23579 35127 23585
rect 35069 23545 35081 23579
rect 35115 23545 35127 23579
rect 35069 23539 35127 23545
rect 36633 23579 36691 23585
rect 36633 23545 36645 23579
rect 36679 23545 36691 23579
rect 36633 23539 36691 23545
rect 37185 23579 37243 23585
rect 37185 23545 37197 23579
rect 37231 23576 37243 23579
rect 37458 23576 37464 23588
rect 37231 23548 37464 23576
rect 37231 23545 37243 23548
rect 37185 23539 37243 23545
rect 29730 23508 29736 23520
rect 24443 23480 24716 23508
rect 29691 23480 29736 23508
rect 24443 23477 24455 23480
rect 24397 23471 24455 23477
rect 29730 23468 29736 23480
rect 29788 23468 29794 23520
rect 30834 23468 30840 23520
rect 30892 23508 30898 23520
rect 34330 23508 34336 23520
rect 30892 23480 34336 23508
rect 30892 23468 30898 23480
rect 34330 23468 34336 23480
rect 34388 23468 34394 23520
rect 34698 23468 34704 23520
rect 34756 23508 34762 23520
rect 35084 23508 35112 23539
rect 35897 23511 35955 23517
rect 35897 23508 35909 23511
rect 34756 23480 35909 23508
rect 34756 23468 34762 23480
rect 35897 23477 35909 23480
rect 35943 23508 35955 23511
rect 36262 23508 36268 23520
rect 35943 23480 36268 23508
rect 35943 23477 35955 23480
rect 35897 23471 35955 23477
rect 36262 23468 36268 23480
rect 36320 23508 36326 23520
rect 36648 23508 36676 23539
rect 37458 23536 37464 23548
rect 37516 23536 37522 23588
rect 38194 23576 38200 23588
rect 38155 23548 38200 23576
rect 38194 23536 38200 23548
rect 38252 23536 38258 23588
rect 39666 23576 39672 23588
rect 39579 23548 39672 23576
rect 39666 23536 39672 23548
rect 39724 23576 39730 23588
rect 40402 23576 40408 23588
rect 39724 23548 40408 23576
rect 39724 23536 39730 23548
rect 40402 23536 40408 23548
rect 40460 23536 40466 23588
rect 40865 23579 40923 23585
rect 40865 23545 40877 23579
rect 40911 23576 40923 23579
rect 41141 23579 41199 23585
rect 41141 23576 41153 23579
rect 40911 23548 41153 23576
rect 40911 23545 40923 23548
rect 40865 23539 40923 23545
rect 41141 23545 41153 23548
rect 41187 23576 41199 23579
rect 41322 23576 41328 23588
rect 41187 23548 41328 23576
rect 41187 23545 41199 23548
rect 41141 23539 41199 23545
rect 41322 23536 41328 23548
rect 41380 23536 41386 23588
rect 41690 23576 41696 23588
rect 41651 23548 41696 23576
rect 41690 23536 41696 23548
rect 41748 23536 41754 23588
rect 43257 23579 43315 23585
rect 43257 23545 43269 23579
rect 43303 23576 43315 23579
rect 43622 23576 43628 23588
rect 43303 23548 43628 23576
rect 43303 23545 43315 23548
rect 43257 23539 43315 23545
rect 39298 23508 39304 23520
rect 36320 23480 36676 23508
rect 39259 23480 39304 23508
rect 36320 23468 36326 23480
rect 39298 23468 39304 23480
rect 39356 23468 39362 23520
rect 42886 23508 42892 23520
rect 42847 23480 42892 23508
rect 42886 23468 42892 23480
rect 42944 23508 42950 23520
rect 43272 23508 43300 23539
rect 43622 23536 43628 23548
rect 43680 23576 43686 23588
rect 44085 23579 44143 23585
rect 44085 23576 44097 23579
rect 43680 23548 44097 23576
rect 43680 23536 43686 23548
rect 44085 23545 44097 23548
rect 44131 23545 44143 23579
rect 44085 23539 44143 23545
rect 42944 23480 43300 23508
rect 42944 23468 42950 23480
rect 44174 23468 44180 23520
rect 44232 23508 44238 23520
rect 44775 23511 44833 23517
rect 44775 23508 44787 23511
rect 44232 23480 44787 23508
rect 44232 23468 44238 23480
rect 44775 23477 44787 23480
rect 44821 23477 44833 23511
rect 44775 23471 44833 23477
rect 1104 23418 48852 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 48852 23418
rect 1104 23344 48852 23366
rect 2498 23304 2504 23316
rect 2459 23276 2504 23304
rect 2498 23264 2504 23276
rect 2556 23264 2562 23316
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 5166 23304 5172 23316
rect 2924 23276 5172 23304
rect 2924 23264 2930 23276
rect 5166 23264 5172 23276
rect 5224 23264 5230 23316
rect 5810 23264 5816 23316
rect 5868 23304 5874 23316
rect 7653 23307 7711 23313
rect 7653 23304 7665 23307
rect 5868 23276 7665 23304
rect 5868 23264 5874 23276
rect 7653 23273 7665 23276
rect 7699 23304 7711 23307
rect 7834 23304 7840 23316
rect 7699 23276 7840 23304
rect 7699 23273 7711 23276
rect 7653 23267 7711 23273
rect 7834 23264 7840 23276
rect 7892 23264 7898 23316
rect 8202 23264 8208 23316
rect 8260 23304 8266 23316
rect 9214 23304 9220 23316
rect 8260 23276 9220 23304
rect 8260 23264 8266 23276
rect 9214 23264 9220 23276
rect 9272 23264 9278 23316
rect 10686 23304 10692 23316
rect 9416 23276 10548 23304
rect 10647 23276 10692 23304
rect 3970 23196 3976 23248
rect 4028 23236 4034 23248
rect 4246 23236 4252 23248
rect 4028 23208 4252 23236
rect 4028 23196 4034 23208
rect 4246 23196 4252 23208
rect 4304 23196 4310 23248
rect 5258 23196 5264 23248
rect 5316 23236 5322 23248
rect 5316 23208 5672 23236
rect 5316 23196 5322 23208
rect 2314 23168 2320 23180
rect 2275 23140 2320 23168
rect 2314 23128 2320 23140
rect 2372 23128 2378 23180
rect 2406 23128 2412 23180
rect 2464 23168 2470 23180
rect 4433 23171 4491 23177
rect 4433 23168 4445 23171
rect 2464 23140 4445 23168
rect 2464 23128 2470 23140
rect 4433 23137 4445 23140
rect 4479 23168 4491 23171
rect 4706 23168 4712 23180
rect 4479 23140 4712 23168
rect 4479 23137 4491 23140
rect 4433 23131 4491 23137
rect 4706 23128 4712 23140
rect 4764 23168 4770 23180
rect 5534 23168 5540 23180
rect 4764 23140 5540 23168
rect 4764 23128 4770 23140
rect 5534 23128 5540 23140
rect 5592 23128 5598 23180
rect 5644 23177 5672 23208
rect 6638 23196 6644 23248
rect 6696 23236 6702 23248
rect 7374 23236 7380 23248
rect 6696 23208 7380 23236
rect 6696 23196 6702 23208
rect 7374 23196 7380 23208
rect 7432 23236 7438 23248
rect 9416 23236 9444 23276
rect 7432 23208 9444 23236
rect 7432 23196 7438 23208
rect 9490 23196 9496 23248
rect 9548 23236 9554 23248
rect 10520 23236 10548 23276
rect 10686 23264 10692 23276
rect 10744 23264 10750 23316
rect 12342 23304 12348 23316
rect 12303 23276 12348 23304
rect 12342 23264 12348 23276
rect 12400 23264 12406 23316
rect 13630 23264 13636 23316
rect 13688 23304 13694 23316
rect 14185 23307 14243 23313
rect 14185 23304 14197 23307
rect 13688 23276 14197 23304
rect 13688 23264 13694 23276
rect 14185 23273 14197 23276
rect 14231 23273 14243 23307
rect 14185 23267 14243 23273
rect 14918 23264 14924 23316
rect 14976 23304 14982 23316
rect 15473 23307 15531 23313
rect 15473 23304 15485 23307
rect 14976 23276 15485 23304
rect 14976 23264 14982 23276
rect 15473 23273 15485 23276
rect 15519 23273 15531 23307
rect 20714 23304 20720 23316
rect 20675 23276 20720 23304
rect 15473 23267 15531 23273
rect 20714 23264 20720 23276
rect 20772 23304 20778 23316
rect 21039 23307 21097 23313
rect 21039 23304 21051 23307
rect 20772 23276 21051 23304
rect 20772 23264 20778 23276
rect 21039 23273 21051 23276
rect 21085 23273 21097 23307
rect 21039 23267 21097 23273
rect 27982 23264 27988 23316
rect 28040 23264 28046 23316
rect 28905 23307 28963 23313
rect 28905 23273 28917 23307
rect 28951 23304 28963 23307
rect 29086 23304 29092 23316
rect 28951 23276 29092 23304
rect 28951 23273 28963 23276
rect 28905 23267 28963 23273
rect 29086 23264 29092 23276
rect 29144 23264 29150 23316
rect 31294 23304 31300 23316
rect 31255 23276 31300 23304
rect 31294 23264 31300 23276
rect 31352 23264 31358 23316
rect 32490 23304 32496 23316
rect 32451 23276 32496 23304
rect 32490 23264 32496 23276
rect 32548 23264 32554 23316
rect 33045 23307 33103 23313
rect 33045 23273 33057 23307
rect 33091 23304 33103 23307
rect 33410 23304 33416 23316
rect 33091 23276 33416 23304
rect 33091 23273 33103 23276
rect 33045 23267 33103 23273
rect 33410 23264 33416 23276
rect 33468 23264 33474 23316
rect 35250 23304 35256 23316
rect 35211 23276 35256 23304
rect 35250 23264 35256 23276
rect 35308 23264 35314 23316
rect 36630 23264 36636 23316
rect 36688 23304 36694 23316
rect 37093 23307 37151 23313
rect 37093 23304 37105 23307
rect 36688 23276 37105 23304
rect 36688 23264 36694 23276
rect 37093 23273 37105 23276
rect 37139 23273 37151 23307
rect 43162 23304 43168 23316
rect 43123 23276 43168 23304
rect 37093 23267 37151 23273
rect 43162 23264 43168 23276
rect 43220 23264 43226 23316
rect 43346 23264 43352 23316
rect 43404 23304 43410 23316
rect 45051 23307 45109 23313
rect 45051 23304 45063 23307
rect 43404 23276 45063 23304
rect 43404 23264 43410 23276
rect 45051 23273 45063 23276
rect 45097 23273 45109 23307
rect 45051 23267 45109 23273
rect 11146 23236 11152 23248
rect 9548 23208 9904 23236
rect 10520 23208 11152 23236
rect 9548 23196 9554 23208
rect 5629 23171 5687 23177
rect 5629 23137 5641 23171
rect 5675 23168 5687 23171
rect 6730 23168 6736 23180
rect 5675 23140 6736 23168
rect 5675 23137 5687 23140
rect 5629 23131 5687 23137
rect 6730 23128 6736 23140
rect 6788 23128 6794 23180
rect 7098 23128 7104 23180
rect 7156 23168 7162 23180
rect 7193 23171 7251 23177
rect 7193 23168 7205 23171
rect 7156 23140 7205 23168
rect 7156 23128 7162 23140
rect 7193 23137 7205 23140
rect 7239 23168 7251 23171
rect 7282 23168 7288 23180
rect 7239 23140 7288 23168
rect 7239 23137 7251 23140
rect 7193 23131 7251 23137
rect 7282 23128 7288 23140
rect 7340 23128 7346 23180
rect 8202 23168 8208 23180
rect 8163 23140 8208 23168
rect 8202 23128 8208 23140
rect 8260 23128 8266 23180
rect 8386 23168 8392 23180
rect 8347 23140 8392 23168
rect 8386 23128 8392 23140
rect 8444 23128 8450 23180
rect 8757 23171 8815 23177
rect 8757 23137 8769 23171
rect 8803 23168 8815 23171
rect 9214 23168 9220 23180
rect 8803 23140 9220 23168
rect 8803 23137 8815 23140
rect 8757 23131 8815 23137
rect 9214 23128 9220 23140
rect 9272 23128 9278 23180
rect 9674 23168 9680 23180
rect 9635 23140 9680 23168
rect 9674 23128 9680 23140
rect 9732 23128 9738 23180
rect 9876 23177 9904 23208
rect 11146 23196 11152 23208
rect 11204 23236 11210 23248
rect 11609 23239 11667 23245
rect 11204 23208 11284 23236
rect 11204 23196 11210 23208
rect 9861 23171 9919 23177
rect 9861 23137 9873 23171
rect 9907 23137 9919 23171
rect 11054 23168 11060 23180
rect 11015 23140 11060 23168
rect 9861 23131 9919 23137
rect 11054 23128 11060 23140
rect 11112 23128 11118 23180
rect 11256 23177 11284 23208
rect 11609 23205 11621 23239
rect 11655 23236 11667 23239
rect 15102 23236 15108 23248
rect 11655 23208 15108 23236
rect 11655 23205 11667 23208
rect 11609 23199 11667 23205
rect 15102 23196 15108 23208
rect 15160 23196 15166 23248
rect 17037 23239 17095 23245
rect 17037 23205 17049 23239
rect 17083 23236 17095 23239
rect 17310 23236 17316 23248
rect 17083 23208 17316 23236
rect 17083 23205 17095 23208
rect 17037 23199 17095 23205
rect 17310 23196 17316 23208
rect 17368 23196 17374 23248
rect 18598 23236 18604 23248
rect 18559 23208 18604 23236
rect 18598 23196 18604 23208
rect 18656 23196 18662 23248
rect 20806 23196 20812 23248
rect 20864 23236 20870 23248
rect 21361 23239 21419 23245
rect 21361 23236 21373 23239
rect 20864 23208 21373 23236
rect 20864 23196 20870 23208
rect 21361 23205 21373 23208
rect 21407 23205 21419 23239
rect 21361 23199 21419 23205
rect 23109 23239 23167 23245
rect 23109 23205 23121 23239
rect 23155 23236 23167 23239
rect 23290 23236 23296 23248
rect 23155 23208 23296 23236
rect 23155 23205 23167 23208
rect 23109 23199 23167 23205
rect 23290 23196 23296 23208
rect 23348 23236 23354 23248
rect 23842 23236 23848 23248
rect 23348 23208 23848 23236
rect 23348 23196 23354 23208
rect 23842 23196 23848 23208
rect 23900 23196 23906 23248
rect 24673 23239 24731 23245
rect 24673 23205 24685 23239
rect 24719 23236 24731 23239
rect 24762 23236 24768 23248
rect 24719 23208 24768 23236
rect 24719 23205 24731 23208
rect 24673 23199 24731 23205
rect 24762 23196 24768 23208
rect 24820 23196 24826 23248
rect 28000 23236 28028 23264
rect 28347 23239 28405 23245
rect 28347 23236 28359 23239
rect 28000 23208 28359 23236
rect 28347 23205 28359 23208
rect 28393 23236 28405 23239
rect 28442 23236 28448 23248
rect 28393 23208 28448 23236
rect 28393 23205 28405 23208
rect 28347 23199 28405 23205
rect 28442 23196 28448 23208
rect 28500 23196 28506 23248
rect 30975 23239 31033 23245
rect 30975 23205 30987 23239
rect 31021 23236 31033 23239
rect 31478 23236 31484 23248
rect 31021 23208 31484 23236
rect 31021 23205 31033 23208
rect 30975 23199 31033 23205
rect 31478 23196 31484 23208
rect 31536 23196 31542 23248
rect 33502 23196 33508 23248
rect 33560 23236 33566 23248
rect 34057 23239 34115 23245
rect 34057 23236 34069 23239
rect 33560 23208 34069 23236
rect 33560 23196 33566 23208
rect 34057 23205 34069 23208
rect 34103 23236 34115 23239
rect 34698 23236 34704 23248
rect 34103 23208 34704 23236
rect 34103 23205 34115 23208
rect 34057 23199 34115 23205
rect 34698 23196 34704 23208
rect 34756 23236 34762 23248
rect 34885 23239 34943 23245
rect 34885 23236 34897 23239
rect 34756 23208 34897 23236
rect 34756 23196 34762 23208
rect 34885 23205 34897 23208
rect 34931 23205 34943 23239
rect 36262 23236 36268 23248
rect 36223 23208 36268 23236
rect 34885 23199 34943 23205
rect 36262 23196 36268 23208
rect 36320 23196 36326 23248
rect 38562 23236 38568 23248
rect 38523 23208 38568 23236
rect 38562 23196 38568 23208
rect 38620 23196 38626 23248
rect 39298 23196 39304 23248
rect 39356 23236 39362 23248
rect 39714 23239 39772 23245
rect 39714 23236 39726 23239
rect 39356 23208 39726 23236
rect 39356 23196 39362 23208
rect 39714 23205 39726 23208
rect 39760 23205 39772 23239
rect 39714 23199 39772 23205
rect 41049 23239 41107 23245
rect 41049 23205 41061 23239
rect 41095 23236 41107 23239
rect 41322 23236 41328 23248
rect 41095 23208 41328 23236
rect 41095 23205 41107 23208
rect 41049 23199 41107 23205
rect 41322 23196 41328 23208
rect 41380 23196 41386 23248
rect 41874 23236 41880 23248
rect 41835 23208 41880 23236
rect 41874 23196 41880 23208
rect 41932 23196 41938 23248
rect 43533 23239 43591 23245
rect 43533 23205 43545 23239
rect 43579 23236 43591 23239
rect 43622 23236 43628 23248
rect 43579 23208 43628 23236
rect 43579 23205 43591 23208
rect 43533 23199 43591 23205
rect 43622 23196 43628 23208
rect 43680 23196 43686 23248
rect 11241 23171 11299 23177
rect 11241 23137 11253 23171
rect 11287 23137 11299 23171
rect 11241 23131 11299 23137
rect 13170 23128 13176 23180
rect 13228 23168 13234 23180
rect 13446 23168 13452 23180
rect 13228 23140 13452 23168
rect 13228 23128 13234 23140
rect 13446 23128 13452 23140
rect 13504 23128 13510 23180
rect 13630 23168 13636 23180
rect 13591 23140 13636 23168
rect 13630 23128 13636 23140
rect 13688 23128 13694 23180
rect 15908 23171 15966 23177
rect 15908 23137 15920 23171
rect 15954 23168 15966 23171
rect 16206 23168 16212 23180
rect 15954 23140 16212 23168
rect 15954 23137 15966 23140
rect 15908 23131 15966 23137
rect 16206 23128 16212 23140
rect 16264 23128 16270 23180
rect 20968 23171 21026 23177
rect 20968 23137 20980 23171
rect 21014 23168 21026 23171
rect 21266 23168 21272 23180
rect 21014 23140 21272 23168
rect 21014 23137 21026 23140
rect 20968 23131 21026 23137
rect 21266 23128 21272 23140
rect 21324 23128 21330 23180
rect 21913 23171 21971 23177
rect 21913 23137 21925 23171
rect 21959 23168 21971 23171
rect 22094 23168 22100 23180
rect 21959 23140 22100 23168
rect 21959 23137 21971 23140
rect 21913 23131 21971 23137
rect 22094 23128 22100 23140
rect 22152 23128 22158 23180
rect 26602 23128 26608 23180
rect 26660 23168 26666 23180
rect 26697 23171 26755 23177
rect 26697 23168 26709 23171
rect 26660 23140 26709 23168
rect 26660 23128 26666 23140
rect 26697 23137 26709 23140
rect 26743 23168 26755 23171
rect 27062 23168 27068 23180
rect 26743 23140 27068 23168
rect 26743 23137 26755 23140
rect 26697 23131 26755 23137
rect 27062 23128 27068 23140
rect 27120 23128 27126 23180
rect 27430 23128 27436 23180
rect 27488 23168 27494 23180
rect 27985 23171 28043 23177
rect 27985 23168 27997 23171
rect 27488 23140 27997 23168
rect 27488 23128 27494 23140
rect 27985 23137 27997 23140
rect 28031 23168 28043 23171
rect 28166 23168 28172 23180
rect 28031 23140 28172 23168
rect 28031 23137 28043 23140
rect 27985 23131 28043 23137
rect 28166 23128 28172 23140
rect 28224 23128 28230 23180
rect 29730 23168 29736 23180
rect 29643 23140 29736 23168
rect 29730 23128 29736 23140
rect 29788 23128 29794 23180
rect 30282 23128 30288 23180
rect 30340 23168 30346 23180
rect 30872 23171 30930 23177
rect 30872 23168 30884 23171
rect 30340 23140 30884 23168
rect 30340 23128 30346 23140
rect 30872 23137 30884 23140
rect 30918 23168 30930 23171
rect 33137 23171 33195 23177
rect 33137 23168 33149 23171
rect 30918 23140 33149 23168
rect 30918 23137 30930 23140
rect 30872 23131 30930 23137
rect 33137 23137 33149 23140
rect 33183 23137 33195 23171
rect 33137 23131 33195 23137
rect 37829 23171 37887 23177
rect 37829 23137 37841 23171
rect 37875 23137 37887 23171
rect 38286 23168 38292 23180
rect 38247 23140 38292 23168
rect 37829 23131 37887 23137
rect 4982 23060 4988 23112
rect 5040 23100 5046 23112
rect 5994 23100 6000 23112
rect 5040 23072 6000 23100
rect 5040 23060 5046 23072
rect 5994 23060 6000 23072
rect 6052 23100 6058 23112
rect 8113 23103 8171 23109
rect 8113 23100 8125 23103
rect 6052 23072 7144 23100
rect 6052 23060 6058 23072
rect 5166 23032 5172 23044
rect 5079 23004 5172 23032
rect 5166 22992 5172 23004
rect 5224 23032 5230 23044
rect 5537 23035 5595 23041
rect 5537 23032 5549 23035
rect 5224 23004 5549 23032
rect 5224 22992 5230 23004
rect 5537 23001 5549 23004
rect 5583 23032 5595 23035
rect 6273 23035 6331 23041
rect 5583 23004 5948 23032
rect 5583 23001 5595 23004
rect 5537 22995 5595 23001
rect 5920 22976 5948 23004
rect 6273 23001 6285 23035
rect 6319 23032 6331 23035
rect 6319 23004 6868 23032
rect 6319 23001 6331 23004
rect 6273 22995 6331 23001
rect 6840 22976 6868 23004
rect 2866 22924 2872 22976
rect 2924 22964 2930 22976
rect 2961 22967 3019 22973
rect 2961 22964 2973 22967
rect 2924 22936 2973 22964
rect 2924 22924 2930 22936
rect 2961 22933 2973 22936
rect 3007 22964 3019 22967
rect 3142 22964 3148 22976
rect 3007 22936 3148 22964
rect 3007 22933 3019 22936
rect 2961 22927 3019 22933
rect 3142 22924 3148 22936
rect 3200 22924 3206 22976
rect 3326 22964 3332 22976
rect 3287 22936 3332 22964
rect 3326 22924 3332 22936
rect 3384 22924 3390 22976
rect 3786 22964 3792 22976
rect 3747 22936 3792 22964
rect 3786 22924 3792 22936
rect 3844 22924 3850 22976
rect 4062 22924 4068 22976
rect 4120 22964 4126 22976
rect 4525 22967 4583 22973
rect 4525 22964 4537 22967
rect 4120 22936 4537 22964
rect 4120 22924 4126 22936
rect 4525 22933 4537 22936
rect 4571 22933 4583 22967
rect 4525 22927 4583 22933
rect 5626 22924 5632 22976
rect 5684 22964 5690 22976
rect 5767 22967 5825 22973
rect 5767 22964 5779 22967
rect 5684 22936 5779 22964
rect 5684 22924 5690 22936
rect 5767 22933 5779 22936
rect 5813 22933 5825 22967
rect 5902 22964 5908 22976
rect 5863 22936 5908 22964
rect 5767 22927 5825 22933
rect 5902 22924 5908 22936
rect 5960 22924 5966 22976
rect 6822 22924 6828 22976
rect 6880 22964 6886 22976
rect 7009 22967 7067 22973
rect 7009 22964 7021 22967
rect 6880 22936 7021 22964
rect 6880 22924 6886 22936
rect 7009 22933 7021 22936
rect 7055 22933 7067 22967
rect 7116 22964 7144 23072
rect 7208 23072 8125 23100
rect 7208 23044 7236 23072
rect 8113 23069 8125 23072
rect 8159 23100 8171 23103
rect 10229 23103 10287 23109
rect 10229 23100 10241 23103
rect 8159 23072 10241 23100
rect 8159 23069 8171 23072
rect 8113 23063 8171 23069
rect 10229 23069 10241 23072
rect 10275 23100 10287 23103
rect 12066 23100 12072 23112
rect 10275 23072 12072 23100
rect 10275 23069 10287 23072
rect 10229 23063 10287 23069
rect 12066 23060 12072 23072
rect 12124 23060 12130 23112
rect 13906 23100 13912 23112
rect 13867 23072 13912 23100
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 16945 23103 17003 23109
rect 16945 23069 16957 23103
rect 16991 23069 17003 23103
rect 16945 23063 17003 23069
rect 7190 22992 7196 23044
rect 7248 22992 7254 23044
rect 7377 23035 7435 23041
rect 7377 23001 7389 23035
rect 7423 23032 7435 23035
rect 9858 23032 9864 23044
rect 7423 23004 9864 23032
rect 7423 23001 7435 23004
rect 7377 22995 7435 23001
rect 9858 22992 9864 23004
rect 9916 22992 9922 23044
rect 15979 23035 16037 23041
rect 15979 23001 15991 23035
rect 16025 23032 16037 23035
rect 16758 23032 16764 23044
rect 16025 23004 16764 23032
rect 16025 23001 16037 23004
rect 15979 22995 16037 23001
rect 16758 22992 16764 23004
rect 16816 23032 16822 23044
rect 16960 23032 16988 23063
rect 18230 23060 18236 23112
rect 18288 23100 18294 23112
rect 18509 23103 18567 23109
rect 18509 23100 18521 23103
rect 18288 23072 18521 23100
rect 18288 23060 18294 23072
rect 18509 23069 18521 23072
rect 18555 23100 18567 23103
rect 18782 23100 18788 23112
rect 18555 23072 18788 23100
rect 18555 23069 18567 23072
rect 18509 23063 18567 23069
rect 18782 23060 18788 23072
rect 18840 23060 18846 23112
rect 23014 23100 23020 23112
rect 22975 23072 23020 23100
rect 23014 23060 23020 23072
rect 23072 23060 23078 23112
rect 23293 23103 23351 23109
rect 23293 23069 23305 23103
rect 23339 23069 23351 23103
rect 24578 23100 24584 23112
rect 24539 23072 24584 23100
rect 23293 23063 23351 23069
rect 16816 23004 16988 23032
rect 17497 23035 17555 23041
rect 16816 22992 16822 23004
rect 17497 23001 17509 23035
rect 17543 23032 17555 23035
rect 17862 23032 17868 23044
rect 17543 23004 17868 23032
rect 17543 23001 17555 23004
rect 17497 22995 17555 23001
rect 17862 22992 17868 23004
rect 17920 23032 17926 23044
rect 19061 23035 19119 23041
rect 19061 23032 19073 23035
rect 17920 23004 19073 23032
rect 17920 22992 17926 23004
rect 19061 23001 19073 23004
rect 19107 23001 19119 23035
rect 19061 22995 19119 23001
rect 21910 22992 21916 23044
rect 21968 23032 21974 23044
rect 23308 23032 23336 23063
rect 24578 23060 24584 23072
rect 24636 23060 24642 23112
rect 24854 23100 24860 23112
rect 24815 23072 24860 23100
rect 24854 23060 24860 23072
rect 24912 23060 24918 23112
rect 27338 23060 27344 23112
rect 27396 23100 27402 23112
rect 29748 23100 29776 23128
rect 32122 23100 32128 23112
rect 27396 23072 29776 23100
rect 32083 23072 32128 23100
rect 27396 23060 27402 23072
rect 32122 23060 32128 23072
rect 32180 23060 32186 23112
rect 33318 23100 33324 23112
rect 33279 23072 33324 23100
rect 33318 23060 33324 23072
rect 33376 23060 33382 23112
rect 33962 23100 33968 23112
rect 33923 23072 33968 23100
rect 33962 23060 33968 23072
rect 34020 23060 34026 23112
rect 34146 23060 34152 23112
rect 34204 23100 34210 23112
rect 34241 23103 34299 23109
rect 34241 23100 34253 23103
rect 34204 23072 34253 23100
rect 34204 23060 34210 23072
rect 34241 23069 34253 23072
rect 34287 23069 34299 23103
rect 34241 23063 34299 23069
rect 34716 23072 35756 23100
rect 25222 23032 25228 23044
rect 21968 23004 25228 23032
rect 21968 22992 21974 23004
rect 25222 22992 25228 23004
rect 25280 22992 25286 23044
rect 26881 23035 26939 23041
rect 26881 23001 26893 23035
rect 26927 23032 26939 23035
rect 26927 23004 28212 23032
rect 26927 23001 26939 23004
rect 26881 22995 26939 23001
rect 8386 22964 8392 22976
rect 7116 22936 8392 22964
rect 7009 22927 7067 22933
rect 8386 22924 8392 22936
rect 8444 22924 8450 22976
rect 18141 22967 18199 22973
rect 18141 22933 18153 22967
rect 18187 22964 18199 22967
rect 18690 22964 18696 22976
rect 18187 22936 18696 22964
rect 18187 22933 18199 22936
rect 18141 22927 18199 22933
rect 18690 22924 18696 22936
rect 18748 22924 18754 22976
rect 20070 22924 20076 22976
rect 20128 22964 20134 22976
rect 22097 22967 22155 22973
rect 22097 22964 22109 22967
rect 20128 22936 22109 22964
rect 20128 22924 20134 22936
rect 22097 22933 22109 22936
rect 22143 22933 22155 22967
rect 27154 22964 27160 22976
rect 27115 22936 27160 22964
rect 22097 22927 22155 22933
rect 27154 22924 27160 22936
rect 27212 22964 27218 22976
rect 27338 22964 27344 22976
rect 27212 22936 27344 22964
rect 27212 22924 27218 22936
rect 27338 22924 27344 22936
rect 27396 22924 27402 22976
rect 28184 22964 28212 23004
rect 28258 22992 28264 23044
rect 28316 23032 28322 23044
rect 29917 23035 29975 23041
rect 29917 23032 29929 23035
rect 28316 23004 29929 23032
rect 28316 22992 28322 23004
rect 29917 23001 29929 23004
rect 29963 23001 29975 23035
rect 34716 23032 34744 23072
rect 29917 22995 29975 23001
rect 30484 23004 34744 23032
rect 30484 22976 30512 23004
rect 34790 22992 34796 23044
rect 34848 23032 34854 23044
rect 35621 23035 35679 23041
rect 35621 23032 35633 23035
rect 34848 23004 35633 23032
rect 34848 22992 34854 23004
rect 35621 23001 35633 23004
rect 35667 23001 35679 23035
rect 35728 23032 35756 23072
rect 35802 23060 35808 23112
rect 35860 23100 35866 23112
rect 36170 23100 36176 23112
rect 35860 23072 36176 23100
rect 35860 23060 35866 23072
rect 36170 23060 36176 23072
rect 36228 23060 36234 23112
rect 37844 23100 37872 23131
rect 38286 23128 38292 23140
rect 38344 23168 38350 23180
rect 38838 23168 38844 23180
rect 38344 23140 38844 23168
rect 38344 23128 38350 23140
rect 38838 23128 38844 23140
rect 38896 23128 38902 23180
rect 44910 23168 44916 23180
rect 44871 23140 44916 23168
rect 44910 23128 44916 23140
rect 44968 23128 44974 23180
rect 38102 23100 38108 23112
rect 36648 23072 38108 23100
rect 36648 23032 36676 23072
rect 38102 23060 38108 23072
rect 38160 23060 38166 23112
rect 39390 23100 39396 23112
rect 39351 23072 39396 23100
rect 39390 23060 39396 23072
rect 39448 23060 39454 23112
rect 40494 23060 40500 23112
rect 40552 23100 40558 23112
rect 40770 23100 40776 23112
rect 40552 23072 40776 23100
rect 40552 23060 40558 23072
rect 40770 23060 40776 23072
rect 40828 23100 40834 23112
rect 41233 23103 41291 23109
rect 41233 23100 41245 23103
rect 40828 23072 41245 23100
rect 40828 23060 40834 23072
rect 41233 23069 41245 23072
rect 41279 23069 41291 23103
rect 41233 23063 41291 23069
rect 41690 23060 41696 23112
rect 41748 23100 41754 23112
rect 42058 23100 42064 23112
rect 41748 23072 42064 23100
rect 41748 23060 41754 23072
rect 42058 23060 42064 23072
rect 42116 23100 42122 23112
rect 43438 23100 43444 23112
rect 42116 23072 42794 23100
rect 43399 23072 43444 23100
rect 42116 23060 42122 23072
rect 35728 23004 36676 23032
rect 36725 23035 36783 23041
rect 35621 22995 35679 23001
rect 36725 23001 36737 23035
rect 36771 23032 36783 23035
rect 36814 23032 36820 23044
rect 36771 23004 36820 23032
rect 36771 23001 36783 23004
rect 36725 22995 36783 23001
rect 36814 22992 36820 23004
rect 36872 22992 36878 23044
rect 40313 23035 40371 23041
rect 40313 23001 40325 23035
rect 40359 23032 40371 23035
rect 42766 23032 42794 23072
rect 43438 23060 43444 23072
rect 43496 23060 43502 23112
rect 43717 23103 43775 23109
rect 43717 23100 43729 23103
rect 43548 23072 43729 23100
rect 43548 23032 43576 23072
rect 43717 23069 43729 23072
rect 43763 23069 43775 23103
rect 43717 23063 43775 23069
rect 40359 23004 41736 23032
rect 42766 23004 43576 23032
rect 40359 23001 40371 23004
rect 40313 22995 40371 23001
rect 28902 22964 28908 22976
rect 28184 22936 28908 22964
rect 28902 22924 28908 22936
rect 28960 22924 28966 22976
rect 29270 22964 29276 22976
rect 29231 22936 29276 22964
rect 29270 22924 29276 22936
rect 29328 22924 29334 22976
rect 30466 22964 30472 22976
rect 30427 22936 30472 22964
rect 30466 22924 30472 22936
rect 30524 22924 30530 22976
rect 33137 22967 33195 22973
rect 33137 22933 33149 22967
rect 33183 22964 33195 22967
rect 37182 22964 37188 22976
rect 33183 22936 37188 22964
rect 33183 22933 33195 22936
rect 33137 22927 33195 22933
rect 37182 22924 37188 22936
rect 37240 22924 37246 22976
rect 41708 22964 41736 23004
rect 42886 22964 42892 22976
rect 41708 22936 42892 22964
rect 42886 22924 42892 22936
rect 42944 22924 42950 22976
rect 1104 22874 48852 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 48852 22874
rect 1104 22800 48852 22822
rect 3970 22760 3976 22772
rect 3931 22732 3976 22760
rect 3970 22720 3976 22732
rect 4028 22720 4034 22772
rect 4341 22763 4399 22769
rect 4341 22729 4353 22763
rect 4387 22760 4399 22763
rect 4706 22760 4712 22772
rect 4387 22732 4712 22760
rect 4387 22729 4399 22732
rect 4341 22723 4399 22729
rect 4706 22720 4712 22732
rect 4764 22720 4770 22772
rect 5994 22720 6000 22772
rect 6052 22760 6058 22772
rect 6365 22763 6423 22769
rect 6365 22760 6377 22763
rect 6052 22732 6377 22760
rect 6052 22720 6058 22732
rect 6365 22729 6377 22732
rect 6411 22729 6423 22763
rect 7006 22760 7012 22772
rect 6967 22732 7012 22760
rect 6365 22723 6423 22729
rect 7006 22720 7012 22732
rect 7064 22720 7070 22772
rect 7282 22760 7288 22772
rect 7243 22732 7288 22760
rect 7282 22720 7288 22732
rect 7340 22720 7346 22772
rect 7834 22760 7840 22772
rect 7795 22732 7840 22760
rect 7834 22720 7840 22732
rect 7892 22720 7898 22772
rect 8202 22760 8208 22772
rect 8163 22732 8208 22760
rect 8202 22720 8208 22732
rect 8260 22720 8266 22772
rect 9490 22720 9496 22772
rect 9548 22760 9554 22772
rect 9769 22763 9827 22769
rect 9769 22760 9781 22763
rect 9548 22732 9781 22760
rect 9548 22720 9554 22732
rect 9769 22729 9781 22732
rect 9815 22729 9827 22763
rect 9769 22723 9827 22729
rect 11146 22720 11152 22772
rect 11204 22760 11210 22772
rect 11425 22763 11483 22769
rect 11425 22760 11437 22763
rect 11204 22732 11437 22760
rect 11204 22720 11210 22732
rect 11425 22729 11437 22732
rect 11471 22729 11483 22763
rect 11425 22723 11483 22729
rect 16025 22763 16083 22769
rect 16025 22729 16037 22763
rect 16071 22760 16083 22763
rect 16206 22760 16212 22772
rect 16071 22732 16212 22760
rect 16071 22729 16083 22732
rect 16025 22723 16083 22729
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 16758 22760 16764 22772
rect 16719 22732 16764 22760
rect 16758 22720 16764 22732
rect 16816 22720 16822 22772
rect 17310 22720 17316 22772
rect 17368 22760 17374 22772
rect 17405 22763 17463 22769
rect 17405 22760 17417 22763
rect 17368 22732 17417 22760
rect 17368 22720 17374 22732
rect 17405 22729 17417 22732
rect 17451 22729 17463 22763
rect 17405 22723 17463 22729
rect 20993 22763 21051 22769
rect 20993 22729 21005 22763
rect 21039 22760 21051 22763
rect 21082 22760 21088 22772
rect 21039 22732 21088 22760
rect 21039 22729 21051 22732
rect 20993 22723 21051 22729
rect 21082 22720 21088 22732
rect 21140 22720 21146 22772
rect 21266 22760 21272 22772
rect 21227 22732 21272 22760
rect 21266 22720 21272 22732
rect 21324 22720 21330 22772
rect 23014 22720 23020 22772
rect 23072 22760 23078 22772
rect 23385 22763 23443 22769
rect 23385 22760 23397 22763
rect 23072 22732 23397 22760
rect 23072 22720 23078 22732
rect 23385 22729 23397 22732
rect 23431 22729 23443 22763
rect 23385 22723 23443 22729
rect 24578 22720 24584 22772
rect 24636 22760 24642 22772
rect 25501 22763 25559 22769
rect 25501 22760 25513 22763
rect 24636 22732 25513 22760
rect 24636 22720 24642 22732
rect 25501 22729 25513 22732
rect 25547 22729 25559 22763
rect 26234 22760 26240 22772
rect 26195 22732 26240 22760
rect 25501 22723 25559 22729
rect 26234 22720 26240 22732
rect 26292 22720 26298 22772
rect 26602 22760 26608 22772
rect 26563 22732 26608 22760
rect 26602 22720 26608 22732
rect 26660 22720 26666 22772
rect 28166 22720 28172 22772
rect 28224 22760 28230 22772
rect 28353 22763 28411 22769
rect 28353 22760 28365 22763
rect 28224 22732 28365 22760
rect 28224 22720 28230 22732
rect 28353 22729 28365 22732
rect 28399 22729 28411 22763
rect 28353 22723 28411 22729
rect 28994 22720 29000 22772
rect 29052 22760 29058 22772
rect 29457 22763 29515 22769
rect 29457 22760 29469 22763
rect 29052 22732 29469 22760
rect 29052 22720 29058 22732
rect 29457 22729 29469 22732
rect 29503 22729 29515 22763
rect 29457 22723 29515 22729
rect 32953 22763 33011 22769
rect 32953 22729 32965 22763
rect 32999 22760 33011 22763
rect 33502 22760 33508 22772
rect 32999 22732 33508 22760
rect 32999 22729 33011 22732
rect 32953 22723 33011 22729
rect 33502 22720 33508 22732
rect 33560 22720 33566 22772
rect 33962 22769 33968 22772
rect 33689 22763 33747 22769
rect 33689 22729 33701 22763
rect 33735 22760 33747 22763
rect 33919 22763 33968 22769
rect 33919 22760 33931 22763
rect 33735 22732 33931 22760
rect 33735 22729 33747 22732
rect 33689 22723 33747 22729
rect 33919 22729 33931 22732
rect 33965 22729 33968 22763
rect 33919 22723 33968 22729
rect 33962 22720 33968 22723
rect 34020 22720 34026 22772
rect 34698 22760 34704 22772
rect 34659 22732 34704 22760
rect 34698 22720 34704 22732
rect 34756 22720 34762 22772
rect 34790 22720 34796 22772
rect 34848 22760 34854 22772
rect 35023 22763 35081 22769
rect 35023 22760 35035 22763
rect 34848 22732 35035 22760
rect 34848 22720 34854 22732
rect 35023 22729 35035 22732
rect 35069 22729 35081 22763
rect 35802 22760 35808 22772
rect 35763 22732 35808 22760
rect 35023 22723 35081 22729
rect 35802 22720 35808 22732
rect 35860 22720 35866 22772
rect 37415 22763 37473 22769
rect 37415 22729 37427 22763
rect 37461 22760 37473 22763
rect 37550 22760 37556 22772
rect 37461 22732 37556 22760
rect 37461 22729 37473 22732
rect 37415 22723 37473 22729
rect 37550 22720 37556 22732
rect 37608 22720 37614 22772
rect 38102 22760 38108 22772
rect 38063 22732 38108 22760
rect 38102 22720 38108 22732
rect 38160 22720 38166 22772
rect 40313 22763 40371 22769
rect 40313 22729 40325 22763
rect 40359 22760 40371 22763
rect 40494 22760 40500 22772
rect 40359 22732 40500 22760
rect 40359 22729 40371 22732
rect 40313 22723 40371 22729
rect 40494 22720 40500 22732
rect 40552 22720 40558 22772
rect 40635 22763 40693 22769
rect 40635 22729 40647 22763
rect 40681 22760 40693 22763
rect 41046 22760 41052 22772
rect 40681 22732 41052 22760
rect 40681 22729 40693 22732
rect 40635 22723 40693 22729
rect 41046 22720 41052 22732
rect 41104 22720 41110 22772
rect 41322 22760 41328 22772
rect 41283 22732 41328 22760
rect 41322 22720 41328 22732
rect 41380 22720 41386 22772
rect 42613 22763 42671 22769
rect 42613 22729 42625 22763
rect 42659 22760 42671 22763
rect 43438 22760 43444 22772
rect 42659 22732 43444 22760
rect 42659 22729 42671 22732
rect 42613 22723 42671 22729
rect 43438 22720 43444 22732
rect 43496 22720 43502 22772
rect 3602 22652 3608 22704
rect 3660 22692 3666 22704
rect 5626 22692 5632 22704
rect 3660 22664 5632 22692
rect 3660 22652 3666 22664
rect 5626 22652 5632 22664
rect 5684 22652 5690 22704
rect 5902 22652 5908 22704
rect 5960 22692 5966 22704
rect 6089 22695 6147 22701
rect 6089 22692 6101 22695
rect 5960 22664 6101 22692
rect 5960 22652 5966 22664
rect 6089 22661 6101 22664
rect 6135 22692 6147 22695
rect 8220 22692 8248 22720
rect 6135 22664 8248 22692
rect 6135 22661 6147 22664
rect 6089 22655 6147 22661
rect 11514 22652 11520 22704
rect 11572 22692 11578 22704
rect 12894 22692 12900 22704
rect 11572 22664 12900 22692
rect 11572 22652 11578 22664
rect 12894 22652 12900 22664
rect 12952 22692 12958 22704
rect 15289 22695 15347 22701
rect 15289 22692 15301 22695
rect 12952 22664 15301 22692
rect 12952 22652 12958 22664
rect 15289 22661 15301 22664
rect 15335 22661 15347 22695
rect 15289 22655 15347 22661
rect 17129 22695 17187 22701
rect 17129 22661 17141 22695
rect 17175 22692 17187 22695
rect 18322 22692 18328 22704
rect 17175 22664 18328 22692
rect 17175 22661 17187 22664
rect 17129 22655 17187 22661
rect 18322 22652 18328 22664
rect 18380 22652 18386 22704
rect 18966 22652 18972 22704
rect 19024 22692 19030 22704
rect 21910 22692 21916 22704
rect 19024 22664 21916 22692
rect 19024 22652 19030 22664
rect 21910 22652 21916 22664
rect 21968 22692 21974 22704
rect 22833 22695 22891 22701
rect 22833 22692 22845 22695
rect 21968 22664 22845 22692
rect 21968 22652 21974 22664
rect 22833 22661 22845 22664
rect 22879 22661 22891 22695
rect 22833 22655 22891 22661
rect 23109 22695 23167 22701
rect 23109 22661 23121 22695
rect 23155 22692 23167 22695
rect 23290 22692 23296 22704
rect 23155 22664 23296 22692
rect 23155 22661 23167 22664
rect 23109 22655 23167 22661
rect 23290 22652 23296 22664
rect 23348 22652 23354 22704
rect 26418 22692 26424 22704
rect 23446 22664 26424 22692
rect 2866 22624 2872 22636
rect 2827 22596 2872 22624
rect 2866 22584 2872 22596
rect 2924 22584 2930 22636
rect 4614 22624 4620 22636
rect 4448 22596 4620 22624
rect 2225 22559 2283 22565
rect 2225 22556 2237 22559
rect 1964 22528 2237 22556
rect 1964 22432 1992 22528
rect 2225 22525 2237 22528
rect 2271 22556 2283 22559
rect 2314 22556 2320 22568
rect 2271 22528 2320 22556
rect 2271 22525 2283 22528
rect 2225 22519 2283 22525
rect 2314 22516 2320 22528
rect 2372 22556 2378 22568
rect 4448 22565 4476 22596
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 9401 22627 9459 22633
rect 9401 22624 9413 22627
rect 8588 22596 9413 22624
rect 3145 22559 3203 22565
rect 3145 22556 3157 22559
rect 2372 22528 3157 22556
rect 2372 22516 2378 22528
rect 3145 22525 3157 22528
rect 3191 22525 3203 22559
rect 3145 22519 3203 22525
rect 4433 22559 4491 22565
rect 4433 22525 4445 22559
rect 4479 22525 4491 22559
rect 4893 22559 4951 22565
rect 4893 22556 4905 22559
rect 4433 22519 4491 22525
rect 4540 22528 4905 22556
rect 3605 22491 3663 22497
rect 3605 22457 3617 22491
rect 3651 22488 3663 22491
rect 3970 22488 3976 22500
rect 3651 22460 3976 22488
rect 3651 22457 3663 22460
rect 3605 22451 3663 22457
rect 3970 22448 3976 22460
rect 4028 22488 4034 22500
rect 4540 22488 4568 22528
rect 4893 22525 4905 22528
rect 4939 22525 4951 22559
rect 6822 22556 6828 22568
rect 6783 22528 6828 22556
rect 4893 22519 4951 22525
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 8110 22516 8116 22568
rect 8168 22556 8174 22568
rect 8588 22565 8616 22596
rect 9401 22593 9413 22596
rect 9447 22593 9459 22627
rect 9401 22587 9459 22593
rect 13265 22627 13323 22633
rect 13265 22593 13277 22627
rect 13311 22624 13323 22627
rect 13722 22624 13728 22636
rect 13311 22596 13728 22624
rect 13311 22593 13323 22596
rect 13265 22587 13323 22593
rect 13722 22584 13728 22596
rect 13780 22624 13786 22636
rect 14734 22624 14740 22636
rect 13780 22596 14740 22624
rect 13780 22584 13786 22596
rect 14734 22584 14740 22596
rect 14792 22584 14798 22636
rect 17865 22627 17923 22633
rect 17865 22624 17877 22627
rect 16960 22596 17877 22624
rect 8573 22559 8631 22565
rect 8573 22556 8585 22559
rect 8168 22528 8585 22556
rect 8168 22516 8174 22528
rect 8573 22525 8585 22528
rect 8619 22525 8631 22559
rect 8573 22519 8631 22525
rect 8757 22559 8815 22565
rect 8757 22525 8769 22559
rect 8803 22525 8815 22559
rect 8757 22519 8815 22525
rect 5166 22488 5172 22500
rect 4028 22460 4568 22488
rect 5127 22460 5172 22488
rect 4028 22448 4034 22460
rect 5166 22448 5172 22460
rect 5224 22448 5230 22500
rect 7834 22448 7840 22500
rect 7892 22488 7898 22500
rect 8772 22488 8800 22519
rect 10686 22516 10692 22568
rect 10744 22556 10750 22568
rect 10781 22559 10839 22565
rect 10781 22556 10793 22559
rect 10744 22528 10793 22556
rect 10744 22516 10750 22528
rect 10781 22525 10793 22528
rect 10827 22525 10839 22559
rect 13354 22556 13360 22568
rect 13315 22528 13360 22556
rect 10781 22519 10839 22525
rect 13354 22516 13360 22528
rect 13412 22556 13418 22568
rect 14553 22559 14611 22565
rect 14553 22556 14565 22559
rect 13412 22528 14565 22556
rect 13412 22516 13418 22528
rect 14553 22525 14565 22528
rect 14599 22525 14611 22559
rect 15102 22556 15108 22568
rect 15063 22528 15108 22556
rect 14553 22519 14611 22525
rect 15102 22516 15108 22528
rect 15160 22556 15166 22568
rect 16960 22565 16988 22596
rect 17865 22593 17877 22596
rect 17911 22624 17923 22627
rect 19242 22624 19248 22636
rect 17911 22596 19248 22624
rect 17911 22593 17923 22596
rect 17865 22587 17923 22593
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 23446 22624 23474 22664
rect 26418 22652 26424 22664
rect 26476 22652 26482 22704
rect 26694 22652 26700 22704
rect 26752 22692 26758 22704
rect 34716 22692 34744 22720
rect 36081 22695 36139 22701
rect 36081 22692 36093 22695
rect 26752 22664 29868 22692
rect 34716 22664 36093 22692
rect 26752 22652 26758 22664
rect 22020 22596 23474 22624
rect 24581 22627 24639 22633
rect 15565 22559 15623 22565
rect 15565 22556 15577 22559
rect 15160 22528 15577 22556
rect 15160 22516 15166 22528
rect 15565 22525 15577 22528
rect 15611 22525 15623 22559
rect 15565 22519 15623 22525
rect 16945 22559 17003 22565
rect 16945 22525 16957 22559
rect 16991 22525 17003 22559
rect 18690 22556 18696 22568
rect 18651 22528 18696 22556
rect 16945 22519 17003 22525
rect 18690 22516 18696 22528
rect 18748 22516 18754 22568
rect 20073 22559 20131 22565
rect 20073 22525 20085 22559
rect 20119 22556 20131 22559
rect 20254 22556 20260 22568
rect 20119 22528 20260 22556
rect 20119 22525 20131 22528
rect 20073 22519 20131 22525
rect 20254 22516 20260 22528
rect 20312 22516 20318 22568
rect 22020 22565 22048 22596
rect 24581 22593 24593 22627
rect 24627 22624 24639 22627
rect 24762 22624 24768 22636
rect 24627 22596 24768 22624
rect 24627 22593 24639 22596
rect 24581 22587 24639 22593
rect 24762 22584 24768 22596
rect 24820 22584 24826 22636
rect 27433 22627 27491 22633
rect 27433 22593 27445 22627
rect 27479 22624 27491 22627
rect 28350 22624 28356 22636
rect 27479 22596 28356 22624
rect 27479 22593 27491 22596
rect 27433 22587 27491 22593
rect 28350 22584 28356 22596
rect 28408 22584 28414 22636
rect 29840 22568 29868 22664
rect 36081 22661 36093 22664
rect 36127 22661 36139 22695
rect 36081 22655 36139 22661
rect 37185 22695 37243 22701
rect 37185 22661 37197 22695
rect 37231 22692 37243 22695
rect 38286 22692 38292 22704
rect 37231 22664 38292 22692
rect 37231 22661 37243 22664
rect 37185 22655 37243 22661
rect 38286 22652 38292 22664
rect 38344 22652 38350 22704
rect 39022 22652 39028 22704
rect 39080 22692 39086 22704
rect 41969 22695 42027 22701
rect 41969 22692 41981 22695
rect 39080 22664 41981 22692
rect 39080 22652 39086 22664
rect 31478 22584 31484 22636
rect 31536 22624 31542 22636
rect 38010 22624 38016 22636
rect 31536 22596 38016 22624
rect 31536 22584 31542 22596
rect 38010 22584 38016 22596
rect 38068 22584 38074 22636
rect 38304 22624 38332 22652
rect 39117 22627 39175 22633
rect 38304 22596 38884 22624
rect 22005 22559 22063 22565
rect 22005 22556 22017 22559
rect 21836 22528 22017 22556
rect 9122 22488 9128 22500
rect 7892 22460 8800 22488
rect 9083 22460 9128 22488
rect 7892 22448 7898 22460
rect 9122 22448 9128 22460
rect 9180 22448 9186 22500
rect 10594 22488 10600 22500
rect 10555 22460 10600 22488
rect 10594 22448 10600 22460
rect 10652 22448 10658 22500
rect 11054 22448 11060 22500
rect 11112 22488 11118 22500
rect 11149 22491 11207 22497
rect 11149 22488 11161 22491
rect 11112 22460 11161 22488
rect 11112 22448 11118 22460
rect 11149 22457 11161 22460
rect 11195 22488 11207 22491
rect 12897 22491 12955 22497
rect 11195 22460 11836 22488
rect 11195 22457 11207 22460
rect 11149 22451 11207 22457
rect 11808 22432 11836 22460
rect 12897 22457 12909 22491
rect 12943 22488 12955 22491
rect 13446 22488 13452 22500
rect 12943 22460 13452 22488
rect 12943 22457 12955 22460
rect 12897 22451 12955 22457
rect 13446 22448 13452 22460
rect 13504 22448 13510 22500
rect 18046 22488 18052 22500
rect 18007 22460 18052 22488
rect 18046 22448 18052 22460
rect 18104 22448 18110 22500
rect 19981 22491 20039 22497
rect 19981 22457 19993 22491
rect 20027 22488 20039 22491
rect 20394 22491 20452 22497
rect 20394 22488 20406 22491
rect 20027 22460 20406 22488
rect 20027 22457 20039 22460
rect 19981 22451 20039 22457
rect 20394 22457 20406 22460
rect 20440 22488 20452 22491
rect 21634 22488 21640 22500
rect 20440 22460 21640 22488
rect 20440 22457 20452 22460
rect 20394 22451 20452 22457
rect 21634 22448 21640 22460
rect 21692 22448 21698 22500
rect 21836 22432 21864 22528
rect 22005 22525 22017 22528
rect 22051 22525 22063 22559
rect 22005 22519 22063 22525
rect 22094 22516 22100 22568
rect 22152 22556 22158 22568
rect 22465 22559 22523 22565
rect 22465 22556 22477 22559
rect 22152 22528 22477 22556
rect 22152 22516 22158 22528
rect 22465 22525 22477 22528
rect 22511 22525 22523 22559
rect 22465 22519 22523 22525
rect 22833 22559 22891 22565
rect 22833 22525 22845 22559
rect 22879 22556 22891 22559
rect 23661 22559 23719 22565
rect 23661 22556 23673 22559
rect 22879 22528 23673 22556
rect 22879 22525 22891 22528
rect 22833 22519 22891 22525
rect 23661 22525 23673 22528
rect 23707 22556 23719 22559
rect 24670 22556 24676 22568
rect 23707 22528 24256 22556
rect 24631 22528 24676 22556
rect 23707 22525 23719 22528
rect 23661 22519 23719 22525
rect 22741 22491 22799 22497
rect 22741 22457 22753 22491
rect 22787 22488 22799 22491
rect 22922 22488 22928 22500
rect 22787 22460 22928 22488
rect 22787 22457 22799 22460
rect 22741 22451 22799 22457
rect 22922 22448 22928 22460
rect 22980 22448 22986 22500
rect 24228 22497 24256 22528
rect 24670 22516 24676 22528
rect 24728 22556 24734 22568
rect 25133 22559 25191 22565
rect 25133 22556 25145 22559
rect 24728 22528 25145 22556
rect 24728 22516 24734 22528
rect 25133 22525 25145 22528
rect 25179 22525 25191 22559
rect 25133 22519 25191 22525
rect 25685 22559 25743 22565
rect 25685 22525 25697 22559
rect 25731 22556 25743 22559
rect 26234 22556 26240 22568
rect 25731 22528 26240 22556
rect 25731 22525 25743 22528
rect 25685 22519 25743 22525
rect 26234 22516 26240 22528
rect 26292 22516 26298 22568
rect 26786 22556 26792 22568
rect 26747 22528 26792 22556
rect 26786 22516 26792 22528
rect 26844 22516 26850 22568
rect 27154 22556 27160 22568
rect 27115 22528 27160 22556
rect 27154 22516 27160 22528
rect 27212 22516 27218 22568
rect 28077 22559 28135 22565
rect 28077 22525 28089 22559
rect 28123 22556 28135 22559
rect 28442 22556 28448 22568
rect 28123 22528 28448 22556
rect 28123 22525 28135 22528
rect 28077 22519 28135 22525
rect 28442 22516 28448 22528
rect 28500 22516 28506 22568
rect 29270 22556 29276 22568
rect 29231 22528 29276 22556
rect 29270 22516 29276 22528
rect 29328 22516 29334 22568
rect 29822 22516 29828 22568
rect 29880 22556 29886 22568
rect 30466 22556 30472 22568
rect 29880 22528 30472 22556
rect 29880 22516 29886 22528
rect 30466 22516 30472 22528
rect 30524 22516 30530 22568
rect 31018 22556 31024 22568
rect 30979 22528 31024 22556
rect 31018 22516 31024 22528
rect 31076 22516 31082 22568
rect 31205 22559 31263 22565
rect 31205 22525 31217 22559
rect 31251 22556 31263 22559
rect 32033 22559 32091 22565
rect 32033 22556 32045 22559
rect 31251 22528 32045 22556
rect 31251 22525 31263 22528
rect 31205 22519 31263 22525
rect 32033 22525 32045 22528
rect 32079 22556 32091 22559
rect 33229 22559 33287 22565
rect 33229 22556 33241 22559
rect 32079 22528 33241 22556
rect 32079 22525 32091 22528
rect 32033 22519 32091 22525
rect 33229 22525 33241 22528
rect 33275 22525 33287 22559
rect 33229 22519 33287 22525
rect 33594 22516 33600 22568
rect 33652 22556 33658 22568
rect 33816 22559 33874 22565
rect 33816 22556 33828 22559
rect 33652 22528 33828 22556
rect 33652 22516 33658 22528
rect 33816 22525 33828 22528
rect 33862 22556 33874 22559
rect 34241 22559 34299 22565
rect 34241 22556 34253 22559
rect 33862 22528 34253 22556
rect 33862 22525 33874 22528
rect 33816 22519 33874 22525
rect 34241 22525 34253 22528
rect 34287 22525 34299 22559
rect 34920 22559 34978 22565
rect 34920 22556 34932 22559
rect 34241 22519 34299 22525
rect 34440 22528 34932 22556
rect 24213 22491 24271 22497
rect 24213 22457 24225 22491
rect 24259 22488 24271 22491
rect 26804 22488 26832 22516
rect 29914 22488 29920 22500
rect 24259 22460 26832 22488
rect 28368 22460 29920 22488
rect 24259 22457 24271 22460
rect 24213 22451 24271 22457
rect 1946 22420 1952 22432
rect 1907 22392 1952 22420
rect 1946 22380 1952 22392
rect 2004 22380 2010 22432
rect 9674 22380 9680 22432
rect 9732 22420 9738 22432
rect 10134 22420 10140 22432
rect 9732 22392 10140 22420
rect 9732 22380 9738 22392
rect 10134 22380 10140 22392
rect 10192 22380 10198 22432
rect 11790 22420 11796 22432
rect 11751 22392 11796 22420
rect 11790 22380 11796 22392
rect 11848 22380 11854 22432
rect 13722 22420 13728 22432
rect 13683 22392 13728 22420
rect 13722 22380 13728 22392
rect 13780 22380 13786 22432
rect 14274 22420 14280 22432
rect 14235 22392 14280 22420
rect 14274 22380 14280 22392
rect 14332 22380 14338 22432
rect 15562 22380 15568 22432
rect 15620 22420 15626 22432
rect 18598 22420 18604 22432
rect 15620 22392 18604 22420
rect 15620 22380 15626 22392
rect 18598 22380 18604 22392
rect 18656 22420 18662 22432
rect 19061 22423 19119 22429
rect 19061 22420 19073 22423
rect 18656 22392 19073 22420
rect 18656 22380 18662 22392
rect 19061 22389 19073 22392
rect 19107 22389 19119 22423
rect 21818 22420 21824 22432
rect 21779 22392 21824 22420
rect 19061 22383 19119 22389
rect 21818 22380 21824 22392
rect 21876 22380 21882 22432
rect 23842 22420 23848 22432
rect 23803 22392 23848 22420
rect 23842 22380 23848 22392
rect 23900 22380 23906 22432
rect 24857 22423 24915 22429
rect 24857 22389 24869 22423
rect 24903 22420 24915 22423
rect 25774 22420 25780 22432
rect 24903 22392 25780 22420
rect 24903 22389 24915 22392
rect 24857 22383 24915 22389
rect 25774 22380 25780 22392
rect 25832 22380 25838 22432
rect 25869 22423 25927 22429
rect 25869 22389 25881 22423
rect 25915 22420 25927 22423
rect 28368 22420 28396 22460
rect 29914 22448 29920 22460
rect 29972 22448 29978 22500
rect 30009 22491 30067 22497
rect 30009 22457 30021 22491
rect 30055 22488 30067 22491
rect 31036 22488 31064 22516
rect 30055 22460 31064 22488
rect 32395 22491 32453 22497
rect 30055 22457 30067 22460
rect 30009 22451 30067 22457
rect 32395 22457 32407 22491
rect 32441 22457 32453 22491
rect 32395 22451 32453 22457
rect 25915 22392 28396 22420
rect 25915 22389 25927 22392
rect 25869 22383 25927 22389
rect 28442 22380 28448 22432
rect 28500 22420 28506 22432
rect 28997 22423 29055 22429
rect 28997 22420 29009 22423
rect 28500 22392 29009 22420
rect 28500 22380 28506 22392
rect 28997 22389 29009 22392
rect 29043 22389 29055 22423
rect 30282 22420 30288 22432
rect 30243 22392 30288 22420
rect 28997 22383 29055 22389
rect 30282 22380 30288 22392
rect 30340 22380 30346 22432
rect 31573 22423 31631 22429
rect 31573 22389 31585 22423
rect 31619 22420 31631 22423
rect 31849 22423 31907 22429
rect 31849 22420 31861 22423
rect 31619 22392 31861 22420
rect 31619 22389 31631 22392
rect 31573 22383 31631 22389
rect 31849 22389 31861 22392
rect 31895 22420 31907 22423
rect 32416 22420 32444 22451
rect 32490 22420 32496 22432
rect 31895 22392 32496 22420
rect 31895 22389 31907 22392
rect 31849 22383 31907 22389
rect 32490 22380 32496 22392
rect 32548 22380 32554 22432
rect 32950 22380 32956 22432
rect 33008 22420 33014 22432
rect 33612 22420 33640 22516
rect 33008 22392 33640 22420
rect 33008 22380 33014 22392
rect 34238 22380 34244 22432
rect 34296 22420 34302 22432
rect 34440 22420 34468 22528
rect 34920 22525 34932 22528
rect 34966 22525 34978 22559
rect 34920 22519 34978 22525
rect 36332 22559 36390 22565
rect 36332 22525 36344 22559
rect 36378 22556 36390 22559
rect 36722 22556 36728 22568
rect 36378 22528 36728 22556
rect 36378 22525 36390 22528
rect 36332 22519 36390 22525
rect 34606 22448 34612 22500
rect 34664 22488 34670 22500
rect 36347 22488 36375 22519
rect 36722 22516 36728 22528
rect 36780 22516 36786 22568
rect 37182 22516 37188 22568
rect 37240 22556 37246 22568
rect 37344 22559 37402 22565
rect 37344 22556 37356 22559
rect 37240 22528 37356 22556
rect 37240 22516 37246 22528
rect 37344 22525 37356 22528
rect 37390 22525 37402 22559
rect 38378 22556 38384 22568
rect 38339 22528 38384 22556
rect 37344 22519 37402 22525
rect 34664 22460 36375 22488
rect 37359 22488 37387 22519
rect 38378 22516 38384 22528
rect 38436 22516 38442 22568
rect 38856 22565 38884 22596
rect 39117 22593 39129 22627
rect 39163 22624 39175 22627
rect 39390 22624 39396 22636
rect 39163 22596 39396 22624
rect 39163 22593 39175 22596
rect 39117 22587 39175 22593
rect 39390 22584 39396 22596
rect 39448 22624 39454 22636
rect 39761 22627 39819 22633
rect 39761 22624 39773 22627
rect 39448 22596 39773 22624
rect 39448 22584 39454 22596
rect 39761 22593 39773 22596
rect 39807 22593 39819 22627
rect 39761 22587 39819 22593
rect 38841 22559 38899 22565
rect 38841 22525 38853 22559
rect 38887 22525 38899 22559
rect 38841 22519 38899 22525
rect 40402 22516 40408 22568
rect 40460 22556 40466 22568
rect 41559 22565 41587 22664
rect 41969 22661 41981 22664
rect 42015 22661 42027 22695
rect 41969 22655 42027 22661
rect 43162 22624 43168 22636
rect 43075 22596 43168 22624
rect 43162 22584 43168 22596
rect 43220 22624 43226 22636
rect 44174 22624 44180 22636
rect 43220 22596 44180 22624
rect 43220 22584 43226 22596
rect 44174 22584 44180 22596
rect 44232 22584 44238 22636
rect 40564 22559 40622 22565
rect 40564 22556 40576 22559
rect 40460 22528 40576 22556
rect 40460 22516 40466 22528
rect 40564 22525 40576 22528
rect 40610 22556 40622 22559
rect 41544 22559 41602 22565
rect 40610 22528 41092 22556
rect 40610 22525 40622 22528
rect 40564 22519 40622 22525
rect 37829 22491 37887 22497
rect 37829 22488 37841 22491
rect 37359 22460 37841 22488
rect 34664 22448 34670 22460
rect 37829 22457 37841 22460
rect 37875 22488 37887 22491
rect 40862 22488 40868 22500
rect 37875 22460 40868 22488
rect 37875 22457 37887 22460
rect 37829 22451 37887 22457
rect 40862 22448 40868 22460
rect 40920 22448 40926 22500
rect 35345 22423 35403 22429
rect 35345 22420 35357 22423
rect 34296 22392 35357 22420
rect 34296 22380 34302 22392
rect 35345 22389 35357 22392
rect 35391 22389 35403 22423
rect 35345 22383 35403 22389
rect 36170 22380 36176 22432
rect 36228 22420 36234 22432
rect 36403 22423 36461 22429
rect 36403 22420 36415 22423
rect 36228 22392 36415 22420
rect 36228 22380 36234 22392
rect 36403 22389 36415 22392
rect 36449 22389 36461 22423
rect 36403 22383 36461 22389
rect 39298 22380 39304 22432
rect 39356 22420 39362 22432
rect 39485 22423 39543 22429
rect 39485 22420 39497 22423
rect 39356 22392 39497 22420
rect 39356 22380 39362 22392
rect 39485 22389 39497 22392
rect 39531 22420 39543 22423
rect 40310 22420 40316 22432
rect 39531 22392 40316 22420
rect 39531 22389 39543 22392
rect 39485 22383 39543 22389
rect 40310 22380 40316 22392
rect 40368 22380 40374 22432
rect 41064 22429 41092 22528
rect 41544 22525 41556 22559
rect 41590 22525 41602 22559
rect 41544 22519 41602 22525
rect 43257 22491 43315 22497
rect 43257 22457 43269 22491
rect 43303 22457 43315 22491
rect 43806 22488 43812 22500
rect 43767 22460 43812 22488
rect 43257 22451 43315 22457
rect 41049 22423 41107 22429
rect 41049 22389 41061 22423
rect 41095 22420 41107 22423
rect 41138 22420 41144 22432
rect 41095 22392 41144 22420
rect 41095 22389 41107 22392
rect 41049 22383 41107 22389
rect 41138 22380 41144 22392
rect 41196 22380 41202 22432
rect 41647 22423 41705 22429
rect 41647 22389 41659 22423
rect 41693 22420 41705 22423
rect 41874 22420 41880 22432
rect 41693 22392 41880 22420
rect 41693 22389 41705 22392
rect 41647 22383 41705 22389
rect 41874 22380 41880 22392
rect 41932 22380 41938 22432
rect 42886 22380 42892 22432
rect 42944 22420 42950 22432
rect 42981 22423 43039 22429
rect 42981 22420 42993 22423
rect 42944 22392 42993 22420
rect 42944 22380 42950 22392
rect 42981 22389 42993 22392
rect 43027 22420 43039 22423
rect 43272 22420 43300 22451
rect 43806 22448 43812 22460
rect 43864 22448 43870 22500
rect 43622 22420 43628 22432
rect 43027 22392 43628 22420
rect 43027 22389 43039 22392
rect 42981 22383 43039 22389
rect 43622 22380 43628 22392
rect 43680 22420 43686 22432
rect 44085 22423 44143 22429
rect 44085 22420 44097 22423
rect 43680 22392 44097 22420
rect 43680 22380 43686 22392
rect 44085 22389 44097 22392
rect 44131 22389 44143 22423
rect 44910 22420 44916 22432
rect 44871 22392 44916 22420
rect 44085 22383 44143 22389
rect 44910 22380 44916 22392
rect 44968 22380 44974 22432
rect 1104 22330 48852 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 48852 22330
rect 1104 22256 48852 22278
rect 4341 22219 4399 22225
rect 4341 22185 4353 22219
rect 4387 22216 4399 22219
rect 4433 22219 4491 22225
rect 4433 22216 4445 22219
rect 4387 22188 4445 22216
rect 4387 22185 4399 22188
rect 4341 22179 4399 22185
rect 4433 22185 4445 22188
rect 4479 22216 4491 22219
rect 4614 22216 4620 22228
rect 4479 22188 4620 22216
rect 4479 22185 4491 22188
rect 4433 22179 4491 22185
rect 4614 22176 4620 22188
rect 4672 22176 4678 22228
rect 5442 22176 5448 22228
rect 5500 22216 5506 22228
rect 5537 22219 5595 22225
rect 5537 22216 5549 22219
rect 5500 22188 5549 22216
rect 5500 22176 5506 22188
rect 5537 22185 5549 22188
rect 5583 22185 5595 22219
rect 5537 22179 5595 22185
rect 6457 22219 6515 22225
rect 6457 22185 6469 22219
rect 6503 22216 6515 22219
rect 6730 22216 6736 22228
rect 6503 22188 6736 22216
rect 6503 22185 6515 22188
rect 6457 22179 6515 22185
rect 6730 22176 6736 22188
rect 6788 22176 6794 22228
rect 8297 22219 8355 22225
rect 8297 22185 8309 22219
rect 8343 22216 8355 22219
rect 8386 22216 8392 22228
rect 8343 22188 8392 22216
rect 8343 22185 8355 22188
rect 8297 22179 8355 22185
rect 8386 22176 8392 22188
rect 8444 22176 8450 22228
rect 8665 22219 8723 22225
rect 8665 22185 8677 22219
rect 8711 22216 8723 22219
rect 9582 22216 9588 22228
rect 8711 22188 9588 22216
rect 8711 22185 8723 22188
rect 8665 22179 8723 22185
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 10686 22216 10692 22228
rect 10647 22188 10692 22216
rect 10686 22176 10692 22188
rect 10744 22176 10750 22228
rect 13906 22176 13912 22228
rect 13964 22216 13970 22228
rect 14001 22219 14059 22225
rect 14001 22216 14013 22219
rect 13964 22188 14013 22216
rect 13964 22176 13970 22188
rect 14001 22185 14013 22188
rect 14047 22185 14059 22219
rect 14001 22179 14059 22185
rect 18690 22176 18696 22228
rect 18748 22216 18754 22228
rect 19475 22219 19533 22225
rect 19475 22216 19487 22219
rect 18748 22188 19487 22216
rect 18748 22176 18754 22188
rect 19475 22185 19487 22188
rect 19521 22185 19533 22219
rect 19475 22179 19533 22185
rect 23293 22219 23351 22225
rect 23293 22185 23305 22219
rect 23339 22216 23351 22219
rect 23474 22216 23480 22228
rect 23339 22188 23480 22216
rect 23339 22185 23351 22188
rect 23293 22179 23351 22185
rect 23474 22176 23480 22188
rect 23532 22176 23538 22228
rect 23845 22219 23903 22225
rect 23845 22185 23857 22219
rect 23891 22216 23903 22219
rect 24581 22219 24639 22225
rect 24581 22216 24593 22219
rect 23891 22188 24593 22216
rect 23891 22185 23903 22188
rect 23845 22179 23903 22185
rect 24581 22185 24593 22188
rect 24627 22216 24639 22219
rect 24762 22216 24768 22228
rect 24627 22188 24768 22216
rect 24627 22185 24639 22188
rect 24581 22179 24639 22185
rect 24762 22176 24768 22188
rect 24820 22216 24826 22228
rect 26786 22216 26792 22228
rect 24820 22188 24900 22216
rect 26747 22188 26792 22216
rect 24820 22176 24826 22188
rect 2777 22151 2835 22157
rect 2777 22117 2789 22151
rect 2823 22148 2835 22151
rect 3786 22148 3792 22160
rect 2823 22120 3792 22148
rect 2823 22117 2835 22120
rect 2777 22111 2835 22117
rect 3786 22108 3792 22120
rect 3844 22108 3850 22160
rect 7101 22151 7159 22157
rect 7101 22117 7113 22151
rect 7147 22148 7159 22151
rect 7190 22148 7196 22160
rect 7147 22120 7196 22148
rect 7147 22117 7159 22120
rect 7101 22111 7159 22117
rect 7190 22108 7196 22120
rect 7248 22108 7254 22160
rect 13354 22148 13360 22160
rect 13315 22120 13360 22148
rect 13354 22108 13360 22120
rect 13412 22108 13418 22160
rect 15194 22108 15200 22160
rect 15252 22148 15258 22160
rect 15473 22151 15531 22157
rect 15473 22148 15485 22151
rect 15252 22120 15485 22148
rect 15252 22108 15258 22120
rect 15473 22117 15485 22120
rect 15519 22148 15531 22151
rect 17310 22148 17316 22160
rect 15519 22120 17316 22148
rect 15519 22117 15531 22120
rect 15473 22111 15531 22117
rect 17310 22108 17316 22120
rect 17368 22108 17374 22160
rect 17862 22148 17868 22160
rect 17823 22120 17868 22148
rect 17862 22108 17868 22120
rect 17920 22108 17926 22160
rect 17957 22151 18015 22157
rect 17957 22117 17969 22151
rect 18003 22148 18015 22151
rect 18046 22148 18052 22160
rect 18003 22120 18052 22148
rect 18003 22117 18015 22120
rect 17957 22111 18015 22117
rect 18046 22108 18052 22120
rect 18104 22108 18110 22160
rect 18782 22148 18788 22160
rect 18743 22120 18788 22148
rect 18782 22108 18788 22120
rect 18840 22108 18846 22160
rect 21082 22148 21088 22160
rect 21043 22120 21088 22148
rect 21082 22108 21088 22120
rect 21140 22108 21146 22160
rect 21637 22151 21695 22157
rect 21637 22117 21649 22151
rect 21683 22148 21695 22151
rect 21726 22148 21732 22160
rect 21683 22120 21732 22148
rect 21683 22117 21695 22120
rect 21637 22111 21695 22117
rect 21726 22108 21732 22120
rect 21784 22108 21790 22160
rect 24872 22157 24900 22188
rect 26786 22176 26792 22188
rect 26844 22176 26850 22228
rect 28534 22176 28540 22228
rect 28592 22216 28598 22228
rect 31110 22216 31116 22228
rect 28592 22188 31116 22216
rect 28592 22176 28598 22188
rect 31110 22176 31116 22188
rect 31168 22176 31174 22228
rect 32907 22219 32965 22225
rect 32907 22185 32919 22219
rect 32953 22216 32965 22219
rect 33318 22216 33324 22228
rect 32953 22188 33324 22216
rect 32953 22185 32965 22188
rect 32907 22179 32965 22185
rect 33318 22176 33324 22188
rect 33376 22176 33382 22228
rect 38378 22216 38384 22228
rect 33888 22188 38384 22216
rect 24857 22151 24915 22157
rect 24857 22117 24869 22151
rect 24903 22117 24915 22151
rect 24857 22111 24915 22117
rect 25774 22108 25780 22160
rect 25832 22148 25838 22160
rect 28718 22148 28724 22160
rect 25832 22120 28724 22148
rect 25832 22108 25838 22120
rect 28718 22108 28724 22120
rect 28776 22108 28782 22160
rect 28813 22151 28871 22157
rect 28813 22117 28825 22151
rect 28859 22148 28871 22151
rect 29270 22148 29276 22160
rect 28859 22120 29276 22148
rect 28859 22117 28871 22120
rect 28813 22111 28871 22117
rect 29270 22108 29276 22120
rect 29328 22108 29334 22160
rect 30374 22108 30380 22160
rect 30432 22148 30438 22160
rect 31205 22151 31263 22157
rect 30432 22120 31156 22148
rect 30432 22108 30438 22120
rect 2130 22080 2136 22092
rect 2091 22052 2136 22080
rect 2130 22040 2136 22052
rect 2188 22040 2194 22092
rect 4062 22040 4068 22092
rect 4120 22080 4126 22092
rect 4157 22083 4215 22089
rect 4157 22080 4169 22083
rect 4120 22052 4169 22080
rect 4120 22040 4126 22052
rect 4157 22049 4169 22052
rect 4203 22049 4215 22083
rect 4157 22043 4215 22049
rect 8294 22040 8300 22092
rect 8352 22080 8358 22092
rect 8481 22083 8539 22089
rect 8481 22080 8493 22083
rect 8352 22052 8493 22080
rect 8352 22040 8358 22052
rect 8481 22049 8493 22052
rect 8527 22049 8539 22083
rect 9674 22080 9680 22092
rect 9635 22052 9680 22080
rect 8481 22043 8539 22049
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 11517 22083 11575 22089
rect 11517 22049 11529 22083
rect 11563 22080 11575 22083
rect 11790 22080 11796 22092
rect 11563 22052 11796 22080
rect 11563 22049 11575 22052
rect 11517 22043 11575 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 12618 22080 12624 22092
rect 12579 22052 12624 22080
rect 12618 22040 12624 22052
rect 12676 22040 12682 22092
rect 13081 22083 13139 22089
rect 13081 22049 13093 22083
rect 13127 22049 13139 22083
rect 13081 22043 13139 22049
rect 14185 22083 14243 22089
rect 14185 22049 14197 22083
rect 14231 22080 14243 22083
rect 14274 22080 14280 22092
rect 14231 22052 14280 22080
rect 14231 22049 14243 22052
rect 14185 22043 14243 22049
rect 5166 22012 5172 22024
rect 5127 21984 5172 22012
rect 5166 21972 5172 21984
rect 5224 21972 5230 22024
rect 7006 22012 7012 22024
rect 6967 21984 7012 22012
rect 7006 21972 7012 21984
rect 7064 21972 7070 22024
rect 13096 21956 13124 22043
rect 14274 22040 14280 22052
rect 14332 22040 14338 22092
rect 19242 22040 19248 22092
rect 19300 22080 19306 22092
rect 19372 22083 19430 22089
rect 19372 22080 19384 22083
rect 19300 22052 19384 22080
rect 19300 22040 19306 22052
rect 19372 22049 19384 22052
rect 19418 22049 19430 22083
rect 26970 22080 26976 22092
rect 19372 22043 19430 22049
rect 26252 22052 26976 22080
rect 15381 22015 15439 22021
rect 15381 22012 15393 22015
rect 14338 21984 15393 22012
rect 3510 21904 3516 21956
rect 3568 21944 3574 21956
rect 6089 21947 6147 21953
rect 6089 21944 6101 21947
rect 3568 21916 6101 21944
rect 3568 21904 3574 21916
rect 6089 21913 6101 21916
rect 6135 21913 6147 21947
rect 7558 21944 7564 21956
rect 7519 21916 7564 21944
rect 6089 21907 6147 21913
rect 7558 21904 7564 21916
rect 7616 21904 7622 21956
rect 9861 21947 9919 21953
rect 9861 21913 9873 21947
rect 9907 21944 9919 21947
rect 10134 21944 10140 21956
rect 9907 21916 10140 21944
rect 9907 21913 9919 21916
rect 9861 21907 9919 21913
rect 10134 21904 10140 21916
rect 10192 21944 10198 21956
rect 11606 21944 11612 21956
rect 10192 21916 11612 21944
rect 10192 21904 10198 21916
rect 11606 21904 11612 21916
rect 11664 21904 11670 21956
rect 13078 21904 13084 21956
rect 13136 21944 13142 21956
rect 13630 21944 13636 21956
rect 13136 21916 13636 21944
rect 13136 21904 13142 21916
rect 13630 21904 13636 21916
rect 13688 21904 13694 21956
rect 14338 21953 14366 21984
rect 15381 21981 15393 21984
rect 15427 22012 15439 22015
rect 16114 22012 16120 22024
rect 15427 21984 16120 22012
rect 15427 21981 15439 21984
rect 15381 21975 15439 21981
rect 16114 21972 16120 21984
rect 16172 21972 16178 22024
rect 18509 22015 18567 22021
rect 18509 21981 18521 22015
rect 18555 22012 18567 22015
rect 18598 22012 18604 22024
rect 18555 21984 18604 22012
rect 18555 21981 18567 21984
rect 18509 21975 18567 21981
rect 18598 21972 18604 21984
rect 18656 21972 18662 22024
rect 20990 22012 20996 22024
rect 20951 21984 20996 22012
rect 20990 21972 20996 21984
rect 21048 21972 21054 22024
rect 22922 22012 22928 22024
rect 22883 21984 22928 22012
rect 22922 21972 22928 21984
rect 22980 21972 22986 22024
rect 24762 22012 24768 22024
rect 24723 21984 24768 22012
rect 24762 21972 24768 21984
rect 24820 21972 24826 22024
rect 25038 22012 25044 22024
rect 24999 21984 25044 22012
rect 25038 21972 25044 21984
rect 25096 21972 25102 22024
rect 14323 21947 14381 21953
rect 14323 21913 14335 21947
rect 14369 21913 14381 21947
rect 14323 21907 14381 21913
rect 15933 21947 15991 21953
rect 15933 21913 15945 21947
rect 15979 21944 15991 21947
rect 16022 21944 16028 21956
rect 15979 21916 16028 21944
rect 15979 21913 15991 21916
rect 15933 21907 15991 21913
rect 16022 21904 16028 21916
rect 16080 21904 16086 21956
rect 19426 21904 19432 21956
rect 19484 21944 19490 21956
rect 26252 21944 26280 22052
rect 26970 22040 26976 22052
rect 27028 22080 27034 22092
rect 27065 22083 27123 22089
rect 27065 22080 27077 22083
rect 27028 22052 27077 22080
rect 27028 22040 27034 22052
rect 27065 22049 27077 22052
rect 27111 22080 27123 22083
rect 27522 22080 27528 22092
rect 27111 22052 27528 22080
rect 27111 22049 27123 22052
rect 27065 22043 27123 22049
rect 27522 22040 27528 22052
rect 27580 22040 27586 22092
rect 28077 22083 28135 22089
rect 28077 22049 28089 22083
rect 28123 22080 28135 22083
rect 29086 22080 29092 22092
rect 28123 22052 29092 22080
rect 28123 22049 28135 22052
rect 28077 22043 28135 22049
rect 29086 22040 29092 22052
rect 29144 22040 29150 22092
rect 30484 22089 30512 22120
rect 30469 22083 30527 22089
rect 30469 22049 30481 22083
rect 30515 22049 30527 22083
rect 31018 22080 31024 22092
rect 30931 22052 31024 22080
rect 30469 22043 30527 22049
rect 31018 22040 31024 22052
rect 31076 22040 31082 22092
rect 31128 22080 31156 22120
rect 31205 22117 31217 22151
rect 31251 22148 31263 22151
rect 32122 22148 32128 22160
rect 31251 22120 32128 22148
rect 31251 22117 31263 22120
rect 31205 22111 31263 22117
rect 32122 22108 32128 22120
rect 32180 22148 32186 22160
rect 32309 22151 32367 22157
rect 32309 22148 32321 22151
rect 32180 22120 32321 22148
rect 32180 22108 32186 22120
rect 32309 22117 32321 22120
rect 32355 22117 32367 22151
rect 33888 22148 33916 22188
rect 38378 22176 38384 22188
rect 38436 22176 38442 22228
rect 41874 22176 41880 22228
rect 41932 22216 41938 22228
rect 42245 22219 42303 22225
rect 42245 22216 42257 22219
rect 41932 22188 42257 22216
rect 41932 22176 41938 22188
rect 42245 22185 42257 22188
rect 42291 22216 42303 22219
rect 42334 22216 42340 22228
rect 42291 22188 42340 22216
rect 42291 22185 42303 22188
rect 42245 22179 42303 22185
rect 42334 22176 42340 22188
rect 42392 22176 42398 22228
rect 43162 22216 43168 22228
rect 43123 22188 43168 22216
rect 43162 22176 43168 22188
rect 43220 22176 43226 22228
rect 32309 22111 32367 22117
rect 32416 22120 33916 22148
rect 33965 22151 34023 22157
rect 32416 22080 32444 22120
rect 33965 22117 33977 22151
rect 34011 22148 34023 22151
rect 34514 22148 34520 22160
rect 34011 22120 34520 22148
rect 34011 22117 34023 22120
rect 33965 22111 34023 22117
rect 34514 22108 34520 22120
rect 34572 22108 34578 22160
rect 35989 22151 36047 22157
rect 35989 22117 36001 22151
rect 36035 22148 36047 22151
rect 36170 22148 36176 22160
rect 36035 22120 36176 22148
rect 36035 22117 36047 22120
rect 35989 22111 36047 22117
rect 36170 22108 36176 22120
rect 36228 22108 36234 22160
rect 36262 22108 36268 22160
rect 36320 22148 36326 22160
rect 41417 22151 41475 22157
rect 36320 22120 36365 22148
rect 36320 22108 36326 22120
rect 41417 22117 41429 22151
rect 41463 22148 41475 22151
rect 41690 22148 41696 22160
rect 41463 22120 41696 22148
rect 41463 22117 41475 22120
rect 41417 22111 41475 22117
rect 41690 22108 41696 22120
rect 41748 22108 41754 22160
rect 31128 22052 32444 22080
rect 32836 22083 32894 22089
rect 32836 22049 32848 22083
rect 32882 22080 32894 22083
rect 33134 22080 33140 22092
rect 32882 22052 33140 22080
rect 32882 22049 32894 22052
rect 32836 22043 32894 22049
rect 33134 22040 33140 22052
rect 33192 22040 33198 22092
rect 37826 22089 37832 22092
rect 37804 22083 37832 22089
rect 37804 22080 37816 22083
rect 37739 22052 37816 22080
rect 37804 22049 37816 22052
rect 37884 22080 37890 22092
rect 38286 22080 38292 22092
rect 37884 22052 38292 22080
rect 37804 22043 37832 22049
rect 37826 22040 37832 22043
rect 37884 22040 37890 22052
rect 38286 22040 38292 22052
rect 38344 22040 38350 22092
rect 38749 22083 38807 22089
rect 38749 22049 38761 22083
rect 38795 22049 38807 22083
rect 39206 22080 39212 22092
rect 39167 22052 39212 22080
rect 38749 22043 38807 22049
rect 28166 22012 28172 22024
rect 19484 21916 26280 21944
rect 26896 21984 28172 22012
rect 19484 21904 19490 21916
rect 2682 21836 2688 21888
rect 2740 21876 2746 21888
rect 4433 21879 4491 21885
rect 4433 21876 4445 21879
rect 2740 21848 4445 21876
rect 2740 21836 2746 21848
rect 4433 21845 4445 21848
rect 4479 21845 4491 21879
rect 4982 21876 4988 21888
rect 4943 21848 4988 21876
rect 4433 21839 4491 21845
rect 4982 21836 4988 21848
rect 5040 21836 5046 21888
rect 10226 21836 10232 21888
rect 10284 21876 10290 21888
rect 10594 21876 10600 21888
rect 10284 21848 10600 21876
rect 10284 21836 10290 21848
rect 10594 21836 10600 21848
rect 10652 21876 10658 21888
rect 10965 21879 11023 21885
rect 10965 21876 10977 21879
rect 10652 21848 10977 21876
rect 10652 21836 10658 21848
rect 10965 21845 10977 21848
rect 11011 21845 11023 21879
rect 10965 21839 11023 21845
rect 11701 21879 11759 21885
rect 11701 21845 11713 21879
rect 11747 21876 11759 21879
rect 13354 21876 13360 21888
rect 11747 21848 13360 21876
rect 11747 21845 11759 21848
rect 11701 21839 11759 21845
rect 13354 21836 13360 21848
rect 13412 21836 13418 21888
rect 20165 21879 20223 21885
rect 20165 21845 20177 21879
rect 20211 21876 20223 21879
rect 20254 21876 20260 21888
rect 20211 21848 20260 21876
rect 20211 21845 20223 21848
rect 20165 21839 20223 21845
rect 20254 21836 20260 21848
rect 20312 21836 20318 21888
rect 22094 21876 22100 21888
rect 22055 21848 22100 21876
rect 22094 21836 22100 21848
rect 22152 21876 22158 21888
rect 22373 21879 22431 21885
rect 22373 21876 22385 21879
rect 22152 21848 22385 21876
rect 22152 21836 22158 21848
rect 22373 21845 22385 21848
rect 22419 21845 22431 21879
rect 22373 21839 22431 21845
rect 25498 21836 25504 21888
rect 25556 21876 25562 21888
rect 25777 21879 25835 21885
rect 25777 21876 25789 21879
rect 25556 21848 25789 21876
rect 25556 21836 25562 21848
rect 25777 21845 25789 21848
rect 25823 21876 25835 21879
rect 26896 21876 26924 21984
rect 28166 21972 28172 21984
rect 28224 21972 28230 22024
rect 28442 22012 28448 22024
rect 28403 21984 28448 22012
rect 28442 21972 28448 21984
rect 28500 21972 28506 22024
rect 30377 22015 30435 22021
rect 30377 21981 30389 22015
rect 30423 22012 30435 22015
rect 31036 22012 31064 22040
rect 33870 22012 33876 22024
rect 30423 21984 33134 22012
rect 33831 21984 33876 22012
rect 30423 21981 30435 21984
rect 30377 21975 30435 21981
rect 27617 21947 27675 21953
rect 27617 21913 27629 21947
rect 27663 21944 27675 21947
rect 29365 21947 29423 21953
rect 27663 21916 28028 21944
rect 27663 21913 27675 21916
rect 27617 21907 27675 21913
rect 28000 21888 28028 21916
rect 29365 21913 29377 21947
rect 29411 21944 29423 21947
rect 29546 21944 29552 21956
rect 29411 21916 29552 21944
rect 29411 21913 29423 21916
rect 29365 21907 29423 21913
rect 29546 21904 29552 21916
rect 29604 21904 29610 21956
rect 33106 21944 33134 21984
rect 33870 21972 33876 21984
rect 33928 21972 33934 22024
rect 34146 22012 34152 22024
rect 34107 21984 34152 22012
rect 34146 21972 34152 21984
rect 34204 21972 34210 22024
rect 36814 22012 36820 22024
rect 36775 21984 36820 22012
rect 36814 21972 36820 21984
rect 36872 21972 36878 22024
rect 38194 21972 38200 22024
rect 38252 22012 38258 22024
rect 38764 22012 38792 22043
rect 39206 22040 39212 22052
rect 39264 22040 39270 22092
rect 42978 22040 42984 22092
rect 43036 22080 43042 22092
rect 43346 22080 43352 22092
rect 43404 22089 43410 22092
rect 43404 22083 43442 22089
rect 43036 22052 43352 22080
rect 43036 22040 43042 22052
rect 43346 22040 43352 22052
rect 43430 22049 43442 22083
rect 43404 22043 43442 22049
rect 44361 22083 44419 22089
rect 44361 22049 44373 22083
rect 44407 22080 44419 22083
rect 44818 22080 44824 22092
rect 44407 22052 44824 22080
rect 44407 22049 44419 22052
rect 44361 22043 44419 22049
rect 43404 22040 43410 22043
rect 44818 22040 44824 22052
rect 44876 22040 44882 22092
rect 39482 22012 39488 22024
rect 38252 21984 38792 22012
rect 39443 21984 39488 22012
rect 38252 21972 38258 21984
rect 39482 21972 39488 21984
rect 39540 21972 39546 22024
rect 41322 22012 41328 22024
rect 41283 21984 41328 22012
rect 41322 21972 41328 21984
rect 41380 21972 41386 22024
rect 41601 22015 41659 22021
rect 41601 21981 41613 22015
rect 41647 22012 41659 22015
rect 41782 22012 41788 22024
rect 41647 21984 41788 22012
rect 41647 21981 41659 21984
rect 41601 21975 41659 21981
rect 40586 21944 40592 21956
rect 33106 21916 40592 21944
rect 40586 21904 40592 21916
rect 40644 21904 40650 21956
rect 40954 21904 40960 21956
rect 41012 21944 41018 21956
rect 41616 21944 41644 21975
rect 41782 21972 41788 21984
rect 41840 22012 41846 22024
rect 43806 22012 43812 22024
rect 41840 21984 43812 22012
rect 41840 21972 41846 21984
rect 43806 21972 43812 21984
rect 43864 21972 43870 22024
rect 43901 22015 43959 22021
rect 43901 21981 43913 22015
rect 43947 22012 43959 22015
rect 43990 22012 43996 22024
rect 43947 21984 43996 22012
rect 43947 21981 43959 21984
rect 43901 21975 43959 21981
rect 43990 21972 43996 21984
rect 44048 21972 44054 22024
rect 41012 21916 41644 21944
rect 43487 21947 43545 21953
rect 41012 21904 41018 21916
rect 43487 21913 43499 21947
rect 43533 21944 43545 21947
rect 43533 21916 43944 21944
rect 43533 21913 43545 21916
rect 43487 21907 43545 21913
rect 43916 21888 43944 21916
rect 25823 21848 26924 21876
rect 27249 21879 27307 21885
rect 25823 21845 25835 21848
rect 25777 21839 25835 21845
rect 27249 21845 27261 21879
rect 27295 21876 27307 21879
rect 27338 21876 27344 21888
rect 27295 21848 27344 21876
rect 27295 21845 27307 21848
rect 27249 21839 27307 21845
rect 27338 21836 27344 21848
rect 27396 21836 27402 21888
rect 27522 21836 27528 21888
rect 27580 21876 27586 21888
rect 27893 21879 27951 21885
rect 27893 21876 27905 21879
rect 27580 21848 27905 21876
rect 27580 21836 27586 21848
rect 27893 21845 27905 21848
rect 27939 21845 27951 21879
rect 27893 21839 27951 21845
rect 27982 21836 27988 21888
rect 28040 21876 28046 21888
rect 28215 21879 28273 21885
rect 28215 21876 28227 21879
rect 28040 21848 28227 21876
rect 28040 21836 28046 21848
rect 28215 21845 28227 21848
rect 28261 21845 28273 21879
rect 28350 21876 28356 21888
rect 28311 21848 28356 21876
rect 28215 21839 28273 21845
rect 28350 21836 28356 21848
rect 28408 21836 28414 21888
rect 29270 21836 29276 21888
rect 29328 21876 29334 21888
rect 29641 21879 29699 21885
rect 29641 21876 29653 21879
rect 29328 21848 29653 21876
rect 29328 21836 29334 21848
rect 29641 21845 29653 21848
rect 29687 21845 29699 21879
rect 35342 21876 35348 21888
rect 35303 21848 35348 21876
rect 29641 21839 29699 21845
rect 35342 21836 35348 21848
rect 35400 21836 35406 21888
rect 36906 21836 36912 21888
rect 36964 21876 36970 21888
rect 37875 21879 37933 21885
rect 37875 21876 37887 21879
rect 36964 21848 37887 21876
rect 36964 21836 36970 21848
rect 37875 21845 37887 21848
rect 37921 21845 37933 21879
rect 40494 21876 40500 21888
rect 40455 21848 40500 21876
rect 37875 21839 37933 21845
rect 40494 21836 40500 21848
rect 40552 21836 40558 21888
rect 43898 21836 43904 21888
rect 43956 21876 43962 21888
rect 44177 21879 44235 21885
rect 44177 21876 44189 21879
rect 43956 21848 44189 21876
rect 43956 21836 43962 21848
rect 44177 21845 44189 21848
rect 44223 21845 44235 21879
rect 44542 21876 44548 21888
rect 44503 21848 44548 21876
rect 44177 21839 44235 21845
rect 44542 21836 44548 21848
rect 44600 21836 44606 21888
rect 1104 21786 48852 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 48852 21786
rect 1104 21712 48852 21734
rect 2501 21675 2559 21681
rect 2501 21641 2513 21675
rect 2547 21672 2559 21675
rect 3326 21672 3332 21684
rect 2547 21644 3332 21672
rect 2547 21641 2559 21644
rect 2501 21635 2559 21641
rect 3326 21632 3332 21644
rect 3384 21632 3390 21684
rect 3510 21672 3516 21684
rect 3471 21644 3516 21672
rect 3510 21632 3516 21644
rect 3568 21632 3574 21684
rect 4062 21672 4068 21684
rect 4023 21644 4068 21672
rect 4062 21632 4068 21644
rect 4120 21632 4126 21684
rect 4525 21675 4583 21681
rect 4525 21641 4537 21675
rect 4571 21672 4583 21675
rect 5442 21672 5448 21684
rect 4571 21644 5448 21672
rect 4571 21641 4583 21644
rect 4525 21635 4583 21641
rect 5442 21632 5448 21644
rect 5500 21672 5506 21684
rect 5813 21675 5871 21681
rect 5813 21672 5825 21675
rect 5500 21644 5825 21672
rect 5500 21632 5506 21644
rect 5813 21641 5825 21644
rect 5859 21641 5871 21675
rect 5813 21635 5871 21641
rect 8021 21675 8079 21681
rect 8021 21641 8033 21675
rect 8067 21672 8079 21675
rect 8294 21672 8300 21684
rect 8067 21644 8300 21672
rect 8067 21641 8079 21644
rect 8021 21635 8079 21641
rect 8294 21632 8300 21644
rect 8352 21632 8358 21684
rect 8386 21632 8392 21684
rect 8444 21672 8450 21684
rect 11790 21672 11796 21684
rect 8444 21644 8489 21672
rect 11751 21644 11796 21672
rect 8444 21632 8450 21644
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 12618 21632 12624 21684
rect 12676 21672 12682 21684
rect 12897 21675 12955 21681
rect 12897 21672 12909 21675
rect 12676 21644 12909 21672
rect 12676 21632 12682 21644
rect 12897 21641 12909 21644
rect 12943 21641 12955 21675
rect 15194 21672 15200 21684
rect 15155 21644 15200 21672
rect 12897 21635 12955 21641
rect 15194 21632 15200 21644
rect 15252 21632 15258 21684
rect 17497 21675 17555 21681
rect 17497 21641 17509 21675
rect 17543 21672 17555 21675
rect 17862 21672 17868 21684
rect 17543 21644 17868 21672
rect 17543 21641 17555 21644
rect 17497 21635 17555 21641
rect 17862 21632 17868 21644
rect 17920 21632 17926 21684
rect 19242 21672 19248 21684
rect 19203 21644 19248 21672
rect 19242 21632 19248 21644
rect 19300 21632 19306 21684
rect 19426 21632 19432 21684
rect 19484 21672 19490 21684
rect 19521 21675 19579 21681
rect 19521 21672 19533 21675
rect 19484 21644 19533 21672
rect 19484 21632 19490 21644
rect 19521 21641 19533 21644
rect 19567 21641 19579 21675
rect 19521 21635 19579 21641
rect 20993 21675 21051 21681
rect 20993 21641 21005 21675
rect 21039 21672 21051 21675
rect 21082 21672 21088 21684
rect 21039 21644 21088 21672
rect 21039 21641 21051 21644
rect 20993 21635 21051 21641
rect 9309 21607 9367 21613
rect 9309 21604 9321 21607
rect 8496 21576 9321 21604
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21536 4675 21539
rect 4982 21536 4988 21548
rect 4663 21508 4988 21536
rect 4663 21505 4675 21508
rect 4617 21499 4675 21505
rect 4982 21496 4988 21508
rect 5040 21496 5046 21548
rect 2130 21468 2136 21480
rect 2043 21440 2136 21468
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 2056 21341 2084 21440
rect 2130 21428 2136 21440
rect 2188 21468 2194 21480
rect 2317 21471 2375 21477
rect 2317 21468 2329 21471
rect 2188 21440 2329 21468
rect 2188 21428 2194 21440
rect 2317 21437 2329 21440
rect 2363 21468 2375 21471
rect 2777 21471 2835 21477
rect 2777 21468 2789 21471
rect 2363 21440 2789 21468
rect 2363 21437 2375 21440
rect 2317 21431 2375 21437
rect 2777 21437 2789 21440
rect 2823 21437 2835 21471
rect 2777 21431 2835 21437
rect 3510 21428 3516 21480
rect 3568 21468 3574 21480
rect 3640 21471 3698 21477
rect 3640 21468 3652 21471
rect 3568 21440 3652 21468
rect 3568 21428 3574 21440
rect 3640 21437 3652 21440
rect 3686 21437 3698 21471
rect 3640 21431 3698 21437
rect 3743 21471 3801 21477
rect 3743 21437 3755 21471
rect 3789 21468 3801 21471
rect 6181 21471 6239 21477
rect 6181 21468 6193 21471
rect 3789 21440 6193 21468
rect 3789 21437 3801 21440
rect 3743 21431 3801 21437
rect 6181 21437 6193 21440
rect 6227 21437 6239 21471
rect 6181 21431 6239 21437
rect 4706 21360 4712 21412
rect 4764 21400 4770 21412
rect 4979 21403 5037 21409
rect 4979 21400 4991 21403
rect 4764 21372 4991 21400
rect 4764 21360 4770 21372
rect 4979 21369 4991 21372
rect 5025 21400 5037 21403
rect 5442 21400 5448 21412
rect 5025 21372 5448 21400
rect 5025 21369 5037 21372
rect 4979 21363 5037 21369
rect 5442 21360 5448 21372
rect 5500 21360 5506 21412
rect 6196 21400 6224 21431
rect 8110 21428 8116 21480
rect 8168 21468 8174 21480
rect 8496 21477 8524 21576
rect 9309 21573 9321 21576
rect 9355 21573 9367 21607
rect 9309 21567 9367 21573
rect 9398 21564 9404 21616
rect 9456 21604 9462 21616
rect 10689 21607 10747 21613
rect 10689 21604 10701 21607
rect 9456 21576 10701 21604
rect 9456 21564 9462 21576
rect 10689 21573 10701 21576
rect 10735 21604 10747 21607
rect 10962 21604 10968 21616
rect 10735 21576 10968 21604
rect 10735 21573 10747 21576
rect 10689 21567 10747 21573
rect 10962 21564 10968 21576
rect 11020 21604 11026 21616
rect 13998 21604 14004 21616
rect 11020 21576 14004 21604
rect 11020 21564 11026 21576
rect 13998 21564 14004 21576
rect 14056 21604 14062 21616
rect 15212 21604 15240 21632
rect 14056 21576 15240 21604
rect 17773 21607 17831 21613
rect 14056 21564 14062 21576
rect 17773 21573 17785 21607
rect 17819 21604 17831 21607
rect 18046 21604 18052 21616
rect 17819 21576 18052 21604
rect 17819 21573 17831 21576
rect 17773 21567 17831 21573
rect 18046 21564 18052 21576
rect 18104 21564 18110 21616
rect 9033 21539 9091 21545
rect 9033 21505 9045 21539
rect 9079 21536 9091 21539
rect 9674 21536 9680 21548
rect 9079 21508 9680 21536
rect 9079 21505 9091 21508
rect 9033 21499 9091 21505
rect 9674 21496 9680 21508
rect 9732 21496 9738 21548
rect 13906 21536 13912 21548
rect 13867 21508 13912 21536
rect 13906 21496 13912 21508
rect 13964 21496 13970 21548
rect 16022 21536 16028 21548
rect 15983 21508 16028 21536
rect 16022 21496 16028 21508
rect 16080 21536 16086 21548
rect 18141 21539 18199 21545
rect 18141 21536 18153 21539
rect 16080 21508 18153 21536
rect 16080 21496 16086 21508
rect 18141 21505 18153 21508
rect 18187 21536 18199 21539
rect 18506 21536 18512 21548
rect 18187 21508 18512 21536
rect 18187 21505 18199 21508
rect 18141 21499 18199 21505
rect 18506 21496 18512 21508
rect 18564 21496 18570 21548
rect 18598 21496 18604 21548
rect 18656 21536 18662 21548
rect 18656 21508 18701 21536
rect 18656 21496 18662 21508
rect 8481 21471 8539 21477
rect 8481 21468 8493 21471
rect 8168 21440 8493 21468
rect 8168 21428 8174 21440
rect 8481 21437 8493 21440
rect 8527 21437 8539 21471
rect 8481 21431 8539 21437
rect 8665 21471 8723 21477
rect 8665 21437 8677 21471
rect 8711 21437 8723 21471
rect 12472 21471 12530 21477
rect 12472 21468 12484 21471
rect 8665 21431 8723 21437
rect 12176 21440 12484 21468
rect 6917 21403 6975 21409
rect 6917 21400 6929 21403
rect 6196 21372 6929 21400
rect 6917 21369 6929 21372
rect 6963 21369 6975 21403
rect 6917 21363 6975 21369
rect 7009 21403 7067 21409
rect 7009 21369 7021 21403
rect 7055 21369 7067 21403
rect 7558 21400 7564 21412
rect 7519 21372 7564 21400
rect 7009 21363 7067 21369
rect 2041 21335 2099 21341
rect 2041 21332 2053 21335
rect 1452 21304 2053 21332
rect 1452 21292 1458 21304
rect 2041 21301 2053 21304
rect 2087 21301 2099 21335
rect 5534 21332 5540 21344
rect 5495 21304 5540 21332
rect 2041 21295 2099 21301
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 6641 21335 6699 21341
rect 6641 21301 6653 21335
rect 6687 21332 6699 21335
rect 6730 21332 6736 21344
rect 6687 21304 6736 21332
rect 6687 21301 6699 21304
rect 6641 21295 6699 21301
rect 6730 21292 6736 21304
rect 6788 21332 6794 21344
rect 7024 21332 7052 21363
rect 7558 21360 7564 21372
rect 7616 21360 7622 21412
rect 8386 21360 8392 21412
rect 8444 21400 8450 21412
rect 8680 21400 8708 21431
rect 8444 21372 8708 21400
rect 10321 21403 10379 21409
rect 8444 21360 8450 21372
rect 10321 21369 10333 21403
rect 10367 21400 10379 21403
rect 10870 21400 10876 21412
rect 10367 21372 10876 21400
rect 10367 21369 10379 21372
rect 10321 21363 10379 21369
rect 10870 21360 10876 21372
rect 10928 21360 10934 21412
rect 10962 21360 10968 21412
rect 11020 21400 11026 21412
rect 11517 21403 11575 21409
rect 11020 21372 11065 21400
rect 11020 21360 11026 21372
rect 11517 21369 11529 21403
rect 11563 21400 11575 21403
rect 12066 21400 12072 21412
rect 11563 21372 12072 21400
rect 11563 21369 11575 21372
rect 11517 21363 11575 21369
rect 12066 21360 12072 21372
rect 12124 21360 12130 21412
rect 12176 21344 12204 21440
rect 12472 21437 12484 21440
rect 12518 21437 12530 21471
rect 12472 21431 12530 21437
rect 13630 21428 13636 21480
rect 13688 21468 13694 21480
rect 13725 21471 13783 21477
rect 13725 21468 13737 21471
rect 13688 21440 13737 21468
rect 13688 21428 13694 21440
rect 13725 21437 13737 21440
rect 13771 21468 13783 21471
rect 19536 21468 19564 21635
rect 21082 21632 21088 21644
rect 21140 21632 21146 21684
rect 21634 21672 21640 21684
rect 21595 21644 21640 21672
rect 21634 21632 21640 21644
rect 21692 21632 21698 21684
rect 22741 21675 22799 21681
rect 22741 21641 22753 21675
rect 22787 21672 22799 21675
rect 23290 21672 23296 21684
rect 22787 21644 23296 21672
rect 22787 21641 22799 21644
rect 22741 21635 22799 21641
rect 23290 21632 23296 21644
rect 23348 21672 23354 21684
rect 23385 21675 23443 21681
rect 23385 21672 23397 21675
rect 23348 21644 23397 21672
rect 23348 21632 23354 21644
rect 23385 21641 23397 21644
rect 23431 21641 23443 21675
rect 25498 21672 25504 21684
rect 25459 21644 25504 21672
rect 23385 21635 23443 21641
rect 25498 21632 25504 21644
rect 25556 21632 25562 21684
rect 25869 21675 25927 21681
rect 25869 21641 25881 21675
rect 25915 21672 25927 21675
rect 25958 21672 25964 21684
rect 25915 21644 25964 21672
rect 25915 21641 25927 21644
rect 25869 21635 25927 21641
rect 25958 21632 25964 21644
rect 26016 21632 26022 21684
rect 26970 21672 26976 21684
rect 26931 21644 26976 21672
rect 26970 21632 26976 21644
rect 27028 21632 27034 21684
rect 27890 21632 27896 21684
rect 27948 21672 27954 21684
rect 27985 21675 28043 21681
rect 27985 21672 27997 21675
rect 27948 21644 27997 21672
rect 27948 21632 27954 21644
rect 27985 21641 27997 21644
rect 28031 21641 28043 21675
rect 27985 21635 28043 21641
rect 28718 21632 28724 21684
rect 28776 21672 28782 21684
rect 31849 21675 31907 21681
rect 31849 21672 31861 21675
rect 28776 21644 31861 21672
rect 28776 21632 28782 21644
rect 31849 21641 31861 21644
rect 31895 21672 31907 21675
rect 31941 21675 31999 21681
rect 31941 21672 31953 21675
rect 31895 21644 31953 21672
rect 31895 21641 31907 21644
rect 31849 21635 31907 21641
rect 31941 21641 31953 21644
rect 31987 21641 31999 21675
rect 33870 21672 33876 21684
rect 31941 21635 31999 21641
rect 33704 21644 33876 21672
rect 21726 21564 21732 21616
rect 21784 21604 21790 21616
rect 27798 21604 27804 21616
rect 21784 21576 24440 21604
rect 27759 21576 27804 21604
rect 21784 21564 21790 21576
rect 20254 21536 20260 21548
rect 20215 21508 20260 21536
rect 20254 21496 20260 21508
rect 20312 21496 20318 21548
rect 22830 21496 22836 21548
rect 22888 21536 22894 21548
rect 24412 21545 24440 21576
rect 27798 21564 27804 21576
rect 27856 21564 27862 21616
rect 29270 21564 29276 21616
rect 29328 21604 29334 21616
rect 29411 21607 29469 21613
rect 29411 21604 29423 21607
rect 29328 21576 29423 21604
rect 29328 21564 29334 21576
rect 29411 21573 29423 21576
rect 29457 21573 29469 21607
rect 29546 21604 29552 21616
rect 29507 21576 29552 21604
rect 29411 21567 29469 21573
rect 29546 21564 29552 21576
rect 29604 21604 29610 21616
rect 31021 21607 31079 21613
rect 31021 21604 31033 21607
rect 29604 21576 31033 21604
rect 29604 21564 29610 21576
rect 31021 21573 31033 21576
rect 31067 21573 31079 21607
rect 31021 21567 31079 21573
rect 24397 21539 24455 21545
rect 22888 21508 23612 21536
rect 22888 21496 22894 21508
rect 19705 21471 19763 21477
rect 19705 21468 19717 21471
rect 13771 21440 13860 21468
rect 19536 21440 19717 21468
rect 13771 21437 13783 21440
rect 13725 21431 13783 21437
rect 12158 21332 12164 21344
rect 6788 21304 7052 21332
rect 12119 21304 12164 21332
rect 6788 21292 6794 21304
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 12250 21292 12256 21344
rect 12308 21332 12314 21344
rect 12575 21335 12633 21341
rect 12575 21332 12587 21335
rect 12308 21304 12587 21332
rect 12308 21292 12314 21304
rect 12575 21301 12587 21304
rect 12621 21301 12633 21335
rect 12575 21295 12633 21301
rect 13078 21292 13084 21344
rect 13136 21332 13142 21344
rect 13265 21335 13323 21341
rect 13265 21332 13277 21335
rect 13136 21304 13277 21332
rect 13136 21292 13142 21304
rect 13265 21301 13277 21304
rect 13311 21301 13323 21335
rect 13832 21332 13860 21440
rect 19705 21437 19717 21440
rect 19751 21437 19763 21471
rect 19705 21431 19763 21437
rect 20070 21428 20076 21480
rect 20128 21468 20134 21480
rect 20165 21471 20223 21477
rect 20165 21468 20177 21471
rect 20128 21440 20177 21468
rect 20128 21428 20134 21440
rect 20165 21437 20177 21440
rect 20211 21437 20223 21471
rect 20165 21431 20223 21437
rect 21361 21471 21419 21477
rect 21361 21437 21373 21471
rect 21407 21468 21419 21471
rect 21726 21468 21732 21480
rect 21407 21440 21732 21468
rect 21407 21437 21419 21440
rect 21361 21431 21419 21437
rect 21726 21428 21732 21440
rect 21784 21468 21790 21480
rect 21821 21471 21879 21477
rect 21821 21468 21833 21471
rect 21784 21440 21833 21468
rect 21784 21428 21790 21440
rect 21821 21437 21833 21440
rect 21867 21437 21879 21471
rect 23474 21468 23480 21480
rect 21821 21431 21879 21437
rect 23032 21440 23480 21468
rect 15746 21400 15752 21412
rect 15707 21372 15752 21400
rect 15746 21360 15752 21372
rect 15804 21360 15810 21412
rect 15841 21403 15899 21409
rect 15841 21369 15853 21403
rect 15887 21369 15899 21403
rect 18230 21400 18236 21412
rect 18191 21372 18236 21400
rect 15841 21363 15899 21369
rect 14277 21335 14335 21341
rect 14277 21332 14289 21335
rect 13832 21304 14289 21332
rect 13265 21295 13323 21301
rect 14277 21301 14289 21304
rect 14323 21301 14335 21335
rect 14826 21332 14832 21344
rect 14787 21304 14832 21332
rect 14277 21295 14335 21301
rect 14826 21292 14832 21304
rect 14884 21292 14890 21344
rect 15562 21332 15568 21344
rect 15523 21304 15568 21332
rect 15562 21292 15568 21304
rect 15620 21332 15626 21344
rect 15856 21332 15884 21363
rect 18230 21360 18236 21372
rect 18288 21360 18294 21412
rect 21634 21360 21640 21412
rect 21692 21400 21698 21412
rect 23032 21409 23060 21440
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 22142 21403 22200 21409
rect 22142 21400 22154 21403
rect 21692 21372 22154 21400
rect 21692 21360 21698 21372
rect 22142 21369 22154 21372
rect 22188 21400 22200 21403
rect 23017 21403 23075 21409
rect 23017 21400 23029 21403
rect 22188 21372 23029 21400
rect 22188 21369 22200 21372
rect 22142 21363 22200 21369
rect 23017 21369 23029 21372
rect 23063 21369 23075 21403
rect 23017 21363 23075 21369
rect 23290 21360 23296 21412
rect 23348 21400 23354 21412
rect 23584 21400 23612 21508
rect 24397 21505 24409 21539
rect 24443 21536 24455 21539
rect 25038 21536 25044 21548
rect 24443 21508 25044 21536
rect 24443 21505 24455 21508
rect 24397 21499 24455 21505
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 25590 21536 25596 21548
rect 25551 21508 25596 21536
rect 25590 21496 25596 21508
rect 25648 21536 25654 21548
rect 26237 21539 26295 21545
rect 26237 21536 26249 21539
rect 25648 21508 26249 21536
rect 25648 21496 25654 21508
rect 26237 21505 26249 21508
rect 26283 21536 26295 21539
rect 26605 21539 26663 21545
rect 26605 21536 26617 21539
rect 26283 21508 26617 21536
rect 26283 21505 26295 21508
rect 26237 21499 26295 21505
rect 26605 21505 26617 21508
rect 26651 21536 26663 21539
rect 27522 21536 27528 21548
rect 26651 21508 27528 21536
rect 26651 21505 26663 21508
rect 26605 21499 26663 21505
rect 27522 21496 27528 21508
rect 27580 21536 27586 21548
rect 27893 21539 27951 21545
rect 27893 21536 27905 21539
rect 27580 21508 27905 21536
rect 27580 21496 27586 21508
rect 27893 21505 27905 21508
rect 27939 21536 27951 21539
rect 28442 21536 28448 21548
rect 27939 21508 28448 21536
rect 27939 21505 27951 21508
rect 27893 21499 27951 21505
rect 28442 21496 28448 21508
rect 28500 21536 28506 21548
rect 29638 21536 29644 21548
rect 28500 21508 29644 21536
rect 28500 21496 28506 21508
rect 29638 21496 29644 21508
rect 29696 21496 29702 21548
rect 30009 21539 30067 21545
rect 30009 21505 30021 21539
rect 30055 21536 30067 21539
rect 33594 21536 33600 21548
rect 30055 21508 33600 21536
rect 30055 21505 30067 21508
rect 30009 21499 30067 21505
rect 33594 21496 33600 21508
rect 33652 21496 33658 21548
rect 33704 21545 33732 21644
rect 33870 21632 33876 21644
rect 33928 21672 33934 21684
rect 34149 21675 34207 21681
rect 34149 21672 34161 21675
rect 33928 21644 34161 21672
rect 33928 21632 33934 21644
rect 34149 21641 34161 21644
rect 34195 21641 34207 21675
rect 43346 21672 43352 21684
rect 43307 21644 43352 21672
rect 34149 21635 34207 21641
rect 43346 21632 43352 21644
rect 43404 21632 43410 21684
rect 37458 21604 37464 21616
rect 37419 21576 37464 21604
rect 37458 21564 37464 21576
rect 37516 21564 37522 21616
rect 43272 21576 44220 21604
rect 43272 21548 43300 21576
rect 33689 21539 33747 21545
rect 33689 21505 33701 21539
rect 33735 21505 33747 21539
rect 35342 21536 35348 21548
rect 35303 21508 35348 21536
rect 33689 21499 33747 21505
rect 35342 21496 35348 21508
rect 35400 21496 35406 21548
rect 35618 21536 35624 21548
rect 35579 21508 35624 21536
rect 35618 21496 35624 21508
rect 35676 21536 35682 21548
rect 36354 21536 36360 21548
rect 35676 21508 36360 21536
rect 35676 21496 35682 21508
rect 36354 21496 36360 21508
rect 36412 21496 36418 21548
rect 36906 21536 36912 21548
rect 36867 21508 36912 21536
rect 36906 21496 36912 21508
rect 36964 21496 36970 21548
rect 39577 21539 39635 21545
rect 39577 21505 39589 21539
rect 39623 21536 39635 21539
rect 40494 21536 40500 21548
rect 39623 21508 40500 21536
rect 39623 21505 39635 21508
rect 39577 21499 39635 21505
rect 40494 21496 40500 21508
rect 40552 21496 40558 21548
rect 42334 21536 42340 21548
rect 42295 21508 42340 21536
rect 42334 21496 42340 21508
rect 42392 21496 42398 21548
rect 42981 21539 43039 21545
rect 42981 21505 42993 21539
rect 43027 21536 43039 21539
rect 43254 21536 43260 21548
rect 43027 21508 43260 21536
rect 43027 21505 43039 21508
rect 42981 21499 43039 21505
rect 43254 21496 43260 21508
rect 43312 21496 43318 21548
rect 43898 21536 43904 21548
rect 43859 21508 43904 21536
rect 43898 21496 43904 21508
rect 43956 21496 43962 21548
rect 44192 21545 44220 21576
rect 44177 21539 44235 21545
rect 44177 21505 44189 21539
rect 44223 21505 44235 21539
rect 44177 21499 44235 21505
rect 25130 21428 25136 21480
rect 25188 21468 25194 21480
rect 25372 21471 25430 21477
rect 25372 21468 25384 21471
rect 25188 21440 25384 21468
rect 25188 21428 25194 21440
rect 25372 21437 25384 21440
rect 25418 21437 25430 21471
rect 25372 21431 25430 21437
rect 27672 21471 27730 21477
rect 27672 21437 27684 21471
rect 27718 21468 27730 21471
rect 27982 21468 27988 21480
rect 27718 21440 27988 21468
rect 27718 21437 27730 21440
rect 27672 21431 27730 21437
rect 27982 21428 27988 21440
rect 28040 21428 28046 21480
rect 28166 21428 28172 21480
rect 28224 21468 28230 21480
rect 30837 21471 30895 21477
rect 30837 21468 30849 21471
rect 28224 21440 30849 21468
rect 28224 21428 28230 21440
rect 30837 21437 30849 21440
rect 30883 21468 30895 21471
rect 31297 21471 31355 21477
rect 31297 21468 31309 21471
rect 30883 21440 31309 21468
rect 30883 21437 30895 21440
rect 30837 21431 30895 21437
rect 31297 21437 31309 21440
rect 31343 21437 31355 21471
rect 31297 21431 31355 21437
rect 31849 21471 31907 21477
rect 31849 21437 31861 21471
rect 31895 21468 31907 21471
rect 32122 21468 32128 21480
rect 31895 21440 32128 21468
rect 31895 21437 31907 21440
rect 31849 21431 31907 21437
rect 32122 21428 32128 21440
rect 32180 21428 32186 21480
rect 32582 21468 32588 21480
rect 32543 21440 32588 21468
rect 32582 21428 32588 21440
rect 32640 21428 32646 21480
rect 37921 21471 37979 21477
rect 37921 21437 37933 21471
rect 37967 21468 37979 21471
rect 38286 21468 38292 21480
rect 37967 21440 38292 21468
rect 37967 21437 37979 21440
rect 37921 21431 37979 21437
rect 38286 21428 38292 21440
rect 38344 21428 38350 21480
rect 38841 21471 38899 21477
rect 38841 21437 38853 21471
rect 38887 21437 38899 21471
rect 38841 21431 38899 21437
rect 23750 21400 23756 21412
rect 23348 21372 23474 21400
rect 23584 21372 23756 21400
rect 23348 21360 23354 21372
rect 15620 21304 15884 21332
rect 23446 21332 23474 21372
rect 23750 21360 23756 21372
rect 23808 21360 23814 21412
rect 23845 21403 23903 21409
rect 23845 21369 23857 21403
rect 23891 21369 23903 21403
rect 23845 21363 23903 21369
rect 23860 21332 23888 21363
rect 24210 21360 24216 21412
rect 24268 21400 24274 21412
rect 24765 21403 24823 21409
rect 24765 21400 24777 21403
rect 24268 21372 24777 21400
rect 24268 21360 24274 21372
rect 24765 21369 24777 21372
rect 24811 21400 24823 21403
rect 25225 21403 25283 21409
rect 25225 21400 25237 21403
rect 24811 21372 25237 21400
rect 24811 21369 24823 21372
rect 24765 21363 24823 21369
rect 25225 21369 25237 21372
rect 25271 21400 25283 21403
rect 26510 21400 26516 21412
rect 25271 21372 26516 21400
rect 25271 21369 25283 21372
rect 25225 21363 25283 21369
rect 26510 21360 26516 21372
rect 26568 21360 26574 21412
rect 27522 21400 27528 21412
rect 27483 21372 27528 21400
rect 27522 21360 27528 21372
rect 27580 21360 27586 21412
rect 29089 21403 29147 21409
rect 29089 21369 29101 21403
rect 29135 21400 29147 21403
rect 29178 21400 29184 21412
rect 29135 21372 29184 21400
rect 29135 21369 29147 21372
rect 29089 21363 29147 21369
rect 29178 21360 29184 21372
rect 29236 21400 29242 21412
rect 29272 21403 29330 21409
rect 29272 21400 29284 21403
rect 29236 21372 29284 21400
rect 29236 21360 29242 21372
rect 29272 21369 29284 21372
rect 29318 21369 29330 21403
rect 29272 21363 29330 21369
rect 30374 21360 30380 21412
rect 30432 21400 30438 21412
rect 30469 21403 30527 21409
rect 30469 21400 30481 21403
rect 30432 21372 30481 21400
rect 30432 21360 30438 21372
rect 30469 21369 30481 21372
rect 30515 21369 30527 21403
rect 32858 21400 32864 21412
rect 32819 21372 32864 21400
rect 30469 21363 30527 21369
rect 32858 21360 32864 21372
rect 32916 21360 32922 21412
rect 33134 21400 33140 21412
rect 33106 21360 33140 21400
rect 33192 21400 33198 21412
rect 33229 21403 33287 21409
rect 33229 21400 33241 21403
rect 33192 21372 33241 21400
rect 33192 21360 33198 21372
rect 33229 21369 33241 21372
rect 33275 21400 33287 21403
rect 35158 21400 35164 21412
rect 33275 21372 35164 21400
rect 33275 21369 33287 21372
rect 33229 21363 33287 21369
rect 35158 21360 35164 21372
rect 35216 21360 35222 21412
rect 35437 21403 35495 21409
rect 35437 21369 35449 21403
rect 35483 21369 35495 21403
rect 35437 21363 35495 21369
rect 37001 21403 37059 21409
rect 37001 21369 37013 21403
rect 37047 21369 37059 21403
rect 37001 21363 37059 21369
rect 25130 21332 25136 21344
rect 23446 21304 23888 21332
rect 25091 21304 25136 21332
rect 15620 21292 15626 21304
rect 25130 21292 25136 21304
rect 25188 21292 25194 21344
rect 27430 21332 27436 21344
rect 27391 21304 27436 21332
rect 27430 21292 27436 21304
rect 27488 21332 27494 21344
rect 27798 21332 27804 21344
rect 27488 21304 27804 21332
rect 27488 21292 27494 21304
rect 27798 21292 27804 21304
rect 27856 21332 27862 21344
rect 28350 21332 28356 21344
rect 27856 21304 28356 21332
rect 27856 21292 27862 21304
rect 28350 21292 28356 21304
rect 28408 21332 28414 21344
rect 28537 21335 28595 21341
rect 28537 21332 28549 21335
rect 28408 21304 28549 21332
rect 28408 21292 28414 21304
rect 28537 21301 28549 21304
rect 28583 21301 28595 21335
rect 28537 21295 28595 21301
rect 31110 21292 31116 21344
rect 31168 21332 31174 21344
rect 31662 21332 31668 21344
rect 31168 21304 31668 21332
rect 31168 21292 31174 21304
rect 31662 21292 31668 21304
rect 31720 21332 31726 21344
rect 33106 21332 33134 21360
rect 34514 21332 34520 21344
rect 31720 21304 33134 21332
rect 34475 21304 34520 21332
rect 31720 21292 31726 21304
rect 34514 21292 34520 21304
rect 34572 21332 34578 21344
rect 35069 21335 35127 21341
rect 35069 21332 35081 21335
rect 34572 21304 35081 21332
rect 34572 21292 34578 21304
rect 35069 21301 35081 21304
rect 35115 21332 35127 21335
rect 35452 21332 35480 21363
rect 36262 21332 36268 21344
rect 35115 21304 36268 21332
rect 35115 21301 35127 21304
rect 35069 21295 35127 21301
rect 36262 21292 36268 21304
rect 36320 21332 36326 21344
rect 36633 21335 36691 21341
rect 36633 21332 36645 21335
rect 36320 21304 36645 21332
rect 36320 21292 36326 21304
rect 36633 21301 36645 21304
rect 36679 21332 36691 21335
rect 37016 21332 37044 21363
rect 37642 21360 37648 21412
rect 37700 21400 37706 21412
rect 38657 21403 38715 21409
rect 38657 21400 38669 21403
rect 37700 21372 38669 21400
rect 37700 21360 37706 21372
rect 38657 21369 38669 21372
rect 38703 21400 38715 21403
rect 38856 21400 38884 21431
rect 39206 21428 39212 21480
rect 39264 21468 39270 21480
rect 39301 21471 39359 21477
rect 39301 21468 39313 21471
rect 39264 21440 39313 21468
rect 39264 21428 39270 21440
rect 39301 21437 39313 21440
rect 39347 21468 39359 21471
rect 39853 21471 39911 21477
rect 39853 21468 39865 21471
rect 39347 21440 39865 21468
rect 39347 21437 39359 21440
rect 39301 21431 39359 21437
rect 39853 21437 39865 21440
rect 39899 21437 39911 21471
rect 39853 21431 39911 21437
rect 40818 21403 40876 21409
rect 40818 21400 40830 21403
rect 38703 21372 38884 21400
rect 40328 21372 40830 21400
rect 38703 21369 38715 21372
rect 38657 21363 38715 21369
rect 40328 21344 40356 21372
rect 40818 21369 40830 21372
rect 40864 21369 40876 21403
rect 40818 21363 40876 21369
rect 42429 21403 42487 21409
rect 42429 21369 42441 21403
rect 42475 21369 42487 21403
rect 43990 21400 43996 21412
rect 43951 21372 43996 21400
rect 42429 21363 42487 21369
rect 36679 21304 37044 21332
rect 36679 21301 36691 21304
rect 36633 21295 36691 21301
rect 38194 21292 38200 21344
rect 38252 21332 38258 21344
rect 38289 21335 38347 21341
rect 38289 21332 38301 21335
rect 38252 21304 38301 21332
rect 38252 21292 38258 21304
rect 38289 21301 38301 21304
rect 38335 21301 38347 21335
rect 40310 21332 40316 21344
rect 40271 21304 40316 21332
rect 38289 21295 38347 21301
rect 40310 21292 40316 21304
rect 40368 21292 40374 21344
rect 41414 21332 41420 21344
rect 41375 21304 41420 21332
rect 41414 21292 41420 21304
rect 41472 21292 41478 21344
rect 41690 21332 41696 21344
rect 41651 21304 41696 21332
rect 41690 21292 41696 21304
rect 41748 21332 41754 21344
rect 42061 21335 42119 21341
rect 42061 21332 42073 21335
rect 41748 21304 42073 21332
rect 41748 21292 41754 21304
rect 42061 21301 42073 21304
rect 42107 21332 42119 21335
rect 42444 21332 42472 21363
rect 43990 21360 43996 21372
rect 44048 21360 44054 21412
rect 44818 21332 44824 21344
rect 42107 21304 42472 21332
rect 44779 21304 44824 21332
rect 42107 21301 42119 21304
rect 42061 21295 42119 21301
rect 44818 21292 44824 21304
rect 44876 21292 44882 21344
rect 1104 21242 48852 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 48852 21242
rect 1104 21168 48852 21190
rect 5166 21128 5172 21140
rect 5127 21100 5172 21128
rect 5166 21088 5172 21100
rect 5224 21088 5230 21140
rect 5951 21131 6009 21137
rect 5951 21097 5963 21131
rect 5997 21128 6009 21131
rect 7006 21128 7012 21140
rect 5997 21100 7012 21128
rect 5997 21097 6009 21100
rect 5951 21091 6009 21097
rect 7006 21088 7012 21100
rect 7064 21128 7070 21140
rect 7285 21131 7343 21137
rect 7285 21128 7297 21131
rect 7064 21100 7297 21128
rect 7064 21088 7070 21100
rect 7285 21097 7297 21100
rect 7331 21097 7343 21131
rect 7285 21091 7343 21097
rect 10597 21131 10655 21137
rect 10597 21097 10609 21131
rect 10643 21128 10655 21131
rect 12158 21128 12164 21140
rect 10643 21100 12164 21128
rect 10643 21097 10655 21100
rect 10597 21091 10655 21097
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 14274 21128 14280 21140
rect 14235 21100 14280 21128
rect 14274 21088 14280 21100
rect 14332 21088 14338 21140
rect 15427 21131 15485 21137
rect 15427 21097 15439 21131
rect 15473 21128 15485 21131
rect 15746 21128 15752 21140
rect 15473 21100 15752 21128
rect 15473 21097 15485 21100
rect 15427 21091 15485 21097
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 16114 21128 16120 21140
rect 16075 21100 16120 21128
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 18506 21128 18512 21140
rect 18467 21100 18512 21128
rect 18506 21088 18512 21100
rect 18564 21088 18570 21140
rect 19797 21131 19855 21137
rect 19797 21097 19809 21131
rect 19843 21128 19855 21131
rect 20070 21128 20076 21140
rect 19843 21100 20076 21128
rect 19843 21097 19855 21100
rect 19797 21091 19855 21097
rect 20070 21088 20076 21100
rect 20128 21088 20134 21140
rect 21726 21128 21732 21140
rect 21687 21100 21732 21128
rect 21726 21088 21732 21100
rect 21784 21088 21790 21140
rect 22922 21128 22928 21140
rect 22883 21100 22928 21128
rect 22922 21088 22928 21100
rect 22980 21088 22986 21140
rect 23750 21128 23756 21140
rect 23711 21100 23756 21128
rect 23750 21088 23756 21100
rect 23808 21088 23814 21140
rect 24397 21131 24455 21137
rect 24397 21097 24409 21131
rect 24443 21128 24455 21131
rect 24762 21128 24768 21140
rect 24443 21100 24768 21128
rect 24443 21097 24455 21100
rect 24397 21091 24455 21097
rect 24762 21088 24768 21100
rect 24820 21128 24826 21140
rect 28215 21131 28273 21137
rect 28215 21128 28227 21131
rect 24820 21100 28227 21128
rect 24820 21088 24826 21100
rect 28215 21097 28227 21100
rect 28261 21097 28273 21131
rect 28215 21091 28273 21097
rect 28810 21088 28816 21140
rect 28868 21128 28874 21140
rect 29733 21131 29791 21137
rect 29733 21128 29745 21131
rect 28868 21100 29745 21128
rect 28868 21088 28874 21100
rect 29733 21097 29745 21100
rect 29779 21097 29791 21131
rect 29733 21091 29791 21097
rect 32401 21131 32459 21137
rect 32401 21097 32413 21131
rect 32447 21128 32459 21131
rect 32582 21128 32588 21140
rect 32447 21100 32588 21128
rect 32447 21097 32459 21100
rect 32401 21091 32459 21097
rect 32582 21088 32588 21100
rect 32640 21088 32646 21140
rect 33321 21131 33379 21137
rect 33321 21128 33333 21131
rect 33106 21100 33333 21128
rect 4801 21063 4859 21069
rect 4801 21029 4813 21063
rect 4847 21060 4859 21063
rect 4982 21060 4988 21072
rect 4847 21032 4988 21060
rect 4847 21029 4859 21032
rect 4801 21023 4859 21029
rect 4982 21020 4988 21032
rect 5040 21020 5046 21072
rect 10039 21063 10097 21069
rect 10039 21029 10051 21063
rect 10085 21060 10097 21063
rect 10778 21060 10784 21072
rect 10085 21032 10784 21060
rect 10085 21029 10097 21032
rect 10039 21023 10097 21029
rect 10778 21020 10784 21032
rect 10836 21020 10842 21072
rect 11606 21060 11612 21072
rect 11567 21032 11612 21060
rect 11606 21020 11612 21032
rect 11664 21020 11670 21072
rect 17310 21060 17316 21072
rect 17271 21032 17316 21060
rect 17310 21020 17316 21032
rect 17368 21020 17374 21072
rect 25593 21063 25651 21069
rect 25593 21029 25605 21063
rect 25639 21060 25651 21063
rect 25866 21060 25872 21072
rect 25639 21032 25872 21060
rect 25639 21029 25651 21032
rect 25593 21023 25651 21029
rect 25866 21020 25872 21032
rect 25924 21020 25930 21072
rect 30101 21063 30159 21069
rect 30101 21060 30113 21063
rect 29104 21032 30113 21060
rect 29104 21004 29132 21032
rect 30101 21029 30113 21032
rect 30147 21029 30159 21063
rect 30101 21023 30159 21029
rect 32490 21020 32496 21072
rect 32548 21060 32554 21072
rect 33106 21060 33134 21100
rect 33321 21097 33333 21100
rect 33367 21097 33379 21131
rect 33321 21091 33379 21097
rect 33873 21131 33931 21137
rect 33873 21097 33885 21131
rect 33919 21128 33931 21131
rect 34514 21128 34520 21140
rect 33919 21100 34520 21128
rect 33919 21097 33931 21100
rect 33873 21091 33931 21097
rect 34514 21088 34520 21100
rect 34572 21088 34578 21140
rect 35115 21131 35173 21137
rect 35115 21097 35127 21131
rect 35161 21128 35173 21131
rect 35342 21128 35348 21140
rect 35161 21100 35348 21128
rect 35161 21097 35173 21100
rect 35115 21091 35173 21097
rect 35342 21088 35348 21100
rect 35400 21088 35406 21140
rect 36906 21088 36912 21140
rect 36964 21128 36970 21140
rect 37001 21131 37059 21137
rect 37001 21128 37013 21131
rect 36964 21100 37013 21128
rect 36964 21088 36970 21100
rect 37001 21097 37013 21100
rect 37047 21097 37059 21131
rect 37001 21091 37059 21097
rect 38703 21131 38761 21137
rect 38703 21097 38715 21131
rect 38749 21128 38761 21131
rect 41141 21131 41199 21137
rect 41141 21128 41153 21131
rect 38749 21100 41153 21128
rect 38749 21097 38761 21100
rect 38703 21091 38761 21097
rect 41141 21097 41153 21100
rect 41187 21128 41199 21131
rect 41322 21128 41328 21140
rect 41187 21100 41328 21128
rect 41187 21097 41199 21100
rect 41141 21091 41199 21097
rect 41322 21088 41328 21100
rect 41380 21088 41386 21140
rect 43990 21128 43996 21140
rect 43548 21100 43996 21128
rect 43548 21072 43576 21100
rect 43990 21088 43996 21100
rect 44048 21088 44054 21140
rect 36170 21060 36176 21072
rect 32548 21032 33134 21060
rect 36131 21032 36176 21060
rect 32548 21020 32554 21032
rect 36170 21020 36176 21032
rect 36228 21020 36234 21072
rect 39117 21063 39175 21069
rect 39117 21029 39129 21063
rect 39163 21060 39175 21063
rect 39206 21060 39212 21072
rect 39163 21032 39212 21060
rect 39163 21029 39175 21032
rect 39117 21023 39175 21029
rect 39206 21020 39212 21032
rect 39264 21020 39270 21072
rect 39939 21063 39997 21069
rect 39939 21029 39951 21063
rect 39985 21060 39997 21063
rect 40310 21060 40316 21072
rect 39985 21032 40316 21060
rect 39985 21029 39997 21032
rect 39939 21023 39997 21029
rect 40310 21020 40316 21032
rect 40368 21020 40374 21072
rect 41046 21020 41052 21072
rect 41104 21060 41110 21072
rect 41509 21063 41567 21069
rect 41509 21060 41521 21063
rect 41104 21032 41521 21060
rect 41104 21020 41110 21032
rect 41509 21029 41521 21032
rect 41555 21060 41567 21063
rect 41690 21060 41696 21072
rect 41555 21032 41696 21060
rect 41555 21029 41567 21032
rect 41509 21023 41567 21029
rect 41690 21020 41696 21032
rect 41748 21020 41754 21072
rect 42058 21060 42064 21072
rect 42019 21032 42064 21060
rect 42058 21020 42064 21032
rect 42116 21020 42122 21072
rect 43530 21060 43536 21072
rect 43443 21032 43536 21060
rect 43530 21020 43536 21032
rect 43588 21020 43594 21072
rect 43806 21020 43812 21072
rect 43864 21060 43870 21072
rect 44085 21063 44143 21069
rect 44085 21060 44097 21063
rect 43864 21032 44097 21060
rect 43864 21020 43870 21032
rect 44085 21029 44097 21032
rect 44131 21029 44143 21063
rect 44085 21023 44143 21029
rect 3878 20952 3884 21004
rect 3936 20992 3942 21004
rect 4065 20995 4123 21001
rect 4065 20992 4077 20995
rect 3936 20964 4077 20992
rect 3936 20952 3942 20964
rect 4065 20961 4077 20964
rect 4111 20961 4123 20995
rect 4614 20992 4620 21004
rect 4575 20964 4620 20992
rect 4065 20955 4123 20961
rect 4614 20952 4620 20964
rect 4672 20952 4678 21004
rect 5534 20952 5540 21004
rect 5592 20992 5598 21004
rect 5848 20995 5906 21001
rect 5848 20992 5860 20995
rect 5592 20964 5860 20992
rect 5592 20952 5598 20964
rect 5848 20961 5860 20964
rect 5894 20961 5906 20995
rect 5848 20955 5906 20961
rect 7098 20952 7104 21004
rect 7156 20992 7162 21004
rect 7742 20992 7748 21004
rect 7156 20964 7748 20992
rect 7156 20952 7162 20964
rect 7742 20952 7748 20964
rect 7800 20952 7806 21004
rect 8202 20992 8208 21004
rect 8163 20964 8208 20992
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 12894 20952 12900 21004
rect 12952 20992 12958 21004
rect 12989 20995 13047 21001
rect 12989 20992 13001 20995
rect 12952 20964 13001 20992
rect 12952 20952 12958 20964
rect 12989 20961 13001 20964
rect 13035 20961 13047 20995
rect 12989 20955 13047 20961
rect 13078 20952 13084 21004
rect 13136 20992 13142 21004
rect 13449 20995 13507 21001
rect 13449 20992 13461 20995
rect 13136 20964 13461 20992
rect 13136 20952 13142 20964
rect 13449 20961 13461 20964
rect 13495 20961 13507 20995
rect 13449 20955 13507 20961
rect 14826 20952 14832 21004
rect 14884 20992 14890 21004
rect 15286 20992 15292 21004
rect 15344 21001 15350 21004
rect 15344 20995 15382 21001
rect 14884 20964 15292 20992
rect 14884 20952 14890 20964
rect 15286 20952 15292 20964
rect 15370 20961 15382 20995
rect 15344 20955 15382 20961
rect 15344 20952 15350 20955
rect 18322 20952 18328 21004
rect 18380 20992 18386 21004
rect 18785 20995 18843 21001
rect 18785 20992 18797 20995
rect 18380 20964 18797 20992
rect 18380 20952 18386 20964
rect 18785 20961 18797 20964
rect 18831 20992 18843 20995
rect 19058 20992 19064 21004
rect 18831 20964 19064 20992
rect 18831 20961 18843 20964
rect 18785 20955 18843 20961
rect 19058 20952 19064 20964
rect 19116 20952 19122 21004
rect 21910 20992 21916 21004
rect 21871 20964 21916 20992
rect 21910 20952 21916 20964
rect 21968 20952 21974 21004
rect 22094 20992 22100 21004
rect 22055 20964 22100 20992
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 23198 20992 23204 21004
rect 23159 20964 23204 20992
rect 23198 20952 23204 20964
rect 23256 20952 23262 21004
rect 24857 20995 24915 21001
rect 24857 20961 24869 20995
rect 24903 20992 24915 20995
rect 25406 20992 25412 21004
rect 24903 20964 25412 20992
rect 24903 20961 24915 20964
rect 24857 20955 24915 20961
rect 25406 20952 25412 20964
rect 25464 20952 25470 21004
rect 26510 20992 26516 21004
rect 26471 20964 26516 20992
rect 26510 20952 26516 20964
rect 26568 20952 26574 21004
rect 27890 20952 27896 21004
rect 27948 20992 27954 21004
rect 28112 20995 28170 21001
rect 28112 20992 28124 20995
rect 27948 20964 28124 20992
rect 27948 20952 27954 20964
rect 28112 20961 28124 20964
rect 28158 20961 28170 20995
rect 29086 20992 29092 21004
rect 29047 20964 29092 20992
rect 28112 20955 28170 20961
rect 29086 20952 29092 20964
rect 29144 20952 29150 21004
rect 30650 20992 30656 21004
rect 30611 20964 30656 20992
rect 30650 20952 30656 20964
rect 30708 20952 30714 21004
rect 32306 20952 32312 21004
rect 32364 20992 32370 21004
rect 32766 20992 32772 21004
rect 32364 20964 32772 20992
rect 32364 20952 32370 20964
rect 32766 20952 32772 20964
rect 32824 20952 32830 21004
rect 32858 20952 32864 21004
rect 32916 20992 32922 21004
rect 32953 20995 33011 21001
rect 32953 20992 32965 20995
rect 32916 20964 32965 20992
rect 32916 20952 32922 20964
rect 32953 20961 32965 20964
rect 32999 20992 33011 20995
rect 33410 20992 33416 21004
rect 32999 20964 33416 20992
rect 32999 20961 33011 20964
rect 32953 20955 33011 20961
rect 33410 20952 33416 20964
rect 33468 20952 33474 21004
rect 35044 20995 35102 21001
rect 35044 20961 35056 20995
rect 35090 20992 35102 20995
rect 35250 20992 35256 21004
rect 35090 20964 35256 20992
rect 35090 20961 35102 20964
rect 35044 20955 35102 20961
rect 35250 20952 35256 20964
rect 35308 20952 35314 21004
rect 39482 20952 39488 21004
rect 39540 20992 39546 21004
rect 39577 20995 39635 21001
rect 39577 20992 39589 20995
rect 39540 20964 39589 20992
rect 39540 20952 39546 20964
rect 39577 20961 39589 20964
rect 39623 20961 39635 20995
rect 39577 20955 39635 20961
rect 44964 20995 45022 21001
rect 44964 20961 44976 20995
rect 45010 20992 45022 20995
rect 45462 20992 45468 21004
rect 45010 20964 45468 20992
rect 45010 20961 45022 20964
rect 44964 20955 45022 20961
rect 45462 20952 45468 20964
rect 45520 20952 45526 21004
rect 8481 20927 8539 20933
rect 8481 20893 8493 20927
rect 8527 20924 8539 20927
rect 9677 20927 9735 20933
rect 9677 20924 9689 20927
rect 8527 20896 9689 20924
rect 8527 20893 8539 20896
rect 8481 20887 8539 20893
rect 9677 20893 9689 20896
rect 9723 20924 9735 20927
rect 10502 20924 10508 20936
rect 9723 20896 10508 20924
rect 9723 20893 9735 20896
rect 9677 20887 9735 20893
rect 10502 20884 10508 20896
rect 10560 20884 10566 20936
rect 11517 20927 11575 20933
rect 11517 20893 11529 20927
rect 11563 20924 11575 20927
rect 12250 20924 12256 20936
rect 11563 20896 12256 20924
rect 11563 20893 11575 20896
rect 11517 20887 11575 20893
rect 12250 20884 12256 20896
rect 12308 20884 12314 20936
rect 13538 20924 13544 20936
rect 13499 20896 13544 20924
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 16942 20884 16948 20936
rect 17000 20924 17006 20936
rect 17221 20927 17279 20933
rect 17221 20924 17233 20927
rect 17000 20896 17233 20924
rect 17000 20884 17006 20896
rect 17221 20893 17233 20896
rect 17267 20893 17279 20927
rect 17221 20887 17279 20893
rect 17865 20927 17923 20933
rect 17865 20893 17877 20927
rect 17911 20924 17923 20927
rect 18966 20924 18972 20936
rect 17911 20896 18972 20924
rect 17911 20893 17923 20896
rect 17865 20887 17923 20893
rect 18966 20884 18972 20896
rect 19024 20884 19030 20936
rect 25004 20927 25062 20933
rect 25004 20893 25016 20927
rect 25050 20924 25062 20927
rect 25130 20924 25136 20936
rect 25050 20896 25136 20924
rect 25050 20893 25062 20896
rect 25004 20887 25062 20893
rect 25130 20884 25136 20896
rect 25188 20884 25194 20936
rect 25225 20927 25283 20933
rect 25225 20893 25237 20927
rect 25271 20924 25283 20927
rect 25590 20924 25596 20936
rect 25271 20896 25596 20924
rect 25271 20893 25283 20896
rect 25225 20887 25283 20893
rect 12066 20856 12072 20868
rect 12027 20828 12072 20856
rect 12066 20816 12072 20828
rect 12124 20816 12130 20868
rect 14553 20859 14611 20865
rect 14553 20856 14565 20859
rect 13786 20828 14565 20856
rect 7006 20788 7012 20800
rect 6967 20760 7012 20788
rect 7006 20748 7012 20760
rect 7064 20748 7070 20800
rect 13354 20748 13360 20800
rect 13412 20788 13418 20800
rect 13786 20788 13814 20828
rect 14553 20825 14565 20828
rect 14599 20825 14611 20859
rect 14553 20819 14611 20825
rect 17954 20816 17960 20868
rect 18012 20856 18018 20868
rect 20625 20859 20683 20865
rect 20625 20856 20637 20859
rect 18012 20828 20637 20856
rect 18012 20816 18018 20828
rect 20625 20825 20637 20828
rect 20671 20856 20683 20859
rect 20990 20856 20996 20868
rect 20671 20828 20996 20856
rect 20671 20825 20683 20828
rect 20625 20819 20683 20825
rect 20990 20816 20996 20828
rect 21048 20816 21054 20868
rect 22094 20816 22100 20868
rect 22152 20856 22158 20868
rect 23385 20859 23443 20865
rect 23385 20856 23397 20859
rect 22152 20828 23397 20856
rect 22152 20816 22158 20828
rect 23385 20825 23397 20828
rect 23431 20825 23443 20859
rect 23385 20819 23443 20825
rect 24302 20816 24308 20868
rect 24360 20856 24366 20868
rect 25240 20856 25268 20887
rect 25590 20884 25596 20896
rect 25648 20884 25654 20936
rect 26881 20927 26939 20933
rect 26881 20924 26893 20927
rect 25884 20896 26893 20924
rect 24360 20828 25268 20856
rect 24360 20816 24366 20828
rect 25884 20800 25912 20896
rect 26881 20893 26893 20896
rect 26927 20924 26939 20927
rect 28810 20924 28816 20936
rect 26927 20896 28816 20924
rect 26927 20893 26939 20896
rect 26881 20887 26939 20893
rect 28810 20884 28816 20896
rect 28868 20924 28874 20936
rect 28905 20927 28963 20933
rect 28905 20924 28917 20927
rect 28868 20896 28917 20924
rect 28868 20884 28874 20896
rect 28905 20893 28917 20896
rect 28951 20924 28963 20927
rect 29457 20927 29515 20933
rect 29457 20924 29469 20927
rect 28951 20896 29469 20924
rect 28951 20893 28963 20896
rect 28905 20887 28963 20893
rect 29457 20893 29469 20896
rect 29503 20893 29515 20927
rect 29457 20887 29515 20893
rect 26329 20859 26387 20865
rect 26329 20825 26341 20859
rect 26375 20856 26387 20859
rect 26973 20859 27031 20865
rect 26973 20856 26985 20859
rect 26375 20828 26985 20856
rect 26375 20825 26387 20828
rect 26329 20819 26387 20825
rect 26973 20825 26985 20828
rect 27019 20856 27031 20859
rect 27062 20856 27068 20868
rect 27019 20828 27068 20856
rect 27019 20825 27031 20828
rect 26973 20819 27031 20825
rect 27062 20816 27068 20828
rect 27120 20816 27126 20868
rect 28994 20816 29000 20868
rect 29052 20856 29058 20868
rect 29270 20865 29276 20868
rect 29236 20859 29276 20865
rect 29236 20856 29248 20859
rect 29052 20828 29248 20856
rect 29052 20816 29058 20828
rect 29236 20825 29248 20828
rect 29236 20819 29276 20825
rect 29270 20816 29276 20819
rect 29328 20816 29334 20868
rect 29472 20856 29500 20887
rect 29546 20884 29552 20936
rect 29604 20924 29610 20936
rect 30469 20927 30527 20933
rect 30469 20924 30481 20927
rect 29604 20896 30481 20924
rect 29604 20884 29610 20896
rect 30469 20893 30481 20896
rect 30515 20893 30527 20927
rect 30469 20887 30527 20893
rect 30558 20884 30564 20936
rect 30616 20924 30622 20936
rect 36078 20924 36084 20936
rect 30616 20896 32489 20924
rect 36039 20896 36084 20924
rect 30616 20884 30622 20896
rect 30837 20859 30895 20865
rect 30837 20856 30849 20859
rect 29472 20828 30849 20856
rect 30837 20825 30849 20828
rect 30883 20856 30895 20859
rect 31018 20856 31024 20868
rect 30883 20828 31024 20856
rect 30883 20825 30895 20828
rect 30837 20819 30895 20825
rect 31018 20816 31024 20828
rect 31076 20856 31082 20868
rect 31113 20859 31171 20865
rect 31113 20856 31125 20859
rect 31076 20828 31125 20856
rect 31076 20816 31082 20828
rect 31113 20825 31125 20828
rect 31159 20825 31171 20859
rect 32461 20856 32489 20896
rect 36078 20884 36084 20896
rect 36136 20884 36142 20936
rect 36354 20924 36360 20936
rect 36315 20896 36360 20924
rect 36354 20884 36360 20896
rect 36412 20884 36418 20936
rect 38194 20924 38200 20936
rect 36556 20896 38200 20924
rect 32766 20856 32772 20868
rect 32461 20828 32772 20856
rect 31113 20819 31171 20825
rect 32766 20816 32772 20828
rect 32824 20856 32830 20868
rect 36556 20856 36584 20896
rect 38194 20884 38200 20896
rect 38252 20884 38258 20936
rect 40770 20884 40776 20936
rect 40828 20924 40834 20936
rect 41417 20927 41475 20933
rect 41417 20924 41429 20927
rect 40828 20896 41429 20924
rect 40828 20884 40834 20896
rect 41417 20893 41429 20896
rect 41463 20893 41475 20927
rect 41417 20887 41475 20893
rect 42610 20884 42616 20936
rect 42668 20924 42674 20936
rect 43441 20927 43499 20933
rect 43441 20924 43453 20927
rect 42668 20896 43453 20924
rect 42668 20884 42674 20896
rect 43441 20893 43453 20896
rect 43487 20924 43499 20927
rect 45051 20927 45109 20933
rect 45051 20924 45063 20927
rect 43487 20896 45063 20924
rect 43487 20893 43499 20896
rect 43441 20887 43499 20893
rect 45051 20893 45063 20896
rect 45097 20893 45109 20927
rect 45051 20887 45109 20893
rect 38470 20856 38476 20868
rect 32824 20828 36584 20856
rect 38431 20828 38476 20856
rect 32824 20816 32830 20828
rect 38470 20816 38476 20828
rect 38528 20816 38534 20868
rect 18230 20788 18236 20800
rect 13412 20760 13814 20788
rect 18191 20760 18236 20788
rect 13412 20748 13418 20760
rect 18230 20748 18236 20760
rect 18288 20788 18294 20800
rect 18969 20791 19027 20797
rect 18969 20788 18981 20791
rect 18288 20760 18981 20788
rect 18288 20748 18294 20760
rect 18969 20757 18981 20760
rect 19015 20757 19027 20791
rect 21266 20788 21272 20800
rect 21227 20760 21272 20788
rect 18969 20751 19027 20757
rect 21266 20748 21272 20760
rect 21324 20748 21330 20800
rect 24765 20791 24823 20797
rect 24765 20757 24777 20791
rect 24811 20788 24823 20791
rect 25133 20791 25191 20797
rect 25133 20788 25145 20791
rect 24811 20760 25145 20788
rect 24811 20757 24823 20760
rect 24765 20751 24823 20757
rect 25133 20757 25145 20760
rect 25179 20788 25191 20791
rect 25498 20788 25504 20800
rect 25179 20760 25504 20788
rect 25179 20757 25191 20760
rect 25133 20751 25191 20757
rect 25498 20748 25504 20760
rect 25556 20748 25562 20800
rect 25866 20788 25872 20800
rect 25827 20760 25872 20788
rect 25866 20748 25872 20760
rect 25924 20748 25930 20800
rect 26602 20748 26608 20800
rect 26660 20797 26666 20800
rect 26660 20791 26709 20797
rect 26660 20757 26663 20791
rect 26697 20757 26709 20791
rect 26786 20788 26792 20800
rect 26747 20760 26792 20788
rect 26660 20751 26709 20757
rect 26660 20748 26666 20751
rect 26786 20748 26792 20760
rect 26844 20748 26850 20800
rect 27614 20788 27620 20800
rect 27575 20760 27620 20788
rect 27614 20748 27620 20760
rect 27672 20748 27678 20800
rect 27982 20788 27988 20800
rect 27943 20760 27988 20788
rect 27982 20748 27988 20760
rect 28040 20748 28046 20800
rect 28629 20791 28687 20797
rect 28629 20757 28641 20791
rect 28675 20788 28687 20791
rect 29086 20788 29092 20800
rect 28675 20760 29092 20788
rect 28675 20757 28687 20760
rect 28629 20751 28687 20757
rect 29086 20748 29092 20760
rect 29144 20748 29150 20800
rect 29362 20788 29368 20800
rect 29323 20760 29368 20788
rect 29362 20748 29368 20760
rect 29420 20748 29426 20800
rect 31573 20791 31631 20797
rect 31573 20757 31585 20791
rect 31619 20788 31631 20791
rect 31938 20788 31944 20800
rect 31619 20760 31944 20788
rect 31619 20757 31631 20760
rect 31573 20751 31631 20757
rect 31938 20748 31944 20760
rect 31996 20748 32002 20800
rect 32122 20748 32128 20800
rect 32180 20788 32186 20800
rect 39298 20788 39304 20800
rect 32180 20760 39304 20788
rect 32180 20748 32186 20760
rect 39298 20748 39304 20760
rect 39356 20748 39362 20800
rect 40497 20791 40555 20797
rect 40497 20757 40509 20791
rect 40543 20788 40555 20791
rect 41046 20788 41052 20800
rect 40543 20760 41052 20788
rect 40543 20757 40555 20760
rect 40497 20751 40555 20757
rect 41046 20748 41052 20760
rect 41104 20748 41110 20800
rect 1104 20698 48852 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 48852 20698
rect 1104 20624 48852 20646
rect 3789 20587 3847 20593
rect 3789 20553 3801 20587
rect 3835 20584 3847 20587
rect 3878 20584 3884 20596
rect 3835 20556 3884 20584
rect 3835 20553 3847 20556
rect 3789 20547 3847 20553
rect 3878 20544 3884 20556
rect 3936 20544 3942 20596
rect 4157 20587 4215 20593
rect 4157 20553 4169 20587
rect 4203 20584 4215 20587
rect 4706 20584 4712 20596
rect 4203 20556 4712 20584
rect 4203 20553 4215 20556
rect 4157 20547 4215 20553
rect 4706 20544 4712 20556
rect 4764 20544 4770 20596
rect 5534 20544 5540 20596
rect 5592 20584 5598 20596
rect 5813 20587 5871 20593
rect 5813 20584 5825 20587
rect 5592 20556 5825 20584
rect 5592 20544 5598 20556
rect 5813 20553 5825 20556
rect 5859 20553 5871 20587
rect 7650 20584 7656 20596
rect 7611 20556 7656 20584
rect 5813 20547 5871 20553
rect 7650 20544 7656 20556
rect 7708 20544 7714 20596
rect 10870 20544 10876 20596
rect 10928 20584 10934 20596
rect 11195 20587 11253 20593
rect 11195 20584 11207 20587
rect 10928 20556 11207 20584
rect 10928 20544 10934 20556
rect 11195 20553 11207 20556
rect 11241 20553 11253 20587
rect 11195 20547 11253 20553
rect 11977 20587 12035 20593
rect 11977 20553 11989 20587
rect 12023 20584 12035 20587
rect 12250 20584 12256 20596
rect 12023 20556 12256 20584
rect 12023 20553 12035 20556
rect 11977 20547 12035 20553
rect 12250 20544 12256 20556
rect 12308 20544 12314 20596
rect 12894 20544 12900 20596
rect 12952 20584 12958 20596
rect 13265 20587 13323 20593
rect 13265 20584 13277 20587
rect 12952 20556 13277 20584
rect 12952 20544 12958 20556
rect 13265 20553 13277 20556
rect 13311 20553 13323 20587
rect 13630 20584 13636 20596
rect 13591 20556 13636 20584
rect 13265 20547 13323 20553
rect 13630 20544 13636 20556
rect 13688 20544 13694 20596
rect 15286 20584 15292 20596
rect 15247 20556 15292 20584
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 19058 20584 19064 20596
rect 19019 20556 19064 20584
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 21085 20587 21143 20593
rect 21085 20553 21097 20587
rect 21131 20584 21143 20587
rect 22094 20584 22100 20596
rect 21131 20556 22100 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 22094 20544 22100 20556
rect 22152 20544 22158 20596
rect 23109 20587 23167 20593
rect 23109 20553 23121 20587
rect 23155 20584 23167 20587
rect 23198 20584 23204 20596
rect 23155 20556 23204 20584
rect 23155 20553 23167 20556
rect 23109 20547 23167 20553
rect 23198 20544 23204 20556
rect 23256 20584 23262 20596
rect 25961 20587 26019 20593
rect 25961 20584 25973 20587
rect 23256 20556 25973 20584
rect 23256 20544 23262 20556
rect 25961 20553 25973 20556
rect 26007 20553 26019 20587
rect 25961 20547 26019 20553
rect 26510 20544 26516 20596
rect 26568 20584 26574 20596
rect 26881 20587 26939 20593
rect 26881 20584 26893 20587
rect 26568 20556 26893 20584
rect 26568 20544 26574 20556
rect 26881 20553 26893 20556
rect 26927 20553 26939 20587
rect 26881 20547 26939 20553
rect 27154 20544 27160 20596
rect 27212 20584 27218 20596
rect 27249 20587 27307 20593
rect 27249 20584 27261 20587
rect 27212 20556 27261 20584
rect 27212 20544 27218 20556
rect 27249 20553 27261 20556
rect 27295 20553 27307 20587
rect 27249 20547 27307 20553
rect 29178 20544 29184 20596
rect 29236 20584 29242 20596
rect 30285 20587 30343 20593
rect 30285 20584 30297 20587
rect 29236 20556 30297 20584
rect 29236 20544 29242 20556
rect 30285 20553 30297 20556
rect 30331 20584 30343 20587
rect 30469 20587 30527 20593
rect 30469 20584 30481 20587
rect 30331 20556 30481 20584
rect 30331 20553 30343 20556
rect 30285 20547 30343 20553
rect 30469 20553 30481 20556
rect 30515 20553 30527 20587
rect 30650 20584 30656 20596
rect 30611 20556 30656 20584
rect 30469 20547 30527 20553
rect 30650 20544 30656 20556
rect 30708 20544 30714 20596
rect 30742 20544 30748 20596
rect 30800 20584 30806 20596
rect 30975 20587 31033 20593
rect 30975 20584 30987 20587
rect 30800 20556 30987 20584
rect 30800 20544 30806 20556
rect 30975 20553 30987 20556
rect 31021 20553 31033 20587
rect 31478 20584 31484 20596
rect 31439 20556 31484 20584
rect 30975 20547 31033 20553
rect 31478 20544 31484 20556
rect 31536 20544 31542 20596
rect 31938 20584 31944 20596
rect 31899 20556 31944 20584
rect 31938 20544 31944 20556
rect 31996 20544 32002 20596
rect 35621 20587 35679 20593
rect 35621 20553 35633 20587
rect 35667 20584 35679 20587
rect 35851 20587 35909 20593
rect 35851 20584 35863 20587
rect 35667 20556 35863 20584
rect 35667 20553 35679 20556
rect 35621 20547 35679 20553
rect 35851 20553 35863 20556
rect 35897 20584 35909 20587
rect 36078 20584 36084 20596
rect 35897 20556 36084 20584
rect 35897 20553 35909 20556
rect 35851 20547 35909 20553
rect 36078 20544 36084 20556
rect 36136 20544 36142 20596
rect 36170 20544 36176 20596
rect 36228 20584 36234 20596
rect 36541 20587 36599 20593
rect 36541 20584 36553 20587
rect 36228 20556 36553 20584
rect 36228 20544 36234 20556
rect 36541 20553 36553 20556
rect 36587 20584 36599 20587
rect 37918 20584 37924 20596
rect 36587 20556 37924 20584
rect 36587 20553 36599 20556
rect 36541 20547 36599 20553
rect 37918 20544 37924 20556
rect 37976 20544 37982 20596
rect 38102 20584 38108 20596
rect 38063 20556 38108 20584
rect 38102 20544 38108 20556
rect 38160 20544 38166 20596
rect 39301 20587 39359 20593
rect 39301 20553 39313 20587
rect 39347 20584 39359 20587
rect 39482 20584 39488 20596
rect 39347 20556 39488 20584
rect 39347 20553 39359 20556
rect 39301 20547 39359 20553
rect 39482 20544 39488 20556
rect 39540 20544 39546 20596
rect 40770 20584 40776 20596
rect 40731 20556 40776 20584
rect 40770 20544 40776 20556
rect 40828 20544 40834 20596
rect 41046 20584 41052 20596
rect 41007 20556 41052 20584
rect 41046 20544 41052 20556
rect 41104 20544 41110 20596
rect 42610 20584 42616 20596
rect 42571 20556 42616 20584
rect 42610 20544 42616 20556
rect 42668 20544 42674 20596
rect 42981 20587 43039 20593
rect 42981 20553 42993 20587
rect 43027 20584 43039 20587
rect 43349 20587 43407 20593
rect 43349 20584 43361 20587
rect 43027 20556 43361 20584
rect 43027 20553 43039 20556
rect 42981 20547 43039 20553
rect 43349 20553 43361 20556
rect 43395 20584 43407 20587
rect 43530 20584 43536 20596
rect 43395 20556 43536 20584
rect 43395 20553 43407 20556
rect 43349 20547 43407 20553
rect 43530 20544 43536 20556
rect 43588 20544 43594 20596
rect 2593 20519 2651 20525
rect 2593 20485 2605 20519
rect 2639 20516 2651 20519
rect 3234 20516 3240 20528
rect 2639 20488 3240 20516
rect 2639 20485 2651 20488
rect 2593 20479 2651 20485
rect 2700 20389 2728 20488
rect 3234 20476 3240 20488
rect 3292 20476 3298 20528
rect 21910 20476 21916 20528
rect 21968 20516 21974 20528
rect 22189 20519 22247 20525
rect 22189 20516 22201 20519
rect 21968 20488 22201 20516
rect 21968 20476 21974 20488
rect 22189 20485 22201 20488
rect 22235 20485 22247 20519
rect 22189 20479 22247 20485
rect 25777 20519 25835 20525
rect 25777 20485 25789 20519
rect 25823 20516 25835 20519
rect 26786 20516 26792 20528
rect 25823 20488 26792 20516
rect 25823 20485 25835 20488
rect 25777 20479 25835 20485
rect 26786 20476 26792 20488
rect 26844 20516 26850 20528
rect 26844 20488 29132 20516
rect 26844 20476 26850 20488
rect 3970 20448 3976 20460
rect 3252 20420 3976 20448
rect 2685 20383 2743 20389
rect 2685 20349 2697 20383
rect 2731 20349 2743 20383
rect 2685 20343 2743 20349
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 3252 20389 3280 20420
rect 3970 20408 3976 20420
rect 4028 20448 4034 20460
rect 4614 20448 4620 20460
rect 4028 20420 4620 20448
rect 4028 20408 4034 20420
rect 4614 20408 4620 20420
rect 4672 20448 4678 20460
rect 4672 20420 5580 20448
rect 4672 20408 4678 20420
rect 3237 20383 3295 20389
rect 3237 20380 3249 20383
rect 2832 20352 3249 20380
rect 2832 20340 2838 20352
rect 3237 20349 3249 20352
rect 3283 20349 3295 20383
rect 3237 20343 3295 20349
rect 3421 20383 3479 20389
rect 3421 20349 3433 20383
rect 3467 20380 3479 20383
rect 3786 20380 3792 20392
rect 3467 20352 3792 20380
rect 3467 20349 3479 20352
rect 3421 20343 3479 20349
rect 3786 20340 3792 20352
rect 3844 20380 3850 20392
rect 4249 20383 4307 20389
rect 4249 20380 4261 20383
rect 3844 20352 4261 20380
rect 3844 20340 3850 20352
rect 4249 20349 4261 20352
rect 4295 20349 4307 20383
rect 4249 20343 4307 20349
rect 4611 20315 4669 20321
rect 4611 20281 4623 20315
rect 4657 20312 4669 20315
rect 4706 20312 4712 20324
rect 4657 20284 4712 20312
rect 4657 20281 4669 20284
rect 4611 20275 4669 20281
rect 4706 20272 4712 20284
rect 4764 20272 4770 20324
rect 5552 20321 5580 20420
rect 6730 20408 6736 20460
rect 6788 20448 6794 20460
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 6788 20420 11529 20448
rect 6788 20408 6794 20420
rect 11517 20417 11529 20420
rect 11563 20448 11575 20451
rect 11606 20448 11612 20460
rect 11563 20420 11612 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 11606 20408 11612 20420
rect 11664 20408 11670 20460
rect 12066 20408 12072 20460
rect 12124 20448 12130 20460
rect 18138 20448 18144 20460
rect 12124 20420 18144 20448
rect 12124 20408 12130 20420
rect 18138 20408 18144 20420
rect 18196 20408 18202 20460
rect 18598 20408 18604 20460
rect 18656 20448 18662 20460
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 18656 20420 19717 20448
rect 18656 20408 18662 20420
rect 19705 20417 19717 20420
rect 19751 20448 19763 20451
rect 20070 20448 20076 20460
rect 19751 20420 20076 20448
rect 19751 20417 19763 20420
rect 19705 20411 19763 20417
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 24210 20448 24216 20460
rect 24171 20420 24216 20448
rect 24210 20408 24216 20420
rect 24268 20408 24274 20460
rect 25866 20448 25872 20460
rect 25827 20420 25872 20448
rect 25866 20408 25872 20420
rect 25924 20448 25930 20460
rect 27525 20451 27583 20457
rect 27525 20448 27537 20451
rect 25924 20420 27537 20448
rect 25924 20408 25930 20420
rect 27525 20417 27537 20420
rect 27571 20417 27583 20451
rect 27525 20411 27583 20417
rect 7650 20340 7656 20392
rect 7708 20380 7714 20392
rect 7745 20383 7803 20389
rect 7745 20380 7757 20383
rect 7708 20352 7757 20380
rect 7708 20340 7714 20352
rect 7745 20349 7757 20352
rect 7791 20349 7803 20383
rect 8202 20380 8208 20392
rect 8115 20352 8208 20380
rect 7745 20343 7803 20349
rect 8202 20340 8208 20352
rect 8260 20380 8266 20392
rect 8481 20383 8539 20389
rect 8260 20352 8432 20380
rect 8260 20340 8266 20352
rect 5537 20315 5595 20321
rect 5537 20281 5549 20315
rect 5583 20312 5595 20315
rect 5718 20312 5724 20324
rect 5583 20284 5724 20312
rect 5583 20281 5595 20284
rect 5537 20275 5595 20281
rect 5718 20272 5724 20284
rect 5776 20312 5782 20324
rect 8294 20312 8300 20324
rect 5776 20284 8300 20312
rect 5776 20272 5782 20284
rect 8294 20272 8300 20284
rect 8352 20272 8358 20324
rect 5166 20244 5172 20256
rect 5127 20216 5172 20244
rect 5166 20204 5172 20216
rect 5224 20204 5230 20256
rect 7285 20247 7343 20253
rect 7285 20213 7297 20247
rect 7331 20244 7343 20247
rect 8404 20244 8432 20352
rect 8481 20349 8493 20383
rect 8527 20380 8539 20383
rect 9306 20380 9312 20392
rect 8527 20352 9312 20380
rect 8527 20349 8539 20352
rect 8481 20343 8539 20349
rect 9306 20340 9312 20352
rect 9364 20340 9370 20392
rect 10229 20383 10287 20389
rect 10229 20349 10241 20383
rect 10275 20380 10287 20383
rect 10873 20383 10931 20389
rect 10873 20380 10885 20383
rect 10275 20352 10885 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 10873 20349 10885 20352
rect 10919 20380 10931 20383
rect 11092 20383 11150 20389
rect 11092 20380 11104 20383
rect 10919 20352 11104 20380
rect 10919 20349 10931 20352
rect 10873 20343 10931 20349
rect 11092 20349 11104 20352
rect 11138 20349 11150 20383
rect 12805 20383 12863 20389
rect 12805 20380 12817 20383
rect 11092 20343 11150 20349
rect 12728 20352 12817 20380
rect 9217 20315 9275 20321
rect 9217 20281 9229 20315
rect 9263 20312 9275 20315
rect 9671 20315 9729 20321
rect 9671 20312 9683 20315
rect 9263 20284 9683 20312
rect 9263 20281 9275 20284
rect 9217 20275 9275 20281
rect 9671 20281 9683 20284
rect 9717 20312 9729 20315
rect 9717 20284 10640 20312
rect 9717 20281 9729 20284
rect 9671 20275 9729 20281
rect 8846 20244 8852 20256
rect 7331 20216 8852 20244
rect 7331 20213 7343 20216
rect 7285 20207 7343 20213
rect 8846 20204 8852 20216
rect 8904 20204 8910 20256
rect 10612 20253 10640 20284
rect 12728 20256 12756 20352
rect 12805 20349 12817 20352
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 13354 20340 13360 20392
rect 13412 20380 13418 20392
rect 13817 20383 13875 20389
rect 13817 20380 13829 20383
rect 13412 20352 13829 20380
rect 13412 20340 13418 20352
rect 13817 20349 13829 20352
rect 13863 20349 13875 20383
rect 13817 20343 13875 20349
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20380 14795 20383
rect 15600 20383 15658 20389
rect 15600 20380 15612 20383
rect 14783 20352 15612 20380
rect 14783 20349 14795 20352
rect 14737 20343 14795 20349
rect 15600 20349 15612 20352
rect 15646 20380 15658 20383
rect 16025 20383 16083 20389
rect 16025 20380 16037 20383
rect 15646 20352 16037 20380
rect 15646 20349 15658 20352
rect 15600 20343 15658 20349
rect 16025 20349 16037 20352
rect 16071 20349 16083 20383
rect 16612 20383 16670 20389
rect 16612 20380 16624 20383
rect 16025 20343 16083 20349
rect 16408 20352 16624 20380
rect 13630 20272 13636 20324
rect 13688 20312 13694 20324
rect 13688 20284 13814 20312
rect 13688 20272 13694 20284
rect 10597 20247 10655 20253
rect 10597 20213 10609 20247
rect 10643 20244 10655 20247
rect 10778 20244 10784 20256
rect 10643 20216 10784 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 10778 20204 10784 20216
rect 10836 20204 10842 20256
rect 12710 20244 12716 20256
rect 12671 20216 12716 20244
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 12986 20244 12992 20256
rect 12947 20216 12992 20244
rect 12986 20204 12992 20216
rect 13044 20204 13050 20256
rect 13786 20244 13814 20284
rect 16408 20256 16436 20352
rect 16612 20349 16624 20352
rect 16658 20349 16670 20383
rect 21266 20380 21272 20392
rect 21227 20352 21272 20380
rect 16612 20343 16670 20349
rect 21266 20340 21272 20352
rect 21324 20340 21330 20392
rect 23014 20340 23020 20392
rect 23072 20380 23078 20392
rect 23385 20383 23443 20389
rect 23385 20380 23397 20383
rect 23072 20352 23397 20380
rect 23072 20340 23078 20352
rect 23385 20349 23397 20352
rect 23431 20380 23443 20383
rect 23845 20383 23903 20389
rect 23845 20380 23857 20383
rect 23431 20352 23857 20380
rect 23431 20349 23443 20352
rect 23385 20343 23443 20349
rect 23845 20349 23857 20352
rect 23891 20349 23903 20383
rect 25648 20383 25706 20389
rect 25648 20380 25660 20383
rect 23845 20343 23903 20349
rect 25332 20352 25660 20380
rect 18230 20312 18236 20324
rect 17788 20284 18236 20312
rect 14185 20247 14243 20253
rect 14185 20244 14197 20247
rect 13786 20216 14197 20244
rect 14185 20213 14197 20216
rect 14231 20213 14243 20247
rect 14185 20207 14243 20213
rect 15470 20204 15476 20256
rect 15528 20244 15534 20256
rect 15703 20247 15761 20253
rect 15703 20244 15715 20247
rect 15528 20216 15715 20244
rect 15528 20204 15534 20216
rect 15703 20213 15715 20216
rect 15749 20213 15761 20247
rect 16390 20244 16396 20256
rect 16351 20216 16396 20244
rect 15703 20207 15761 20213
rect 16390 20204 16396 20216
rect 16448 20204 16454 20256
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 16715 20247 16773 20253
rect 16715 20244 16727 20247
rect 16632 20216 16727 20244
rect 16632 20204 16638 20216
rect 16715 20213 16727 20216
rect 16761 20213 16773 20247
rect 16715 20207 16773 20213
rect 17221 20247 17279 20253
rect 17221 20213 17233 20247
rect 17267 20244 17279 20247
rect 17310 20244 17316 20256
rect 17267 20216 17316 20244
rect 17267 20213 17279 20216
rect 17221 20207 17279 20213
rect 17310 20204 17316 20216
rect 17368 20244 17374 20256
rect 17788 20253 17816 20284
rect 18230 20272 18236 20284
rect 18288 20272 18294 20324
rect 18782 20312 18788 20324
rect 18743 20284 18788 20312
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 19797 20315 19855 20321
rect 19797 20281 19809 20315
rect 19843 20281 19855 20315
rect 20346 20312 20352 20324
rect 20307 20284 20352 20312
rect 19797 20275 19855 20281
rect 17773 20247 17831 20253
rect 17773 20244 17785 20247
rect 17368 20216 17785 20244
rect 17368 20204 17374 20216
rect 17773 20213 17785 20216
rect 17819 20213 17831 20247
rect 17773 20207 17831 20213
rect 19426 20204 19432 20256
rect 19484 20244 19490 20256
rect 19521 20247 19579 20253
rect 19521 20244 19533 20247
rect 19484 20216 19533 20244
rect 19484 20204 19490 20216
rect 19521 20213 19533 20216
rect 19567 20244 19579 20247
rect 19812 20244 19840 20275
rect 20346 20272 20352 20284
rect 20404 20272 20410 20324
rect 21177 20315 21235 20321
rect 21177 20312 21189 20315
rect 20456 20284 21189 20312
rect 20456 20244 20484 20284
rect 21177 20281 21189 20284
rect 21223 20281 21235 20315
rect 21177 20275 21235 20281
rect 23661 20315 23719 20321
rect 23661 20281 23673 20315
rect 23707 20312 23719 20315
rect 24489 20315 24547 20321
rect 24489 20312 24501 20315
rect 23707 20284 24501 20312
rect 23707 20281 23719 20284
rect 23661 20275 23719 20281
rect 24489 20281 24501 20284
rect 24535 20281 24547 20315
rect 24489 20275 24547 20281
rect 19567 20216 20484 20244
rect 19567 20213 19579 20216
rect 19521 20207 19579 20213
rect 22646 20204 22652 20256
rect 22704 20244 22710 20256
rect 23676 20244 23704 20275
rect 22704 20216 23704 20244
rect 24949 20247 25007 20253
rect 22704 20204 22710 20216
rect 24949 20213 24961 20247
rect 24995 20244 25007 20247
rect 25130 20244 25136 20256
rect 24995 20216 25136 20244
rect 24995 20213 25007 20216
rect 24949 20207 25007 20213
rect 25130 20204 25136 20216
rect 25188 20244 25194 20256
rect 25332 20253 25360 20352
rect 25648 20349 25660 20352
rect 25694 20380 25706 20383
rect 26513 20383 26571 20389
rect 26513 20380 26525 20383
rect 25694 20352 26525 20380
rect 25694 20349 25706 20352
rect 25648 20343 25706 20349
rect 26513 20349 26525 20352
rect 26559 20380 26571 20383
rect 26602 20380 26608 20392
rect 26559 20352 26608 20380
rect 26559 20349 26571 20352
rect 26513 20343 26571 20349
rect 26602 20340 26608 20352
rect 26660 20340 26666 20392
rect 27062 20380 27068 20392
rect 27023 20352 27068 20380
rect 27062 20340 27068 20352
rect 27120 20340 27126 20392
rect 28169 20383 28227 20389
rect 28169 20349 28181 20383
rect 28215 20380 28227 20383
rect 28718 20380 28724 20392
rect 28215 20352 28724 20380
rect 28215 20349 28227 20352
rect 28169 20343 28227 20349
rect 28718 20340 28724 20352
rect 28776 20340 28782 20392
rect 29104 20380 29132 20488
rect 29270 20476 29276 20528
rect 29328 20516 29334 20528
rect 29411 20519 29469 20525
rect 29411 20516 29423 20519
rect 29328 20488 29423 20516
rect 29328 20476 29334 20488
rect 29411 20485 29423 20488
rect 29457 20485 29469 20519
rect 29411 20479 29469 20485
rect 29546 20476 29552 20528
rect 29604 20516 29610 20528
rect 31110 20516 31116 20528
rect 29604 20488 31116 20516
rect 29604 20476 29610 20488
rect 31110 20476 31116 20488
rect 31168 20476 31174 20528
rect 31294 20476 31300 20528
rect 31352 20516 31358 20528
rect 33778 20516 33784 20528
rect 31352 20488 33784 20516
rect 31352 20476 31358 20488
rect 33778 20476 33784 20488
rect 33836 20476 33842 20528
rect 37645 20519 37703 20525
rect 37645 20485 37657 20519
rect 37691 20516 37703 20519
rect 39022 20516 39028 20528
rect 37691 20488 39028 20516
rect 37691 20485 37703 20488
rect 37645 20479 37703 20485
rect 39022 20476 39028 20488
rect 39080 20476 39086 20528
rect 29564 20380 29592 20476
rect 29638 20408 29644 20460
rect 29696 20448 29702 20460
rect 33137 20451 33195 20457
rect 29696 20420 30144 20448
rect 29696 20408 29702 20420
rect 29104 20352 29592 20380
rect 25406 20272 25412 20324
rect 25464 20312 25470 20324
rect 25501 20315 25559 20321
rect 25501 20312 25513 20315
rect 25464 20284 25513 20312
rect 25464 20272 25470 20284
rect 25501 20281 25513 20284
rect 25547 20281 25559 20315
rect 28997 20315 29055 20321
rect 28997 20312 29009 20315
rect 25501 20275 25559 20281
rect 28368 20284 29009 20312
rect 25317 20247 25375 20253
rect 25317 20244 25329 20247
rect 25188 20216 25329 20244
rect 25188 20204 25194 20216
rect 25317 20213 25329 20216
rect 25363 20213 25375 20247
rect 25317 20207 25375 20213
rect 26326 20204 26332 20256
rect 26384 20244 26390 20256
rect 27890 20244 27896 20256
rect 26384 20216 27896 20244
rect 26384 20204 26390 20216
rect 27890 20204 27896 20216
rect 27948 20244 27954 20256
rect 27985 20247 28043 20253
rect 27985 20244 27997 20247
rect 27948 20216 27997 20244
rect 27948 20204 27954 20216
rect 27985 20213 27997 20216
rect 28031 20213 28043 20247
rect 27985 20207 28043 20213
rect 28258 20204 28264 20256
rect 28316 20244 28322 20256
rect 28368 20253 28396 20284
rect 28997 20281 29009 20284
rect 29043 20281 29055 20315
rect 28997 20275 29055 20281
rect 29086 20272 29092 20324
rect 29144 20312 29150 20324
rect 29273 20315 29331 20321
rect 29273 20312 29285 20315
rect 29144 20284 29285 20312
rect 29144 20272 29150 20284
rect 29273 20281 29285 20284
rect 29319 20281 29331 20315
rect 29564 20312 29592 20352
rect 29638 20312 29644 20324
rect 29564 20284 29644 20312
rect 29273 20275 29331 20281
rect 29638 20272 29644 20284
rect 29696 20272 29702 20324
rect 30006 20312 30012 20324
rect 29967 20284 30012 20312
rect 30006 20272 30012 20284
rect 30064 20272 30070 20324
rect 28353 20247 28411 20253
rect 28353 20244 28365 20247
rect 28316 20216 28365 20244
rect 28316 20204 28322 20216
rect 28353 20213 28365 20216
rect 28399 20213 28411 20247
rect 28718 20244 28724 20256
rect 28679 20216 28724 20244
rect 28353 20207 28411 20213
rect 28718 20204 28724 20216
rect 28776 20204 28782 20256
rect 30116 20244 30144 20420
rect 33137 20417 33149 20451
rect 33183 20448 33195 20451
rect 34146 20448 34152 20460
rect 33183 20420 34152 20448
rect 33183 20417 33195 20420
rect 33137 20411 33195 20417
rect 34146 20408 34152 20420
rect 34204 20408 34210 20460
rect 38470 20448 38476 20460
rect 36188 20420 38476 20448
rect 30469 20383 30527 20389
rect 30469 20349 30481 20383
rect 30515 20380 30527 20383
rect 30837 20383 30895 20389
rect 30837 20380 30849 20383
rect 30515 20352 30849 20380
rect 30515 20349 30527 20352
rect 30469 20343 30527 20349
rect 30837 20349 30849 20352
rect 30883 20349 30895 20383
rect 30837 20343 30895 20349
rect 31018 20340 31024 20392
rect 31076 20380 31082 20392
rect 31176 20383 31234 20389
rect 31176 20380 31188 20383
rect 31076 20352 31188 20380
rect 31076 20340 31082 20352
rect 31176 20349 31188 20352
rect 31222 20349 31234 20383
rect 31176 20343 31234 20349
rect 31665 20383 31723 20389
rect 31665 20349 31677 20383
rect 31711 20380 31723 20383
rect 32217 20383 32275 20389
rect 32217 20380 32229 20383
rect 31711 20352 32229 20380
rect 31711 20349 31723 20352
rect 31665 20343 31723 20349
rect 32217 20349 32229 20352
rect 32263 20349 32275 20383
rect 32217 20343 32275 20349
rect 35780 20383 35838 20389
rect 35780 20349 35792 20383
rect 35826 20380 35838 20383
rect 35894 20380 35900 20392
rect 35826 20352 35900 20380
rect 35826 20349 35838 20352
rect 35780 20343 35838 20349
rect 35894 20340 35900 20352
rect 35952 20380 35958 20392
rect 36078 20380 36084 20392
rect 35952 20352 36084 20380
rect 35952 20340 35958 20352
rect 36078 20340 36084 20352
rect 36136 20380 36142 20392
rect 36188 20389 36216 20420
rect 38470 20408 38476 20420
rect 38528 20448 38534 20460
rect 38565 20451 38623 20457
rect 38565 20448 38577 20451
rect 38528 20420 38577 20448
rect 38528 20408 38534 20420
rect 38565 20417 38577 20420
rect 38611 20417 38623 20451
rect 38565 20411 38623 20417
rect 39531 20451 39589 20457
rect 39531 20417 39543 20451
rect 39577 20448 39589 20451
rect 40788 20448 40816 20544
rect 42058 20476 42064 20528
rect 42116 20516 42122 20528
rect 42794 20516 42800 20528
rect 42116 20488 42800 20516
rect 42116 20476 42122 20488
rect 42794 20476 42800 20488
rect 42852 20516 42858 20528
rect 44085 20519 44143 20525
rect 44085 20516 44097 20519
rect 42852 20488 44097 20516
rect 42852 20476 42858 20488
rect 44085 20485 44097 20488
rect 44131 20485 44143 20519
rect 44085 20479 44143 20485
rect 39577 20420 40816 20448
rect 43533 20451 43591 20457
rect 39577 20417 39589 20420
rect 39531 20411 39589 20417
rect 43533 20417 43545 20451
rect 43579 20448 43591 20451
rect 44450 20448 44456 20460
rect 43579 20420 44456 20448
rect 43579 20417 43591 20420
rect 43533 20411 43591 20417
rect 44450 20408 44456 20420
rect 44508 20408 44514 20460
rect 45462 20448 45468 20460
rect 45423 20420 45468 20448
rect 45462 20408 45468 20420
rect 45520 20408 45526 20460
rect 36998 20389 37004 20392
rect 36173 20383 36231 20389
rect 36173 20380 36185 20383
rect 36136 20352 36185 20380
rect 36136 20340 36142 20352
rect 36173 20349 36185 20352
rect 36219 20349 36231 20383
rect 36976 20383 37004 20389
rect 36976 20380 36988 20383
rect 36911 20352 36988 20380
rect 36173 20343 36231 20349
rect 36976 20349 36988 20352
rect 37056 20380 37062 20392
rect 37369 20383 37427 20389
rect 37369 20380 37381 20383
rect 37056 20352 37381 20380
rect 36976 20343 37004 20349
rect 36998 20340 37004 20343
rect 37056 20340 37062 20352
rect 37369 20349 37381 20352
rect 37415 20380 37427 20383
rect 37645 20383 37703 20389
rect 37645 20380 37657 20383
rect 37415 20352 37657 20380
rect 37415 20349 37427 20352
rect 37369 20343 37427 20349
rect 37645 20349 37657 20352
rect 37691 20349 37703 20383
rect 37645 20343 37703 20349
rect 37921 20383 37979 20389
rect 37921 20349 37933 20383
rect 37967 20349 37979 20383
rect 37921 20343 37979 20349
rect 39444 20383 39502 20389
rect 39444 20349 39456 20383
rect 39490 20380 39502 20383
rect 39490 20349 39503 20380
rect 39444 20343 39503 20349
rect 33229 20315 33287 20321
rect 33229 20281 33241 20315
rect 33275 20281 33287 20315
rect 33778 20312 33784 20324
rect 33739 20284 33784 20312
rect 33229 20275 33287 20281
rect 31665 20247 31723 20253
rect 31665 20244 31677 20247
rect 30116 20216 31677 20244
rect 31665 20213 31677 20216
rect 31711 20213 31723 20247
rect 31665 20207 31723 20213
rect 32490 20204 32496 20256
rect 32548 20244 32554 20256
rect 32861 20247 32919 20253
rect 32861 20244 32873 20247
rect 32548 20216 32873 20244
rect 32548 20204 32554 20216
rect 32861 20213 32873 20216
rect 32907 20213 32919 20247
rect 32861 20207 32919 20213
rect 32950 20204 32956 20256
rect 33008 20244 33014 20256
rect 33244 20244 33272 20275
rect 33778 20272 33784 20284
rect 33836 20272 33842 20324
rect 34057 20247 34115 20253
rect 34057 20244 34069 20247
rect 33008 20216 34069 20244
rect 33008 20204 33014 20216
rect 34057 20213 34069 20216
rect 34103 20213 34115 20247
rect 35158 20244 35164 20256
rect 35119 20216 35164 20244
rect 34057 20207 34115 20213
rect 35158 20204 35164 20216
rect 35216 20204 35222 20256
rect 37047 20247 37105 20253
rect 37047 20213 37059 20247
rect 37093 20244 37105 20247
rect 37274 20244 37280 20256
rect 37093 20216 37280 20244
rect 37093 20213 37105 20216
rect 37047 20207 37105 20213
rect 37274 20204 37280 20216
rect 37332 20204 37338 20256
rect 37734 20244 37740 20256
rect 37695 20216 37740 20244
rect 37734 20204 37740 20216
rect 37792 20244 37798 20256
rect 37936 20244 37964 20343
rect 38470 20272 38476 20324
rect 38528 20312 38534 20324
rect 39475 20312 39503 20343
rect 40221 20315 40279 20321
rect 40221 20312 40233 20315
rect 38528 20284 40233 20312
rect 38528 20272 38534 20284
rect 40221 20281 40233 20284
rect 40267 20281 40279 20315
rect 40221 20275 40279 20281
rect 40954 20272 40960 20324
rect 41012 20312 41018 20324
rect 41325 20315 41383 20321
rect 41325 20312 41337 20315
rect 41012 20284 41337 20312
rect 41012 20272 41018 20284
rect 41325 20281 41337 20284
rect 41371 20281 41383 20315
rect 41325 20275 41383 20281
rect 41414 20272 41420 20324
rect 41472 20312 41478 20324
rect 41966 20312 41972 20324
rect 41472 20284 41517 20312
rect 41927 20284 41972 20312
rect 41472 20272 41478 20284
rect 41966 20272 41972 20284
rect 42024 20272 42030 20324
rect 43530 20272 43536 20324
rect 43588 20312 43594 20324
rect 43625 20315 43683 20321
rect 43625 20312 43637 20315
rect 43588 20284 43637 20312
rect 43588 20272 43594 20284
rect 43625 20281 43637 20284
rect 43671 20281 43683 20315
rect 43625 20275 43683 20281
rect 37792 20216 37964 20244
rect 39945 20247 40003 20253
rect 37792 20204 37798 20216
rect 39945 20213 39957 20247
rect 39991 20244 40003 20247
rect 40310 20244 40316 20256
rect 39991 20216 40316 20244
rect 39991 20213 40003 20216
rect 39945 20207 40003 20213
rect 40310 20204 40316 20216
rect 40368 20204 40374 20256
rect 45002 20244 45008 20256
rect 44963 20216 45008 20244
rect 45002 20204 45008 20216
rect 45060 20204 45066 20256
rect 1104 20154 48852 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 48852 20154
rect 1104 20080 48852 20102
rect 2774 20040 2780 20052
rect 2735 20012 2780 20040
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 3786 20040 3792 20052
rect 3747 20012 3792 20040
rect 3786 20000 3792 20012
rect 3844 20000 3850 20052
rect 4706 20040 4712 20052
rect 4667 20012 4712 20040
rect 4706 20000 4712 20012
rect 4764 20000 4770 20052
rect 7742 20040 7748 20052
rect 7703 20012 7748 20040
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 8294 20040 8300 20052
rect 8255 20012 8300 20040
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 9306 20040 9312 20052
rect 9267 20012 9312 20040
rect 9306 20000 9312 20012
rect 9364 20000 9370 20052
rect 10502 20040 10508 20052
rect 10463 20012 10508 20040
rect 10502 20000 10508 20012
rect 10560 20000 10566 20052
rect 13262 20000 13268 20052
rect 13320 20040 13326 20052
rect 13630 20040 13636 20052
rect 13320 20012 13636 20040
rect 13320 20000 13326 20012
rect 13630 20000 13636 20012
rect 13688 20040 13694 20052
rect 13817 20043 13875 20049
rect 13817 20040 13829 20043
rect 13688 20012 13829 20040
rect 13688 20000 13694 20012
rect 13817 20009 13829 20012
rect 13863 20009 13875 20043
rect 13817 20003 13875 20009
rect 14369 20043 14427 20049
rect 14369 20009 14381 20043
rect 14415 20040 14427 20043
rect 16390 20040 16396 20052
rect 14415 20012 16396 20040
rect 14415 20009 14427 20012
rect 14369 20003 14427 20009
rect 16390 20000 16396 20012
rect 16448 20000 16454 20052
rect 16942 20040 16948 20052
rect 16903 20012 16948 20040
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 18138 20040 18144 20052
rect 18099 20012 18144 20040
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 20070 20040 20076 20052
rect 20031 20012 20076 20040
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 26329 20043 26387 20049
rect 26329 20009 26341 20043
rect 26375 20040 26387 20043
rect 26786 20040 26792 20052
rect 26375 20012 26792 20040
rect 26375 20009 26387 20012
rect 26329 20003 26387 20009
rect 26786 20000 26792 20012
rect 26844 20040 26850 20052
rect 27157 20043 27215 20049
rect 27157 20040 27169 20043
rect 26844 20012 27169 20040
rect 26844 20000 26850 20012
rect 27157 20009 27169 20012
rect 27203 20009 27215 20043
rect 27157 20003 27215 20009
rect 27522 20000 27528 20052
rect 27580 20040 27586 20052
rect 27617 20043 27675 20049
rect 27617 20040 27629 20043
rect 27580 20012 27629 20040
rect 27580 20000 27586 20012
rect 27617 20009 27629 20012
rect 27663 20040 27675 20043
rect 28074 20040 28080 20052
rect 27663 20012 28080 20040
rect 27663 20009 27675 20012
rect 27617 20003 27675 20009
rect 28074 20000 28080 20012
rect 28132 20000 28138 20052
rect 28810 20040 28816 20052
rect 28771 20012 28816 20040
rect 28810 20000 28816 20012
rect 28868 20000 28874 20052
rect 28994 20000 29000 20052
rect 29052 20040 29058 20052
rect 30742 20040 30748 20052
rect 29052 20012 30748 20040
rect 29052 20000 29058 20012
rect 6730 19972 6736 19984
rect 6691 19944 6736 19972
rect 6730 19932 6736 19944
rect 6788 19932 6794 19984
rect 10318 19932 10324 19984
rect 10376 19972 10382 19984
rect 12621 19975 12679 19981
rect 10376 19944 11928 19972
rect 10376 19932 10382 19944
rect 11900 19916 11928 19944
rect 12621 19941 12633 19975
rect 12667 19972 12679 19975
rect 13354 19972 13360 19984
rect 12667 19944 13360 19972
rect 12667 19941 12679 19944
rect 12621 19935 12679 19941
rect 13354 19932 13360 19944
rect 13412 19932 13418 19984
rect 15470 19972 15476 19984
rect 15431 19944 15476 19972
rect 15470 19932 15476 19944
rect 15528 19932 15534 19984
rect 15562 19932 15568 19984
rect 15620 19972 15626 19984
rect 17313 19975 17371 19981
rect 15620 19944 15665 19972
rect 15620 19932 15626 19944
rect 17313 19941 17325 19975
rect 17359 19972 17371 19975
rect 18046 19972 18052 19984
rect 17359 19944 18052 19972
rect 17359 19941 17371 19944
rect 17313 19935 17371 19941
rect 18046 19932 18052 19944
rect 18104 19972 18110 19984
rect 18877 19975 18935 19981
rect 18877 19972 18889 19975
rect 18104 19944 18889 19972
rect 18104 19932 18110 19944
rect 18877 19941 18889 19944
rect 18923 19941 18935 19975
rect 18877 19935 18935 19941
rect 25498 19932 25504 19984
rect 25556 19972 25562 19984
rect 25593 19975 25651 19981
rect 25593 19972 25605 19975
rect 25556 19944 25605 19972
rect 25556 19932 25562 19944
rect 25593 19941 25605 19944
rect 25639 19941 25651 19975
rect 27430 19972 27436 19984
rect 25593 19935 25651 19941
rect 26620 19944 27436 19972
rect 3028 19907 3086 19913
rect 3028 19873 3040 19907
rect 3074 19904 3086 19907
rect 3786 19904 3792 19916
rect 3074 19876 3792 19904
rect 3074 19873 3086 19876
rect 3028 19867 3086 19873
rect 3786 19864 3792 19876
rect 3844 19864 3850 19916
rect 7926 19864 7932 19916
rect 7984 19904 7990 19916
rect 8113 19907 8171 19913
rect 8113 19904 8125 19907
rect 7984 19876 8125 19904
rect 7984 19864 7990 19876
rect 8113 19873 8125 19876
rect 8159 19904 8171 19907
rect 8846 19904 8852 19916
rect 8159 19876 8852 19904
rect 8159 19873 8171 19876
rect 8113 19867 8171 19873
rect 8846 19864 8852 19876
rect 8904 19864 8910 19916
rect 9122 19864 9128 19916
rect 9180 19904 9186 19916
rect 9674 19904 9680 19916
rect 9180 19876 9680 19904
rect 9180 19864 9186 19876
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 10940 19907 10998 19913
rect 10940 19873 10952 19907
rect 10986 19904 10998 19907
rect 11054 19904 11060 19916
rect 10986 19876 11060 19904
rect 10986 19873 10998 19876
rect 10940 19867 10998 19873
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 11882 19904 11888 19916
rect 11795 19876 11888 19904
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 12342 19904 12348 19916
rect 12303 19876 12348 19904
rect 12342 19864 12348 19876
rect 12400 19904 12406 19916
rect 12986 19904 12992 19916
rect 12400 19876 12992 19904
rect 12400 19864 12406 19876
rect 12986 19864 12992 19876
rect 13044 19864 13050 19916
rect 13449 19907 13507 19913
rect 13449 19873 13461 19907
rect 13495 19904 13507 19907
rect 13538 19904 13544 19916
rect 13495 19876 13544 19904
rect 13495 19873 13507 19876
rect 13449 19867 13507 19873
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 20990 19904 20996 19916
rect 20951 19876 20996 19904
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 22741 19907 22799 19913
rect 22741 19904 22753 19907
rect 22664 19876 22753 19904
rect 22664 19848 22692 19876
rect 22741 19873 22753 19876
rect 22787 19873 22799 19907
rect 22741 19867 22799 19873
rect 23198 19864 23204 19916
rect 23256 19904 23262 19916
rect 23293 19907 23351 19913
rect 23293 19904 23305 19907
rect 23256 19876 23305 19904
rect 23256 19864 23262 19876
rect 23293 19873 23305 19876
rect 23339 19873 23351 19907
rect 25314 19904 25320 19916
rect 25275 19876 25320 19904
rect 23293 19867 23351 19873
rect 25314 19864 25320 19876
rect 25372 19904 25378 19916
rect 26620 19904 26648 19944
rect 27430 19932 27436 19944
rect 27488 19972 27494 19984
rect 28258 19972 28264 19984
rect 27488 19944 28264 19972
rect 27488 19932 27494 19944
rect 28258 19932 28264 19944
rect 28316 19932 28322 19984
rect 29178 19932 29184 19984
rect 29236 19972 29242 19984
rect 29273 19975 29331 19981
rect 29273 19972 29285 19975
rect 29236 19944 29285 19972
rect 29236 19932 29242 19944
rect 29273 19941 29285 19944
rect 29319 19941 29331 19975
rect 29273 19935 29331 19941
rect 29435 19916 29463 20012
rect 30742 20000 30748 20012
rect 30800 20040 30806 20052
rect 31570 20040 31576 20052
rect 30800 20012 31576 20040
rect 30800 20000 30806 20012
rect 31570 20000 31576 20012
rect 31628 20040 31634 20052
rect 31757 20043 31815 20049
rect 31757 20040 31769 20043
rect 31628 20012 31769 20040
rect 31628 20000 31634 20012
rect 31757 20009 31769 20012
rect 31803 20040 31815 20043
rect 31938 20040 31944 20052
rect 31803 20012 31944 20040
rect 31803 20009 31815 20012
rect 31757 20003 31815 20009
rect 31938 20000 31944 20012
rect 31996 20000 32002 20052
rect 32490 20000 32496 20052
rect 32548 20040 32554 20052
rect 32585 20043 32643 20049
rect 32585 20040 32597 20043
rect 32548 20012 32597 20040
rect 32548 20000 32554 20012
rect 32585 20009 32597 20012
rect 32631 20009 32643 20043
rect 33410 20040 33416 20052
rect 33371 20012 33416 20040
rect 32585 20003 32643 20009
rect 33410 20000 33416 20012
rect 33468 20000 33474 20052
rect 33873 20043 33931 20049
rect 33873 20009 33885 20043
rect 33919 20040 33931 20043
rect 34054 20040 34060 20052
rect 33919 20012 34060 20040
rect 33919 20009 33931 20012
rect 33873 20003 33931 20009
rect 34054 20000 34060 20012
rect 34112 20000 34118 20052
rect 40954 20040 40960 20052
rect 40915 20012 40960 20040
rect 40954 20000 40960 20012
rect 41012 20000 41018 20052
rect 41325 20043 41383 20049
rect 41325 20009 41337 20043
rect 41371 20040 41383 20043
rect 41414 20040 41420 20052
rect 41371 20012 41420 20040
rect 41371 20009 41383 20012
rect 41325 20003 41383 20009
rect 41414 20000 41420 20012
rect 41472 20000 41478 20052
rect 43714 20040 43720 20052
rect 43548 20012 43720 20040
rect 31110 19932 31116 19984
rect 31168 19972 31174 19984
rect 31389 19975 31447 19981
rect 31389 19972 31401 19975
rect 31168 19944 31401 19972
rect 31168 19932 31174 19944
rect 31389 19941 31401 19944
rect 31435 19941 31447 19975
rect 33594 19972 33600 19984
rect 31389 19935 31447 19941
rect 33152 19944 33600 19972
rect 25372 19876 26648 19904
rect 26697 19907 26755 19913
rect 25372 19864 25378 19876
rect 26697 19873 26709 19907
rect 26743 19904 26755 19907
rect 27246 19904 27252 19916
rect 26743 19876 27252 19904
rect 26743 19873 26755 19876
rect 26697 19867 26755 19873
rect 27246 19864 27252 19876
rect 27304 19864 27310 19916
rect 27985 19907 28043 19913
rect 27985 19873 27997 19907
rect 28031 19873 28043 19907
rect 27985 19867 28043 19873
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19836 4399 19839
rect 4614 19836 4620 19848
rect 4387 19808 4620 19836
rect 4387 19805 4399 19808
rect 4341 19799 4399 19805
rect 4614 19796 4620 19808
rect 4672 19836 4678 19848
rect 5534 19836 5540 19848
rect 4672 19808 5540 19836
rect 4672 19796 4678 19808
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 6641 19839 6699 19845
rect 6641 19805 6653 19839
rect 6687 19805 6699 19839
rect 6641 19799 6699 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19836 7343 19839
rect 7558 19836 7564 19848
rect 7331 19808 7564 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 3099 19771 3157 19777
rect 3099 19737 3111 19771
rect 3145 19768 3157 19771
rect 6546 19768 6552 19780
rect 3145 19740 6552 19768
rect 3145 19737 3157 19740
rect 3099 19731 3157 19737
rect 6546 19728 6552 19740
rect 6604 19768 6610 19780
rect 6656 19768 6684 19799
rect 7558 19796 7564 19808
rect 7616 19796 7622 19848
rect 16114 19836 16120 19848
rect 16075 19808 16120 19836
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 16942 19796 16948 19848
rect 17000 19836 17006 19848
rect 17221 19839 17279 19845
rect 17221 19836 17233 19839
rect 17000 19808 17233 19836
rect 17000 19796 17006 19808
rect 17221 19805 17233 19808
rect 17267 19805 17279 19839
rect 18598 19836 18604 19848
rect 17221 19799 17279 19805
rect 17512 19808 18604 19836
rect 6604 19740 6684 19768
rect 9861 19771 9919 19777
rect 6604 19728 6610 19740
rect 9861 19737 9873 19771
rect 9907 19768 9919 19771
rect 10226 19768 10232 19780
rect 9907 19740 10232 19768
rect 9907 19737 9919 19740
rect 9861 19731 9919 19737
rect 10226 19728 10232 19740
rect 10284 19728 10290 19780
rect 16132 19768 16160 19796
rect 17512 19768 17540 19808
rect 18598 19796 18604 19808
rect 18656 19836 18662 19848
rect 18785 19839 18843 19845
rect 18785 19836 18797 19839
rect 18656 19808 18797 19836
rect 18656 19796 18662 19808
rect 18785 19805 18797 19808
rect 18831 19805 18843 19839
rect 18785 19799 18843 19805
rect 18966 19796 18972 19848
rect 19024 19836 19030 19848
rect 19061 19839 19119 19845
rect 19061 19836 19073 19839
rect 19024 19808 19073 19836
rect 19024 19796 19030 19808
rect 19061 19805 19073 19808
rect 19107 19805 19119 19839
rect 19061 19799 19119 19805
rect 22646 19796 22652 19848
rect 22704 19796 22710 19848
rect 23109 19839 23167 19845
rect 23109 19805 23121 19839
rect 23155 19836 23167 19839
rect 28000 19836 28028 19867
rect 28074 19864 28080 19916
rect 28132 19904 28138 19916
rect 28353 19907 28411 19913
rect 28132 19876 28177 19904
rect 28132 19864 28138 19876
rect 28353 19873 28365 19907
rect 28399 19904 28411 19907
rect 28534 19904 28540 19916
rect 28399 19876 28540 19904
rect 28399 19873 28411 19876
rect 28353 19867 28411 19873
rect 28534 19864 28540 19876
rect 28592 19864 28598 19916
rect 29435 19913 29460 19916
rect 29420 19907 29460 19913
rect 29420 19904 29432 19907
rect 29367 19876 29432 19904
rect 29420 19873 29432 19876
rect 29420 19867 29460 19873
rect 29454 19864 29460 19867
rect 29512 19864 29518 19916
rect 30904 19907 30962 19913
rect 30904 19873 30916 19907
rect 30950 19904 30962 19907
rect 31018 19904 31024 19916
rect 30950 19876 31024 19904
rect 30950 19873 30962 19876
rect 30904 19867 30962 19873
rect 31018 19864 31024 19876
rect 31076 19904 31082 19916
rect 31294 19904 31300 19916
rect 31076 19876 31300 19904
rect 31076 19864 31082 19876
rect 31294 19864 31300 19876
rect 31352 19864 31358 19916
rect 33152 19913 33180 19944
rect 33594 19932 33600 19944
rect 33652 19972 33658 19984
rect 34149 19975 34207 19981
rect 34149 19972 34161 19975
rect 33652 19944 34161 19972
rect 33652 19932 33658 19944
rect 34149 19941 34161 19944
rect 34195 19941 34207 19975
rect 36262 19972 36268 19984
rect 36223 19944 36268 19972
rect 34149 19935 34207 19941
rect 36262 19932 36268 19944
rect 36320 19932 36326 19984
rect 37274 19932 37280 19984
rect 37332 19972 37338 19984
rect 37826 19972 37832 19984
rect 37332 19944 37832 19972
rect 37332 19932 37338 19944
rect 37826 19932 37832 19944
rect 37884 19932 37890 19984
rect 37918 19932 37924 19984
rect 37976 19972 37982 19984
rect 37976 19944 38021 19972
rect 37976 19932 37982 19944
rect 39206 19932 39212 19984
rect 39264 19972 39270 19984
rect 41782 19972 41788 19984
rect 39264 19944 39804 19972
rect 41743 19944 41788 19972
rect 39264 19932 39270 19944
rect 33137 19907 33195 19913
rect 33137 19873 33149 19907
rect 33183 19873 33195 19907
rect 39298 19904 39304 19916
rect 39259 19876 39304 19904
rect 33137 19867 33195 19873
rect 39298 19864 39304 19876
rect 39356 19864 39362 19916
rect 39776 19913 39804 19944
rect 41782 19932 41788 19944
rect 41840 19932 41846 19984
rect 43548 19981 43576 20012
rect 43714 20000 43720 20012
rect 43772 20040 43778 20052
rect 45002 20040 45008 20052
rect 43772 20012 45008 20040
rect 43772 20000 43778 20012
rect 45002 20000 45008 20012
rect 45060 20000 45066 20052
rect 43533 19975 43591 19981
rect 43533 19941 43545 19975
rect 43579 19941 43591 19975
rect 43533 19935 43591 19941
rect 43622 19932 43628 19984
rect 43680 19972 43686 19984
rect 43680 19944 43725 19972
rect 43680 19932 43686 19944
rect 44450 19932 44456 19984
rect 44508 19972 44514 19984
rect 45143 19975 45201 19981
rect 45143 19972 45155 19975
rect 44508 19944 45155 19972
rect 44508 19932 44514 19944
rect 45143 19941 45155 19944
rect 45189 19941 45201 19975
rect 45143 19935 45201 19941
rect 39761 19907 39819 19913
rect 39761 19873 39773 19907
rect 39807 19873 39819 19907
rect 45002 19904 45008 19916
rect 44963 19876 45008 19904
rect 39761 19867 39819 19873
rect 45002 19864 45008 19876
rect 45060 19864 45066 19916
rect 28442 19836 28448 19848
rect 23155 19808 23474 19836
rect 28000 19808 28448 19836
rect 23155 19805 23167 19808
rect 23109 19799 23167 19805
rect 16132 19740 17540 19768
rect 17773 19771 17831 19777
rect 17773 19737 17785 19771
rect 17819 19768 17831 19771
rect 17862 19768 17868 19780
rect 17819 19740 17868 19768
rect 17819 19737 17831 19740
rect 17773 19731 17831 19737
rect 17862 19728 17868 19740
rect 17920 19728 17926 19780
rect 23446 19768 23474 19808
rect 28442 19796 28448 19808
rect 28500 19796 28506 19848
rect 28810 19796 28816 19848
rect 28868 19836 28874 19848
rect 29641 19839 29699 19845
rect 29641 19836 29653 19839
rect 28868 19808 29653 19836
rect 28868 19796 28874 19808
rect 29641 19805 29653 19808
rect 29687 19836 29699 19839
rect 29730 19836 29736 19848
rect 29687 19808 29736 19836
rect 29687 19805 29699 19808
rect 29641 19799 29699 19805
rect 29730 19796 29736 19808
rect 29788 19836 29794 19848
rect 30285 19839 30343 19845
rect 30285 19836 30297 19839
rect 29788 19808 30297 19836
rect 29788 19796 29794 19808
rect 30285 19805 30297 19808
rect 30331 19805 30343 19839
rect 32214 19836 32220 19848
rect 32175 19808 32220 19836
rect 30285 19799 30343 19805
rect 32214 19796 32220 19808
rect 32272 19796 32278 19848
rect 34057 19839 34115 19845
rect 34057 19805 34069 19839
rect 34103 19836 34115 19839
rect 34790 19836 34796 19848
rect 34103 19808 34796 19836
rect 34103 19805 34115 19808
rect 34057 19799 34115 19805
rect 34790 19796 34796 19808
rect 34848 19836 34854 19848
rect 35618 19836 35624 19848
rect 34848 19808 35624 19836
rect 34848 19796 34854 19808
rect 35618 19796 35624 19808
rect 35676 19796 35682 19848
rect 36170 19836 36176 19848
rect 36131 19808 36176 19836
rect 36170 19796 36176 19808
rect 36228 19796 36234 19848
rect 36814 19836 36820 19848
rect 36775 19808 36820 19836
rect 36814 19796 36820 19808
rect 36872 19796 36878 19848
rect 37458 19796 37464 19848
rect 37516 19836 37522 19848
rect 38105 19839 38163 19845
rect 38105 19836 38117 19839
rect 37516 19808 38117 19836
rect 37516 19796 37522 19808
rect 38105 19805 38117 19808
rect 38151 19805 38163 19839
rect 38105 19799 38163 19805
rect 40037 19839 40095 19845
rect 40037 19805 40049 19839
rect 40083 19836 40095 19839
rect 41506 19836 41512 19848
rect 40083 19808 41512 19836
rect 40083 19805 40095 19808
rect 40037 19799 40095 19805
rect 41506 19796 41512 19808
rect 41564 19796 41570 19848
rect 41693 19839 41751 19845
rect 41693 19805 41705 19839
rect 41739 19805 41751 19839
rect 41966 19836 41972 19848
rect 41927 19808 41972 19836
rect 41693 19799 41751 19805
rect 24765 19771 24823 19777
rect 24765 19768 24777 19771
rect 23446 19740 24777 19768
rect 24765 19737 24777 19740
rect 24811 19768 24823 19771
rect 29917 19771 29975 19777
rect 24811 19740 25452 19768
rect 24811 19737 24823 19740
rect 24765 19731 24823 19737
rect 25424 19712 25452 19740
rect 29917 19737 29929 19771
rect 29963 19768 29975 19771
rect 33226 19768 33232 19780
rect 29963 19740 33232 19768
rect 29963 19737 29975 19740
rect 29917 19731 29975 19737
rect 33226 19728 33232 19740
rect 33284 19728 33290 19780
rect 33778 19728 33784 19780
rect 33836 19768 33842 19780
rect 34609 19771 34667 19777
rect 34609 19768 34621 19771
rect 33836 19740 34621 19768
rect 33836 19728 33842 19740
rect 34609 19737 34621 19740
rect 34655 19768 34667 19771
rect 36832 19768 36860 19796
rect 34655 19740 36860 19768
rect 34655 19737 34667 19740
rect 34609 19731 34667 19737
rect 4062 19660 4068 19712
rect 4120 19700 4126 19712
rect 4798 19700 4804 19712
rect 4120 19672 4804 19700
rect 4120 19660 4126 19672
rect 4798 19660 4804 19672
rect 4856 19660 4862 19712
rect 5258 19700 5264 19712
rect 5219 19672 5264 19700
rect 5258 19660 5264 19672
rect 5316 19660 5322 19712
rect 6362 19700 6368 19712
rect 6323 19672 6368 19700
rect 6362 19660 6368 19672
rect 6420 19660 6426 19712
rect 8846 19660 8852 19712
rect 8904 19700 8910 19712
rect 10137 19703 10195 19709
rect 10137 19700 10149 19703
rect 8904 19672 10149 19700
rect 8904 19660 8910 19672
rect 10137 19669 10149 19672
rect 10183 19700 10195 19703
rect 10502 19700 10508 19712
rect 10183 19672 10508 19700
rect 10183 19669 10195 19672
rect 10137 19663 10195 19669
rect 10502 19660 10508 19672
rect 10560 19660 10566 19712
rect 11011 19703 11069 19709
rect 11011 19669 11023 19703
rect 11057 19700 11069 19703
rect 12434 19700 12440 19712
rect 11057 19672 12440 19700
rect 11057 19669 11069 19672
rect 11011 19663 11069 19669
rect 12434 19660 12440 19672
rect 12492 19660 12498 19712
rect 19702 19700 19708 19712
rect 19663 19672 19708 19700
rect 19702 19660 19708 19672
rect 19760 19660 19766 19712
rect 21174 19700 21180 19712
rect 21135 19672 21180 19700
rect 21174 19660 21180 19672
rect 21232 19660 21238 19712
rect 24302 19700 24308 19712
rect 24263 19672 24308 19700
rect 24302 19660 24308 19672
rect 24360 19660 24366 19712
rect 25406 19660 25412 19712
rect 25464 19700 25470 19712
rect 25869 19703 25927 19709
rect 25869 19700 25881 19703
rect 25464 19672 25881 19700
rect 25464 19660 25470 19672
rect 25869 19669 25881 19672
rect 25915 19669 25927 19703
rect 26878 19700 26884 19712
rect 26839 19672 26884 19700
rect 25869 19663 25927 19669
rect 26878 19660 26884 19672
rect 26936 19660 26942 19712
rect 29086 19700 29092 19712
rect 29047 19672 29092 19700
rect 29086 19660 29092 19672
rect 29144 19660 29150 19712
rect 29362 19660 29368 19712
rect 29420 19700 29426 19712
rect 29549 19703 29607 19709
rect 29549 19700 29561 19703
rect 29420 19672 29561 19700
rect 29420 19660 29426 19672
rect 29549 19669 29561 19672
rect 29595 19669 29607 19703
rect 29549 19663 29607 19669
rect 30742 19660 30748 19712
rect 30800 19700 30806 19712
rect 30975 19703 31033 19709
rect 30975 19700 30987 19703
rect 30800 19672 30987 19700
rect 30800 19660 30806 19672
rect 30975 19669 30987 19672
rect 31021 19669 31033 19703
rect 30975 19663 31033 19669
rect 34422 19660 34428 19712
rect 34480 19700 34486 19712
rect 35069 19703 35127 19709
rect 35069 19700 35081 19703
rect 34480 19672 35081 19700
rect 34480 19660 34486 19672
rect 35069 19669 35081 19672
rect 35115 19669 35127 19703
rect 35069 19663 35127 19669
rect 36170 19660 36176 19712
rect 36228 19700 36234 19712
rect 37476 19700 37504 19796
rect 41708 19768 41736 19799
rect 41966 19796 41972 19808
rect 42024 19796 42030 19848
rect 42886 19796 42892 19848
rect 42944 19836 42950 19848
rect 43806 19836 43812 19848
rect 42944 19808 43812 19836
rect 42944 19796 42950 19808
rect 43806 19796 43812 19808
rect 43864 19796 43870 19848
rect 42058 19768 42064 19780
rect 41708 19740 42064 19768
rect 42058 19728 42064 19740
rect 42116 19728 42122 19780
rect 40494 19700 40500 19712
rect 36228 19672 37504 19700
rect 40455 19672 40500 19700
rect 36228 19660 36234 19672
rect 40494 19660 40500 19672
rect 40552 19660 40558 19712
rect 40586 19660 40592 19712
rect 40644 19700 40650 19712
rect 41874 19700 41880 19712
rect 40644 19672 41880 19700
rect 40644 19660 40650 19672
rect 41874 19660 41880 19672
rect 41932 19700 41938 19712
rect 44542 19700 44548 19712
rect 41932 19672 44548 19700
rect 41932 19660 41938 19672
rect 44542 19660 44548 19672
rect 44600 19660 44606 19712
rect 1104 19610 48852 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 48852 19610
rect 1104 19536 48852 19558
rect 3786 19496 3792 19508
rect 3747 19468 3792 19496
rect 3786 19456 3792 19468
rect 3844 19496 3850 19508
rect 5166 19496 5172 19508
rect 3844 19468 5172 19496
rect 3844 19456 3850 19468
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 5534 19496 5540 19508
rect 5495 19468 5540 19496
rect 5534 19456 5540 19468
rect 5592 19456 5598 19508
rect 6273 19499 6331 19505
rect 6273 19465 6285 19499
rect 6319 19496 6331 19499
rect 7006 19496 7012 19508
rect 6319 19468 7012 19496
rect 6319 19465 6331 19468
rect 6273 19459 6331 19465
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 7926 19496 7932 19508
rect 7887 19468 7932 19496
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 9674 19496 9680 19508
rect 9635 19468 9680 19496
rect 9674 19456 9680 19468
rect 9732 19456 9738 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19496 11575 19499
rect 12342 19496 12348 19508
rect 11563 19468 12348 19496
rect 11563 19465 11575 19468
rect 11517 19459 11575 19465
rect 12342 19456 12348 19468
rect 12400 19456 12406 19508
rect 13354 19456 13360 19508
rect 13412 19496 13418 19508
rect 13449 19499 13507 19505
rect 13449 19496 13461 19499
rect 13412 19468 13461 19496
rect 13412 19456 13418 19468
rect 13449 19465 13461 19468
rect 13495 19465 13507 19499
rect 13449 19459 13507 19465
rect 13909 19499 13967 19505
rect 13909 19465 13921 19499
rect 13955 19496 13967 19499
rect 13998 19496 14004 19508
rect 13955 19468 14004 19496
rect 13955 19465 13967 19468
rect 13909 19459 13967 19465
rect 13998 19456 14004 19468
rect 14056 19456 14062 19508
rect 15105 19499 15163 19505
rect 15105 19465 15117 19499
rect 15151 19496 15163 19499
rect 15470 19496 15476 19508
rect 15151 19468 15476 19496
rect 15151 19465 15163 19468
rect 15105 19459 15163 19465
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 16574 19496 16580 19508
rect 16535 19468 16580 19496
rect 16574 19456 16580 19468
rect 16632 19456 16638 19508
rect 17221 19499 17279 19505
rect 17221 19465 17233 19499
rect 17267 19496 17279 19499
rect 17865 19499 17923 19505
rect 17865 19496 17877 19499
rect 17267 19468 17877 19496
rect 17267 19465 17279 19468
rect 17221 19459 17279 19465
rect 17865 19465 17877 19468
rect 17911 19496 17923 19499
rect 18046 19496 18052 19508
rect 17911 19468 18052 19496
rect 17911 19465 17923 19468
rect 17865 19459 17923 19465
rect 18046 19456 18052 19468
rect 18104 19496 18110 19508
rect 18230 19496 18236 19508
rect 18104 19468 18236 19496
rect 18104 19456 18110 19468
rect 18230 19456 18236 19468
rect 18288 19496 18294 19508
rect 19061 19499 19119 19505
rect 19061 19496 19073 19499
rect 18288 19468 19073 19496
rect 18288 19456 18294 19468
rect 19061 19465 19073 19468
rect 19107 19465 19119 19499
rect 19061 19459 19119 19465
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19496 20775 19499
rect 20990 19496 20996 19508
rect 20763 19468 20996 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 21085 19499 21143 19505
rect 21085 19465 21097 19499
rect 21131 19496 21143 19499
rect 21174 19496 21180 19508
rect 21131 19468 21180 19496
rect 21131 19465 21143 19468
rect 21085 19459 21143 19465
rect 21174 19456 21180 19468
rect 21232 19456 21238 19508
rect 22646 19456 22652 19508
rect 22704 19496 22710 19508
rect 22741 19499 22799 19505
rect 22741 19496 22753 19499
rect 22704 19468 22753 19496
rect 22704 19456 22710 19468
rect 22741 19465 22753 19468
rect 22787 19465 22799 19499
rect 22741 19459 22799 19465
rect 27246 19456 27252 19508
rect 27304 19496 27310 19508
rect 27341 19499 27399 19505
rect 27341 19496 27353 19499
rect 27304 19468 27353 19496
rect 27304 19456 27310 19468
rect 27341 19465 27353 19468
rect 27387 19465 27399 19499
rect 27341 19459 27399 19465
rect 28258 19456 28264 19508
rect 28316 19496 28322 19508
rect 28997 19499 29055 19505
rect 28997 19496 29009 19499
rect 28316 19468 29009 19496
rect 28316 19456 28322 19468
rect 28997 19465 29009 19468
rect 29043 19496 29055 19499
rect 29362 19496 29368 19508
rect 29043 19468 29368 19496
rect 29043 19465 29055 19468
rect 28997 19459 29055 19465
rect 29362 19456 29368 19468
rect 29420 19456 29426 19508
rect 29454 19456 29460 19508
rect 29512 19505 29518 19508
rect 29512 19499 29561 19505
rect 29512 19465 29515 19499
rect 29549 19465 29561 19499
rect 29638 19496 29644 19508
rect 29599 19468 29644 19496
rect 29512 19459 29561 19465
rect 29512 19456 29518 19459
rect 29638 19456 29644 19468
rect 29696 19456 29702 19508
rect 30837 19499 30895 19505
rect 30837 19465 30849 19499
rect 30883 19496 30895 19499
rect 30926 19496 30932 19508
rect 30883 19468 30932 19496
rect 30883 19465 30895 19468
rect 30837 19459 30895 19465
rect 30926 19456 30932 19468
rect 30984 19456 30990 19508
rect 32861 19499 32919 19505
rect 32861 19465 32873 19499
rect 32907 19496 32919 19499
rect 32950 19496 32956 19508
rect 32907 19468 32956 19496
rect 32907 19465 32919 19468
rect 32861 19459 32919 19465
rect 32950 19456 32956 19468
rect 33008 19456 33014 19508
rect 33594 19496 33600 19508
rect 33555 19468 33600 19496
rect 33594 19456 33600 19468
rect 33652 19456 33658 19508
rect 35989 19499 36047 19505
rect 35989 19465 36001 19499
rect 36035 19496 36047 19499
rect 36262 19496 36268 19508
rect 36035 19468 36268 19496
rect 36035 19465 36047 19468
rect 35989 19459 36047 19465
rect 36262 19456 36268 19468
rect 36320 19456 36326 19508
rect 37642 19496 37648 19508
rect 36740 19468 37648 19496
rect 4249 19431 4307 19437
rect 4249 19397 4261 19431
rect 4295 19428 4307 19431
rect 4706 19428 4712 19440
rect 4295 19400 4712 19428
rect 4295 19397 4307 19400
rect 4249 19391 4307 19397
rect 4706 19388 4712 19400
rect 4764 19388 4770 19440
rect 6641 19431 6699 19437
rect 6641 19397 6653 19431
rect 6687 19428 6699 19431
rect 6730 19428 6736 19440
rect 6687 19400 6736 19428
rect 6687 19397 6699 19400
rect 6641 19391 6699 19397
rect 6730 19388 6736 19400
rect 6788 19388 6794 19440
rect 11882 19428 11888 19440
rect 11843 19400 11888 19428
rect 11882 19388 11888 19400
rect 11940 19388 11946 19440
rect 13265 19431 13323 19437
rect 13265 19397 13277 19431
rect 13311 19428 13323 19431
rect 15381 19431 15439 19437
rect 15381 19428 15393 19431
rect 13311 19400 15393 19428
rect 13311 19397 13323 19400
rect 13265 19391 13323 19397
rect 15381 19397 15393 19400
rect 15427 19428 15439 19431
rect 15562 19428 15568 19440
rect 15427 19400 15568 19428
rect 15427 19397 15439 19400
rect 15381 19391 15439 19397
rect 15562 19388 15568 19400
rect 15620 19388 15626 19440
rect 16114 19388 16120 19440
rect 16172 19428 16178 19440
rect 16209 19431 16267 19437
rect 16209 19428 16221 19431
rect 16172 19400 16221 19428
rect 16172 19388 16178 19400
rect 16209 19397 16221 19400
rect 16255 19397 16267 19431
rect 16209 19391 16267 19397
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 2958 19360 2964 19372
rect 2731 19332 2964 19360
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 2792 19301 2820 19332
rect 2958 19320 2964 19332
rect 3016 19320 3022 19372
rect 8846 19360 8852 19372
rect 8807 19332 8852 19360
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 12710 19360 12716 19372
rect 10520 19332 12716 19360
rect 10520 19304 10548 19332
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 14369 19363 14427 19369
rect 14369 19360 14381 19363
rect 13786 19332 14381 19360
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19261 2835 19295
rect 2777 19255 2835 19261
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 3237 19295 3295 19301
rect 3237 19292 3249 19295
rect 2924 19264 3249 19292
rect 2924 19252 2930 19264
rect 3237 19261 3249 19264
rect 3283 19261 3295 19295
rect 3237 19255 3295 19261
rect 3513 19295 3571 19301
rect 3513 19261 3525 19295
rect 3559 19292 3571 19295
rect 4338 19292 4344 19304
rect 3559 19264 4344 19292
rect 3559 19261 3571 19264
rect 3513 19255 3571 19261
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 9582 19252 9588 19304
rect 9640 19292 9646 19304
rect 9950 19292 9956 19304
rect 9640 19264 9956 19292
rect 9640 19252 9646 19264
rect 9950 19252 9956 19264
rect 10008 19252 10014 19304
rect 10502 19292 10508 19304
rect 10415 19264 10508 19292
rect 10502 19252 10508 19264
rect 10560 19252 10566 19304
rect 11606 19252 11612 19304
rect 11664 19292 11670 19304
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 11664 19264 12173 19292
rect 11664 19252 11670 19264
rect 12161 19261 12173 19264
rect 12207 19261 12219 19295
rect 12161 19255 12219 19261
rect 6362 19184 6368 19236
rect 6420 19224 6426 19236
rect 6917 19227 6975 19233
rect 6917 19224 6929 19227
rect 6420 19196 6929 19224
rect 6420 19184 6426 19196
rect 6917 19193 6929 19196
rect 6963 19193 6975 19227
rect 6917 19187 6975 19193
rect 7006 19184 7012 19236
rect 7064 19224 7070 19236
rect 7558 19224 7564 19236
rect 7064 19196 7157 19224
rect 7519 19196 7564 19224
rect 7064 19184 7070 19196
rect 7558 19184 7564 19196
rect 7616 19184 7622 19236
rect 8294 19184 8300 19236
rect 8352 19224 8358 19236
rect 8481 19227 8539 19233
rect 8481 19224 8493 19227
rect 8352 19196 8493 19224
rect 8352 19184 8358 19196
rect 8481 19193 8493 19196
rect 8527 19193 8539 19227
rect 8481 19187 8539 19193
rect 8573 19227 8631 19233
rect 8573 19193 8585 19227
rect 8619 19224 8631 19227
rect 9398 19224 9404 19236
rect 8619 19196 9404 19224
rect 8619 19193 8631 19196
rect 8573 19187 8631 19193
rect 4706 19156 4712 19168
rect 4667 19128 4712 19156
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 5261 19159 5319 19165
rect 5261 19125 5273 19159
rect 5307 19156 5319 19159
rect 5442 19156 5448 19168
rect 5307 19128 5448 19156
rect 5307 19125 5319 19128
rect 5261 19119 5319 19125
rect 5442 19116 5448 19128
rect 5500 19116 5506 19168
rect 7024 19156 7052 19184
rect 8205 19159 8263 19165
rect 8205 19156 8217 19159
rect 7024 19128 8217 19156
rect 8205 19125 8217 19128
rect 8251 19156 8263 19159
rect 8588 19156 8616 19187
rect 9398 19184 9404 19196
rect 9456 19184 9462 19236
rect 10686 19224 10692 19236
rect 10647 19196 10692 19224
rect 10686 19184 10692 19196
rect 10744 19184 10750 19236
rect 11054 19156 11060 19168
rect 8251 19128 8616 19156
rect 11015 19128 11060 19156
rect 8251 19125 8263 19128
rect 8205 19119 8263 19125
rect 11054 19116 11060 19128
rect 11112 19116 11118 19168
rect 12176 19156 12204 19255
rect 12250 19184 12256 19236
rect 12308 19224 12314 19236
rect 12529 19227 12587 19233
rect 12529 19224 12541 19227
rect 12308 19196 12541 19224
rect 12308 19184 12314 19196
rect 12529 19193 12541 19196
rect 12575 19193 12587 19227
rect 12529 19187 12587 19193
rect 12621 19227 12679 19233
rect 12621 19193 12633 19227
rect 12667 19193 12679 19227
rect 12621 19187 12679 19193
rect 13173 19227 13231 19233
rect 13173 19193 13185 19227
rect 13219 19224 13231 19227
rect 13786 19224 13814 19332
rect 14369 19329 14381 19332
rect 14415 19360 14427 19363
rect 15657 19363 15715 19369
rect 14415 19332 15516 19360
rect 14415 19329 14427 19332
rect 14369 19323 14427 19329
rect 14090 19224 14096 19236
rect 13219 19196 13814 19224
rect 14051 19196 14096 19224
rect 13219 19193 13231 19196
rect 13173 19187 13231 19193
rect 12636 19156 12664 19187
rect 14090 19184 14096 19196
rect 14148 19184 14154 19236
rect 14185 19227 14243 19233
rect 14185 19193 14197 19227
rect 14231 19193 14243 19227
rect 14185 19187 14243 19193
rect 13265 19159 13323 19165
rect 13265 19156 13277 19159
rect 12176 19128 13277 19156
rect 13265 19125 13277 19128
rect 13311 19125 13323 19159
rect 13265 19119 13323 19125
rect 13998 19116 14004 19168
rect 14056 19156 14062 19168
rect 14200 19156 14228 19187
rect 14056 19128 14228 19156
rect 15488 19156 15516 19332
rect 15657 19329 15669 19363
rect 15703 19360 15715 19363
rect 16592 19360 16620 19456
rect 18966 19388 18972 19440
rect 19024 19428 19030 19440
rect 26786 19428 26792 19440
rect 19024 19400 21312 19428
rect 19024 19388 19030 19400
rect 18782 19360 18788 19372
rect 15703 19332 16620 19360
rect 18743 19332 18788 19360
rect 15703 19329 15715 19332
rect 15657 19323 15715 19329
rect 18782 19320 18788 19332
rect 18840 19360 18846 19372
rect 19702 19360 19708 19372
rect 18840 19332 19708 19360
rect 18840 19320 18846 19332
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 20346 19360 20352 19372
rect 20307 19332 20352 19360
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 21284 19369 21312 19400
rect 25332 19400 26792 19428
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 21358 19360 21364 19372
rect 21315 19332 21364 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 21358 19320 21364 19332
rect 21416 19320 21422 19372
rect 21542 19360 21548 19372
rect 21503 19332 21548 19360
rect 21542 19320 21548 19332
rect 21600 19320 21606 19372
rect 23937 19363 23995 19369
rect 23937 19329 23949 19363
rect 23983 19360 23995 19363
rect 24210 19360 24216 19372
rect 23983 19332 24216 19360
rect 23983 19329 23995 19332
rect 23937 19323 23995 19329
rect 24210 19320 24216 19332
rect 24268 19360 24274 19372
rect 25332 19369 25360 19400
rect 26786 19388 26792 19400
rect 26844 19428 26850 19440
rect 30650 19428 30656 19440
rect 26844 19400 30656 19428
rect 26844 19388 26850 19400
rect 30650 19388 30656 19400
rect 30708 19388 30714 19440
rect 32122 19388 32128 19440
rect 32180 19428 32186 19440
rect 36740 19428 36768 19468
rect 37642 19456 37648 19468
rect 37700 19456 37706 19508
rect 37826 19456 37832 19508
rect 37884 19496 37890 19508
rect 38197 19499 38255 19505
rect 38197 19496 38209 19499
rect 37884 19468 38209 19496
rect 37884 19456 37890 19468
rect 38197 19465 38209 19468
rect 38243 19465 38255 19499
rect 38197 19459 38255 19465
rect 39298 19456 39304 19508
rect 39356 19496 39362 19508
rect 39853 19499 39911 19505
rect 39853 19496 39865 19499
rect 39356 19468 39865 19496
rect 39356 19456 39362 19468
rect 39853 19465 39865 19468
rect 39899 19465 39911 19499
rect 39853 19459 39911 19465
rect 41417 19499 41475 19505
rect 41417 19465 41429 19499
rect 41463 19496 41475 19499
rect 41782 19496 41788 19508
rect 41463 19468 41788 19496
rect 41463 19465 41475 19468
rect 41417 19459 41475 19465
rect 41782 19456 41788 19468
rect 41840 19456 41846 19508
rect 43349 19499 43407 19505
rect 43349 19465 43361 19499
rect 43395 19496 43407 19499
rect 43530 19496 43536 19508
rect 43395 19468 43536 19496
rect 43395 19465 43407 19468
rect 43349 19459 43407 19465
rect 43530 19456 43536 19468
rect 43588 19456 43594 19508
rect 43714 19496 43720 19508
rect 43675 19468 43720 19496
rect 43714 19456 43720 19468
rect 43772 19456 43778 19508
rect 32180 19400 36768 19428
rect 32180 19388 32186 19400
rect 36814 19388 36820 19440
rect 36872 19428 36878 19440
rect 37461 19431 37519 19437
rect 37461 19428 37473 19431
rect 36872 19400 37473 19428
rect 36872 19388 36878 19400
rect 37461 19397 37473 19400
rect 37507 19397 37519 19431
rect 37918 19428 37924 19440
rect 37879 19400 37924 19428
rect 37461 19391 37519 19397
rect 37918 19388 37924 19400
rect 37976 19388 37982 19440
rect 43548 19428 43576 19456
rect 43993 19431 44051 19437
rect 43993 19428 44005 19431
rect 43548 19400 44005 19428
rect 43993 19397 44005 19400
rect 44039 19397 44051 19431
rect 43993 19391 44051 19397
rect 25317 19363 25375 19369
rect 25317 19360 25329 19363
rect 24268 19332 25329 19360
rect 24268 19320 24274 19332
rect 25317 19329 25329 19332
rect 25363 19329 25375 19363
rect 29730 19360 29736 19372
rect 29691 19332 29736 19360
rect 25317 19323 25375 19329
rect 29730 19320 29736 19332
rect 29788 19320 29794 19372
rect 32306 19320 32312 19372
rect 32364 19320 32370 19372
rect 39577 19363 39635 19369
rect 39577 19329 39589 19363
rect 39623 19360 39635 19363
rect 40494 19360 40500 19372
rect 39623 19332 40500 19360
rect 39623 19329 39635 19332
rect 39577 19323 39635 19329
rect 40494 19320 40500 19332
rect 40552 19320 40558 19372
rect 41506 19320 41512 19372
rect 41564 19360 41570 19372
rect 42426 19360 42432 19372
rect 41564 19332 42432 19360
rect 41564 19320 41570 19332
rect 42426 19320 42432 19332
rect 42484 19320 42490 19372
rect 24673 19295 24731 19301
rect 24673 19292 24685 19295
rect 24412 19264 24685 19292
rect 15746 19224 15752 19236
rect 15707 19196 15752 19224
rect 15746 19184 15752 19196
rect 15804 19184 15810 19236
rect 18138 19224 18144 19236
rect 16224 19196 18144 19224
rect 16224 19156 16252 19196
rect 18138 19184 18144 19196
rect 18196 19184 18202 19236
rect 18230 19184 18236 19236
rect 18288 19224 18294 19236
rect 19521 19227 19579 19233
rect 18288 19196 18333 19224
rect 18288 19184 18294 19196
rect 19521 19193 19533 19227
rect 19567 19224 19579 19227
rect 19797 19227 19855 19233
rect 19797 19224 19809 19227
rect 19567 19196 19809 19224
rect 19567 19193 19579 19196
rect 19521 19187 19579 19193
rect 19797 19193 19809 19196
rect 19843 19193 19855 19227
rect 19797 19187 19855 19193
rect 21361 19227 21419 19233
rect 21361 19193 21373 19227
rect 21407 19193 21419 19227
rect 21361 19187 21419 19193
rect 15488 19128 16252 19156
rect 19812 19156 19840 19187
rect 21174 19156 21180 19168
rect 19812 19128 21180 19156
rect 14056 19116 14062 19128
rect 21174 19116 21180 19128
rect 21232 19156 21238 19168
rect 21376 19156 21404 19187
rect 24412 19168 24440 19264
rect 24673 19261 24685 19264
rect 24719 19292 24731 19295
rect 26329 19295 26387 19301
rect 26329 19292 26341 19295
rect 24719 19264 26341 19292
rect 24719 19261 24731 19264
rect 24673 19255 24731 19261
rect 26329 19261 26341 19264
rect 26375 19292 26387 19295
rect 26973 19295 27031 19301
rect 26973 19292 26985 19295
rect 26375 19264 26985 19292
rect 26375 19261 26387 19264
rect 26329 19255 26387 19261
rect 26973 19261 26985 19264
rect 27019 19261 27031 19295
rect 27522 19292 27528 19304
rect 27483 19264 27528 19292
rect 26973 19255 27031 19261
rect 27522 19252 27528 19264
rect 27580 19252 27586 19304
rect 27706 19252 27712 19304
rect 27764 19292 27770 19304
rect 29086 19292 29092 19304
rect 27764 19264 29092 19292
rect 27764 19252 27770 19264
rect 29086 19252 29092 19264
rect 29144 19292 29150 19304
rect 29365 19295 29423 19301
rect 29365 19292 29377 19295
rect 29144 19264 29377 19292
rect 29144 19252 29150 19264
rect 29365 19261 29377 19264
rect 29411 19292 29423 19295
rect 30377 19295 30435 19301
rect 30377 19292 30389 19295
rect 29411 19264 30389 19292
rect 29411 19261 29423 19264
rect 29365 19255 29423 19261
rect 30377 19261 30389 19264
rect 30423 19261 30435 19295
rect 30377 19255 30435 19261
rect 30837 19295 30895 19301
rect 30837 19261 30849 19295
rect 30883 19292 30895 19295
rect 30926 19292 30932 19304
rect 30984 19301 30990 19304
rect 30984 19295 31022 19301
rect 30883 19264 30932 19292
rect 30883 19261 30895 19264
rect 30837 19255 30895 19261
rect 30926 19252 30932 19264
rect 31010 19261 31022 19295
rect 31938 19292 31944 19304
rect 31899 19264 31944 19292
rect 30984 19255 31022 19261
rect 30984 19252 30990 19255
rect 31938 19252 31944 19264
rect 31996 19252 32002 19304
rect 32324 19292 32352 19320
rect 32950 19292 32956 19304
rect 32324 19264 32956 19292
rect 32950 19252 32956 19264
rect 33008 19292 33014 19304
rect 33756 19295 33814 19301
rect 33756 19292 33768 19295
rect 33008 19264 33768 19292
rect 33008 19252 33014 19264
rect 33756 19261 33768 19264
rect 33802 19292 33814 19295
rect 34149 19295 34207 19301
rect 34149 19292 34161 19295
rect 33802 19264 34161 19292
rect 33802 19261 33814 19264
rect 33756 19255 33814 19261
rect 34149 19261 34161 19264
rect 34195 19261 34207 19295
rect 34149 19255 34207 19261
rect 34422 19252 34428 19304
rect 34480 19292 34486 19304
rect 35069 19295 35127 19301
rect 35069 19292 35081 19295
rect 34480 19264 35081 19292
rect 34480 19252 34486 19264
rect 35069 19261 35081 19264
rect 35115 19261 35127 19295
rect 35069 19255 35127 19261
rect 37550 19252 37556 19304
rect 37608 19292 37614 19304
rect 38749 19295 38807 19301
rect 38749 19292 38761 19295
rect 37608 19264 38761 19292
rect 37608 19252 37614 19264
rect 38749 19261 38761 19264
rect 38795 19292 38807 19295
rect 38841 19295 38899 19301
rect 38841 19292 38853 19295
rect 38795 19264 38853 19292
rect 38795 19261 38807 19264
rect 38749 19255 38807 19261
rect 38841 19261 38853 19264
rect 38887 19261 38899 19295
rect 38841 19255 38899 19261
rect 39206 19252 39212 19304
rect 39264 19292 39270 19304
rect 39301 19295 39359 19301
rect 39301 19292 39313 19295
rect 39264 19264 39313 19292
rect 39264 19252 39270 19264
rect 39301 19261 39313 19264
rect 39347 19261 39359 19295
rect 39301 19255 39359 19261
rect 26053 19227 26111 19233
rect 26053 19193 26065 19227
rect 26099 19224 26111 19227
rect 26142 19224 26148 19236
rect 26099 19196 26148 19224
rect 26099 19193 26111 19196
rect 26053 19187 26111 19193
rect 26142 19184 26148 19196
rect 26200 19184 26206 19236
rect 30098 19224 30104 19236
rect 30059 19196 30104 19224
rect 30098 19184 30104 19196
rect 30156 19184 30162 19236
rect 32030 19184 32036 19236
rect 32088 19224 32094 19236
rect 32262 19227 32320 19233
rect 32262 19224 32274 19227
rect 32088 19196 32274 19224
rect 32088 19184 32094 19196
rect 32262 19193 32274 19196
rect 32308 19224 32320 19227
rect 32490 19224 32496 19236
rect 32308 19196 32496 19224
rect 32308 19193 32320 19196
rect 32262 19187 32320 19193
rect 32490 19184 32496 19196
rect 32548 19224 32554 19236
rect 34609 19227 34667 19233
rect 34609 19224 34621 19227
rect 32548 19196 34621 19224
rect 32548 19184 32554 19196
rect 34609 19193 34621 19196
rect 34655 19224 34667 19227
rect 35342 19224 35348 19236
rect 34655 19196 35348 19224
rect 34655 19193 34667 19196
rect 34609 19187 34667 19193
rect 35342 19184 35348 19196
rect 35400 19233 35406 19236
rect 35400 19227 35448 19233
rect 35400 19193 35402 19227
rect 35436 19193 35448 19227
rect 36906 19224 36912 19236
rect 36867 19196 36912 19224
rect 35400 19187 35448 19193
rect 35400 19184 35406 19187
rect 36906 19184 36912 19196
rect 36964 19184 36970 19236
rect 37001 19227 37059 19233
rect 37001 19193 37013 19227
rect 37047 19193 37059 19227
rect 37001 19187 37059 19193
rect 40818 19227 40876 19233
rect 40818 19193 40830 19227
rect 40864 19193 40876 19227
rect 40818 19187 40876 19193
rect 42750 19227 42808 19233
rect 42750 19193 42762 19227
rect 42796 19193 42808 19227
rect 42750 19187 42808 19193
rect 23106 19156 23112 19168
rect 21232 19128 21404 19156
rect 23067 19128 23112 19156
rect 21232 19116 21238 19128
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 24394 19156 24400 19168
rect 24355 19128 24400 19156
rect 24394 19116 24400 19128
rect 24452 19116 24458 19168
rect 25314 19116 25320 19168
rect 25372 19156 25378 19168
rect 25593 19159 25651 19165
rect 25593 19156 25605 19159
rect 25372 19128 25605 19156
rect 25372 19116 25378 19128
rect 25593 19125 25605 19128
rect 25639 19125 25651 19159
rect 26418 19156 26424 19168
rect 26379 19128 26424 19156
rect 25593 19119 25651 19125
rect 26418 19116 26424 19128
rect 26476 19116 26482 19168
rect 27522 19116 27528 19168
rect 27580 19156 27586 19168
rect 27709 19159 27767 19165
rect 27709 19156 27721 19159
rect 27580 19128 27721 19156
rect 27580 19116 27586 19128
rect 27709 19125 27721 19128
rect 27755 19125 27767 19159
rect 27982 19156 27988 19168
rect 27943 19128 27988 19156
rect 27709 19119 27767 19125
rect 27982 19116 27988 19128
rect 28040 19116 28046 19168
rect 28442 19156 28448 19168
rect 28403 19128 28448 19156
rect 28442 19116 28448 19128
rect 28500 19116 28506 19168
rect 31067 19159 31125 19165
rect 31067 19125 31079 19159
rect 31113 19156 31125 19159
rect 31294 19156 31300 19168
rect 31113 19128 31300 19156
rect 31113 19125 31125 19128
rect 31067 19119 31125 19125
rect 31294 19116 31300 19128
rect 31352 19116 31358 19168
rect 31386 19116 31392 19168
rect 31444 19156 31450 19168
rect 31757 19159 31815 19165
rect 31757 19156 31769 19159
rect 31444 19128 31769 19156
rect 31444 19116 31450 19128
rect 31757 19125 31769 19128
rect 31803 19125 31815 19159
rect 31757 19119 31815 19125
rect 32398 19116 32404 19168
rect 32456 19156 32462 19168
rect 33137 19159 33195 19165
rect 33137 19156 33149 19159
rect 32456 19128 33149 19156
rect 32456 19116 32462 19128
rect 33137 19125 33149 19128
rect 33183 19125 33195 19159
rect 33137 19119 33195 19125
rect 33318 19116 33324 19168
rect 33376 19156 33382 19168
rect 33827 19159 33885 19165
rect 33827 19156 33839 19159
rect 33376 19128 33839 19156
rect 33376 19116 33382 19128
rect 33827 19125 33839 19128
rect 33873 19125 33885 19159
rect 36630 19156 36636 19168
rect 36591 19128 36636 19156
rect 33827 19119 33885 19125
rect 36630 19116 36636 19128
rect 36688 19156 36694 19168
rect 37016 19156 37044 19187
rect 40310 19156 40316 19168
rect 36688 19128 37044 19156
rect 40271 19128 40316 19156
rect 36688 19116 36694 19128
rect 40310 19116 40316 19128
rect 40368 19156 40374 19168
rect 40833 19156 40861 19187
rect 42245 19159 42303 19165
rect 42245 19156 42257 19159
rect 40368 19128 42257 19156
rect 40368 19116 40374 19128
rect 42245 19125 42257 19128
rect 42291 19156 42303 19159
rect 42765 19156 42793 19187
rect 42291 19128 42793 19156
rect 42291 19125 42303 19128
rect 42245 19119 42303 19125
rect 43438 19116 43444 19168
rect 43496 19156 43502 19168
rect 43990 19156 43996 19168
rect 43496 19128 43996 19156
rect 43496 19116 43502 19128
rect 43990 19116 43996 19128
rect 44048 19156 44054 19168
rect 45002 19156 45008 19168
rect 44048 19128 45008 19156
rect 44048 19116 44054 19128
rect 45002 19116 45008 19128
rect 45060 19116 45066 19168
rect 1104 19066 48852 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 48852 19066
rect 1104 18992 48852 19014
rect 2866 18952 2872 18964
rect 2827 18924 2872 18952
rect 2866 18912 2872 18924
rect 2924 18912 2930 18964
rect 4338 18912 4344 18964
rect 4396 18952 4402 18964
rect 4709 18955 4767 18961
rect 4709 18952 4721 18955
rect 4396 18924 4721 18952
rect 4396 18912 4402 18924
rect 4709 18921 4721 18924
rect 4755 18921 4767 18955
rect 6546 18952 6552 18964
rect 6507 18924 6552 18952
rect 4709 18915 4767 18921
rect 6546 18912 6552 18924
rect 6604 18912 6610 18964
rect 7098 18912 7104 18964
rect 7156 18952 7162 18964
rect 7193 18955 7251 18961
rect 7193 18952 7205 18955
rect 7156 18924 7205 18952
rect 7156 18912 7162 18924
rect 7193 18921 7205 18924
rect 7239 18921 7251 18955
rect 9950 18952 9956 18964
rect 9911 18924 9956 18952
rect 7193 18915 7251 18921
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10870 18952 10876 18964
rect 10831 18924 10876 18952
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 12161 18955 12219 18961
rect 12161 18921 12173 18955
rect 12207 18952 12219 18955
rect 12250 18952 12256 18964
rect 12207 18924 12256 18952
rect 12207 18921 12219 18924
rect 12161 18915 12219 18921
rect 12250 18912 12256 18924
rect 12308 18912 12314 18964
rect 13538 18952 13544 18964
rect 13499 18924 13544 18952
rect 13538 18912 13544 18924
rect 13596 18912 13602 18964
rect 14090 18952 14096 18964
rect 14051 18924 14096 18952
rect 14090 18912 14096 18924
rect 14148 18912 14154 18964
rect 14366 18952 14372 18964
rect 14327 18924 14372 18952
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 16255 18955 16313 18961
rect 16255 18921 16267 18955
rect 16301 18952 16313 18955
rect 17954 18952 17960 18964
rect 16301 18924 17960 18952
rect 16301 18921 16313 18924
rect 16255 18915 16313 18921
rect 17954 18912 17960 18924
rect 18012 18912 18018 18964
rect 18138 18952 18144 18964
rect 18099 18924 18144 18952
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 18598 18912 18604 18964
rect 18656 18952 18662 18964
rect 18693 18955 18751 18961
rect 18693 18952 18705 18955
rect 18656 18924 18705 18952
rect 18656 18912 18662 18924
rect 18693 18921 18705 18924
rect 18739 18921 18751 18955
rect 18693 18915 18751 18921
rect 20990 18912 20996 18964
rect 21048 18952 21054 18964
rect 21177 18955 21235 18961
rect 21177 18952 21189 18955
rect 21048 18924 21189 18952
rect 21048 18912 21054 18924
rect 21177 18921 21189 18924
rect 21223 18921 21235 18955
rect 21358 18952 21364 18964
rect 21319 18924 21364 18952
rect 21177 18915 21235 18921
rect 21358 18912 21364 18924
rect 21416 18912 21422 18964
rect 25593 18955 25651 18961
rect 25593 18921 25605 18955
rect 25639 18952 25651 18955
rect 27614 18952 27620 18964
rect 25639 18924 27620 18952
rect 25639 18921 25651 18924
rect 25593 18915 25651 18921
rect 27614 18912 27620 18924
rect 27672 18952 27678 18964
rect 29270 18952 29276 18964
rect 27672 18924 29276 18952
rect 27672 18912 27678 18924
rect 10888 18884 10916 18912
rect 12574 18887 12632 18893
rect 12574 18884 12586 18887
rect 10888 18856 12586 18884
rect 12574 18853 12586 18856
rect 12620 18884 12632 18887
rect 13262 18884 13268 18896
rect 12620 18856 13268 18884
rect 12620 18853 12632 18856
rect 12574 18847 12632 18853
rect 13262 18844 13268 18856
rect 13320 18844 13326 18896
rect 13998 18844 14004 18896
rect 14056 18884 14062 18896
rect 15565 18887 15623 18893
rect 15565 18884 15577 18887
rect 14056 18856 15577 18884
rect 14056 18844 14062 18856
rect 15565 18853 15577 18856
rect 15611 18884 15623 18887
rect 15746 18884 15752 18896
rect 15611 18856 15752 18884
rect 15611 18853 15623 18856
rect 15565 18847 15623 18853
rect 15746 18844 15752 18856
rect 15804 18844 15810 18896
rect 17218 18884 17224 18896
rect 17179 18856 17224 18884
rect 17218 18844 17224 18856
rect 17276 18844 17282 18896
rect 17310 18844 17316 18896
rect 17368 18884 17374 18896
rect 17862 18884 17868 18896
rect 17368 18856 17413 18884
rect 17823 18856 17868 18884
rect 17368 18844 17374 18856
rect 17862 18844 17868 18856
rect 17920 18884 17926 18896
rect 19334 18884 19340 18896
rect 17920 18856 19340 18884
rect 17920 18844 17926 18856
rect 19334 18844 19340 18856
rect 19392 18844 19398 18896
rect 19426 18844 19432 18896
rect 19484 18884 19490 18896
rect 19981 18887 20039 18893
rect 19484 18856 19529 18884
rect 19484 18844 19490 18856
rect 19981 18853 19993 18887
rect 20027 18884 20039 18887
rect 20530 18884 20536 18896
rect 20027 18856 20536 18884
rect 20027 18853 20039 18856
rect 19981 18847 20039 18853
rect 20530 18844 20536 18856
rect 20588 18884 20594 18896
rect 21542 18884 21548 18896
rect 20588 18856 21548 18884
rect 20588 18844 20594 18856
rect 21542 18844 21548 18856
rect 21600 18844 21606 18896
rect 23014 18884 23020 18896
rect 22975 18856 23020 18884
rect 23014 18844 23020 18856
rect 23072 18844 23078 18896
rect 28184 18893 28212 18924
rect 29270 18912 29276 18924
rect 29328 18912 29334 18964
rect 29638 18912 29644 18964
rect 29696 18952 29702 18964
rect 30561 18955 30619 18961
rect 30561 18952 30573 18955
rect 29696 18924 30573 18952
rect 29696 18912 29702 18924
rect 30561 18921 30573 18924
rect 30607 18921 30619 18955
rect 31570 18952 31576 18964
rect 31531 18924 31576 18952
rect 30561 18915 30619 18921
rect 31570 18912 31576 18924
rect 31628 18912 31634 18964
rect 32214 18952 32220 18964
rect 32175 18924 32220 18952
rect 32214 18912 32220 18924
rect 32272 18912 32278 18964
rect 33594 18912 33600 18964
rect 33652 18952 33658 18964
rect 34790 18952 34796 18964
rect 33652 18924 33732 18952
rect 34751 18924 34796 18952
rect 33652 18912 33658 18924
rect 28169 18887 28227 18893
rect 28169 18853 28181 18887
rect 28215 18853 28227 18887
rect 28169 18847 28227 18853
rect 28902 18844 28908 18896
rect 28960 18884 28966 18896
rect 28960 18856 31385 18884
rect 28960 18844 28966 18856
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 4706 18816 4712 18828
rect 4479 18788 4712 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 5074 18776 5080 18828
rect 5132 18816 5138 18828
rect 5261 18819 5319 18825
rect 5261 18816 5273 18819
rect 5132 18788 5273 18816
rect 5132 18776 5138 18788
rect 5261 18785 5273 18788
rect 5307 18785 5319 18819
rect 5718 18816 5724 18828
rect 5679 18788 5724 18816
rect 5261 18779 5319 18785
rect 5718 18776 5724 18788
rect 5776 18776 5782 18828
rect 7745 18819 7803 18825
rect 7745 18785 7757 18819
rect 7791 18816 7803 18819
rect 8570 18816 8576 18828
rect 8628 18825 8634 18828
rect 8628 18819 8666 18825
rect 7791 18788 8576 18816
rect 7791 18785 7803 18788
rect 7745 18779 7803 18785
rect 8570 18776 8576 18788
rect 8654 18785 8666 18819
rect 8628 18779 8666 18785
rect 8628 18776 8634 18779
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 13173 18819 13231 18825
rect 13173 18816 13185 18819
rect 11112 18788 13185 18816
rect 11112 18776 11118 18788
rect 13173 18785 13185 18788
rect 13219 18785 13231 18819
rect 13173 18779 13231 18785
rect 14185 18819 14243 18825
rect 14185 18785 14197 18819
rect 14231 18816 14243 18819
rect 14366 18816 14372 18828
rect 14231 18788 14372 18816
rect 14231 18785 14243 18788
rect 14185 18779 14243 18785
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 16184 18819 16242 18825
rect 16184 18785 16196 18819
rect 16230 18816 16242 18819
rect 16758 18816 16764 18828
rect 16230 18788 16764 18816
rect 16230 18785 16242 18788
rect 16184 18779 16242 18785
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 20968 18819 21026 18825
rect 20968 18785 20980 18819
rect 21014 18816 21026 18819
rect 21726 18816 21732 18828
rect 21014 18788 21732 18816
rect 21014 18785 21026 18788
rect 20968 18779 21026 18785
rect 21726 18776 21732 18788
rect 21784 18776 21790 18828
rect 22925 18819 22983 18825
rect 22925 18785 22937 18819
rect 22971 18785 22983 18819
rect 22925 18779 22983 18785
rect 23385 18819 23443 18825
rect 23385 18785 23397 18819
rect 23431 18816 23443 18819
rect 23658 18816 23664 18828
rect 23431 18788 23664 18816
rect 23431 18785 23443 18788
rect 23385 18779 23443 18785
rect 5997 18751 6055 18757
rect 5997 18717 6009 18751
rect 6043 18748 6055 18751
rect 6825 18751 6883 18757
rect 6825 18748 6837 18751
rect 6043 18720 6837 18748
rect 6043 18717 6055 18720
rect 5997 18711 6055 18717
rect 6825 18717 6837 18720
rect 6871 18748 6883 18751
rect 7374 18748 7380 18760
rect 6871 18720 7380 18748
rect 6871 18717 6883 18720
rect 6825 18711 6883 18717
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 10410 18708 10416 18760
rect 10468 18748 10474 18760
rect 10505 18751 10563 18757
rect 10505 18748 10517 18751
rect 10468 18720 10517 18748
rect 10468 18708 10474 18720
rect 10505 18717 10517 18720
rect 10551 18717 10563 18751
rect 10505 18711 10563 18717
rect 10686 18708 10692 18760
rect 10744 18748 10750 18760
rect 12253 18751 12311 18757
rect 12253 18748 12265 18751
rect 10744 18720 12265 18748
rect 10744 18708 10750 18720
rect 12253 18717 12265 18720
rect 12299 18748 12311 18751
rect 13446 18748 13452 18760
rect 12299 18720 13452 18748
rect 12299 18717 12311 18720
rect 12253 18711 12311 18717
rect 13446 18708 13452 18720
rect 13504 18708 13510 18760
rect 22940 18748 22968 18779
rect 23658 18776 23664 18788
rect 23716 18816 23722 18828
rect 23845 18819 23903 18825
rect 23845 18816 23857 18819
rect 23716 18788 23857 18816
rect 23716 18776 23722 18788
rect 23845 18785 23857 18788
rect 23891 18816 23903 18819
rect 24949 18819 25007 18825
rect 24949 18816 24961 18819
rect 23891 18788 24961 18816
rect 23891 18785 23903 18788
rect 23845 18779 23903 18785
rect 24949 18785 24961 18788
rect 24995 18816 25007 18819
rect 25406 18816 25412 18828
rect 24995 18788 25412 18816
rect 24995 18785 25007 18788
rect 24949 18779 25007 18785
rect 25406 18776 25412 18788
rect 25464 18776 25470 18828
rect 26602 18816 26608 18828
rect 26563 18788 26608 18816
rect 26602 18776 26608 18788
rect 26660 18776 26666 18828
rect 28316 18819 28374 18825
rect 28316 18785 28328 18819
rect 28362 18816 28374 18819
rect 28626 18816 28632 18828
rect 28362 18788 28632 18816
rect 28362 18785 28374 18788
rect 28316 18779 28374 18785
rect 23014 18748 23020 18760
rect 22940 18720 23020 18748
rect 23014 18708 23020 18720
rect 23072 18708 23078 18760
rect 24210 18748 24216 18760
rect 24171 18720 24216 18748
rect 24210 18708 24216 18720
rect 24268 18708 24274 18760
rect 26970 18748 26976 18760
rect 26931 18720 26976 18748
rect 26970 18708 26976 18720
rect 27028 18708 27034 18760
rect 27709 18751 27767 18757
rect 27709 18717 27721 18751
rect 27755 18748 27767 18751
rect 28331 18748 28359 18779
rect 28626 18776 28632 18788
rect 28684 18776 28690 18828
rect 29800 18819 29858 18825
rect 29800 18785 29812 18819
rect 29846 18816 29858 18819
rect 30282 18816 30288 18828
rect 29846 18788 30288 18816
rect 29846 18785 29858 18788
rect 29800 18779 29858 18785
rect 30282 18776 30288 18788
rect 30340 18776 30346 18828
rect 31021 18819 31079 18825
rect 31021 18785 31033 18819
rect 31067 18816 31079 18819
rect 31110 18816 31116 18828
rect 31067 18788 31116 18816
rect 31067 18785 31079 18788
rect 31021 18779 31079 18785
rect 31110 18776 31116 18788
rect 31168 18776 31174 18828
rect 31357 18816 31385 18856
rect 32122 18816 32128 18828
rect 31357 18788 32128 18816
rect 32122 18776 32128 18788
rect 32180 18776 32186 18828
rect 32214 18776 32220 18828
rect 32272 18816 32278 18828
rect 32398 18816 32404 18828
rect 32272 18788 32404 18816
rect 32272 18776 32278 18788
rect 32398 18776 32404 18788
rect 32456 18776 32462 18828
rect 32582 18816 32588 18828
rect 32543 18788 32588 18816
rect 32582 18776 32588 18788
rect 32640 18816 32646 18828
rect 33704 18825 33732 18924
rect 34790 18912 34796 18924
rect 34848 18912 34854 18964
rect 36173 18955 36231 18961
rect 36173 18921 36185 18955
rect 36219 18952 36231 18955
rect 36630 18952 36636 18964
rect 36219 18924 36636 18952
rect 36219 18921 36231 18924
rect 36173 18915 36231 18921
rect 36630 18912 36636 18924
rect 36688 18912 36694 18964
rect 38933 18955 38991 18961
rect 38933 18921 38945 18955
rect 38979 18952 38991 18955
rect 39206 18952 39212 18964
rect 38979 18924 39212 18952
rect 38979 18921 38991 18924
rect 38933 18915 38991 18921
rect 39206 18912 39212 18924
rect 39264 18952 39270 18964
rect 39301 18955 39359 18961
rect 39301 18952 39313 18955
rect 39264 18924 39313 18952
rect 39264 18912 39270 18924
rect 39301 18921 39313 18924
rect 39347 18921 39359 18955
rect 39301 18915 39359 18921
rect 41693 18955 41751 18961
rect 41693 18921 41705 18955
rect 41739 18952 41751 18955
rect 42794 18952 42800 18964
rect 41739 18924 42800 18952
rect 41739 18921 41751 18924
rect 41693 18915 41751 18921
rect 42794 18912 42800 18924
rect 42852 18912 42858 18964
rect 34422 18884 34428 18896
rect 34383 18856 34428 18884
rect 34422 18844 34428 18856
rect 34480 18844 34486 18896
rect 35342 18844 35348 18896
rect 35400 18884 35406 18896
rect 35574 18887 35632 18893
rect 35574 18884 35586 18887
rect 35400 18856 35586 18884
rect 35400 18844 35406 18856
rect 35574 18853 35586 18856
rect 35620 18853 35632 18887
rect 37918 18884 37924 18896
rect 37879 18856 37924 18884
rect 35574 18847 35632 18853
rect 37918 18844 37924 18856
rect 37976 18844 37982 18896
rect 40310 18844 40316 18896
rect 40368 18884 40374 18896
rect 40542 18887 40600 18893
rect 40542 18884 40554 18887
rect 40368 18856 40554 18884
rect 40368 18844 40374 18856
rect 40542 18853 40554 18856
rect 40588 18853 40600 18887
rect 42426 18884 42432 18896
rect 42387 18856 42432 18884
rect 40542 18847 40600 18853
rect 42426 18844 42432 18856
rect 42484 18844 42490 18896
rect 43530 18884 43536 18896
rect 43491 18856 43536 18884
rect 43530 18844 43536 18856
rect 43588 18844 43594 18896
rect 33689 18819 33747 18825
rect 32640 18788 33364 18816
rect 32640 18776 32646 18788
rect 28534 18748 28540 18760
rect 27755 18720 28359 18748
rect 28495 18720 28540 18748
rect 27755 18717 27767 18720
rect 27709 18711 27767 18717
rect 28534 18708 28540 18720
rect 28592 18708 28598 18760
rect 28905 18751 28963 18757
rect 28905 18717 28917 18751
rect 28951 18748 28963 18751
rect 32306 18748 32312 18760
rect 28951 18720 32312 18748
rect 28951 18717 28963 18720
rect 28905 18711 28963 18717
rect 32306 18708 32312 18720
rect 32364 18708 32370 18760
rect 33336 18757 33364 18788
rect 33689 18785 33701 18819
rect 33735 18785 33747 18819
rect 33689 18779 33747 18785
rect 34241 18819 34299 18825
rect 34241 18785 34253 18819
rect 34287 18816 34299 18819
rect 34698 18816 34704 18828
rect 34287 18788 34704 18816
rect 34287 18785 34299 18788
rect 34241 18779 34299 18785
rect 33321 18751 33379 18757
rect 33321 18717 33333 18751
rect 33367 18748 33379 18751
rect 34256 18748 34284 18779
rect 34698 18776 34704 18788
rect 34756 18776 34762 18828
rect 36170 18776 36176 18828
rect 36228 18816 36234 18828
rect 36449 18819 36507 18825
rect 36449 18816 36461 18819
rect 36228 18788 36461 18816
rect 36228 18776 36234 18788
rect 36449 18785 36461 18788
rect 36495 18785 36507 18819
rect 36449 18779 36507 18785
rect 41874 18776 41880 18828
rect 41932 18816 41938 18828
rect 41969 18819 42027 18825
rect 41969 18816 41981 18819
rect 41932 18788 41981 18816
rect 41932 18776 41938 18788
rect 41969 18785 41981 18788
rect 42015 18785 42027 18819
rect 41969 18779 42027 18785
rect 33367 18720 34284 18748
rect 35253 18751 35311 18757
rect 33367 18717 33379 18720
rect 33321 18711 33379 18717
rect 35253 18717 35265 18751
rect 35299 18717 35311 18751
rect 35253 18711 35311 18717
rect 37829 18751 37887 18757
rect 37829 18717 37841 18751
rect 37875 18748 37887 18751
rect 37918 18748 37924 18760
rect 37875 18720 37924 18748
rect 37875 18717 37887 18720
rect 37829 18711 37887 18717
rect 12434 18640 12440 18692
rect 12492 18680 12498 18692
rect 14090 18680 14096 18692
rect 12492 18652 14096 18680
rect 12492 18640 12498 18652
rect 14090 18640 14096 18652
rect 14148 18640 14154 18692
rect 24010 18683 24068 18689
rect 24010 18649 24022 18683
rect 24056 18680 24068 18683
rect 26329 18683 26387 18689
rect 24056 18652 25176 18680
rect 24056 18649 24068 18652
rect 24010 18643 24068 18649
rect 25148 18624 25176 18652
rect 26329 18649 26341 18683
rect 26375 18680 26387 18683
rect 26418 18680 26424 18692
rect 26375 18652 26424 18680
rect 26375 18649 26387 18652
rect 26329 18643 26387 18649
rect 26418 18640 26424 18652
rect 26476 18680 26482 18692
rect 26770 18683 26828 18689
rect 26770 18680 26782 18683
rect 26476 18652 26782 18680
rect 26476 18640 26482 18652
rect 26770 18649 26782 18652
rect 26816 18680 26828 18683
rect 31159 18683 31217 18689
rect 26816 18652 30236 18680
rect 26816 18649 26828 18652
rect 26770 18643 26828 18649
rect 30208 18624 30236 18652
rect 31159 18649 31171 18683
rect 31205 18680 31217 18683
rect 32214 18680 32220 18692
rect 31205 18652 32220 18680
rect 31205 18649 31217 18652
rect 31159 18643 31217 18649
rect 32214 18640 32220 18652
rect 32272 18640 32278 18692
rect 35268 18624 35296 18711
rect 37918 18708 37924 18720
rect 37976 18708 37982 18760
rect 40221 18751 40279 18757
rect 40221 18748 40233 18751
rect 40052 18720 40233 18748
rect 36906 18680 36912 18692
rect 36819 18652 36912 18680
rect 36906 18640 36912 18652
rect 36964 18680 36970 18692
rect 38381 18683 38439 18689
rect 38381 18680 38393 18683
rect 36964 18652 38393 18680
rect 36964 18640 36970 18652
rect 38381 18649 38393 18652
rect 38427 18649 38439 18683
rect 38381 18643 38439 18649
rect 7190 18572 7196 18624
rect 7248 18612 7254 18624
rect 8294 18612 8300 18624
rect 7248 18584 8300 18612
rect 7248 18572 7254 18584
rect 8294 18572 8300 18584
rect 8352 18612 8358 18624
rect 8389 18615 8447 18621
rect 8389 18612 8401 18615
rect 8352 18584 8401 18612
rect 8352 18572 8358 18584
rect 8389 18581 8401 18584
rect 8435 18581 8447 18615
rect 8389 18575 8447 18581
rect 8478 18572 8484 18624
rect 8536 18612 8542 18624
rect 8711 18615 8769 18621
rect 8711 18612 8723 18615
rect 8536 18584 8723 18612
rect 8536 18572 8542 18584
rect 8711 18581 8723 18584
rect 8757 18581 8769 18615
rect 8711 18575 8769 18581
rect 11238 18572 11244 18624
rect 11296 18612 11302 18624
rect 11425 18615 11483 18621
rect 11425 18612 11437 18615
rect 11296 18584 11437 18612
rect 11296 18572 11302 18584
rect 11425 18581 11437 18584
rect 11471 18581 11483 18615
rect 16022 18612 16028 18624
rect 15983 18584 16028 18612
rect 11425 18575 11483 18581
rect 16022 18572 16028 18584
rect 16080 18572 16086 18624
rect 16942 18612 16948 18624
rect 16903 18584 16948 18612
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 23750 18612 23756 18624
rect 23711 18584 23756 18612
rect 23750 18572 23756 18584
rect 23808 18612 23814 18624
rect 24121 18615 24179 18621
rect 24121 18612 24133 18615
rect 23808 18584 24133 18612
rect 23808 18572 23814 18584
rect 24121 18581 24133 18584
rect 24167 18581 24179 18615
rect 24302 18612 24308 18624
rect 24263 18584 24308 18612
rect 24121 18575 24179 18581
rect 24302 18572 24308 18584
rect 24360 18572 24366 18624
rect 25130 18572 25136 18624
rect 25188 18612 25194 18624
rect 25225 18615 25283 18621
rect 25225 18612 25237 18615
rect 25188 18584 25237 18612
rect 25188 18572 25194 18584
rect 25225 18581 25237 18584
rect 25271 18581 25283 18615
rect 26878 18612 26884 18624
rect 26839 18584 26884 18612
rect 25225 18575 25283 18581
rect 26878 18572 26884 18584
rect 26936 18572 26942 18624
rect 27062 18612 27068 18624
rect 27023 18584 27068 18612
rect 27062 18572 27068 18584
rect 27120 18572 27126 18624
rect 28077 18615 28135 18621
rect 28077 18581 28089 18615
rect 28123 18612 28135 18615
rect 28442 18612 28448 18624
rect 28123 18584 28448 18612
rect 28123 18581 28135 18584
rect 28077 18575 28135 18581
rect 28442 18572 28448 18584
rect 28500 18572 28506 18624
rect 29362 18572 29368 18624
rect 29420 18612 29426 18624
rect 29871 18615 29929 18621
rect 29871 18612 29883 18615
rect 29420 18584 29883 18612
rect 29420 18572 29426 18584
rect 29871 18581 29883 18584
rect 29917 18581 29929 18615
rect 30190 18612 30196 18624
rect 30151 18584 30196 18612
rect 29871 18575 29929 18581
rect 30190 18572 30196 18584
rect 30248 18572 30254 18624
rect 31938 18612 31944 18624
rect 31899 18584 31944 18612
rect 31938 18572 31944 18584
rect 31996 18572 32002 18624
rect 35161 18615 35219 18621
rect 35161 18581 35173 18615
rect 35207 18612 35219 18615
rect 35250 18612 35256 18624
rect 35207 18584 35256 18612
rect 35207 18581 35219 18584
rect 35161 18575 35219 18581
rect 35250 18572 35256 18584
rect 35308 18572 35314 18624
rect 39574 18572 39580 18624
rect 39632 18612 39638 18624
rect 40052 18621 40080 18720
rect 40221 18717 40233 18720
rect 40267 18717 40279 18751
rect 40221 18711 40279 18717
rect 43254 18708 43260 18760
rect 43312 18748 43318 18760
rect 43441 18751 43499 18757
rect 43441 18748 43453 18751
rect 43312 18720 43453 18748
rect 43312 18708 43318 18720
rect 43441 18717 43453 18720
rect 43487 18717 43499 18751
rect 43714 18748 43720 18760
rect 43675 18720 43720 18748
rect 43441 18711 43499 18717
rect 43714 18708 43720 18720
rect 43772 18708 43778 18760
rect 41141 18683 41199 18689
rect 41141 18649 41153 18683
rect 41187 18680 41199 18683
rect 42334 18680 42340 18692
rect 41187 18652 42340 18680
rect 41187 18649 41199 18652
rect 41141 18643 41199 18649
rect 42334 18640 42340 18652
rect 42392 18640 42398 18692
rect 40037 18615 40095 18621
rect 40037 18612 40049 18615
rect 39632 18584 40049 18612
rect 39632 18572 39638 18584
rect 40037 18581 40049 18584
rect 40083 18581 40095 18615
rect 40037 18575 40095 18581
rect 40126 18572 40132 18624
rect 40184 18612 40190 18624
rect 42153 18615 42211 18621
rect 42153 18612 42165 18615
rect 40184 18584 42165 18612
rect 40184 18572 40190 18584
rect 42153 18581 42165 18584
rect 42199 18581 42211 18615
rect 42153 18575 42211 18581
rect 1104 18522 48852 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 48852 18522
rect 1104 18448 48852 18470
rect 5074 18368 5080 18420
rect 5132 18408 5138 18420
rect 5261 18411 5319 18417
rect 5261 18408 5273 18411
rect 5132 18380 5273 18408
rect 5132 18368 5138 18380
rect 5261 18377 5273 18380
rect 5307 18377 5319 18411
rect 5261 18371 5319 18377
rect 5859 18411 5917 18417
rect 5859 18377 5871 18411
rect 5905 18408 5917 18411
rect 7190 18408 7196 18420
rect 5905 18380 7196 18408
rect 5905 18377 5917 18380
rect 5859 18371 5917 18377
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 7374 18408 7380 18420
rect 7335 18380 7380 18408
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 9585 18411 9643 18417
rect 9585 18377 9597 18411
rect 9631 18408 9643 18411
rect 9766 18408 9772 18420
rect 9631 18380 9772 18408
rect 9631 18377 9643 18380
rect 9585 18371 9643 18377
rect 9766 18368 9772 18380
rect 9824 18368 9830 18420
rect 11238 18408 11244 18420
rect 11199 18380 11244 18408
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 13446 18408 13452 18420
rect 13407 18380 13452 18408
rect 13446 18368 13452 18380
rect 13504 18368 13510 18420
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 13872 18380 13917 18408
rect 13872 18368 13878 18380
rect 14458 18368 14464 18420
rect 14516 18408 14522 18420
rect 15749 18411 15807 18417
rect 15749 18408 15761 18411
rect 14516 18380 15761 18408
rect 14516 18368 14522 18380
rect 15749 18377 15761 18380
rect 15795 18408 15807 18411
rect 15930 18408 15936 18420
rect 15795 18380 15936 18408
rect 15795 18377 15807 18380
rect 15749 18371 15807 18377
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 17310 18408 17316 18420
rect 17271 18380 17316 18408
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 19426 18408 19432 18420
rect 19387 18380 19432 18408
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 19797 18411 19855 18417
rect 19797 18377 19809 18411
rect 19843 18408 19855 18411
rect 21266 18408 21272 18420
rect 19843 18380 21272 18408
rect 19843 18377 19855 18380
rect 19797 18371 19855 18377
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 24121 18411 24179 18417
rect 24121 18408 24133 18411
rect 23446 18380 24133 18408
rect 4985 18343 5043 18349
rect 4985 18309 4997 18343
rect 5031 18340 5043 18343
rect 5718 18340 5724 18352
rect 5031 18312 5724 18340
rect 5031 18309 5043 18312
rect 4985 18303 5043 18309
rect 4525 18275 4583 18281
rect 4525 18241 4537 18275
rect 4571 18272 4583 18275
rect 4614 18272 4620 18284
rect 4571 18244 4620 18272
rect 4571 18241 4583 18244
rect 4525 18235 4583 18241
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 3697 18207 3755 18213
rect 3697 18173 3709 18207
rect 3743 18204 3755 18207
rect 4062 18204 4068 18216
rect 3743 18176 4068 18204
rect 3743 18173 3755 18176
rect 3697 18167 3755 18173
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 4341 18207 4399 18213
rect 4341 18204 4353 18207
rect 4251 18176 4353 18204
rect 4341 18173 4353 18176
rect 4387 18204 4399 18207
rect 5000 18204 5028 18303
rect 5718 18300 5724 18312
rect 5776 18300 5782 18352
rect 6730 18300 6736 18352
rect 6788 18340 6794 18352
rect 7929 18343 7987 18349
rect 7929 18340 7941 18343
rect 6788 18312 7941 18340
rect 6788 18300 6794 18312
rect 7929 18309 7941 18312
rect 7975 18309 7987 18343
rect 23446 18340 23474 18380
rect 24121 18377 24133 18380
rect 24167 18377 24179 18411
rect 26329 18411 26387 18417
rect 26329 18408 26341 18411
rect 24121 18371 24179 18377
rect 25240 18380 26341 18408
rect 7929 18303 7987 18309
rect 19444 18312 23474 18340
rect 4387 18176 5028 18204
rect 4387 18173 4399 18176
rect 4341 18167 4399 18173
rect 5442 18164 5448 18216
rect 5500 18204 5506 18216
rect 5756 18207 5814 18213
rect 5756 18204 5768 18207
rect 5500 18176 5768 18204
rect 5500 18164 5506 18176
rect 5756 18173 5768 18176
rect 5802 18204 5814 18207
rect 6181 18207 6239 18213
rect 6181 18204 6193 18207
rect 5802 18176 6193 18204
rect 5802 18173 5814 18176
rect 5756 18167 5814 18173
rect 6181 18173 6193 18176
rect 6227 18173 6239 18207
rect 6181 18167 6239 18173
rect 7944 18136 7972 18303
rect 19444 18284 19472 18312
rect 23750 18300 23756 18352
rect 23808 18340 23814 18352
rect 23937 18343 23995 18349
rect 23937 18340 23949 18343
rect 23808 18312 23949 18340
rect 23808 18300 23814 18312
rect 23937 18309 23949 18312
rect 23983 18340 23995 18343
rect 24762 18340 24768 18352
rect 23983 18312 24768 18340
rect 23983 18309 23995 18312
rect 23937 18303 23995 18309
rect 24762 18300 24768 18312
rect 24820 18300 24826 18352
rect 8205 18275 8263 18281
rect 8205 18241 8217 18275
rect 8251 18272 8263 18275
rect 8478 18272 8484 18284
rect 8251 18244 8484 18272
rect 8251 18241 8263 18244
rect 8205 18235 8263 18241
rect 8478 18232 8484 18244
rect 8536 18232 8542 18284
rect 8846 18272 8852 18284
rect 8807 18244 8852 18272
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 9217 18275 9275 18281
rect 9217 18241 9229 18275
rect 9263 18272 9275 18275
rect 11471 18275 11529 18281
rect 9263 18244 10272 18272
rect 9263 18241 9275 18244
rect 9217 18235 9275 18241
rect 9766 18204 9772 18216
rect 9727 18176 9772 18204
rect 9766 18164 9772 18176
rect 9824 18164 9830 18216
rect 10244 18213 10272 18244
rect 11471 18241 11483 18275
rect 11517 18272 11529 18275
rect 12250 18272 12256 18284
rect 11517 18244 12256 18272
rect 11517 18241 11529 18244
rect 11471 18235 11529 18241
rect 12250 18232 12256 18244
rect 12308 18232 12314 18284
rect 14936 18244 16068 18272
rect 10229 18207 10287 18213
rect 10229 18173 10241 18207
rect 10275 18204 10287 18207
rect 10502 18204 10508 18216
rect 10275 18176 10508 18204
rect 10275 18173 10287 18176
rect 10229 18167 10287 18173
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 11238 18164 11244 18216
rect 11296 18204 11302 18216
rect 11368 18207 11426 18213
rect 11368 18204 11380 18207
rect 11296 18176 11380 18204
rect 11296 18164 11302 18176
rect 11368 18173 11380 18176
rect 11414 18173 11426 18207
rect 11368 18167 11426 18173
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 12618 18204 12624 18216
rect 11931 18176 12624 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 12894 18204 12900 18216
rect 12855 18176 12900 18204
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 13814 18164 13820 18216
rect 13872 18204 13878 18216
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 13872 18176 14381 18204
rect 13872 18164 13878 18176
rect 14369 18173 14381 18176
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 14642 18164 14648 18216
rect 14700 18204 14706 18216
rect 14936 18213 14964 18244
rect 16040 18216 16068 18244
rect 19426 18232 19432 18284
rect 19484 18232 19490 18284
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 19628 18244 20177 18272
rect 14921 18207 14979 18213
rect 14921 18204 14933 18207
rect 14700 18176 14933 18204
rect 14700 18164 14706 18176
rect 14921 18173 14933 18176
rect 14967 18173 14979 18207
rect 15930 18204 15936 18216
rect 15891 18176 15936 18204
rect 14921 18167 14979 18173
rect 15930 18164 15936 18176
rect 15988 18164 15994 18216
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 19628 18213 19656 18244
rect 20165 18241 20177 18244
rect 20211 18272 20223 18275
rect 21726 18272 21732 18284
rect 20211 18244 21732 18272
rect 20211 18241 20223 18244
rect 20165 18235 20223 18241
rect 21726 18232 21732 18244
rect 21784 18232 21790 18284
rect 23474 18232 23480 18284
rect 23532 18272 23538 18284
rect 24029 18275 24087 18281
rect 24029 18272 24041 18275
rect 23532 18244 24041 18272
rect 23532 18232 23538 18244
rect 24029 18241 24041 18244
rect 24075 18272 24087 18275
rect 24394 18272 24400 18284
rect 24075 18244 24400 18272
rect 24075 18241 24087 18244
rect 24029 18235 24087 18241
rect 24394 18232 24400 18244
rect 24452 18272 24458 18284
rect 25038 18272 25044 18284
rect 24452 18244 25044 18272
rect 24452 18232 24458 18244
rect 25038 18232 25044 18244
rect 25096 18232 25102 18284
rect 25240 18216 25268 18380
rect 26329 18377 26341 18380
rect 26375 18408 26387 18411
rect 26510 18408 26516 18420
rect 26375 18380 26516 18408
rect 26375 18377 26387 18380
rect 26329 18371 26387 18377
rect 26510 18368 26516 18380
rect 26568 18368 26574 18420
rect 26878 18368 26884 18420
rect 26936 18408 26942 18420
rect 27065 18411 27123 18417
rect 27065 18408 27077 18411
rect 26936 18380 27077 18408
rect 26936 18368 26942 18380
rect 27065 18377 27077 18380
rect 27111 18408 27123 18411
rect 27893 18411 27951 18417
rect 27893 18408 27905 18411
rect 27111 18380 27905 18408
rect 27111 18377 27123 18380
rect 27065 18371 27123 18377
rect 27893 18377 27905 18380
rect 27939 18408 27951 18411
rect 28442 18408 28448 18420
rect 27939 18380 28448 18408
rect 27939 18377 27951 18380
rect 27893 18371 27951 18377
rect 28442 18368 28448 18380
rect 28500 18368 28506 18420
rect 29438 18411 29496 18417
rect 29438 18377 29450 18411
rect 29484 18408 29496 18411
rect 30190 18408 30196 18420
rect 29484 18380 30196 18408
rect 29484 18377 29496 18380
rect 29438 18371 29496 18377
rect 30190 18368 30196 18380
rect 30248 18368 30254 18420
rect 30282 18368 30288 18420
rect 30340 18408 30346 18420
rect 33502 18408 33508 18420
rect 30340 18380 33508 18408
rect 30340 18368 30346 18380
rect 33502 18368 33508 18380
rect 33560 18368 33566 18420
rect 33594 18368 33600 18420
rect 33652 18408 33658 18420
rect 34241 18411 34299 18417
rect 34241 18408 34253 18411
rect 33652 18380 34253 18408
rect 33652 18368 33658 18380
rect 34241 18377 34253 18380
rect 34287 18377 34299 18411
rect 35342 18408 35348 18420
rect 35303 18380 35348 18408
rect 34241 18371 34299 18377
rect 25314 18300 25320 18352
rect 25372 18340 25378 18352
rect 25501 18343 25559 18349
rect 25501 18340 25513 18343
rect 25372 18312 25513 18340
rect 25372 18300 25378 18312
rect 25501 18309 25513 18312
rect 25547 18309 25559 18343
rect 25501 18303 25559 18309
rect 28629 18343 28687 18349
rect 28629 18309 28641 18343
rect 28675 18340 28687 18343
rect 28997 18343 29055 18349
rect 28997 18340 29009 18343
rect 28675 18312 29009 18340
rect 28675 18309 28687 18312
rect 28629 18303 28687 18309
rect 28997 18309 29009 18312
rect 29043 18309 29055 18343
rect 29546 18340 29552 18352
rect 29507 18312 29552 18340
rect 28997 18303 29055 18309
rect 25593 18275 25651 18281
rect 25593 18272 25605 18275
rect 25516 18244 25605 18272
rect 16393 18207 16451 18213
rect 16393 18204 16405 18207
rect 16080 18176 16405 18204
rect 16080 18164 16086 18176
rect 16393 18173 16405 18176
rect 16439 18173 16451 18207
rect 16393 18167 16451 18173
rect 18325 18207 18383 18213
rect 18325 18173 18337 18207
rect 18371 18204 18383 18207
rect 19613 18207 19671 18213
rect 18371 18176 18552 18204
rect 18371 18173 18383 18176
rect 18325 18167 18383 18173
rect 8297 18139 8355 18145
rect 8297 18136 8309 18139
rect 7944 18108 8309 18136
rect 8297 18105 8309 18108
rect 8343 18105 8355 18139
rect 10410 18136 10416 18148
rect 10371 18108 10416 18136
rect 8297 18099 8355 18105
rect 10410 18096 10416 18108
rect 10468 18096 10474 18148
rect 13170 18136 13176 18148
rect 13131 18108 13176 18136
rect 13170 18096 13176 18108
rect 13228 18096 13234 18148
rect 15105 18139 15163 18145
rect 15105 18105 15117 18139
rect 15151 18136 15163 18139
rect 15286 18136 15292 18148
rect 15151 18108 15292 18136
rect 15151 18105 15163 18108
rect 15105 18099 15163 18105
rect 15286 18096 15292 18108
rect 15344 18096 15350 18148
rect 17773 18139 17831 18145
rect 17773 18105 17785 18139
rect 17819 18136 17831 18139
rect 18141 18139 18199 18145
rect 18141 18136 18153 18139
rect 17819 18108 18153 18136
rect 17819 18105 17831 18108
rect 17773 18099 17831 18105
rect 18141 18105 18153 18108
rect 18187 18136 18199 18139
rect 18230 18136 18236 18148
rect 18187 18108 18236 18136
rect 18187 18105 18199 18108
rect 18141 18099 18199 18105
rect 18230 18096 18236 18108
rect 18288 18096 18294 18148
rect 18524 18080 18552 18176
rect 19613 18173 19625 18207
rect 19659 18173 19671 18207
rect 19613 18167 19671 18173
rect 20717 18207 20775 18213
rect 20717 18173 20729 18207
rect 20763 18173 20775 18207
rect 22224 18207 22282 18213
rect 22224 18204 22236 18207
rect 20717 18167 20775 18173
rect 22020 18176 22236 18204
rect 20622 18136 20628 18148
rect 20583 18108 20628 18136
rect 20622 18096 20628 18108
rect 20680 18096 20686 18148
rect 7098 18068 7104 18080
rect 7059 18040 7104 18068
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 10318 18028 10324 18080
rect 10376 18068 10382 18080
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 10376 18040 10701 18068
rect 10376 18028 10382 18040
rect 10689 18037 10701 18040
rect 10735 18068 10747 18071
rect 10870 18068 10876 18080
rect 10735 18040 10876 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 10870 18028 10876 18040
rect 10928 18068 10934 18080
rect 12161 18071 12219 18077
rect 12161 18068 12173 18071
rect 10928 18040 12173 18068
rect 10928 18028 10934 18040
rect 12161 18037 12173 18040
rect 12207 18037 12219 18071
rect 12161 18031 12219 18037
rect 14277 18071 14335 18077
rect 14277 18037 14289 18071
rect 14323 18068 14335 18071
rect 14366 18068 14372 18080
rect 14323 18040 14372 18068
rect 14323 18037 14335 18040
rect 14277 18031 14335 18037
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 16206 18068 16212 18080
rect 16167 18040 16212 18068
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 16758 18028 16764 18080
rect 16816 18068 16822 18080
rect 16945 18071 17003 18077
rect 16945 18068 16957 18071
rect 16816 18040 16957 18068
rect 16816 18028 16822 18040
rect 16945 18037 16957 18040
rect 16991 18037 17003 18071
rect 16945 18031 17003 18037
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 18417 18071 18475 18077
rect 18417 18068 18429 18071
rect 17920 18040 18429 18068
rect 17920 18028 17926 18040
rect 18417 18037 18429 18040
rect 18463 18037 18475 18071
rect 18417 18031 18475 18037
rect 18506 18028 18512 18080
rect 18564 18068 18570 18080
rect 18969 18071 19027 18077
rect 18969 18068 18981 18071
rect 18564 18040 18981 18068
rect 18564 18028 18570 18040
rect 18969 18037 18981 18040
rect 19015 18037 19027 18071
rect 20438 18068 20444 18080
rect 20399 18040 20444 18068
rect 18969 18031 19027 18037
rect 20438 18028 20444 18040
rect 20496 18068 20502 18080
rect 20732 18068 20760 18167
rect 22020 18080 22048 18176
rect 22224 18173 22236 18176
rect 22270 18173 22282 18207
rect 23808 18207 23866 18213
rect 23808 18204 23820 18207
rect 22224 18167 22282 18173
rect 23216 18176 23820 18204
rect 23216 18080 23244 18176
rect 23808 18173 23820 18176
rect 23854 18173 23866 18207
rect 25222 18204 25228 18216
rect 25135 18176 25228 18204
rect 23808 18167 23866 18173
rect 25222 18164 25228 18176
rect 25280 18164 25286 18216
rect 25372 18207 25430 18213
rect 25372 18173 25384 18207
rect 25418 18173 25430 18207
rect 25372 18167 25430 18173
rect 23658 18136 23664 18148
rect 23619 18108 23664 18136
rect 23658 18096 23664 18108
rect 23716 18096 23722 18148
rect 25130 18096 25136 18148
rect 25188 18136 25194 18148
rect 25387 18136 25415 18167
rect 25188 18108 25415 18136
rect 25188 18096 25194 18108
rect 22002 18068 22008 18080
rect 20496 18040 20760 18068
rect 21963 18040 22008 18068
rect 20496 18028 20502 18040
rect 22002 18028 22008 18040
rect 22060 18028 22066 18080
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 22327 18071 22385 18077
rect 22327 18068 22339 18071
rect 22152 18040 22339 18068
rect 22152 18028 22158 18040
rect 22327 18037 22339 18040
rect 22373 18037 22385 18071
rect 22327 18031 22385 18037
rect 22741 18071 22799 18077
rect 22741 18037 22753 18071
rect 22787 18068 22799 18071
rect 23014 18068 23020 18080
rect 22787 18040 23020 18068
rect 22787 18037 22799 18040
rect 22741 18031 22799 18037
rect 23014 18028 23020 18040
rect 23072 18028 23078 18080
rect 23109 18071 23167 18077
rect 23109 18037 23121 18071
rect 23155 18068 23167 18071
rect 23198 18068 23204 18080
rect 23155 18040 23204 18068
rect 23155 18037 23167 18040
rect 23109 18031 23167 18037
rect 23198 18028 23204 18040
rect 23256 18028 23262 18080
rect 24762 18068 24768 18080
rect 24723 18040 24768 18068
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 25038 18068 25044 18080
rect 24999 18040 25044 18068
rect 25038 18028 25044 18040
rect 25096 18068 25102 18080
rect 25516 18068 25544 18244
rect 25593 18241 25605 18244
rect 25639 18241 25651 18275
rect 25593 18235 25651 18241
rect 26970 18232 26976 18284
rect 27028 18272 27034 18284
rect 27982 18272 27988 18284
rect 27028 18244 27988 18272
rect 27028 18232 27034 18244
rect 27982 18232 27988 18244
rect 28040 18272 28046 18284
rect 28534 18272 28540 18284
rect 28040 18244 28540 18272
rect 28040 18232 28046 18244
rect 28534 18232 28540 18244
rect 28592 18272 28598 18284
rect 28644 18272 28672 18303
rect 28592 18244 28672 18272
rect 29012 18272 29040 18303
rect 29546 18300 29552 18312
rect 29604 18300 29610 18352
rect 31110 18340 31116 18352
rect 31023 18312 31116 18340
rect 31110 18300 31116 18312
rect 31168 18340 31174 18352
rect 34054 18340 34060 18352
rect 31168 18312 34060 18340
rect 31168 18300 31174 18312
rect 34054 18300 34060 18312
rect 34112 18300 34118 18352
rect 34256 18340 34284 18371
rect 35342 18368 35348 18380
rect 35400 18368 35406 18420
rect 36449 18411 36507 18417
rect 36449 18377 36461 18411
rect 36495 18408 36507 18411
rect 37093 18411 37151 18417
rect 37093 18408 37105 18411
rect 36495 18380 37105 18408
rect 36495 18377 36507 18380
rect 36449 18371 36507 18377
rect 37093 18377 37105 18380
rect 37139 18408 37151 18411
rect 37826 18408 37832 18420
rect 37139 18380 37832 18408
rect 37139 18377 37151 18380
rect 37093 18371 37151 18377
rect 37826 18368 37832 18380
rect 37884 18368 37890 18420
rect 38102 18368 38108 18420
rect 38160 18408 38166 18420
rect 39298 18408 39304 18420
rect 38160 18380 39304 18408
rect 38160 18368 38166 18380
rect 39298 18368 39304 18380
rect 39356 18368 39362 18420
rect 41874 18368 41880 18420
rect 41932 18408 41938 18420
rect 41969 18411 42027 18417
rect 41969 18408 41981 18411
rect 41932 18380 41981 18408
rect 41932 18368 41938 18380
rect 41969 18377 41981 18380
rect 42015 18377 42027 18411
rect 43441 18411 43499 18417
rect 43441 18408 43453 18411
rect 41969 18371 42027 18377
rect 42766 18380 43453 18408
rect 40034 18340 40040 18352
rect 34256 18312 40040 18340
rect 40034 18300 40040 18312
rect 40092 18300 40098 18352
rect 41417 18343 41475 18349
rect 41417 18309 41429 18343
rect 41463 18340 41475 18343
rect 42766 18340 42794 18380
rect 43441 18377 43453 18380
rect 43487 18408 43499 18411
rect 43530 18408 43536 18420
rect 43487 18380 43536 18408
rect 43487 18377 43499 18380
rect 43441 18371 43499 18377
rect 43530 18368 43536 18380
rect 43588 18368 43594 18420
rect 41463 18312 42794 18340
rect 41463 18309 41475 18312
rect 41417 18303 41475 18309
rect 43254 18300 43260 18352
rect 43312 18340 43318 18352
rect 43809 18343 43867 18349
rect 43809 18340 43821 18343
rect 43312 18312 43821 18340
rect 43312 18300 43318 18312
rect 43809 18309 43821 18312
rect 43855 18309 43867 18343
rect 43809 18303 43867 18309
rect 29641 18275 29699 18281
rect 29641 18272 29653 18275
rect 29012 18244 29653 18272
rect 28592 18232 28598 18244
rect 29641 18241 29653 18244
rect 29687 18241 29699 18275
rect 29641 18235 29699 18241
rect 29914 18232 29920 18284
rect 29972 18272 29978 18284
rect 31938 18272 31944 18284
rect 29972 18244 31432 18272
rect 31899 18244 31944 18272
rect 29972 18232 29978 18244
rect 27154 18164 27160 18216
rect 27212 18204 27218 18216
rect 27764 18207 27822 18213
rect 27764 18204 27776 18207
rect 27212 18176 27776 18204
rect 27212 18164 27218 18176
rect 27764 18173 27776 18176
rect 27810 18204 27822 18207
rect 28626 18204 28632 18216
rect 27810 18176 28632 18204
rect 27810 18173 27822 18176
rect 27764 18167 27822 18173
rect 28626 18164 28632 18176
rect 28684 18164 28690 18216
rect 29270 18204 29276 18216
rect 29231 18176 29276 18204
rect 29270 18164 29276 18176
rect 29328 18204 29334 18216
rect 31404 18213 31432 18244
rect 31938 18232 31944 18244
rect 31996 18232 32002 18284
rect 33042 18232 33048 18284
rect 33100 18272 33106 18284
rect 34146 18272 34152 18284
rect 33100 18244 34152 18272
rect 33100 18232 33106 18244
rect 34146 18232 34152 18244
rect 34204 18232 34210 18284
rect 38381 18275 38439 18281
rect 38381 18241 38393 18275
rect 38427 18272 38439 18275
rect 39574 18272 39580 18284
rect 38427 18244 39252 18272
rect 39535 18244 39580 18272
rect 38427 18241 38439 18244
rect 38381 18235 38439 18241
rect 39224 18216 39252 18244
rect 39574 18232 39580 18244
rect 39632 18232 39638 18284
rect 42334 18232 42340 18284
rect 42392 18272 42398 18284
rect 42794 18272 42800 18284
rect 42392 18244 42800 18272
rect 42392 18232 42398 18244
rect 42794 18232 42800 18244
rect 42852 18232 42858 18284
rect 42981 18275 43039 18281
rect 42981 18241 42993 18275
rect 43027 18272 43039 18275
rect 43714 18272 43720 18284
rect 43027 18244 43720 18272
rect 43027 18241 43039 18244
rect 42981 18235 43039 18241
rect 30653 18207 30711 18213
rect 30653 18204 30665 18207
rect 29328 18176 30665 18204
rect 29328 18164 29334 18176
rect 30653 18173 30665 18176
rect 30699 18173 30711 18207
rect 30653 18167 30711 18173
rect 31389 18207 31447 18213
rect 31389 18173 31401 18207
rect 31435 18204 31447 18207
rect 31478 18204 31484 18216
rect 31435 18176 31484 18204
rect 31435 18173 31447 18176
rect 31389 18167 31447 18173
rect 31478 18164 31484 18176
rect 31536 18164 31542 18216
rect 31846 18204 31852 18216
rect 31807 18176 31852 18204
rect 31846 18164 31852 18176
rect 31904 18164 31910 18216
rect 33229 18207 33287 18213
rect 33229 18173 33241 18207
rect 33275 18173 33287 18207
rect 33229 18167 33287 18173
rect 33781 18207 33839 18213
rect 33781 18173 33793 18207
rect 33827 18173 33839 18207
rect 33781 18167 33839 18173
rect 33965 18207 34023 18213
rect 33965 18173 33977 18207
rect 34011 18204 34023 18207
rect 35529 18207 35587 18213
rect 35529 18204 35541 18207
rect 34011 18176 35541 18204
rect 34011 18173 34023 18176
rect 33965 18167 34023 18173
rect 35529 18173 35541 18176
rect 35575 18204 35587 18207
rect 36725 18207 36783 18213
rect 36725 18204 36737 18207
rect 35575 18176 36737 18204
rect 35575 18173 35587 18176
rect 35529 18167 35587 18173
rect 36725 18173 36737 18176
rect 36771 18173 36783 18207
rect 36725 18167 36783 18173
rect 37328 18207 37386 18213
rect 37328 18173 37340 18207
rect 37374 18204 37386 18207
rect 37374 18173 37387 18204
rect 37328 18167 37387 18173
rect 26694 18096 26700 18148
rect 26752 18136 26758 18148
rect 27614 18136 27620 18148
rect 26752 18108 27620 18136
rect 26752 18096 26758 18108
rect 27614 18096 27620 18108
rect 27672 18096 27678 18148
rect 28353 18139 28411 18145
rect 28353 18105 28365 18139
rect 28399 18136 28411 18139
rect 29178 18136 29184 18148
rect 28399 18108 29184 18136
rect 28399 18105 28411 18108
rect 28353 18099 28411 18105
rect 29178 18096 29184 18108
rect 29236 18096 29242 18148
rect 31110 18136 31116 18148
rect 29288 18108 31116 18136
rect 25866 18068 25872 18080
rect 25096 18040 25544 18068
rect 25827 18040 25872 18068
rect 25096 18028 25102 18040
rect 25866 18028 25872 18040
rect 25924 18028 25930 18080
rect 26234 18028 26240 18080
rect 26292 18068 26298 18080
rect 26605 18071 26663 18077
rect 26605 18068 26617 18071
rect 26292 18040 26617 18068
rect 26292 18028 26298 18040
rect 26605 18037 26617 18040
rect 26651 18068 26663 18071
rect 26970 18068 26976 18080
rect 26651 18040 26976 18068
rect 26651 18037 26663 18040
rect 26605 18031 26663 18037
rect 26970 18028 26976 18040
rect 27028 18068 27034 18080
rect 27433 18071 27491 18077
rect 27433 18068 27445 18071
rect 27028 18040 27445 18068
rect 27028 18028 27034 18040
rect 27433 18037 27445 18040
rect 27479 18037 27491 18071
rect 27433 18031 27491 18037
rect 27890 18028 27896 18080
rect 27948 18068 27954 18080
rect 29288 18068 29316 18108
rect 31110 18096 31116 18108
rect 31168 18096 31174 18148
rect 32674 18096 32680 18148
rect 32732 18136 32738 18148
rect 33042 18136 33048 18148
rect 32732 18108 33048 18136
rect 32732 18096 32738 18108
rect 33042 18096 33048 18108
rect 33100 18136 33106 18148
rect 33244 18136 33272 18167
rect 33100 18108 33272 18136
rect 33796 18136 33824 18167
rect 33796 18108 34744 18136
rect 33100 18096 33106 18108
rect 34716 18080 34744 18108
rect 35342 18096 35348 18148
rect 35400 18136 35406 18148
rect 35802 18136 35808 18148
rect 35400 18108 35808 18136
rect 35400 18096 35406 18108
rect 35802 18096 35808 18108
rect 35860 18145 35866 18148
rect 35860 18139 35908 18145
rect 35860 18105 35862 18139
rect 35896 18105 35908 18139
rect 35860 18099 35908 18105
rect 35860 18096 35866 18099
rect 29914 18068 29920 18080
rect 27948 18040 29316 18068
rect 29875 18040 29920 18068
rect 27948 18028 27954 18040
rect 29914 18028 29920 18040
rect 29972 18028 29978 18080
rect 30282 18068 30288 18080
rect 30243 18040 30288 18068
rect 30282 18028 30288 18040
rect 30340 18028 30346 18080
rect 32398 18028 32404 18080
rect 32456 18068 32462 18080
rect 32493 18071 32551 18077
rect 32493 18068 32505 18071
rect 32456 18040 32505 18068
rect 32456 18028 32462 18040
rect 32493 18037 32505 18040
rect 32539 18068 32551 18071
rect 32766 18068 32772 18080
rect 32539 18040 32772 18068
rect 32539 18037 32551 18040
rect 32493 18031 32551 18037
rect 32766 18028 32772 18040
rect 32824 18028 32830 18080
rect 34698 18068 34704 18080
rect 34659 18040 34704 18068
rect 34698 18028 34704 18040
rect 34756 18028 34762 18080
rect 37359 18068 37387 18167
rect 38654 18164 38660 18216
rect 38712 18204 38718 18216
rect 38841 18207 38899 18213
rect 38841 18204 38853 18207
rect 38712 18176 38853 18204
rect 38712 18164 38718 18176
rect 38841 18173 38853 18176
rect 38887 18204 38899 18207
rect 39022 18204 39028 18216
rect 38887 18176 39028 18204
rect 38887 18173 38899 18176
rect 38841 18167 38899 18173
rect 39022 18164 39028 18176
rect 39080 18164 39086 18216
rect 39206 18164 39212 18216
rect 39264 18204 39270 18216
rect 39301 18207 39359 18213
rect 39301 18204 39313 18207
rect 39264 18176 39313 18204
rect 39264 18164 39270 18176
rect 39301 18173 39313 18176
rect 39347 18173 39359 18207
rect 40494 18204 40500 18216
rect 40455 18176 40500 18204
rect 39301 18167 39359 18173
rect 40494 18164 40500 18176
rect 40552 18164 40558 18216
rect 37415 18139 37473 18145
rect 37415 18105 37427 18139
rect 37461 18136 37473 18139
rect 37918 18136 37924 18148
rect 37461 18108 37924 18136
rect 37461 18105 37473 18108
rect 37415 18099 37473 18105
rect 37918 18096 37924 18108
rect 37976 18096 37982 18148
rect 40818 18139 40876 18145
rect 40818 18105 40830 18139
rect 40864 18105 40876 18139
rect 42334 18136 42340 18148
rect 42295 18108 42340 18136
rect 40818 18099 40876 18105
rect 37642 18068 37648 18080
rect 37359 18040 37648 18068
rect 37642 18028 37648 18040
rect 37700 18068 37706 18080
rect 37737 18071 37795 18077
rect 37737 18068 37749 18071
rect 37700 18040 37749 18068
rect 37700 18028 37706 18040
rect 37737 18037 37749 18040
rect 37783 18068 37795 18071
rect 38470 18068 38476 18080
rect 37783 18040 38476 18068
rect 37783 18037 37795 18040
rect 37737 18031 37795 18037
rect 38470 18028 38476 18040
rect 38528 18028 38534 18080
rect 38654 18068 38660 18080
rect 38615 18040 38660 18068
rect 38654 18028 38660 18040
rect 38712 18028 38718 18080
rect 39666 18028 39672 18080
rect 39724 18068 39730 18080
rect 39853 18071 39911 18077
rect 39853 18068 39865 18071
rect 39724 18040 39865 18068
rect 39724 18028 39730 18040
rect 39853 18037 39865 18040
rect 39899 18068 39911 18071
rect 40221 18071 40279 18077
rect 40221 18068 40233 18071
rect 39899 18040 40233 18068
rect 39899 18037 39911 18040
rect 39853 18031 39911 18037
rect 40221 18037 40233 18040
rect 40267 18068 40279 18071
rect 40310 18068 40316 18080
rect 40267 18040 40316 18068
rect 40267 18037 40279 18040
rect 40221 18031 40279 18037
rect 40310 18028 40316 18040
rect 40368 18068 40374 18080
rect 40833 18068 40861 18099
rect 42334 18096 42340 18108
rect 42392 18096 42398 18148
rect 42426 18096 42432 18148
rect 42484 18136 42490 18148
rect 42484 18108 42529 18136
rect 42484 18096 42490 18108
rect 40368 18040 40861 18068
rect 40368 18028 40374 18040
rect 42058 18028 42064 18080
rect 42116 18068 42122 18080
rect 42996 18068 43024 18235
rect 43714 18232 43720 18244
rect 43772 18232 43778 18284
rect 42116 18040 43024 18068
rect 42116 18028 42122 18040
rect 1104 17978 48852 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 48852 17978
rect 1104 17904 48852 17926
rect 2866 17824 2872 17876
rect 2924 17864 2930 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 2924 17836 3801 17864
rect 2924 17824 2930 17836
rect 3789 17833 3801 17836
rect 3835 17833 3847 17867
rect 3789 17827 3847 17833
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4157 17867 4215 17873
rect 4157 17864 4169 17867
rect 4120 17836 4169 17864
rect 4120 17824 4126 17836
rect 4157 17833 4169 17836
rect 4203 17833 4215 17867
rect 4157 17827 4215 17833
rect 5767 17867 5825 17873
rect 5767 17833 5779 17867
rect 5813 17864 5825 17867
rect 6362 17864 6368 17876
rect 5813 17836 6368 17864
rect 5813 17833 5825 17836
rect 5767 17827 5825 17833
rect 6362 17824 6368 17836
rect 6420 17824 6426 17876
rect 8205 17867 8263 17873
rect 8205 17833 8217 17867
rect 8251 17864 8263 17867
rect 8478 17864 8484 17876
rect 8251 17836 8484 17864
rect 8251 17833 8263 17836
rect 8205 17827 8263 17833
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 8570 17824 8576 17876
rect 8628 17864 8634 17876
rect 9766 17864 9772 17876
rect 8628 17836 8673 17864
rect 9727 17836 9772 17864
rect 8628 17824 8634 17836
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 10410 17824 10416 17876
rect 10468 17864 10474 17876
rect 10689 17867 10747 17873
rect 10689 17864 10701 17867
rect 10468 17836 10701 17864
rect 10468 17824 10474 17836
rect 10689 17833 10701 17836
rect 10735 17833 10747 17867
rect 11790 17864 11796 17876
rect 11751 17836 11796 17864
rect 10689 17827 10747 17833
rect 11790 17824 11796 17836
rect 11848 17824 11854 17876
rect 14642 17864 14648 17876
rect 14603 17836 14648 17864
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 15654 17864 15660 17876
rect 15615 17836 15660 17864
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 17497 17867 17555 17873
rect 17497 17864 17509 17867
rect 17276 17836 17509 17864
rect 17276 17824 17282 17836
rect 17497 17833 17509 17836
rect 17543 17833 17555 17867
rect 17497 17827 17555 17833
rect 17678 17824 17684 17876
rect 17736 17864 17742 17876
rect 18325 17867 18383 17873
rect 18325 17864 18337 17867
rect 17736 17836 18337 17864
rect 17736 17824 17742 17836
rect 18325 17833 18337 17836
rect 18371 17833 18383 17867
rect 19334 17864 19340 17876
rect 19295 17836 19340 17864
rect 18325 17827 18383 17833
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 19444 17836 19717 17864
rect 7742 17796 7748 17808
rect 7392 17768 7748 17796
rect 3786 17688 3792 17740
rect 3844 17728 3850 17740
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 3844 17700 4077 17728
rect 3844 17688 3850 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 4614 17728 4620 17740
rect 4575 17700 4620 17728
rect 4065 17691 4123 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 5258 17688 5264 17740
rect 5316 17728 5322 17740
rect 7392 17737 7420 17768
rect 7742 17756 7748 17768
rect 7800 17756 7806 17808
rect 12802 17796 12808 17808
rect 11992 17768 12808 17796
rect 11992 17740 12020 17768
rect 12802 17756 12808 17768
rect 12860 17756 12866 17808
rect 5664 17731 5722 17737
rect 5664 17728 5676 17731
rect 5316 17700 5676 17728
rect 5316 17688 5322 17700
rect 5664 17697 5676 17700
rect 5710 17697 5722 17731
rect 5664 17691 5722 17697
rect 7377 17731 7435 17737
rect 7377 17697 7389 17731
rect 7423 17697 7435 17731
rect 7558 17728 7564 17740
rect 7519 17700 7564 17728
rect 7377 17691 7435 17697
rect 7558 17688 7564 17700
rect 7616 17688 7622 17740
rect 9950 17728 9956 17740
rect 9911 17700 9956 17728
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 10134 17728 10140 17740
rect 10095 17700 10140 17728
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 11974 17728 11980 17740
rect 11887 17700 11980 17728
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 12158 17728 12164 17740
rect 12119 17700 12164 17728
rect 12158 17688 12164 17700
rect 12216 17728 12222 17740
rect 12713 17731 12771 17737
rect 12713 17728 12725 17731
rect 12216 17700 12725 17728
rect 12216 17688 12222 17700
rect 12713 17697 12725 17700
rect 12759 17728 12771 17731
rect 12894 17728 12900 17740
rect 12759 17700 12900 17728
rect 12759 17697 12771 17700
rect 12713 17691 12771 17697
rect 12894 17688 12900 17700
rect 12952 17688 12958 17740
rect 13538 17728 13544 17740
rect 13499 17700 13544 17728
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 14093 17731 14151 17737
rect 14093 17697 14105 17731
rect 14139 17728 14151 17731
rect 14182 17728 14188 17740
rect 14139 17700 14188 17728
rect 14139 17697 14151 17700
rect 14093 17691 14151 17697
rect 14182 17688 14188 17700
rect 14240 17728 14246 17740
rect 14660 17728 14688 17824
rect 18874 17756 18880 17808
rect 18932 17796 18938 17808
rect 19444 17796 19472 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 19705 17827 19763 17833
rect 22833 17867 22891 17873
rect 22833 17833 22845 17867
rect 22879 17864 22891 17867
rect 24673 17867 24731 17873
rect 24673 17864 24685 17867
rect 22879 17836 24685 17864
rect 22879 17833 22891 17836
rect 22833 17827 22891 17833
rect 24673 17833 24685 17836
rect 24719 17864 24731 17867
rect 25130 17864 25136 17876
rect 24719 17836 25136 17864
rect 24719 17833 24731 17836
rect 24673 17827 24731 17833
rect 25130 17824 25136 17836
rect 25188 17824 25194 17876
rect 25314 17864 25320 17876
rect 25275 17836 25320 17864
rect 25314 17824 25320 17836
rect 25372 17824 25378 17876
rect 25406 17824 25412 17876
rect 25464 17864 25470 17876
rect 25869 17867 25927 17873
rect 25869 17864 25881 17867
rect 25464 17836 25881 17864
rect 25464 17824 25470 17836
rect 25869 17833 25881 17836
rect 25915 17833 25927 17867
rect 25869 17827 25927 17833
rect 27709 17867 27767 17873
rect 27709 17833 27721 17867
rect 27755 17864 27767 17867
rect 28442 17864 28448 17876
rect 27755 17836 28448 17864
rect 27755 17833 27767 17836
rect 27709 17827 27767 17833
rect 28442 17824 28448 17836
rect 28500 17864 28506 17876
rect 29365 17867 29423 17873
rect 29365 17864 29377 17867
rect 28500 17836 29377 17864
rect 28500 17824 28506 17836
rect 21082 17796 21088 17808
rect 18932 17768 19472 17796
rect 21043 17768 21088 17796
rect 18932 17756 18938 17768
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 23198 17796 23204 17808
rect 22664 17768 23204 17796
rect 14240 17700 14688 17728
rect 14240 17688 14246 17700
rect 16850 17688 16856 17740
rect 16908 17728 16914 17740
rect 17037 17731 17095 17737
rect 17037 17728 17049 17731
rect 16908 17700 17049 17728
rect 16908 17688 16914 17700
rect 17037 17697 17049 17700
rect 17083 17728 17095 17731
rect 17862 17728 17868 17740
rect 17083 17700 17868 17728
rect 17083 17697 17095 17700
rect 17037 17691 17095 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 18049 17731 18107 17737
rect 18049 17728 18061 17731
rect 18012 17700 18061 17728
rect 18012 17688 18018 17700
rect 18049 17697 18061 17700
rect 18095 17697 18107 17731
rect 18049 17691 18107 17697
rect 18233 17731 18291 17737
rect 18233 17697 18245 17731
rect 18279 17728 18291 17731
rect 18506 17728 18512 17740
rect 18279 17700 18512 17728
rect 18279 17697 18291 17700
rect 18233 17691 18291 17697
rect 18506 17688 18512 17700
rect 18564 17688 18570 17740
rect 19426 17728 19432 17740
rect 19387 17700 19432 17728
rect 19426 17688 19432 17700
rect 19484 17688 19490 17740
rect 19610 17728 19616 17740
rect 19571 17700 19616 17728
rect 19610 17688 19616 17700
rect 19668 17688 19674 17740
rect 22664 17737 22692 17768
rect 23198 17756 23204 17768
rect 23256 17756 23262 17808
rect 24762 17756 24768 17808
rect 24820 17796 24826 17808
rect 27065 17799 27123 17805
rect 24820 17768 26188 17796
rect 24820 17756 24826 17768
rect 26160 17740 26188 17768
rect 27065 17765 27077 17799
rect 27111 17796 27123 17799
rect 27154 17796 27160 17808
rect 27111 17768 27160 17796
rect 27111 17765 27123 17768
rect 27065 17759 27123 17765
rect 27154 17756 27160 17768
rect 27212 17756 27218 17808
rect 28736 17805 28764 17836
rect 29365 17833 29377 17836
rect 29411 17864 29423 17867
rect 29546 17864 29552 17876
rect 29411 17836 29552 17864
rect 29411 17833 29423 17836
rect 29365 17827 29423 17833
rect 29546 17824 29552 17836
rect 29604 17824 29610 17876
rect 31018 17864 31024 17876
rect 30979 17836 31024 17864
rect 31018 17824 31024 17836
rect 31076 17824 31082 17876
rect 31478 17864 31484 17876
rect 31439 17836 31484 17864
rect 31478 17824 31484 17836
rect 31536 17824 31542 17876
rect 31846 17864 31852 17876
rect 31759 17836 31852 17864
rect 31846 17824 31852 17836
rect 31904 17864 31910 17876
rect 32582 17864 32588 17876
rect 31904 17836 32588 17864
rect 31904 17824 31910 17836
rect 32582 17824 32588 17836
rect 32640 17864 32646 17876
rect 32769 17867 32827 17873
rect 32769 17864 32781 17867
rect 32640 17836 32781 17864
rect 32640 17824 32646 17836
rect 32769 17833 32781 17836
rect 32815 17833 32827 17867
rect 32769 17827 32827 17833
rect 35161 17867 35219 17873
rect 35161 17833 35173 17867
rect 35207 17864 35219 17867
rect 35250 17864 35256 17876
rect 35207 17836 35256 17864
rect 35207 17833 35219 17836
rect 35161 17827 35219 17833
rect 35250 17824 35256 17836
rect 35308 17824 35314 17876
rect 35802 17824 35808 17876
rect 35860 17864 35866 17876
rect 35897 17867 35955 17873
rect 35897 17864 35909 17867
rect 35860 17836 35909 17864
rect 35860 17824 35866 17836
rect 35897 17833 35909 17836
rect 35943 17833 35955 17867
rect 37918 17864 37924 17876
rect 37879 17836 37924 17864
rect 35897 17827 35955 17833
rect 37918 17824 37924 17836
rect 37976 17824 37982 17876
rect 40126 17864 40132 17876
rect 38672 17836 40132 17864
rect 28721 17799 28779 17805
rect 28721 17765 28733 17799
rect 28767 17765 28779 17799
rect 28721 17759 28779 17765
rect 28902 17756 28908 17808
rect 28960 17796 28966 17808
rect 28960 17768 33134 17796
rect 28960 17756 28966 17768
rect 22649 17731 22707 17737
rect 22649 17697 22661 17731
rect 22695 17697 22707 17731
rect 22649 17691 22707 17697
rect 23569 17731 23627 17737
rect 23569 17697 23581 17731
rect 23615 17728 23627 17731
rect 23661 17731 23719 17737
rect 23661 17728 23673 17731
rect 23615 17700 23673 17728
rect 23615 17697 23627 17700
rect 23569 17691 23627 17697
rect 23661 17697 23673 17700
rect 23707 17728 23719 17731
rect 25222 17728 25228 17740
rect 23707 17700 25228 17728
rect 23707 17697 23719 17700
rect 23661 17691 23719 17697
rect 25222 17688 25228 17700
rect 25280 17728 25286 17740
rect 25409 17731 25467 17737
rect 25409 17728 25421 17731
rect 25280 17700 25421 17728
rect 25280 17688 25286 17700
rect 25409 17697 25421 17700
rect 25455 17697 25467 17731
rect 25409 17691 25467 17697
rect 26142 17688 26148 17740
rect 26200 17728 26206 17740
rect 26510 17728 26516 17740
rect 26200 17700 26516 17728
rect 26200 17688 26206 17700
rect 26510 17688 26516 17700
rect 26568 17688 26574 17740
rect 26697 17731 26755 17737
rect 26697 17697 26709 17731
rect 26743 17728 26755 17731
rect 26786 17728 26792 17740
rect 26743 17700 26792 17728
rect 26743 17697 26755 17700
rect 26697 17691 26755 17697
rect 26786 17688 26792 17700
rect 26844 17688 26850 17740
rect 27890 17688 27896 17740
rect 27948 17728 27954 17740
rect 28077 17731 28135 17737
rect 28077 17728 28089 17731
rect 27948 17700 28089 17728
rect 27948 17688 27954 17700
rect 28077 17697 28089 17700
rect 28123 17697 28135 17731
rect 29638 17728 29644 17740
rect 29599 17700 29644 17728
rect 28077 17691 28135 17697
rect 29638 17688 29644 17700
rect 29696 17688 29702 17740
rect 30006 17728 30012 17740
rect 29967 17700 30012 17728
rect 30006 17688 30012 17700
rect 30064 17688 30070 17740
rect 32306 17728 32312 17740
rect 32267 17700 32312 17728
rect 32306 17688 32312 17700
rect 32364 17688 32370 17740
rect 33106 17728 33134 17768
rect 34698 17756 34704 17808
rect 34756 17796 34762 17808
rect 38672 17796 38700 17836
rect 40126 17824 40132 17836
rect 40184 17824 40190 17876
rect 40405 17867 40463 17873
rect 40405 17833 40417 17867
rect 40451 17864 40463 17867
rect 40494 17864 40500 17876
rect 40451 17836 40500 17864
rect 40451 17833 40463 17836
rect 40405 17827 40463 17833
rect 40494 17824 40500 17836
rect 40552 17864 40558 17876
rect 41141 17867 41199 17873
rect 41141 17864 41153 17867
rect 40552 17836 41153 17864
rect 40552 17824 40558 17836
rect 41141 17833 41153 17836
rect 41187 17833 41199 17867
rect 41141 17827 41199 17833
rect 42334 17824 42340 17876
rect 42392 17864 42398 17876
rect 42613 17867 42671 17873
rect 42613 17864 42625 17867
rect 42392 17836 42625 17864
rect 42392 17824 42398 17836
rect 42613 17833 42625 17836
rect 42659 17833 42671 17867
rect 42613 17827 42671 17833
rect 34756 17768 38700 17796
rect 34756 17756 34762 17768
rect 33410 17728 33416 17740
rect 33106 17700 33416 17728
rect 33410 17688 33416 17700
rect 33468 17728 33474 17740
rect 33597 17731 33655 17737
rect 33597 17728 33609 17731
rect 33468 17700 33609 17728
rect 33468 17688 33474 17700
rect 33597 17697 33609 17700
rect 33643 17697 33655 17731
rect 33778 17728 33784 17740
rect 33739 17700 33784 17728
rect 33597 17691 33655 17697
rect 7009 17663 7067 17669
rect 7009 17629 7021 17663
rect 7055 17660 7067 17663
rect 7576 17660 7604 17688
rect 7742 17660 7748 17672
rect 7055 17632 7604 17660
rect 7703 17632 7748 17660
rect 7055 17629 7067 17632
rect 7009 17623 7067 17629
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 14274 17660 14280 17672
rect 14235 17632 14280 17660
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 15286 17660 15292 17672
rect 15247 17632 15292 17660
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 20346 17620 20352 17672
rect 20404 17660 20410 17672
rect 20990 17660 20996 17672
rect 20404 17632 20996 17660
rect 20404 17620 20410 17632
rect 20990 17620 20996 17632
rect 21048 17620 21054 17672
rect 21174 17620 21180 17672
rect 21232 17660 21238 17672
rect 21269 17663 21327 17669
rect 21269 17660 21281 17663
rect 21232 17632 21281 17660
rect 21232 17620 21238 17632
rect 21269 17629 21281 17632
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 23201 17663 23259 17669
rect 23201 17629 23213 17663
rect 23247 17660 23259 17663
rect 24026 17660 24032 17672
rect 23247 17632 24032 17660
rect 23247 17629 23259 17632
rect 23201 17623 23259 17629
rect 24026 17620 24032 17632
rect 24084 17620 24090 17672
rect 30098 17620 30104 17672
rect 30156 17660 30162 17672
rect 30285 17663 30343 17669
rect 30285 17660 30297 17663
rect 30156 17632 30297 17660
rect 30156 17620 30162 17632
rect 30285 17629 30297 17632
rect 30331 17660 30343 17663
rect 30561 17663 30619 17669
rect 30561 17660 30573 17663
rect 30331 17632 30573 17660
rect 30331 17629 30343 17632
rect 30285 17623 30343 17629
rect 30561 17629 30573 17632
rect 30607 17629 30619 17663
rect 33612 17660 33640 17691
rect 33778 17688 33784 17700
rect 33836 17688 33842 17740
rect 35452 17737 35480 17768
rect 39206 17756 39212 17808
rect 39264 17796 39270 17808
rect 39264 17768 40632 17796
rect 39264 17756 39270 17768
rect 35161 17731 35219 17737
rect 35161 17697 35173 17731
rect 35207 17728 35219 17731
rect 35437 17731 35495 17737
rect 35207 17700 35388 17728
rect 35207 17697 35219 17700
rect 35161 17691 35219 17697
rect 35360 17672 35388 17700
rect 35437 17697 35449 17731
rect 35483 17697 35495 17731
rect 35437 17691 35495 17697
rect 36262 17688 36268 17740
rect 36320 17728 36326 17740
rect 36484 17731 36542 17737
rect 36484 17728 36496 17731
rect 36320 17700 36496 17728
rect 36320 17688 36326 17700
rect 36484 17697 36496 17700
rect 36530 17697 36542 17731
rect 36484 17691 36542 17697
rect 38378 17688 38384 17740
rect 38436 17728 38442 17740
rect 38565 17731 38623 17737
rect 38565 17728 38577 17731
rect 38436 17700 38577 17728
rect 38436 17688 38442 17700
rect 38565 17697 38577 17700
rect 38611 17728 38623 17731
rect 38838 17728 38844 17740
rect 38611 17700 38844 17728
rect 38611 17697 38623 17700
rect 38565 17691 38623 17697
rect 38838 17688 38844 17700
rect 38896 17688 38902 17740
rect 39117 17731 39175 17737
rect 39117 17697 39129 17731
rect 39163 17728 39175 17731
rect 39482 17728 39488 17740
rect 39163 17700 39488 17728
rect 39163 17697 39175 17700
rect 39117 17691 39175 17697
rect 39482 17688 39488 17700
rect 39540 17688 39546 17740
rect 40034 17688 40040 17740
rect 40092 17728 40098 17740
rect 40604 17737 40632 17768
rect 40129 17731 40187 17737
rect 40129 17728 40141 17731
rect 40092 17700 40141 17728
rect 40092 17688 40098 17700
rect 40129 17697 40141 17700
rect 40175 17697 40187 17731
rect 40129 17691 40187 17697
rect 40589 17731 40647 17737
rect 40589 17697 40601 17731
rect 40635 17697 40647 17731
rect 40589 17691 40647 17697
rect 41760 17731 41818 17737
rect 41760 17697 41772 17731
rect 41806 17728 41818 17731
rect 41966 17728 41972 17740
rect 41806 17700 41972 17728
rect 41806 17697 41818 17700
rect 41760 17691 41818 17697
rect 41966 17688 41972 17700
rect 42024 17688 42030 17740
rect 42337 17731 42395 17737
rect 42337 17697 42349 17731
rect 42383 17728 42395 17731
rect 42426 17728 42432 17740
rect 42383 17700 42432 17728
rect 42383 17697 42395 17700
rect 42337 17691 42395 17697
rect 42426 17688 42432 17700
rect 42484 17688 42490 17740
rect 34057 17663 34115 17669
rect 33612 17632 34008 17660
rect 30561 17623 30619 17629
rect 12710 17552 12716 17604
rect 12768 17592 12774 17604
rect 17221 17595 17279 17601
rect 17221 17592 17233 17595
rect 12768 17564 17233 17592
rect 12768 17552 12774 17564
rect 17221 17561 17233 17564
rect 17267 17561 17279 17595
rect 17221 17555 17279 17561
rect 18230 17552 18236 17604
rect 18288 17592 18294 17604
rect 19334 17592 19340 17604
rect 18288 17564 19340 17592
rect 18288 17552 18294 17564
rect 19334 17552 19340 17564
rect 19392 17592 19398 17604
rect 24121 17595 24179 17601
rect 24121 17592 24133 17595
rect 19392 17564 24133 17592
rect 19392 17552 19398 17564
rect 24121 17561 24133 17564
rect 24167 17561 24179 17595
rect 24121 17555 24179 17561
rect 25593 17595 25651 17601
rect 25593 17561 25605 17595
rect 25639 17592 25651 17595
rect 26237 17595 26295 17601
rect 26237 17592 26249 17595
rect 25639 17564 26249 17592
rect 25639 17561 25651 17564
rect 25593 17555 25651 17561
rect 26237 17561 26249 17564
rect 26283 17592 26295 17595
rect 26602 17592 26608 17604
rect 26283 17564 26608 17592
rect 26283 17561 26295 17564
rect 26237 17555 26295 17561
rect 26602 17552 26608 17564
rect 26660 17552 26666 17604
rect 30926 17552 30932 17604
rect 30984 17592 30990 17604
rect 33980 17592 34008 17632
rect 34057 17629 34069 17663
rect 34103 17660 34115 17663
rect 35250 17660 35256 17672
rect 34103 17632 35256 17660
rect 34103 17629 34115 17632
rect 34057 17623 34115 17629
rect 35250 17620 35256 17632
rect 35308 17620 35314 17672
rect 35342 17620 35348 17672
rect 35400 17660 35406 17672
rect 37550 17660 37556 17672
rect 35400 17632 37556 17660
rect 35400 17620 35406 17632
rect 37550 17620 37556 17632
rect 37608 17620 37614 17672
rect 39301 17663 39359 17669
rect 39301 17629 39313 17663
rect 39347 17660 39359 17663
rect 42058 17660 42064 17672
rect 39347 17632 42064 17660
rect 39347 17629 39359 17632
rect 39301 17623 39359 17629
rect 42058 17620 42064 17632
rect 42116 17620 42122 17672
rect 38378 17592 38384 17604
rect 30984 17564 33870 17592
rect 33980 17564 38384 17592
rect 30984 17552 30990 17564
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 16209 17527 16267 17533
rect 16209 17524 16221 17527
rect 14700 17496 16221 17524
rect 14700 17484 14706 17496
rect 16209 17493 16221 17496
rect 16255 17493 16267 17527
rect 16209 17487 16267 17493
rect 18138 17484 18144 17536
rect 18196 17524 18202 17536
rect 22002 17524 22008 17536
rect 18196 17496 22008 17524
rect 18196 17484 18202 17496
rect 22002 17484 22008 17496
rect 22060 17484 22066 17536
rect 23198 17484 23204 17536
rect 23256 17524 23262 17536
rect 23808 17527 23866 17533
rect 23808 17524 23820 17527
rect 23256 17496 23820 17524
rect 23256 17484 23262 17496
rect 23808 17493 23820 17496
rect 23854 17493 23866 17527
rect 23934 17524 23940 17536
rect 23895 17496 23940 17524
rect 23808 17487 23866 17493
rect 23934 17484 23940 17496
rect 23992 17484 23998 17536
rect 32490 17524 32496 17536
rect 32451 17496 32496 17524
rect 32490 17484 32496 17496
rect 32548 17484 32554 17536
rect 33842 17524 33870 17564
rect 38378 17552 38384 17564
rect 38436 17552 38442 17604
rect 34330 17524 34336 17536
rect 33842 17496 34336 17524
rect 34330 17484 34336 17496
rect 34388 17484 34394 17536
rect 36587 17527 36645 17533
rect 36587 17493 36599 17527
rect 36633 17524 36645 17527
rect 36722 17524 36728 17536
rect 36633 17496 36728 17524
rect 36633 17493 36645 17496
rect 36587 17487 36645 17493
rect 36722 17484 36728 17496
rect 36780 17484 36786 17536
rect 36906 17524 36912 17536
rect 36867 17496 36912 17524
rect 36906 17484 36912 17496
rect 36964 17484 36970 17536
rect 37366 17484 37372 17536
rect 37424 17524 37430 17536
rect 41831 17527 41889 17533
rect 41831 17524 41843 17527
rect 37424 17496 41843 17524
rect 37424 17484 37430 17496
rect 41831 17493 41843 17496
rect 41877 17493 41889 17527
rect 41831 17487 41889 17493
rect 1104 17434 48852 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 48852 17434
rect 1104 17360 48852 17382
rect 2958 17280 2964 17332
rect 3016 17320 3022 17332
rect 3605 17323 3663 17329
rect 3605 17320 3617 17323
rect 3016 17292 3617 17320
rect 3016 17280 3022 17292
rect 3605 17289 3617 17292
rect 3651 17320 3663 17323
rect 3786 17320 3792 17332
rect 3651 17292 3792 17320
rect 3651 17289 3663 17292
rect 3605 17283 3663 17289
rect 3786 17280 3792 17292
rect 3844 17280 3850 17332
rect 3970 17320 3976 17332
rect 3931 17292 3976 17320
rect 3970 17280 3976 17292
rect 4028 17280 4034 17332
rect 5258 17280 5264 17332
rect 5316 17320 5322 17332
rect 5537 17323 5595 17329
rect 5537 17320 5549 17323
rect 5316 17292 5549 17320
rect 5316 17280 5322 17292
rect 5537 17289 5549 17292
rect 5583 17289 5595 17323
rect 5537 17283 5595 17289
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 7929 17323 7987 17329
rect 7929 17320 7941 17323
rect 7892 17292 7941 17320
rect 7892 17280 7898 17292
rect 7929 17289 7941 17292
rect 7975 17289 7987 17323
rect 7929 17283 7987 17289
rect 9950 17280 9956 17332
rect 10008 17320 10014 17332
rect 10321 17323 10379 17329
rect 10321 17320 10333 17323
rect 10008 17292 10333 17320
rect 10008 17280 10014 17292
rect 10321 17289 10333 17292
rect 10367 17289 10379 17323
rect 10321 17283 10379 17289
rect 11425 17323 11483 17329
rect 11425 17289 11437 17323
rect 11471 17320 11483 17323
rect 12158 17320 12164 17332
rect 11471 17292 12164 17320
rect 11471 17289 11483 17292
rect 11425 17283 11483 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 13538 17320 13544 17332
rect 13499 17292 13544 17320
rect 13538 17280 13544 17292
rect 13596 17280 13602 17332
rect 14182 17320 14188 17332
rect 14143 17292 14188 17320
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 16206 17280 16212 17332
rect 16264 17320 16270 17332
rect 16393 17323 16451 17329
rect 16393 17320 16405 17323
rect 16264 17292 16405 17320
rect 16264 17280 16270 17292
rect 16393 17289 16405 17292
rect 16439 17289 16451 17323
rect 16850 17320 16856 17332
rect 16811 17292 16856 17320
rect 16393 17283 16451 17289
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 19337 17323 19395 17329
rect 19337 17320 19349 17323
rect 18248 17292 19349 17320
rect 11793 17255 11851 17261
rect 11793 17221 11805 17255
rect 11839 17252 11851 17255
rect 11974 17252 11980 17264
rect 11839 17224 11980 17252
rect 11839 17221 11851 17224
rect 11793 17215 11851 17221
rect 11974 17212 11980 17224
rect 12032 17212 12038 17264
rect 6641 17187 6699 17193
rect 6641 17153 6653 17187
rect 6687 17184 6699 17187
rect 7650 17184 7656 17196
rect 6687 17156 7656 17184
rect 6687 17153 6699 17156
rect 6641 17147 6699 17153
rect 3970 17076 3976 17128
rect 4028 17116 4034 17128
rect 4157 17119 4215 17125
rect 4157 17116 4169 17119
rect 4028 17088 4169 17116
rect 4028 17076 4034 17088
rect 4157 17085 4169 17088
rect 4203 17085 4215 17119
rect 4614 17116 4620 17128
rect 4575 17088 4620 17116
rect 4157 17079 4215 17085
rect 4614 17076 4620 17088
rect 4672 17116 4678 17128
rect 7208 17125 7236 17156
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 12176 17184 12204 17280
rect 15197 17187 15255 17193
rect 12176 17156 12940 17184
rect 5169 17119 5227 17125
rect 5169 17116 5181 17119
rect 4672 17088 5181 17116
rect 4672 17076 4678 17088
rect 5169 17085 5181 17088
rect 5215 17085 5227 17119
rect 5169 17079 5227 17085
rect 5721 17119 5779 17125
rect 5721 17085 5733 17119
rect 5767 17116 5779 17119
rect 7193 17119 7251 17125
rect 5767 17088 6316 17116
rect 5767 17085 5779 17088
rect 5721 17079 5779 17085
rect 4798 17008 4804 17060
rect 4856 17048 4862 17060
rect 4893 17051 4951 17057
rect 4893 17048 4905 17051
rect 4856 17020 4905 17048
rect 4856 17008 4862 17020
rect 4893 17017 4905 17020
rect 4939 17017 4951 17051
rect 4893 17011 4951 17017
rect 3234 16980 3240 16992
rect 3195 16952 3240 16980
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 5184 16980 5212 17079
rect 6288 17057 6316 17088
rect 7193 17085 7205 17119
rect 7239 17085 7251 17119
rect 7193 17079 7251 17085
rect 7469 17119 7527 17125
rect 7469 17085 7481 17119
rect 7515 17116 7527 17119
rect 7558 17116 7564 17128
rect 7515 17088 7564 17116
rect 7515 17085 7527 17088
rect 7469 17079 7527 17085
rect 6273 17051 6331 17057
rect 6273 17017 6285 17051
rect 6319 17048 6331 17051
rect 7484 17048 7512 17079
rect 7558 17076 7564 17088
rect 7616 17116 7622 17128
rect 9217 17119 9275 17125
rect 7616 17088 8892 17116
rect 7616 17076 7622 17088
rect 7650 17048 7656 17060
rect 6319 17020 7512 17048
rect 7611 17020 7656 17048
rect 6319 17017 6331 17020
rect 6273 17011 6331 17017
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 8864 17057 8892 17088
rect 9217 17085 9229 17119
rect 9263 17116 9275 17119
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 9263 17088 9597 17116
rect 9263 17085 9275 17088
rect 9217 17079 9275 17085
rect 9585 17085 9597 17088
rect 9631 17116 9643 17119
rect 9674 17116 9680 17128
rect 9631 17088 9680 17116
rect 9631 17085 9643 17088
rect 9585 17079 9643 17085
rect 9674 17076 9680 17088
rect 9732 17076 9738 17128
rect 9861 17119 9919 17125
rect 9861 17085 9873 17119
rect 9907 17085 9919 17119
rect 10778 17116 10784 17128
rect 10691 17088 10784 17116
rect 9861 17079 9919 17085
rect 8849 17051 8907 17057
rect 8849 17017 8861 17051
rect 8895 17048 8907 17051
rect 9398 17048 9404 17060
rect 8895 17020 9404 17048
rect 8895 17017 8907 17020
rect 8849 17011 8907 17017
rect 9398 17008 9404 17020
rect 9456 17048 9462 17060
rect 9876 17048 9904 17079
rect 10778 17076 10784 17088
rect 10836 17116 10842 17128
rect 10908 17119 10966 17125
rect 10908 17116 10920 17119
rect 10836 17088 10920 17116
rect 10836 17076 10842 17088
rect 10908 17085 10920 17088
rect 10954 17085 10966 17119
rect 10908 17079 10966 17085
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 12912 17125 12940 17156
rect 15197 17153 15209 17187
rect 15243 17184 15255 17187
rect 16224 17184 16252 17280
rect 18248 17184 18276 17292
rect 19337 17289 19349 17292
rect 19383 17320 19395 17323
rect 19426 17320 19432 17332
rect 19383 17292 19432 17320
rect 19383 17289 19395 17292
rect 19337 17283 19395 17289
rect 19426 17280 19432 17292
rect 19484 17280 19490 17332
rect 21082 17280 21088 17332
rect 21140 17320 21146 17332
rect 21453 17323 21511 17329
rect 21453 17320 21465 17323
rect 21140 17292 21465 17320
rect 21140 17280 21146 17292
rect 21453 17289 21465 17292
rect 21499 17289 21511 17323
rect 21453 17283 21511 17289
rect 22738 17280 22744 17332
rect 22796 17320 22802 17332
rect 23198 17320 23204 17332
rect 22796 17292 23204 17320
rect 22796 17280 22802 17292
rect 23198 17280 23204 17292
rect 23256 17320 23262 17332
rect 23477 17323 23535 17329
rect 23477 17320 23489 17323
rect 23256 17292 23489 17320
rect 23256 17280 23262 17292
rect 23477 17289 23489 17292
rect 23523 17320 23535 17323
rect 24581 17323 24639 17329
rect 24581 17320 24593 17323
rect 23523 17292 24593 17320
rect 23523 17289 23535 17292
rect 23477 17283 23535 17289
rect 24581 17289 24593 17292
rect 24627 17289 24639 17323
rect 24581 17283 24639 17289
rect 25222 17280 25228 17332
rect 25280 17320 25286 17332
rect 25501 17323 25559 17329
rect 25501 17320 25513 17323
rect 25280 17292 25513 17320
rect 25280 17280 25286 17292
rect 25501 17289 25513 17292
rect 25547 17289 25559 17323
rect 25501 17283 25559 17289
rect 26237 17323 26295 17329
rect 26237 17289 26249 17323
rect 26283 17320 26295 17323
rect 26786 17320 26792 17332
rect 26283 17292 26792 17320
rect 26283 17289 26295 17292
rect 26237 17283 26295 17289
rect 26786 17280 26792 17292
rect 26844 17280 26850 17332
rect 28626 17320 28632 17332
rect 28587 17292 28632 17320
rect 28626 17280 28632 17292
rect 28684 17280 28690 17332
rect 29089 17323 29147 17329
rect 29089 17289 29101 17323
rect 29135 17320 29147 17323
rect 29270 17320 29276 17332
rect 29135 17292 29276 17320
rect 29135 17289 29147 17292
rect 29089 17283 29147 17289
rect 29270 17280 29276 17292
rect 29328 17280 29334 17332
rect 32490 17280 32496 17332
rect 32548 17320 32554 17332
rect 33134 17320 33140 17332
rect 32548 17292 33140 17320
rect 32548 17280 32554 17292
rect 33134 17280 33140 17292
rect 33192 17320 33198 17332
rect 33321 17323 33379 17329
rect 33321 17320 33333 17323
rect 33192 17292 33333 17320
rect 33192 17280 33198 17292
rect 33321 17289 33333 17292
rect 33367 17320 33379 17323
rect 33778 17320 33784 17332
rect 33367 17292 33784 17320
rect 33367 17289 33379 17292
rect 33321 17283 33379 17289
rect 33778 17280 33784 17292
rect 33836 17280 33842 17332
rect 34698 17320 34704 17332
rect 34659 17292 34704 17320
rect 34698 17280 34704 17292
rect 34756 17280 34762 17332
rect 34790 17280 34796 17332
rect 34848 17320 34854 17332
rect 35161 17323 35219 17329
rect 35161 17320 35173 17323
rect 34848 17292 35173 17320
rect 34848 17280 34854 17292
rect 35161 17289 35173 17292
rect 35207 17320 35219 17323
rect 35342 17320 35348 17332
rect 35207 17292 35348 17320
rect 35207 17289 35219 17292
rect 35161 17283 35219 17289
rect 35342 17280 35348 17292
rect 35400 17280 35406 17332
rect 36280 17292 40678 17320
rect 36280 17264 36308 17292
rect 19150 17212 19156 17264
rect 19208 17252 19214 17264
rect 19567 17255 19625 17261
rect 19567 17252 19579 17255
rect 19208 17224 19579 17252
rect 19208 17212 19214 17224
rect 19567 17221 19579 17224
rect 19613 17221 19625 17255
rect 19567 17215 19625 17221
rect 20990 17212 20996 17264
rect 21048 17252 21054 17264
rect 21821 17255 21879 17261
rect 21821 17252 21833 17255
rect 21048 17224 21833 17252
rect 21048 17212 21054 17224
rect 21821 17221 21833 17224
rect 21867 17221 21879 17255
rect 23934 17252 23940 17264
rect 23847 17224 23940 17252
rect 21821 17215 21879 17221
rect 23934 17212 23940 17224
rect 23992 17252 23998 17264
rect 24762 17252 24768 17264
rect 23992 17224 24768 17252
rect 23992 17212 23998 17224
rect 24762 17212 24768 17224
rect 24820 17212 24826 17264
rect 32306 17212 32312 17264
rect 32364 17252 32370 17264
rect 32861 17255 32919 17261
rect 32861 17252 32873 17255
rect 32364 17224 32873 17252
rect 32364 17212 32370 17224
rect 32861 17221 32873 17224
rect 32907 17221 32919 17255
rect 32861 17215 32919 17221
rect 32950 17212 32956 17264
rect 33008 17252 33014 17264
rect 33045 17255 33103 17261
rect 33045 17252 33057 17255
rect 33008 17224 33057 17252
rect 33008 17212 33014 17224
rect 33045 17221 33057 17224
rect 33091 17252 33103 17255
rect 36262 17252 36268 17264
rect 33091 17224 36268 17252
rect 33091 17221 33103 17224
rect 33045 17215 33103 17221
rect 36262 17212 36268 17224
rect 36320 17212 36326 17264
rect 36630 17212 36636 17264
rect 36688 17252 36694 17264
rect 37829 17255 37887 17261
rect 37829 17252 37841 17255
rect 36688 17224 37841 17252
rect 36688 17212 36694 17224
rect 37829 17221 37841 17224
rect 37875 17252 37887 17255
rect 38194 17252 38200 17264
rect 37875 17224 38200 17252
rect 37875 17221 37887 17224
rect 37829 17215 37887 17221
rect 38194 17212 38200 17224
rect 38252 17212 38258 17264
rect 38838 17212 38844 17264
rect 38896 17252 38902 17264
rect 39025 17255 39083 17261
rect 39025 17252 39037 17255
rect 38896 17224 39037 17252
rect 38896 17212 38902 17224
rect 39025 17221 39037 17224
rect 39071 17221 39083 17255
rect 39025 17215 39083 17221
rect 39206 17212 39212 17264
rect 39264 17252 39270 17264
rect 39761 17255 39819 17261
rect 39761 17252 39773 17255
rect 39264 17224 39773 17252
rect 39264 17212 39270 17224
rect 39761 17221 39773 17224
rect 39807 17221 39819 17255
rect 39761 17215 39819 17221
rect 40034 17212 40040 17264
rect 40092 17252 40098 17264
rect 40129 17255 40187 17261
rect 40129 17252 40141 17255
rect 40092 17224 40141 17252
rect 40092 17212 40098 17224
rect 40129 17221 40141 17224
rect 40175 17221 40187 17255
rect 40129 17215 40187 17221
rect 20530 17184 20536 17196
rect 15243 17156 16252 17184
rect 18064 17156 18276 17184
rect 20491 17156 20536 17184
rect 15243 17153 15255 17156
rect 15197 17147 15255 17153
rect 12161 17119 12219 17125
rect 12161 17116 12173 17119
rect 11940 17088 12173 17116
rect 11940 17076 11946 17088
rect 12161 17085 12173 17088
rect 12207 17116 12219 17119
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12207 17088 12449 17116
rect 12207 17085 12219 17088
rect 12161 17079 12219 17085
rect 12437 17085 12449 17088
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17116 12955 17119
rect 12986 17116 12992 17128
rect 12943 17088 12992 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 12986 17076 12992 17088
rect 13044 17076 13050 17128
rect 13998 17116 14004 17128
rect 13096 17088 14004 17116
rect 10134 17048 10140 17060
rect 9456 17020 10140 17048
rect 9456 17008 9462 17020
rect 10134 17008 10140 17020
rect 10192 17048 10198 17060
rect 13096 17048 13124 17088
rect 13998 17076 14004 17088
rect 14056 17076 14062 17128
rect 18064 17125 18092 17156
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 21174 17184 21180 17196
rect 21135 17156 21180 17184
rect 21174 17144 21180 17156
rect 21232 17144 21238 17196
rect 26694 17184 26700 17196
rect 26607 17156 26700 17184
rect 16945 17119 17003 17125
rect 16945 17085 16957 17119
rect 16991 17116 17003 17119
rect 18049 17119 18107 17125
rect 16991 17088 17540 17116
rect 16991 17085 17003 17088
rect 16945 17079 17003 17085
rect 15518 17051 15576 17057
rect 15518 17048 15530 17051
rect 10192 17020 13124 17048
rect 15028 17020 15530 17048
rect 10192 17008 10198 17020
rect 5905 16983 5963 16989
rect 5905 16980 5917 16983
rect 5184 16952 5917 16980
rect 5905 16949 5917 16952
rect 5951 16980 5963 16983
rect 6086 16980 6092 16992
rect 5951 16952 6092 16980
rect 5951 16949 5963 16952
rect 5905 16943 5963 16949
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 9582 16980 9588 16992
rect 9543 16952 9588 16980
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 10870 16940 10876 16992
rect 10928 16980 10934 16992
rect 11011 16983 11069 16989
rect 11011 16980 11023 16983
rect 10928 16952 11023 16980
rect 10928 16940 10934 16952
rect 11011 16949 11023 16952
rect 11057 16949 11069 16983
rect 12526 16980 12532 16992
rect 12487 16952 12532 16980
rect 11011 16943 11069 16949
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 14550 16940 14556 16992
rect 14608 16980 14614 16992
rect 15028 16989 15056 17020
rect 15518 17017 15530 17020
rect 15564 17048 15576 17051
rect 15654 17048 15660 17060
rect 15564 17020 15660 17048
rect 15564 17017 15576 17020
rect 15518 17011 15576 17017
rect 15654 17008 15660 17020
rect 15712 17008 15718 17060
rect 17512 16992 17540 17088
rect 18049 17085 18061 17119
rect 18095 17085 18107 17119
rect 18230 17116 18236 17128
rect 18191 17088 18236 17116
rect 18049 17079 18107 17085
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 19496 17119 19554 17125
rect 19496 17085 19508 17119
rect 19542 17116 19554 17119
rect 19886 17116 19892 17128
rect 19542 17088 19892 17116
rect 19542 17085 19554 17088
rect 19496 17079 19554 17085
rect 19886 17076 19892 17088
rect 19944 17076 19950 17128
rect 22332 17119 22390 17125
rect 22332 17085 22344 17119
rect 22378 17116 22390 17119
rect 22830 17116 22836 17128
rect 22378 17088 22836 17116
rect 22378 17085 22390 17088
rect 22332 17079 22390 17085
rect 22830 17076 22836 17088
rect 22888 17076 22894 17128
rect 24486 17116 24492 17128
rect 24447 17088 24492 17116
rect 24486 17076 24492 17088
rect 24544 17116 24550 17128
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24544 17088 25145 17116
rect 24544 17076 24550 17088
rect 25133 17085 25145 17088
rect 25179 17116 25191 17119
rect 26234 17116 26240 17128
rect 25179 17088 26240 17116
rect 25179 17085 25191 17088
rect 25133 17079 25191 17085
rect 26234 17076 26240 17088
rect 26292 17076 26298 17128
rect 26620 17125 26648 17156
rect 26694 17144 26700 17156
rect 26752 17184 26758 17196
rect 29638 17184 29644 17196
rect 26752 17156 29644 17184
rect 26752 17144 26758 17156
rect 29638 17144 29644 17156
rect 29696 17144 29702 17196
rect 30098 17184 30104 17196
rect 30059 17156 30104 17184
rect 30098 17144 30104 17156
rect 30156 17144 30162 17196
rect 31938 17184 31944 17196
rect 31851 17156 31944 17184
rect 31938 17144 31944 17156
rect 31996 17184 32002 17196
rect 33318 17184 33324 17196
rect 31996 17156 33324 17184
rect 31996 17144 32002 17156
rect 33318 17144 33324 17156
rect 33376 17144 33382 17196
rect 35575 17187 35633 17193
rect 35575 17153 35587 17187
rect 35621 17184 35633 17187
rect 36541 17187 36599 17193
rect 36541 17184 36553 17187
rect 35621 17156 36553 17184
rect 35621 17153 35633 17156
rect 35575 17147 35633 17153
rect 36541 17153 36553 17156
rect 36587 17184 36599 17187
rect 36906 17184 36912 17196
rect 36587 17156 36912 17184
rect 36587 17153 36599 17156
rect 36541 17147 36599 17153
rect 36906 17144 36912 17156
rect 36964 17144 36970 17196
rect 38470 17184 38476 17196
rect 38431 17156 38476 17184
rect 38470 17144 38476 17156
rect 38528 17144 38534 17196
rect 26605 17119 26663 17125
rect 26605 17085 26617 17119
rect 26651 17085 26663 17119
rect 26605 17079 26663 17085
rect 26881 17119 26939 17125
rect 26881 17085 26893 17119
rect 26927 17116 26939 17119
rect 27154 17116 27160 17128
rect 26927 17088 27160 17116
rect 26927 17085 26939 17088
rect 26881 17079 26939 17085
rect 27154 17076 27160 17088
rect 27212 17076 27218 17128
rect 28169 17119 28227 17125
rect 28169 17085 28181 17119
rect 28215 17116 28227 17119
rect 28258 17116 28264 17128
rect 28215 17088 28264 17116
rect 28215 17085 28227 17088
rect 28169 17079 28227 17085
rect 28258 17076 28264 17088
rect 28316 17116 28322 17128
rect 29914 17116 29920 17128
rect 28316 17088 29920 17116
rect 28316 17076 28322 17088
rect 29914 17076 29920 17088
rect 29972 17076 29978 17128
rect 32674 17076 32680 17128
rect 32732 17116 32738 17128
rect 33045 17119 33103 17125
rect 33045 17116 33057 17119
rect 32732 17088 33057 17116
rect 32732 17076 32738 17088
rect 33045 17085 33057 17088
rect 33091 17085 33103 17119
rect 33045 17079 33103 17085
rect 33226 17076 33232 17128
rect 33284 17116 33290 17128
rect 33464 17119 33522 17125
rect 33464 17116 33476 17119
rect 33284 17088 33476 17116
rect 33284 17076 33290 17088
rect 33464 17085 33476 17088
rect 33510 17116 33522 17119
rect 40564 17119 40622 17125
rect 33510 17088 34008 17116
rect 33510 17085 33522 17088
rect 33464 17079 33522 17085
rect 19610 17008 19616 17060
rect 19668 17008 19674 17060
rect 20622 17008 20628 17060
rect 20680 17048 20686 17060
rect 22419 17051 22477 17057
rect 20680 17020 20725 17048
rect 20680 17008 20686 17020
rect 22419 17017 22431 17051
rect 22465 17048 22477 17051
rect 24118 17048 24124 17060
rect 22465 17020 24124 17048
rect 22465 17017 22477 17020
rect 22419 17011 22477 17017
rect 24118 17008 24124 17020
rect 24176 17008 24182 17060
rect 24302 17048 24308 17060
rect 24263 17020 24308 17048
rect 24302 17008 24308 17020
rect 24360 17008 24366 17060
rect 26510 17008 26516 17060
rect 26568 17048 26574 17060
rect 27433 17051 27491 17057
rect 27433 17048 27445 17051
rect 26568 17020 27445 17048
rect 26568 17008 26574 17020
rect 27433 17017 27445 17020
rect 27479 17048 27491 17051
rect 28534 17048 28540 17060
rect 27479 17020 28540 17048
rect 27479 17017 27491 17020
rect 27433 17011 27491 17017
rect 28534 17008 28540 17020
rect 28592 17008 28598 17060
rect 30422 17051 30480 17057
rect 30422 17048 30434 17051
rect 30300 17020 30434 17048
rect 14645 16983 14703 16989
rect 14645 16980 14657 16983
rect 14608 16952 14657 16980
rect 14608 16940 14614 16952
rect 14645 16949 14657 16952
rect 14691 16980 14703 16983
rect 15013 16983 15071 16989
rect 15013 16980 15025 16983
rect 14691 16952 15025 16980
rect 14691 16949 14703 16952
rect 14645 16943 14703 16949
rect 15013 16949 15025 16952
rect 15059 16949 15071 16983
rect 16114 16980 16120 16992
rect 16075 16952 16120 16980
rect 15013 16943 15071 16949
rect 16114 16940 16120 16952
rect 16172 16940 16178 16992
rect 16206 16940 16212 16992
rect 16264 16980 16270 16992
rect 17129 16983 17187 16989
rect 17129 16980 17141 16983
rect 16264 16952 17141 16980
rect 16264 16940 16270 16952
rect 17129 16949 17141 16952
rect 17175 16949 17187 16983
rect 17494 16980 17500 16992
rect 17455 16952 17500 16980
rect 17129 16943 17187 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 17862 16980 17868 16992
rect 17823 16952 17868 16980
rect 17862 16940 17868 16952
rect 17920 16940 17926 16992
rect 18322 16980 18328 16992
rect 18283 16952 18328 16980
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 18506 16940 18512 16992
rect 18564 16980 18570 16992
rect 18877 16983 18935 16989
rect 18877 16980 18889 16983
rect 18564 16952 18889 16980
rect 18564 16940 18570 16952
rect 18877 16949 18889 16952
rect 18923 16980 18935 16983
rect 19628 16980 19656 17008
rect 19889 16983 19947 16989
rect 19889 16980 19901 16983
rect 18923 16952 19901 16980
rect 18923 16949 18935 16952
rect 18877 16943 18935 16949
rect 19889 16949 19901 16952
rect 19935 16949 19947 16983
rect 19889 16943 19947 16949
rect 20349 16983 20407 16989
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 20640 16980 20668 17008
rect 30300 16992 30328 17020
rect 30422 17017 30434 17020
rect 30468 17048 30480 17051
rect 31386 17048 31392 17060
rect 30468 17020 31392 17048
rect 30468 17017 30480 17020
rect 30422 17011 30480 17017
rect 31386 17008 31392 17020
rect 31444 17048 31450 17060
rect 31754 17048 31760 17060
rect 31444 17020 31760 17048
rect 31444 17008 31450 17020
rect 31754 17008 31760 17020
rect 31812 17008 31818 17060
rect 32033 17051 32091 17057
rect 32033 17017 32045 17051
rect 32079 17017 32091 17051
rect 32582 17048 32588 17060
rect 32543 17020 32588 17048
rect 32033 17011 32091 17017
rect 26418 16980 26424 16992
rect 20395 16952 20668 16980
rect 26379 16952 26424 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 26418 16940 26424 16952
rect 26476 16940 26482 16992
rect 27890 16940 27896 16992
rect 27948 16980 27954 16992
rect 27985 16983 28043 16989
rect 27985 16980 27997 16983
rect 27948 16952 27997 16980
rect 27948 16940 27954 16952
rect 27985 16949 27997 16952
rect 28031 16949 28043 16983
rect 28350 16980 28356 16992
rect 28311 16952 28356 16980
rect 27985 16943 28043 16949
rect 28350 16940 28356 16952
rect 28408 16940 28414 16992
rect 29638 16980 29644 16992
rect 29599 16952 29644 16980
rect 29638 16940 29644 16952
rect 29696 16940 29702 16992
rect 30009 16983 30067 16989
rect 30009 16949 30021 16983
rect 30055 16980 30067 16983
rect 30282 16980 30288 16992
rect 30055 16952 30288 16980
rect 30055 16949 30067 16952
rect 30009 16943 30067 16949
rect 30282 16940 30288 16952
rect 30340 16940 30346 16992
rect 31021 16983 31079 16989
rect 31021 16949 31033 16983
rect 31067 16980 31079 16983
rect 31665 16983 31723 16989
rect 31665 16980 31677 16983
rect 31067 16952 31677 16980
rect 31067 16949 31079 16952
rect 31021 16943 31079 16949
rect 31665 16949 31677 16952
rect 31711 16980 31723 16983
rect 32048 16980 32076 17011
rect 32582 17008 32588 17020
rect 32640 17008 32646 17060
rect 33551 17051 33609 17057
rect 33551 17048 33563 17051
rect 33106 17020 33563 17048
rect 32306 16980 32312 16992
rect 31711 16952 32312 16980
rect 31711 16949 31723 16952
rect 31665 16943 31723 16949
rect 32306 16940 32312 16952
rect 32364 16940 32370 16992
rect 32950 16940 32956 16992
rect 33008 16980 33014 16992
rect 33106 16980 33134 17020
rect 33551 17017 33563 17020
rect 33597 17017 33609 17051
rect 33551 17011 33609 17017
rect 33980 16989 34008 17088
rect 40564 17085 40576 17119
rect 40610 17085 40622 17119
rect 40650 17116 40678 17292
rect 41966 17280 41972 17332
rect 42024 17320 42030 17332
rect 42337 17323 42395 17329
rect 42337 17320 42349 17323
rect 42024 17292 42349 17320
rect 42024 17280 42030 17292
rect 42337 17289 42349 17292
rect 42383 17289 42395 17323
rect 42337 17283 42395 17289
rect 41544 17119 41602 17125
rect 41544 17116 41556 17119
rect 40650 17088 41556 17116
rect 40564 17079 40622 17085
rect 41544 17085 41556 17088
rect 41590 17116 41602 17119
rect 41969 17119 42027 17125
rect 41969 17116 41981 17119
rect 41590 17088 41981 17116
rect 41590 17085 41602 17088
rect 41544 17079 41602 17085
rect 41969 17085 41981 17088
rect 42015 17085 42027 17119
rect 41969 17079 42027 17085
rect 43140 17119 43198 17125
rect 43140 17085 43152 17119
rect 43186 17116 43198 17119
rect 43530 17116 43536 17128
rect 43186 17088 43536 17116
rect 43186 17085 43198 17088
rect 43140 17079 43198 17085
rect 34330 17008 34336 17060
rect 34388 17048 34394 17060
rect 35345 17051 35403 17057
rect 35345 17048 35357 17051
rect 34388 17020 35357 17048
rect 34388 17008 34394 17020
rect 35345 17017 35357 17020
rect 35391 17048 35403 17051
rect 35986 17048 35992 17060
rect 35391 17020 35992 17048
rect 35391 17017 35403 17020
rect 35345 17011 35403 17017
rect 35986 17008 35992 17020
rect 36044 17008 36050 17060
rect 36630 17048 36636 17060
rect 36591 17020 36636 17048
rect 36630 17008 36636 17020
rect 36688 17008 36694 17060
rect 37182 17048 37188 17060
rect 37143 17020 37188 17048
rect 37182 17008 37188 17020
rect 37240 17008 37246 17060
rect 38105 17051 38163 17057
rect 38105 17048 38117 17051
rect 37476 17020 38117 17048
rect 33008 16952 33134 16980
rect 33965 16983 34023 16989
rect 33008 16940 33014 16952
rect 33965 16949 33977 16983
rect 34011 16980 34023 16983
rect 34606 16980 34612 16992
rect 34011 16952 34612 16980
rect 34011 16949 34023 16952
rect 33965 16943 34023 16949
rect 34606 16940 34612 16952
rect 34664 16940 34670 16992
rect 36446 16940 36452 16992
rect 36504 16980 36510 16992
rect 37476 16989 37504 17020
rect 38105 17017 38117 17020
rect 38151 17017 38163 17051
rect 38105 17011 38163 17017
rect 38194 17008 38200 17060
rect 38252 17048 38258 17060
rect 38252 17020 38297 17048
rect 38252 17008 38258 17020
rect 38562 17008 38568 17060
rect 38620 17048 38626 17060
rect 40579 17048 40607 17079
rect 43530 17076 43536 17088
rect 43588 17076 43594 17128
rect 38620 17020 40816 17048
rect 38620 17008 38626 17020
rect 37461 16983 37519 16989
rect 37461 16980 37473 16983
rect 36504 16952 37473 16980
rect 36504 16940 36510 16952
rect 37461 16949 37473 16952
rect 37507 16949 37519 16983
rect 39482 16980 39488 16992
rect 39443 16952 39488 16980
rect 37461 16943 37519 16949
rect 39482 16940 39488 16952
rect 39540 16940 39546 16992
rect 40310 16940 40316 16992
rect 40368 16980 40374 16992
rect 40635 16983 40693 16989
rect 40635 16980 40647 16983
rect 40368 16952 40647 16980
rect 40368 16940 40374 16952
rect 40635 16949 40647 16952
rect 40681 16949 40693 16983
rect 40788 16980 40816 17020
rect 40862 17008 40868 17060
rect 40920 17048 40926 17060
rect 41647 17051 41705 17057
rect 41647 17048 41659 17051
rect 40920 17020 41659 17048
rect 40920 17008 40926 17020
rect 41647 17017 41659 17020
rect 41693 17017 41705 17051
rect 41647 17011 41705 17017
rect 40957 16983 41015 16989
rect 40957 16980 40969 16983
rect 40788 16952 40969 16980
rect 40635 16943 40693 16949
rect 40957 16949 40969 16952
rect 41003 16980 41015 16983
rect 41138 16980 41144 16992
rect 41003 16952 41144 16980
rect 41003 16949 41015 16952
rect 40957 16943 41015 16949
rect 41138 16940 41144 16952
rect 41196 16940 41202 16992
rect 43211 16983 43269 16989
rect 43211 16949 43223 16983
rect 43257 16980 43269 16983
rect 44082 16980 44088 16992
rect 43257 16952 44088 16980
rect 43257 16949 43269 16952
rect 43211 16943 43269 16949
rect 44082 16940 44088 16952
rect 44140 16940 44146 16992
rect 1104 16890 48852 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 48852 16890
rect 1104 16816 48852 16838
rect 7561 16779 7619 16785
rect 7561 16745 7573 16779
rect 7607 16776 7619 16779
rect 7650 16776 7656 16788
rect 7607 16748 7656 16776
rect 7607 16745 7619 16748
rect 7561 16739 7619 16745
rect 7650 16736 7656 16748
rect 7708 16736 7714 16788
rect 9398 16776 9404 16788
rect 9359 16748 9404 16776
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 10778 16776 10784 16788
rect 10739 16748 10784 16776
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 12158 16776 12164 16788
rect 12119 16748 12164 16776
rect 12158 16736 12164 16748
rect 12216 16736 12222 16788
rect 12986 16776 12992 16788
rect 12947 16748 12992 16776
rect 12986 16736 12992 16748
rect 13044 16776 13050 16788
rect 13541 16779 13599 16785
rect 13541 16776 13553 16779
rect 13044 16748 13553 16776
rect 13044 16736 13050 16748
rect 13541 16745 13553 16748
rect 13587 16745 13599 16779
rect 13541 16739 13599 16745
rect 7098 16668 7104 16720
rect 7156 16708 7162 16720
rect 8015 16711 8073 16717
rect 8015 16708 8027 16711
rect 7156 16680 8027 16708
rect 7156 16668 7162 16680
rect 8015 16677 8027 16680
rect 8061 16708 8073 16711
rect 9490 16708 9496 16720
rect 8061 16680 9496 16708
rect 8061 16677 8073 16680
rect 8015 16671 8073 16677
rect 9490 16668 9496 16680
rect 9548 16708 9554 16720
rect 10223 16711 10281 16717
rect 10223 16708 10235 16711
rect 9548 16680 10235 16708
rect 9548 16668 9554 16680
rect 10223 16677 10235 16680
rect 10269 16708 10281 16711
rect 10318 16708 10324 16720
rect 10269 16680 10324 16708
rect 10269 16677 10281 16680
rect 10223 16671 10281 16677
rect 10318 16668 10324 16680
rect 10376 16668 10382 16720
rect 13556 16708 13584 16739
rect 14182 16736 14188 16788
rect 14240 16736 14246 16788
rect 15286 16736 15292 16788
rect 15344 16776 15350 16788
rect 15933 16779 15991 16785
rect 15933 16776 15945 16779
rect 15344 16748 15945 16776
rect 15344 16736 15350 16748
rect 15933 16745 15945 16748
rect 15979 16745 15991 16779
rect 15933 16739 15991 16745
rect 18141 16779 18199 16785
rect 18141 16745 18153 16779
rect 18187 16776 18199 16779
rect 18230 16776 18236 16788
rect 18187 16748 18236 16776
rect 18187 16745 18199 16748
rect 18141 16739 18199 16745
rect 18230 16736 18236 16748
rect 18288 16776 18294 16788
rect 19426 16776 19432 16788
rect 18288 16748 18368 16776
rect 19387 16748 19432 16776
rect 18288 16736 18294 16748
rect 14200 16708 14228 16736
rect 17494 16708 17500 16720
rect 13556 16680 14228 16708
rect 17455 16680 17500 16708
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 18340 16717 18368 16748
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 20530 16776 20536 16788
rect 20491 16748 20536 16776
rect 20530 16736 20536 16748
rect 20588 16736 20594 16788
rect 21082 16736 21088 16788
rect 21140 16776 21146 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 21140 16748 21189 16776
rect 21140 16736 21146 16748
rect 21177 16745 21189 16748
rect 21223 16745 21235 16779
rect 22738 16776 22744 16788
rect 22699 16748 22744 16776
rect 21177 16739 21235 16745
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 26602 16776 26608 16788
rect 26563 16748 26608 16776
rect 26602 16736 26608 16748
rect 26660 16736 26666 16788
rect 27614 16776 27620 16788
rect 27575 16748 27620 16776
rect 27614 16736 27620 16748
rect 27672 16736 27678 16788
rect 28258 16776 28264 16788
rect 28219 16748 28264 16776
rect 28258 16736 28264 16748
rect 28316 16736 28322 16788
rect 29365 16779 29423 16785
rect 29365 16745 29377 16779
rect 29411 16776 29423 16779
rect 29730 16776 29736 16788
rect 29411 16748 29736 16776
rect 29411 16745 29423 16748
rect 29365 16739 29423 16745
rect 18325 16711 18383 16717
rect 18325 16677 18337 16711
rect 18371 16677 18383 16711
rect 23198 16708 23204 16720
rect 23159 16680 23204 16708
rect 18325 16671 18383 16677
rect 23198 16668 23204 16680
rect 23256 16668 23262 16720
rect 26237 16711 26295 16717
rect 26237 16677 26249 16711
rect 26283 16708 26295 16711
rect 26694 16708 26700 16720
rect 26283 16680 26700 16708
rect 26283 16677 26295 16680
rect 26237 16671 26295 16677
rect 26694 16668 26700 16680
rect 26752 16668 26758 16720
rect 27246 16708 27252 16720
rect 26804 16680 27252 16708
rect 2682 16640 2688 16652
rect 2643 16612 2688 16640
rect 2682 16600 2688 16612
rect 2740 16600 2746 16652
rect 2961 16643 3019 16649
rect 2961 16609 2973 16643
rect 3007 16640 3019 16643
rect 3234 16640 3240 16652
rect 3007 16612 3240 16640
rect 3007 16609 3019 16612
rect 2961 16603 3019 16609
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 3326 16600 3332 16652
rect 3384 16640 3390 16652
rect 3970 16640 3976 16652
rect 3384 16612 3976 16640
rect 3384 16600 3390 16612
rect 3970 16600 3976 16612
rect 4028 16640 4034 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 4028 16612 4077 16640
rect 4028 16600 4034 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4614 16640 4620 16652
rect 4575 16612 4620 16640
rect 4065 16603 4123 16609
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 5074 16600 5080 16652
rect 5132 16640 5138 16652
rect 5629 16643 5687 16649
rect 5629 16640 5641 16643
rect 5132 16612 5641 16640
rect 5132 16600 5138 16612
rect 5629 16609 5641 16612
rect 5675 16640 5687 16643
rect 5902 16640 5908 16652
rect 5675 16612 5908 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 5902 16600 5908 16612
rect 5960 16600 5966 16652
rect 6086 16640 6092 16652
rect 6047 16612 6092 16640
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16640 7251 16643
rect 7558 16640 7564 16652
rect 7239 16612 7564 16640
rect 7239 16609 7251 16612
rect 7193 16603 7251 16609
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16640 7711 16643
rect 7742 16640 7748 16652
rect 7699 16612 7748 16640
rect 7699 16609 7711 16612
rect 7653 16603 7711 16609
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9824 16612 9873 16640
rect 9824 16600 9830 16612
rect 9861 16609 9873 16612
rect 9907 16609 9919 16643
rect 11790 16640 11796 16652
rect 11751 16612 11796 16640
rect 9861 16603 9919 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 14252 16643 14310 16649
rect 14252 16640 14264 16643
rect 13872 16612 14264 16640
rect 13872 16600 13878 16612
rect 14252 16609 14264 16612
rect 14298 16640 14310 16643
rect 14642 16640 14648 16652
rect 14298 16612 14648 16640
rect 14298 16609 14310 16612
rect 14252 16603 14310 16609
rect 14642 16600 14648 16612
rect 14700 16600 14706 16652
rect 15562 16649 15568 16652
rect 15540 16643 15568 16649
rect 15540 16640 15552 16643
rect 15475 16612 15552 16640
rect 15540 16609 15552 16612
rect 15620 16640 15626 16652
rect 16114 16640 16120 16652
rect 15620 16612 16120 16640
rect 15540 16603 15568 16609
rect 15562 16600 15568 16603
rect 15620 16600 15626 16612
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 17129 16643 17187 16649
rect 17129 16609 17141 16643
rect 17175 16640 17187 16643
rect 18506 16640 18512 16652
rect 17175 16612 18512 16640
rect 17175 16609 17187 16612
rect 17129 16603 17187 16609
rect 3142 16572 3148 16584
rect 3103 16544 3148 16572
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 4801 16575 4859 16581
rect 4801 16541 4813 16575
rect 4847 16572 4859 16575
rect 4890 16572 4896 16584
rect 4847 16544 4896 16572
rect 4847 16541 4859 16544
rect 4801 16535 4859 16541
rect 4890 16532 4896 16544
rect 4948 16532 4954 16584
rect 6362 16572 6368 16584
rect 6323 16544 6368 16572
rect 6362 16532 6368 16544
rect 6420 16532 6426 16584
rect 13998 16532 14004 16584
rect 14056 16572 14062 16584
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 14056 16544 14105 16572
rect 14056 16532 14062 16544
rect 14093 16541 14105 16544
rect 14139 16572 14151 16575
rect 16206 16572 16212 16584
rect 14139 16544 16212 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 16960 16572 16988 16603
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 21082 16600 21088 16652
rect 21140 16640 21146 16652
rect 21545 16643 21603 16649
rect 21545 16640 21557 16643
rect 21140 16612 21557 16640
rect 21140 16600 21146 16612
rect 21545 16609 21557 16612
rect 21591 16640 21603 16643
rect 22094 16640 22100 16652
rect 21591 16612 22100 16640
rect 21591 16609 21603 16612
rect 21545 16603 21603 16609
rect 22094 16600 22100 16612
rect 22152 16600 22158 16652
rect 24486 16640 24492 16652
rect 24447 16612 24492 16640
rect 24486 16600 24492 16612
rect 24544 16640 24550 16652
rect 26326 16640 26332 16652
rect 24544 16612 26332 16640
rect 24544 16600 24550 16612
rect 26326 16600 26332 16612
rect 26384 16600 26390 16652
rect 26804 16649 26832 16680
rect 27246 16668 27252 16680
rect 27304 16708 27310 16720
rect 28902 16708 28908 16720
rect 27304 16680 28908 16708
rect 27304 16668 27310 16680
rect 28902 16668 28908 16680
rect 28960 16668 28966 16720
rect 26789 16643 26847 16649
rect 26789 16609 26801 16643
rect 26835 16609 26847 16643
rect 26789 16603 26847 16609
rect 27065 16643 27123 16649
rect 27065 16609 27077 16643
rect 27111 16640 27123 16643
rect 27154 16640 27160 16652
rect 27111 16612 27160 16640
rect 27111 16609 27123 16612
rect 27065 16603 27123 16609
rect 18046 16572 18052 16584
rect 16960 16544 18052 16572
rect 18046 16532 18052 16544
rect 18104 16532 18110 16584
rect 19886 16572 19892 16584
rect 19799 16544 19892 16572
rect 19886 16532 19892 16544
rect 19944 16572 19950 16584
rect 21174 16572 21180 16584
rect 19944 16544 21180 16572
rect 19944 16532 19950 16544
rect 21174 16532 21180 16544
rect 21232 16532 21238 16584
rect 22554 16532 22560 16584
rect 22612 16572 22618 16584
rect 23109 16575 23167 16581
rect 23109 16572 23121 16575
rect 22612 16544 23121 16572
rect 22612 16532 22618 16544
rect 23109 16541 23121 16544
rect 23155 16572 23167 16575
rect 24719 16575 24777 16581
rect 24719 16572 24731 16575
rect 23155 16544 24731 16572
rect 23155 16541 23167 16544
rect 23109 16535 23167 16541
rect 24719 16541 24731 16544
rect 24765 16541 24777 16575
rect 24719 16535 24777 16541
rect 25961 16575 26019 16581
rect 25961 16541 25973 16575
rect 26007 16572 26019 16575
rect 27080 16572 27108 16603
rect 27154 16600 27160 16612
rect 27212 16600 27218 16652
rect 28350 16600 28356 16652
rect 28408 16640 28414 16652
rect 28813 16643 28871 16649
rect 28813 16640 28825 16643
rect 28408 16612 28825 16640
rect 28408 16600 28414 16612
rect 28813 16609 28825 16612
rect 28859 16640 28871 16643
rect 29380 16640 29408 16739
rect 29730 16736 29736 16748
rect 29788 16776 29794 16788
rect 30006 16776 30012 16788
rect 29788 16748 30012 16776
rect 29788 16736 29794 16748
rect 30006 16736 30012 16748
rect 30064 16736 30070 16788
rect 31294 16736 31300 16788
rect 31352 16776 31358 16788
rect 31389 16779 31447 16785
rect 31389 16776 31401 16779
rect 31352 16748 31401 16776
rect 31352 16736 31358 16748
rect 31389 16745 31401 16748
rect 31435 16745 31447 16779
rect 31938 16776 31944 16788
rect 31899 16748 31944 16776
rect 31389 16739 31447 16745
rect 31938 16736 31944 16748
rect 31996 16736 32002 16788
rect 33410 16776 33416 16788
rect 33371 16748 33416 16776
rect 33410 16736 33416 16748
rect 33468 16736 33474 16788
rect 34330 16776 34336 16788
rect 34291 16748 34336 16776
rect 34330 16736 34336 16748
rect 34388 16736 34394 16788
rect 40310 16776 40316 16788
rect 40271 16748 40316 16776
rect 40310 16736 40316 16748
rect 40368 16736 40374 16788
rect 45051 16779 45109 16785
rect 45051 16776 45063 16779
rect 43456 16748 45063 16776
rect 30282 16668 30288 16720
rect 30340 16708 30346 16720
rect 30514 16711 30572 16717
rect 30514 16708 30526 16711
rect 30340 16680 30526 16708
rect 30340 16668 30346 16680
rect 30514 16677 30526 16680
rect 30560 16677 30572 16711
rect 32214 16708 32220 16720
rect 32175 16680 32220 16708
rect 30514 16671 30572 16677
rect 32214 16668 32220 16680
rect 32272 16668 32278 16720
rect 32306 16668 32312 16720
rect 32364 16708 32370 16720
rect 36075 16711 36133 16717
rect 32364 16680 32409 16708
rect 32364 16668 32370 16680
rect 36075 16677 36087 16711
rect 36121 16708 36133 16711
rect 36170 16708 36176 16720
rect 36121 16680 36176 16708
rect 36121 16677 36133 16680
rect 36075 16671 36133 16677
rect 36170 16668 36176 16680
rect 36228 16668 36234 16720
rect 36722 16668 36728 16720
rect 36780 16708 36786 16720
rect 37458 16708 37464 16720
rect 36780 16680 37464 16708
rect 36780 16668 36786 16680
rect 37458 16668 37464 16680
rect 37516 16708 37522 16720
rect 37829 16711 37887 16717
rect 37829 16708 37841 16711
rect 37516 16680 37841 16708
rect 37516 16668 37522 16680
rect 37829 16677 37841 16680
rect 37875 16677 37887 16711
rect 37829 16671 37887 16677
rect 37921 16711 37979 16717
rect 37921 16677 37933 16711
rect 37967 16708 37979 16711
rect 38010 16708 38016 16720
rect 37967 16680 38016 16708
rect 37967 16677 37979 16680
rect 37921 16671 37979 16677
rect 38010 16668 38016 16680
rect 38068 16668 38074 16720
rect 38470 16708 38476 16720
rect 38431 16680 38476 16708
rect 38470 16668 38476 16680
rect 38528 16668 38534 16720
rect 40681 16711 40739 16717
rect 40681 16677 40693 16711
rect 40727 16708 40739 16711
rect 40862 16708 40868 16720
rect 40727 16680 40868 16708
rect 40727 16677 40739 16680
rect 40681 16671 40739 16677
rect 40862 16668 40868 16680
rect 40920 16668 40926 16720
rect 40957 16711 41015 16717
rect 40957 16677 40969 16711
rect 41003 16708 41015 16711
rect 41046 16708 41052 16720
rect 41003 16680 41052 16708
rect 41003 16677 41015 16680
rect 40957 16671 41015 16677
rect 41046 16668 41052 16680
rect 41104 16668 41110 16720
rect 43162 16668 43168 16720
rect 43220 16708 43226 16720
rect 43456 16717 43484 16748
rect 45051 16745 45063 16748
rect 45097 16745 45109 16779
rect 45051 16739 45109 16745
rect 43441 16711 43499 16717
rect 43441 16708 43453 16711
rect 43220 16680 43453 16708
rect 43220 16668 43226 16680
rect 43441 16677 43453 16680
rect 43487 16677 43499 16711
rect 43441 16671 43499 16677
rect 43533 16711 43591 16717
rect 43533 16677 43545 16711
rect 43579 16708 43591 16711
rect 43622 16708 43628 16720
rect 43579 16680 43628 16708
rect 43579 16677 43591 16680
rect 43533 16671 43591 16677
rect 43622 16668 43628 16680
rect 43680 16668 43686 16720
rect 28859 16612 29408 16640
rect 28859 16609 28871 16612
rect 28813 16603 28871 16609
rect 35250 16600 35256 16652
rect 35308 16640 35314 16652
rect 35713 16643 35771 16649
rect 35713 16640 35725 16643
rect 35308 16612 35725 16640
rect 35308 16600 35314 16612
rect 35713 16609 35725 16612
rect 35759 16609 35771 16643
rect 39298 16640 39304 16652
rect 39259 16612 39304 16640
rect 35713 16603 35771 16609
rect 39298 16600 39304 16612
rect 39356 16600 39362 16652
rect 44913 16643 44971 16649
rect 44913 16609 44925 16643
rect 44959 16640 44971 16643
rect 45002 16640 45008 16652
rect 44959 16612 45008 16640
rect 44959 16609 44971 16612
rect 44913 16603 44971 16609
rect 45002 16600 45008 16612
rect 45060 16600 45066 16652
rect 30190 16572 30196 16584
rect 26007 16544 27108 16572
rect 30151 16544 30196 16572
rect 26007 16541 26019 16544
rect 25961 16535 26019 16541
rect 30190 16532 30196 16544
rect 30248 16532 30254 16584
rect 32490 16572 32496 16584
rect 32451 16544 32496 16572
rect 32490 16532 32496 16544
rect 32548 16532 32554 16584
rect 33962 16572 33968 16584
rect 33923 16544 33968 16572
rect 33962 16532 33968 16544
rect 34020 16532 34026 16584
rect 43717 16575 43775 16581
rect 43717 16572 43729 16575
rect 43548 16544 43729 16572
rect 23566 16464 23572 16516
rect 23624 16504 23630 16516
rect 23661 16507 23719 16513
rect 23661 16504 23673 16507
rect 23624 16476 23673 16504
rect 23624 16464 23630 16476
rect 23661 16473 23673 16476
rect 23707 16473 23719 16507
rect 23661 16467 23719 16473
rect 24302 16464 24308 16516
rect 24360 16504 24366 16516
rect 24397 16507 24455 16513
rect 24397 16504 24409 16507
rect 24360 16476 24409 16504
rect 24360 16464 24366 16476
rect 24397 16473 24409 16476
rect 24443 16504 24455 16507
rect 27890 16504 27896 16516
rect 24443 16476 27896 16504
rect 24443 16473 24455 16476
rect 24397 16467 24455 16473
rect 27890 16464 27896 16476
rect 27948 16464 27954 16516
rect 41417 16507 41475 16513
rect 41417 16473 41429 16507
rect 41463 16504 41475 16507
rect 42242 16504 42248 16516
rect 41463 16476 42248 16504
rect 41463 16473 41475 16476
rect 41417 16467 41475 16473
rect 42242 16464 42248 16476
rect 42300 16504 42306 16516
rect 43548 16504 43576 16544
rect 43717 16541 43729 16544
rect 43763 16541 43775 16575
rect 43717 16535 43775 16541
rect 42300 16476 43576 16504
rect 42300 16464 42306 16476
rect 8570 16436 8576 16448
rect 8531 16408 8576 16436
rect 8570 16396 8576 16408
rect 8628 16396 8634 16448
rect 12710 16436 12716 16448
rect 12671 16408 12716 16436
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 14323 16439 14381 16445
rect 14323 16405 14335 16439
rect 14369 16436 14381 16439
rect 15470 16436 15476 16448
rect 14369 16408 15476 16436
rect 14369 16405 14381 16408
rect 14323 16399 14381 16405
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15611 16439 15669 16445
rect 15611 16405 15623 16439
rect 15657 16436 15669 16439
rect 15838 16436 15844 16448
rect 15657 16408 15844 16436
rect 15657 16405 15669 16408
rect 15611 16399 15669 16405
rect 15838 16396 15844 16408
rect 15896 16396 15902 16448
rect 22094 16436 22100 16448
rect 22055 16408 22100 16436
rect 22094 16396 22100 16408
rect 22152 16396 22158 16448
rect 28994 16436 29000 16448
rect 28955 16408 29000 16436
rect 28994 16396 29000 16408
rect 29052 16396 29058 16448
rect 31110 16436 31116 16448
rect 31071 16408 31116 16436
rect 31110 16396 31116 16408
rect 31168 16396 31174 16448
rect 34885 16439 34943 16445
rect 34885 16405 34897 16439
rect 34931 16436 34943 16439
rect 36354 16436 36360 16448
rect 34931 16408 36360 16436
rect 34931 16405 34943 16408
rect 34885 16399 34943 16405
rect 36354 16396 36360 16408
rect 36412 16396 36418 16448
rect 36630 16436 36636 16448
rect 36591 16408 36636 16436
rect 36630 16396 36636 16408
rect 36688 16436 36694 16448
rect 36909 16439 36967 16445
rect 36909 16436 36921 16439
rect 36688 16408 36921 16436
rect 36688 16396 36694 16408
rect 36909 16405 36921 16408
rect 36955 16405 36967 16439
rect 39482 16436 39488 16448
rect 39443 16408 39488 16436
rect 36909 16399 36967 16405
rect 39482 16396 39488 16408
rect 39540 16396 39546 16448
rect 1104 16346 48852 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 48852 16346
rect 1104 16272 48852 16294
rect 2501 16235 2559 16241
rect 2501 16201 2513 16235
rect 2547 16232 2559 16235
rect 2682 16232 2688 16244
rect 2547 16204 2688 16232
rect 2547 16201 2559 16204
rect 2501 16195 2559 16201
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 2869 16235 2927 16241
rect 2869 16201 2881 16235
rect 2915 16232 2927 16235
rect 3234 16232 3240 16244
rect 2915 16204 3240 16232
rect 2915 16201 2927 16204
rect 2869 16195 2927 16201
rect 3234 16192 3240 16204
rect 3292 16232 3298 16244
rect 3694 16232 3700 16244
rect 3292 16204 3700 16232
rect 3292 16192 3298 16204
rect 3694 16192 3700 16204
rect 3752 16192 3758 16244
rect 3970 16192 3976 16244
rect 4028 16232 4034 16244
rect 4065 16235 4123 16241
rect 4065 16232 4077 16235
rect 4028 16204 4077 16232
rect 4028 16192 4034 16204
rect 4065 16201 4077 16204
rect 4111 16201 4123 16235
rect 5902 16232 5908 16244
rect 5863 16204 5908 16232
rect 4065 16195 4123 16201
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 6086 16192 6092 16244
rect 6144 16232 6150 16244
rect 6273 16235 6331 16241
rect 6273 16232 6285 16235
rect 6144 16204 6285 16232
rect 6144 16192 6150 16204
rect 6273 16201 6285 16204
rect 6319 16201 6331 16235
rect 6273 16195 6331 16201
rect 7101 16235 7159 16241
rect 7101 16201 7113 16235
rect 7147 16232 7159 16235
rect 7742 16232 7748 16244
rect 7147 16204 7748 16232
rect 7147 16201 7159 16204
rect 7101 16195 7159 16201
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 15562 16232 15568 16244
rect 13872 16204 13917 16232
rect 15523 16204 15568 16232
rect 13872 16192 13878 16204
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 17129 16235 17187 16241
rect 17129 16201 17141 16235
rect 17175 16232 17187 16235
rect 20438 16232 20444 16244
rect 17175 16204 20444 16232
rect 17175 16201 17187 16204
rect 17129 16195 17187 16201
rect 20438 16192 20444 16204
rect 20496 16192 20502 16244
rect 21082 16232 21088 16244
rect 21043 16204 21088 16232
rect 21082 16192 21088 16204
rect 21140 16192 21146 16244
rect 23109 16235 23167 16241
rect 23109 16201 23121 16235
rect 23155 16232 23167 16235
rect 23198 16232 23204 16244
rect 23155 16204 23204 16232
rect 23155 16201 23167 16204
rect 23109 16195 23167 16201
rect 23198 16192 23204 16204
rect 23256 16192 23262 16244
rect 23293 16235 23351 16241
rect 23293 16201 23305 16235
rect 23339 16232 23351 16235
rect 25866 16232 25872 16244
rect 23339 16204 25872 16232
rect 23339 16201 23351 16204
rect 23293 16195 23351 16201
rect 25866 16192 25872 16204
rect 25924 16192 25930 16244
rect 27246 16232 27252 16244
rect 27207 16204 27252 16232
rect 27246 16192 27252 16204
rect 27304 16192 27310 16244
rect 28902 16192 28908 16244
rect 28960 16232 28966 16244
rect 28997 16235 29055 16241
rect 28997 16232 29009 16235
rect 28960 16204 29009 16232
rect 28960 16192 28966 16204
rect 28997 16201 29009 16204
rect 29043 16201 29055 16235
rect 28997 16195 29055 16201
rect 17865 16167 17923 16173
rect 17865 16133 17877 16167
rect 17911 16164 17923 16167
rect 18046 16164 18052 16176
rect 17911 16136 18052 16164
rect 17911 16133 17923 16136
rect 17865 16127 17923 16133
rect 18046 16124 18052 16136
rect 18104 16124 18110 16176
rect 22649 16167 22707 16173
rect 22649 16133 22661 16167
rect 22695 16164 22707 16167
rect 23566 16164 23572 16176
rect 22695 16136 23572 16164
rect 22695 16133 22707 16136
rect 22649 16127 22707 16133
rect 23566 16124 23572 16136
rect 23624 16124 23630 16176
rect 24486 16124 24492 16176
rect 24544 16164 24550 16176
rect 24673 16167 24731 16173
rect 24673 16164 24685 16167
rect 24544 16136 24685 16164
rect 24544 16124 24550 16136
rect 24673 16133 24685 16136
rect 24719 16133 24731 16167
rect 24673 16127 24731 16133
rect 3142 16056 3148 16108
rect 3200 16096 3206 16108
rect 7561 16099 7619 16105
rect 3200 16068 4154 16096
rect 3200 16056 3206 16068
rect 4126 16028 4154 16068
rect 7561 16065 7573 16099
rect 7607 16096 7619 16099
rect 7650 16096 7656 16108
rect 7607 16068 7656 16096
rect 7607 16065 7619 16068
rect 7561 16059 7619 16065
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 9582 16096 9588 16108
rect 9495 16068 9588 16096
rect 9582 16056 9588 16068
rect 9640 16096 9646 16108
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 9640 16068 10793 16096
rect 9640 16056 9646 16068
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 12437 16099 12495 16105
rect 12437 16065 12449 16099
rect 12483 16096 12495 16099
rect 12526 16096 12532 16108
rect 12483 16068 12532 16096
rect 12483 16065 12495 16068
rect 12437 16059 12495 16065
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 14274 16096 14280 16108
rect 14235 16068 14280 16096
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 17497 16099 17555 16105
rect 17497 16065 17509 16099
rect 17543 16096 17555 16099
rect 18417 16099 18475 16105
rect 18417 16096 18429 16099
rect 17543 16068 18429 16096
rect 17543 16065 17555 16068
rect 17497 16059 17555 16065
rect 18417 16065 18429 16068
rect 18463 16096 18475 16099
rect 18506 16096 18512 16108
rect 18463 16068 18512 16096
rect 18463 16065 18475 16068
rect 18417 16059 18475 16065
rect 18506 16056 18512 16068
rect 18564 16056 18570 16108
rect 19705 16099 19763 16105
rect 19705 16065 19717 16099
rect 19751 16096 19763 16099
rect 23293 16099 23351 16105
rect 23293 16096 23305 16099
rect 19751 16068 23305 16096
rect 19751 16065 19763 16068
rect 19705 16059 19763 16065
rect 23293 16065 23305 16068
rect 23339 16065 23351 16099
rect 23293 16059 23351 16065
rect 25961 16099 26019 16105
rect 25961 16065 25973 16099
rect 26007 16096 26019 16099
rect 26050 16096 26056 16108
rect 26007 16068 26056 16096
rect 26007 16065 26019 16068
rect 25961 16059 26019 16065
rect 4706 16028 4712 16040
rect 4126 16000 4712 16028
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 16028 10563 16031
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 10551 16000 11161 16028
rect 10551 15997 10563 16000
rect 10505 15991 10563 15997
rect 11149 15997 11161 16000
rect 11195 16028 11207 16031
rect 11368 16031 11426 16037
rect 11368 16028 11380 16031
rect 11195 16000 11380 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11368 15997 11380 16000
rect 11414 15997 11426 16031
rect 11368 15991 11426 15997
rect 16853 16031 16911 16037
rect 16853 15997 16865 16031
rect 16899 16028 16911 16031
rect 16945 16031 17003 16037
rect 16945 16028 16957 16031
rect 16899 16000 16957 16028
rect 16899 15997 16911 16000
rect 16853 15991 16911 15997
rect 16945 15997 16957 16000
rect 16991 16028 17003 16031
rect 18138 16028 18144 16040
rect 16991 16000 18144 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 18138 15988 18144 16000
rect 18196 15988 18202 16040
rect 18230 15988 18236 16040
rect 18288 16028 18294 16040
rect 18969 16031 19027 16037
rect 18969 16028 18981 16031
rect 18288 16000 18981 16028
rect 18288 15988 18294 16000
rect 18969 15997 18981 16000
rect 19015 15997 19027 16031
rect 18969 15991 19027 15997
rect 6454 15960 6460 15972
rect 5092 15932 6460 15960
rect 4617 15895 4675 15901
rect 4617 15861 4629 15895
rect 4663 15892 4675 15895
rect 4982 15892 4988 15904
rect 4663 15864 4988 15892
rect 4663 15861 4675 15864
rect 4617 15855 4675 15861
rect 4982 15852 4988 15864
rect 5040 15892 5046 15904
rect 5092 15901 5120 15932
rect 6454 15920 6460 15932
rect 6512 15920 6518 15972
rect 7469 15963 7527 15969
rect 7469 15929 7481 15963
rect 7515 15960 7527 15963
rect 7650 15960 7656 15972
rect 7515 15932 7656 15960
rect 7515 15929 7527 15932
rect 7469 15923 7527 15929
rect 7650 15920 7656 15932
rect 7708 15960 7714 15972
rect 7923 15963 7981 15969
rect 7923 15960 7935 15963
rect 7708 15932 7935 15960
rect 7708 15920 7714 15932
rect 7923 15929 7935 15932
rect 7969 15960 7981 15963
rect 9125 15963 9183 15969
rect 9125 15960 9137 15963
rect 7969 15932 9137 15960
rect 7969 15929 7981 15932
rect 7923 15923 7981 15929
rect 9125 15929 9137 15932
rect 9171 15960 9183 15963
rect 9490 15960 9496 15972
rect 9171 15932 9496 15960
rect 9171 15929 9183 15932
rect 9125 15923 9183 15929
rect 9490 15920 9496 15932
rect 9548 15960 9554 15972
rect 9906 15963 9964 15969
rect 9906 15960 9918 15963
rect 9548 15932 9918 15960
rect 9548 15920 9554 15932
rect 9906 15929 9918 15932
rect 9952 15929 9964 15963
rect 9906 15923 9964 15929
rect 10318 15920 10324 15972
rect 10376 15960 10382 15972
rect 11885 15963 11943 15969
rect 11885 15960 11897 15963
rect 10376 15932 11897 15960
rect 10376 15920 10382 15932
rect 11885 15929 11897 15932
rect 11931 15960 11943 15963
rect 12158 15960 12164 15972
rect 11931 15932 12164 15960
rect 11931 15929 11943 15932
rect 11885 15923 11943 15929
rect 12158 15920 12164 15932
rect 12216 15960 12222 15972
rect 12799 15963 12857 15969
rect 12799 15960 12811 15963
rect 12216 15932 12811 15960
rect 12216 15920 12222 15932
rect 12799 15929 12811 15932
rect 12845 15960 12857 15963
rect 13538 15960 13544 15972
rect 12845 15932 13544 15960
rect 12845 15929 12857 15932
rect 12799 15923 12857 15929
rect 13538 15920 13544 15932
rect 13596 15960 13602 15972
rect 14093 15963 14151 15969
rect 14093 15960 14105 15963
rect 13596 15932 14105 15960
rect 13596 15920 13602 15932
rect 14093 15929 14105 15932
rect 14139 15960 14151 15963
rect 14550 15960 14556 15972
rect 14139 15932 14556 15960
rect 14139 15929 14151 15932
rect 14093 15923 14151 15929
rect 14550 15920 14556 15932
rect 14608 15969 14614 15972
rect 14608 15963 14656 15969
rect 14608 15929 14610 15963
rect 14644 15929 14656 15963
rect 14608 15923 14656 15929
rect 14608 15920 14614 15923
rect 17862 15920 17868 15972
rect 17920 15960 17926 15972
rect 18785 15963 18843 15969
rect 18785 15960 18797 15963
rect 17920 15932 18797 15960
rect 17920 15920 17926 15932
rect 18785 15929 18797 15932
rect 18831 15960 18843 15963
rect 19720 15960 19748 16059
rect 26050 16056 26056 16068
rect 26108 16096 26114 16108
rect 26418 16096 26424 16108
rect 26108 16068 26424 16096
rect 26108 16056 26114 16068
rect 26418 16056 26424 16068
rect 26476 16056 26482 16108
rect 26510 16056 26516 16108
rect 26568 16096 26574 16108
rect 28626 16096 28632 16108
rect 26568 16068 28632 16096
rect 26568 16056 26574 16068
rect 19886 15988 19892 16040
rect 19944 16028 19950 16040
rect 20165 16031 20223 16037
rect 20165 16028 20177 16031
rect 19944 16000 20177 16028
rect 19944 15988 19950 16000
rect 20165 15997 20177 16000
rect 20211 16028 20223 16031
rect 20625 16031 20683 16037
rect 20625 16028 20637 16031
rect 20211 16000 20637 16028
rect 20211 15997 20223 16000
rect 20165 15991 20223 15997
rect 20625 15997 20637 16000
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 23308 16000 23520 16028
rect 18831 15932 19748 15960
rect 18831 15929 18843 15932
rect 18785 15923 18843 15929
rect 20898 15920 20904 15972
rect 20956 15960 20962 15972
rect 22094 15960 22100 15972
rect 20956 15932 22100 15960
rect 20956 15920 20962 15932
rect 22094 15920 22100 15932
rect 22152 15920 22158 15972
rect 22189 15963 22247 15969
rect 22189 15929 22201 15963
rect 22235 15960 22247 15963
rect 23308 15960 23336 16000
rect 23492 15969 23520 16000
rect 27154 15988 27160 16040
rect 27212 16028 27218 16040
rect 28219 16037 28247 16068
rect 28626 16056 28632 16068
rect 28684 16056 28690 16108
rect 27525 16031 27583 16037
rect 27525 16028 27537 16031
rect 27212 16000 27537 16028
rect 27212 15988 27218 16000
rect 27525 15997 27537 16000
rect 27571 15997 27583 16031
rect 27525 15991 27583 15997
rect 28204 16031 28262 16037
rect 28204 15997 28216 16031
rect 28250 15997 28262 16031
rect 29012 16028 29040 16195
rect 31110 16192 31116 16244
rect 31168 16232 31174 16244
rect 31205 16235 31263 16241
rect 31205 16232 31217 16235
rect 31168 16204 31217 16232
rect 31168 16192 31174 16204
rect 31205 16201 31217 16204
rect 31251 16232 31263 16235
rect 31570 16232 31576 16244
rect 31251 16204 31576 16232
rect 31251 16201 31263 16204
rect 31205 16195 31263 16201
rect 31570 16192 31576 16204
rect 31628 16192 31634 16244
rect 32306 16192 32312 16244
rect 32364 16232 32370 16244
rect 32401 16235 32459 16241
rect 32401 16232 32413 16235
rect 32364 16204 32413 16232
rect 32364 16192 32370 16204
rect 32401 16201 32413 16204
rect 32447 16201 32459 16235
rect 32401 16195 32459 16201
rect 33134 16192 33140 16244
rect 33192 16232 33198 16244
rect 35250 16232 35256 16244
rect 33192 16204 33237 16232
rect 35211 16204 35256 16232
rect 33192 16192 33198 16204
rect 35250 16192 35256 16204
rect 35308 16192 35314 16244
rect 36170 16192 36176 16244
rect 36228 16232 36234 16244
rect 38381 16235 38439 16241
rect 38381 16232 38393 16235
rect 36228 16204 38393 16232
rect 36228 16192 36234 16204
rect 38381 16201 38393 16204
rect 38427 16232 38439 16235
rect 38473 16235 38531 16241
rect 38473 16232 38485 16235
rect 38427 16204 38485 16232
rect 38427 16201 38439 16204
rect 38381 16195 38439 16201
rect 38473 16201 38485 16204
rect 38519 16201 38531 16235
rect 38473 16195 38531 16201
rect 39298 16192 39304 16244
rect 39356 16232 39362 16244
rect 39853 16235 39911 16241
rect 39853 16232 39865 16235
rect 39356 16204 39865 16232
rect 39356 16192 39362 16204
rect 39853 16201 39865 16204
rect 39899 16201 39911 16235
rect 39853 16195 39911 16201
rect 29638 16124 29644 16176
rect 29696 16164 29702 16176
rect 29696 16136 32622 16164
rect 29696 16124 29702 16136
rect 30009 16099 30067 16105
rect 30009 16065 30021 16099
rect 30055 16096 30067 16099
rect 30190 16096 30196 16108
rect 30055 16068 30196 16096
rect 30055 16065 30067 16068
rect 30009 16059 30067 16065
rect 30190 16056 30196 16068
rect 30248 16096 30254 16108
rect 30653 16099 30711 16105
rect 30653 16096 30665 16099
rect 30248 16068 30665 16096
rect 30248 16056 30254 16068
rect 30653 16065 30665 16068
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 31294 16056 31300 16108
rect 31352 16096 31358 16108
rect 31481 16099 31539 16105
rect 31481 16096 31493 16099
rect 31352 16068 31493 16096
rect 31352 16056 31358 16068
rect 31481 16065 31493 16068
rect 31527 16065 31539 16099
rect 31481 16059 31539 16065
rect 32125 16099 32183 16105
rect 32125 16065 32137 16099
rect 32171 16096 32183 16099
rect 32306 16096 32312 16108
rect 32171 16068 32312 16096
rect 32171 16065 32183 16068
rect 32125 16059 32183 16065
rect 32306 16056 32312 16068
rect 32364 16096 32370 16108
rect 32490 16096 32496 16108
rect 32364 16068 32496 16096
rect 32364 16056 32370 16068
rect 32490 16056 32496 16068
rect 32548 16056 32554 16108
rect 29273 16031 29331 16037
rect 29273 16028 29285 16031
rect 29012 16000 29285 16028
rect 28204 15991 28262 15997
rect 29273 15997 29285 16000
rect 29319 15997 29331 16031
rect 29730 16028 29736 16040
rect 29691 16000 29736 16028
rect 29273 15991 29331 15997
rect 29730 15988 29736 16000
rect 29788 15988 29794 16040
rect 32594 16028 32622 16136
rect 33152 16096 33180 16192
rect 38562 16164 38568 16176
rect 36648 16136 38568 16164
rect 33962 16096 33968 16108
rect 33152 16068 33732 16096
rect 33875 16068 33968 16096
rect 33502 16028 33508 16040
rect 32594 16000 33508 16028
rect 33502 15988 33508 16000
rect 33560 15988 33566 16040
rect 33704 16037 33732 16068
rect 33962 16056 33968 16068
rect 34020 16096 34026 16108
rect 34609 16099 34667 16105
rect 34609 16096 34621 16099
rect 34020 16068 34621 16096
rect 34020 16056 34026 16068
rect 34609 16065 34621 16068
rect 34655 16065 34667 16099
rect 34609 16059 34667 16065
rect 36357 16099 36415 16105
rect 36357 16065 36369 16099
rect 36403 16096 36415 16099
rect 36648 16096 36676 16136
rect 38562 16124 38568 16136
rect 38620 16124 38626 16176
rect 41325 16167 41383 16173
rect 41325 16133 41337 16167
rect 41371 16164 41383 16167
rect 42150 16164 42156 16176
rect 41371 16136 42156 16164
rect 41371 16133 41383 16136
rect 41325 16127 41383 16133
rect 42150 16124 42156 16136
rect 42208 16164 42214 16176
rect 42208 16136 44404 16164
rect 42208 16124 42214 16136
rect 37182 16096 37188 16108
rect 36403 16068 36676 16096
rect 37143 16068 37188 16096
rect 36403 16065 36415 16068
rect 36357 16059 36415 16065
rect 33689 16031 33747 16037
rect 33689 15997 33701 16031
rect 33735 15997 33747 16031
rect 33689 15991 33747 15997
rect 34054 15988 34060 16040
rect 34112 16028 34118 16040
rect 35488 16031 35546 16037
rect 35488 16028 35500 16031
rect 34112 16000 35500 16028
rect 34112 15988 34118 16000
rect 35488 15997 35500 16000
rect 35534 16028 35546 16031
rect 36372 16028 36400 16059
rect 37182 16056 37188 16068
rect 37240 16056 37246 16108
rect 40310 16056 40316 16108
rect 40368 16096 40374 16108
rect 40773 16099 40831 16105
rect 40773 16096 40785 16099
rect 40368 16068 40785 16096
rect 40368 16056 40374 16068
rect 40773 16065 40785 16068
rect 40819 16065 40831 16099
rect 40773 16059 40831 16065
rect 42058 16056 42064 16108
rect 42116 16096 42122 16108
rect 42245 16099 42303 16105
rect 42245 16096 42257 16099
rect 42116 16068 42257 16096
rect 42116 16056 42122 16068
rect 42245 16065 42257 16068
rect 42291 16065 42303 16099
rect 44082 16096 44088 16108
rect 44043 16068 44088 16096
rect 42245 16059 42303 16065
rect 44082 16056 44088 16068
rect 44140 16056 44146 16108
rect 44376 16105 44404 16136
rect 44361 16099 44419 16105
rect 44361 16065 44373 16099
rect 44407 16065 44419 16099
rect 44361 16059 44419 16065
rect 35534 16000 36400 16028
rect 38197 16031 38255 16037
rect 35534 15997 35546 16000
rect 35488 15991 35546 15997
rect 38197 15997 38209 16031
rect 38243 16028 38255 16031
rect 38562 16028 38568 16040
rect 38243 16000 38568 16028
rect 38243 15997 38255 16000
rect 38197 15991 38255 15997
rect 38562 15988 38568 16000
rect 38620 16028 38626 16040
rect 38657 16031 38715 16037
rect 38657 16028 38669 16031
rect 38620 16000 38669 16028
rect 38620 15988 38626 16000
rect 38657 15997 38669 16000
rect 38703 15997 38715 16031
rect 38657 15991 38715 15997
rect 39577 16031 39635 16037
rect 39577 15997 39589 16031
rect 39623 16028 39635 16031
rect 40221 16031 40279 16037
rect 40221 16028 40233 16031
rect 39623 16000 40233 16028
rect 39623 15997 39635 16000
rect 39577 15991 39635 15997
rect 40221 15997 40233 16000
rect 40267 15997 40279 16031
rect 40221 15991 40279 15997
rect 22235 15932 23336 15960
rect 23477 15963 23535 15969
rect 22235 15929 22247 15932
rect 22189 15923 22247 15929
rect 23477 15929 23489 15963
rect 23523 15929 23535 15963
rect 23750 15960 23756 15972
rect 23711 15932 23756 15960
rect 23477 15923 23535 15929
rect 5077 15895 5135 15901
rect 5077 15892 5089 15895
rect 5040 15864 5089 15892
rect 5040 15852 5046 15864
rect 5077 15861 5089 15864
rect 5123 15861 5135 15895
rect 5077 15855 5135 15861
rect 5629 15895 5687 15901
rect 5629 15861 5641 15895
rect 5675 15892 5687 15895
rect 5810 15892 5816 15904
rect 5675 15864 5816 15892
rect 5675 15861 5687 15864
rect 5629 15855 5687 15861
rect 5810 15852 5816 15864
rect 5868 15852 5874 15904
rect 8478 15892 8484 15904
rect 8439 15864 8484 15892
rect 8478 15852 8484 15864
rect 8536 15852 8542 15904
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 11471 15895 11529 15901
rect 11471 15892 11483 15895
rect 10560 15864 11483 15892
rect 10560 15852 10566 15864
rect 11471 15861 11483 15864
rect 11517 15861 11529 15895
rect 11471 15855 11529 15861
rect 12250 15852 12256 15904
rect 12308 15892 12314 15904
rect 13357 15895 13415 15901
rect 13357 15892 13369 15895
rect 12308 15864 13369 15892
rect 12308 15852 12314 15864
rect 13357 15861 13369 15864
rect 13403 15861 13415 15895
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 13357 15855 13415 15861
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 19058 15892 19064 15904
rect 19019 15864 19064 15892
rect 19058 15852 19064 15864
rect 19116 15852 19122 15904
rect 20162 15852 20168 15904
rect 20220 15892 20226 15904
rect 20349 15895 20407 15901
rect 20349 15892 20361 15895
rect 20220 15864 20361 15892
rect 20220 15852 20226 15864
rect 20349 15861 20361 15864
rect 20395 15861 20407 15895
rect 20349 15855 20407 15861
rect 21913 15895 21971 15901
rect 21913 15861 21925 15895
rect 21959 15892 21971 15895
rect 22204 15892 22232 15923
rect 21959 15864 22232 15892
rect 23492 15892 23520 15923
rect 23750 15920 23756 15932
rect 23808 15920 23814 15972
rect 23842 15920 23848 15972
rect 23900 15960 23906 15972
rect 24397 15963 24455 15969
rect 23900 15932 23945 15960
rect 23900 15920 23906 15932
rect 24397 15929 24409 15963
rect 24443 15960 24455 15963
rect 24578 15960 24584 15972
rect 24443 15932 24584 15960
rect 24443 15929 24455 15932
rect 24397 15923 24455 15929
rect 24578 15920 24584 15932
rect 24636 15920 24642 15972
rect 26326 15969 26332 15972
rect 25869 15963 25927 15969
rect 25869 15929 25881 15963
rect 25915 15960 25927 15963
rect 26282 15963 26332 15969
rect 26282 15960 26294 15963
rect 25915 15932 26294 15960
rect 25915 15929 25927 15932
rect 25869 15923 25927 15929
rect 26282 15929 26294 15932
rect 26328 15929 26332 15963
rect 26282 15923 26332 15929
rect 26326 15920 26332 15923
rect 26384 15920 26390 15972
rect 28307 15963 28365 15969
rect 28307 15929 28319 15963
rect 28353 15960 28365 15963
rect 31478 15960 31484 15972
rect 28353 15932 31484 15960
rect 28353 15929 28365 15932
rect 28307 15923 28365 15929
rect 31478 15920 31484 15932
rect 31536 15920 31542 15972
rect 31570 15920 31576 15972
rect 31628 15960 31634 15972
rect 31628 15932 31673 15960
rect 31628 15920 31634 15932
rect 31754 15920 31760 15972
rect 31812 15960 31818 15972
rect 34241 15963 34299 15969
rect 34241 15960 34253 15963
rect 31812 15932 34253 15960
rect 31812 15920 31818 15932
rect 34241 15929 34253 15932
rect 34287 15960 34299 15963
rect 34330 15960 34336 15972
rect 34287 15932 34336 15960
rect 34287 15929 34299 15932
rect 34241 15923 34299 15929
rect 34330 15920 34336 15932
rect 34388 15920 34394 15972
rect 35575 15963 35633 15969
rect 35575 15929 35587 15963
rect 35621 15960 35633 15963
rect 36538 15960 36544 15972
rect 35621 15932 36544 15960
rect 35621 15929 35633 15932
rect 35575 15923 35633 15929
rect 36538 15920 36544 15932
rect 36596 15920 36602 15972
rect 36633 15963 36691 15969
rect 36633 15929 36645 15963
rect 36679 15929 36691 15963
rect 36633 15923 36691 15929
rect 38381 15963 38439 15969
rect 38381 15929 38393 15963
rect 38427 15960 38439 15963
rect 39019 15963 39077 15969
rect 39019 15960 39031 15963
rect 38427 15932 39031 15960
rect 38427 15929 38439 15932
rect 38381 15923 38439 15929
rect 39019 15929 39031 15932
rect 39065 15960 39077 15963
rect 39666 15960 39672 15972
rect 39065 15932 39672 15960
rect 39065 15929 39077 15932
rect 39019 15923 39077 15929
rect 23860 15892 23888 15920
rect 23492 15864 23888 15892
rect 21959 15861 21971 15864
rect 21913 15855 21971 15861
rect 25314 15852 25320 15904
rect 25372 15892 25378 15904
rect 26881 15895 26939 15901
rect 26881 15892 26893 15895
rect 25372 15864 26893 15892
rect 25372 15852 25378 15864
rect 26881 15861 26893 15864
rect 26927 15861 26939 15895
rect 30282 15892 30288 15904
rect 30243 15864 30288 15892
rect 26881 15855 26939 15861
rect 30282 15852 30288 15864
rect 30340 15852 30346 15904
rect 34348 15892 34376 15920
rect 34514 15892 34520 15904
rect 34348 15864 34520 15892
rect 34514 15852 34520 15864
rect 34572 15892 34578 15904
rect 35897 15895 35955 15901
rect 35897 15892 35909 15895
rect 34572 15864 35909 15892
rect 34572 15852 34578 15864
rect 35897 15861 35909 15864
rect 35943 15892 35955 15895
rect 36170 15892 36176 15904
rect 35943 15864 36176 15892
rect 35943 15861 35955 15864
rect 35897 15855 35955 15861
rect 36170 15852 36176 15864
rect 36228 15852 36234 15904
rect 36354 15852 36360 15904
rect 36412 15892 36418 15904
rect 36648 15892 36676 15923
rect 39666 15920 39672 15932
rect 39724 15920 39730 15972
rect 40236 15960 40264 15991
rect 40310 15960 40316 15972
rect 40223 15932 40316 15960
rect 40310 15920 40316 15932
rect 40368 15960 40374 15972
rect 40865 15963 40923 15969
rect 40865 15960 40877 15963
rect 40368 15932 40877 15960
rect 40368 15920 40374 15932
rect 40865 15929 40877 15932
rect 40911 15960 40923 15963
rect 41046 15960 41052 15972
rect 40911 15932 41052 15960
rect 40911 15929 40923 15932
rect 40865 15923 40923 15929
rect 41046 15920 41052 15932
rect 41104 15920 41110 15972
rect 44177 15963 44235 15969
rect 44177 15929 44189 15963
rect 44223 15929 44235 15963
rect 44177 15923 44235 15929
rect 37461 15895 37519 15901
rect 37461 15892 37473 15895
rect 36412 15864 37473 15892
rect 36412 15852 36418 15864
rect 37461 15861 37473 15864
rect 37507 15892 37519 15895
rect 37826 15892 37832 15904
rect 37507 15864 37832 15892
rect 37507 15861 37519 15864
rect 37461 15855 37519 15861
rect 37826 15852 37832 15864
rect 37884 15892 37890 15904
rect 38010 15892 38016 15904
rect 37884 15864 38016 15892
rect 37884 15852 37890 15864
rect 38010 15852 38016 15864
rect 38068 15852 38074 15904
rect 41064 15892 41092 15920
rect 41693 15895 41751 15901
rect 41693 15892 41705 15895
rect 41064 15864 41705 15892
rect 41693 15861 41705 15864
rect 41739 15861 41751 15895
rect 41693 15855 41751 15861
rect 42153 15895 42211 15901
rect 42153 15861 42165 15895
rect 42199 15892 42211 15895
rect 42610 15892 42616 15904
rect 42199 15864 42616 15892
rect 42199 15861 42211 15864
rect 42153 15855 42211 15861
rect 42610 15852 42616 15864
rect 42668 15852 42674 15904
rect 43165 15895 43223 15901
rect 43165 15861 43177 15895
rect 43211 15892 43223 15895
rect 43533 15895 43591 15901
rect 43533 15892 43545 15895
rect 43211 15864 43545 15892
rect 43211 15861 43223 15864
rect 43165 15855 43223 15861
rect 43533 15861 43545 15864
rect 43579 15892 43591 15895
rect 43622 15892 43628 15904
rect 43579 15864 43628 15892
rect 43579 15861 43591 15864
rect 43533 15855 43591 15861
rect 43622 15852 43628 15864
rect 43680 15892 43686 15904
rect 43809 15895 43867 15901
rect 43809 15892 43821 15895
rect 43680 15864 43821 15892
rect 43680 15852 43686 15864
rect 43809 15861 43821 15864
rect 43855 15892 43867 15895
rect 44192 15892 44220 15923
rect 45002 15892 45008 15904
rect 43855 15864 44220 15892
rect 44963 15864 45008 15892
rect 43855 15861 43867 15864
rect 43809 15855 43867 15861
rect 45002 15852 45008 15864
rect 45060 15852 45066 15904
rect 1104 15802 48852 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 48852 15802
rect 1104 15728 48852 15750
rect 4706 15648 4712 15700
rect 4764 15688 4770 15700
rect 5077 15691 5135 15697
rect 5077 15688 5089 15691
rect 4764 15660 5089 15688
rect 4764 15648 4770 15660
rect 5077 15657 5089 15660
rect 5123 15657 5135 15691
rect 7650 15688 7656 15700
rect 7611 15660 7656 15688
rect 5077 15651 5135 15657
rect 7650 15648 7656 15660
rect 7708 15648 7714 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 9766 15688 9772 15700
rect 9539 15660 9772 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9766 15648 9772 15660
rect 9824 15648 9830 15700
rect 10781 15691 10839 15697
rect 10781 15657 10793 15691
rect 10827 15688 10839 15691
rect 10870 15688 10876 15700
rect 10827 15660 10876 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 11790 15688 11796 15700
rect 11751 15660 11796 15688
rect 11790 15648 11796 15660
rect 11848 15648 11854 15700
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 12897 15691 12955 15697
rect 12897 15688 12909 15691
rect 12584 15660 12909 15688
rect 12584 15648 12590 15660
rect 12897 15657 12909 15660
rect 12943 15657 12955 15691
rect 14274 15688 14280 15700
rect 14235 15660 14280 15688
rect 12897 15651 12955 15657
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 22554 15688 22560 15700
rect 22515 15660 22560 15688
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 23750 15688 23756 15700
rect 23711 15660 23756 15688
rect 23750 15648 23756 15660
rect 23808 15648 23814 15700
rect 26050 15688 26056 15700
rect 26011 15660 26056 15688
rect 26050 15648 26056 15660
rect 26108 15648 26114 15700
rect 28905 15691 28963 15697
rect 28905 15657 28917 15691
rect 28951 15688 28963 15691
rect 29730 15688 29736 15700
rect 28951 15660 29736 15688
rect 28951 15657 28963 15660
rect 28905 15651 28963 15657
rect 29730 15648 29736 15660
rect 29788 15648 29794 15700
rect 31941 15691 31999 15697
rect 31941 15657 31953 15691
rect 31987 15688 31999 15691
rect 32214 15688 32220 15700
rect 31987 15660 32220 15688
rect 31987 15657 31999 15660
rect 31941 15651 31999 15657
rect 32214 15648 32220 15660
rect 32272 15648 32278 15700
rect 35299 15691 35357 15697
rect 35299 15657 35311 15691
rect 35345 15688 35357 15691
rect 36446 15688 36452 15700
rect 35345 15660 36452 15688
rect 35345 15657 35357 15660
rect 35299 15651 35357 15657
rect 36446 15648 36452 15660
rect 36504 15648 36510 15700
rect 36538 15648 36544 15700
rect 36596 15688 36602 15700
rect 37001 15691 37059 15697
rect 37001 15688 37013 15691
rect 36596 15660 37013 15688
rect 36596 15648 36602 15660
rect 37001 15657 37013 15660
rect 37047 15657 37059 15691
rect 37458 15688 37464 15700
rect 37419 15660 37464 15688
rect 37001 15651 37059 15657
rect 37458 15648 37464 15660
rect 37516 15648 37522 15700
rect 37826 15648 37832 15700
rect 37884 15688 37890 15700
rect 37921 15691 37979 15697
rect 37921 15688 37933 15691
rect 37884 15660 37933 15688
rect 37884 15648 37890 15660
rect 37921 15657 37933 15660
rect 37967 15657 37979 15691
rect 38562 15688 38568 15700
rect 38523 15660 38568 15688
rect 37921 15651 37979 15657
rect 38562 15648 38568 15660
rect 38620 15648 38626 15700
rect 42058 15648 42064 15700
rect 42116 15688 42122 15700
rect 42245 15691 42303 15697
rect 42245 15688 42257 15691
rect 42116 15660 42257 15688
rect 42116 15648 42122 15660
rect 42245 15657 42257 15660
rect 42291 15657 42303 15691
rect 43162 15688 43168 15700
rect 43123 15660 43168 15688
rect 42245 15651 42303 15657
rect 43162 15648 43168 15660
rect 43220 15648 43226 15700
rect 44082 15648 44088 15700
rect 44140 15688 44146 15700
rect 44361 15691 44419 15697
rect 44361 15688 44373 15691
rect 44140 15660 44373 15688
rect 44140 15648 44146 15660
rect 44361 15657 44373 15660
rect 44407 15657 44419 15691
rect 44361 15651 44419 15657
rect 3694 15580 3700 15632
rect 3752 15620 3758 15632
rect 4614 15620 4620 15632
rect 3752 15592 4620 15620
rect 3752 15580 3758 15592
rect 3878 15512 3884 15564
rect 3936 15552 3942 15564
rect 4540 15561 4568 15592
rect 4614 15580 4620 15592
rect 4672 15580 4678 15632
rect 6454 15580 6460 15632
rect 6512 15620 6518 15632
rect 6727 15623 6785 15629
rect 6727 15620 6739 15623
rect 6512 15592 6739 15620
rect 6512 15580 6518 15592
rect 6727 15589 6739 15592
rect 6773 15620 6785 15623
rect 7668 15620 7696 15648
rect 9858 15620 9864 15632
rect 6773 15592 7696 15620
rect 9819 15592 9864 15620
rect 6773 15589 6785 15592
rect 6727 15583 6785 15589
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 13443 15623 13501 15629
rect 13443 15589 13455 15623
rect 13489 15620 13501 15623
rect 13538 15620 13544 15632
rect 13489 15592 13544 15620
rect 13489 15589 13501 15592
rect 13443 15583 13501 15589
rect 13538 15580 13544 15592
rect 13596 15580 13602 15632
rect 15838 15620 15844 15632
rect 15799 15592 15844 15620
rect 15838 15580 15844 15592
rect 15896 15580 15902 15632
rect 15930 15580 15936 15632
rect 15988 15620 15994 15632
rect 17957 15623 18015 15629
rect 15988 15592 16033 15620
rect 15988 15580 15994 15592
rect 17957 15589 17969 15623
rect 18003 15620 18015 15623
rect 18046 15620 18052 15632
rect 18003 15592 18052 15620
rect 18003 15589 18015 15592
rect 17957 15583 18015 15589
rect 18046 15580 18052 15592
rect 18104 15580 18110 15632
rect 19886 15620 19892 15632
rect 18800 15592 19564 15620
rect 19847 15592 19892 15620
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 3936 15524 4077 15552
rect 3936 15512 3942 15524
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15521 4583 15555
rect 6362 15552 6368 15564
rect 6323 15524 6368 15552
rect 4525 15515 4583 15521
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 8180 15555 8238 15561
rect 8180 15521 8192 15555
rect 8226 15552 8238 15555
rect 8478 15552 8484 15564
rect 8226 15524 8484 15552
rect 8226 15521 8238 15524
rect 8180 15515 8238 15521
rect 8478 15512 8484 15524
rect 8536 15512 8542 15564
rect 12136 15555 12194 15561
rect 12136 15521 12148 15555
rect 12182 15552 12194 15555
rect 12250 15552 12256 15564
rect 12182 15524 12256 15552
rect 12182 15521 12194 15524
rect 12136 15515 12194 15521
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15552 13139 15555
rect 13170 15552 13176 15564
rect 13127 15524 13176 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 13170 15512 13176 15524
rect 13228 15512 13234 15564
rect 18141 15555 18199 15561
rect 18141 15521 18153 15555
rect 18187 15552 18199 15555
rect 18230 15552 18236 15564
rect 18187 15524 18236 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 18230 15512 18236 15524
rect 18288 15552 18294 15564
rect 18598 15552 18604 15564
rect 18288 15524 18604 15552
rect 18288 15512 18294 15524
rect 18598 15512 18604 15524
rect 18656 15552 18662 15564
rect 18800 15561 18828 15592
rect 18785 15555 18843 15561
rect 18785 15552 18797 15555
rect 18656 15524 18797 15552
rect 18656 15512 18662 15524
rect 18785 15521 18797 15524
rect 18831 15521 18843 15555
rect 19334 15552 19340 15564
rect 19295 15524 19340 15552
rect 18785 15515 18843 15521
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 19536 15561 19564 15592
rect 19886 15580 19892 15592
rect 19944 15580 19950 15632
rect 22833 15623 22891 15629
rect 22833 15589 22845 15623
rect 22879 15620 22891 15623
rect 23198 15620 23204 15632
rect 22879 15592 23204 15620
rect 22879 15589 22891 15592
rect 22833 15583 22891 15589
rect 23198 15580 23204 15592
rect 23256 15580 23262 15632
rect 24118 15580 24124 15632
rect 24176 15620 24182 15632
rect 24305 15623 24363 15629
rect 24305 15620 24317 15623
rect 24176 15592 24317 15620
rect 24176 15580 24182 15592
rect 24305 15589 24317 15592
rect 24351 15589 24363 15623
rect 24305 15583 24363 15589
rect 24397 15623 24455 15629
rect 24397 15589 24409 15623
rect 24443 15620 24455 15623
rect 25314 15620 25320 15632
rect 24443 15592 25320 15620
rect 24443 15589 24455 15592
rect 24397 15583 24455 15589
rect 25314 15580 25320 15592
rect 25372 15580 25378 15632
rect 26326 15580 26332 15632
rect 26384 15620 26390 15632
rect 26834 15623 26892 15629
rect 26834 15620 26846 15623
rect 26384 15592 26846 15620
rect 26384 15580 26390 15592
rect 26834 15589 26846 15592
rect 26880 15589 26892 15623
rect 29270 15620 29276 15632
rect 29231 15592 29276 15620
rect 26834 15583 26892 15589
rect 29270 15580 29276 15592
rect 29328 15580 29334 15632
rect 31570 15580 31576 15632
rect 31628 15620 31634 15632
rect 32030 15620 32036 15632
rect 31628 15592 32036 15620
rect 31628 15580 31634 15592
rect 32030 15580 32036 15592
rect 32088 15620 32094 15632
rect 32309 15623 32367 15629
rect 32309 15620 32321 15623
rect 32088 15592 32321 15620
rect 32088 15580 32094 15592
rect 32309 15589 32321 15592
rect 32355 15589 32367 15623
rect 32309 15583 32367 15589
rect 32582 15580 32588 15632
rect 32640 15620 32646 15632
rect 32861 15623 32919 15629
rect 32861 15620 32873 15623
rect 32640 15592 32873 15620
rect 32640 15580 32646 15592
rect 32861 15589 32873 15592
rect 32907 15589 32919 15623
rect 41046 15620 41052 15632
rect 41007 15592 41052 15620
rect 32861 15583 32919 15589
rect 41046 15580 41052 15592
rect 41104 15580 41110 15632
rect 43533 15623 43591 15629
rect 43533 15589 43545 15623
rect 43579 15620 43591 15623
rect 43622 15620 43628 15632
rect 43579 15592 43628 15620
rect 43579 15589 43591 15592
rect 43533 15583 43591 15589
rect 43622 15580 43628 15592
rect 43680 15580 43686 15632
rect 19521 15555 19579 15561
rect 19521 15521 19533 15555
rect 19567 15521 19579 15555
rect 19521 15515 19579 15521
rect 21637 15555 21695 15561
rect 21637 15521 21649 15555
rect 21683 15552 21695 15555
rect 21726 15552 21732 15564
rect 21683 15524 21732 15552
rect 21683 15521 21695 15524
rect 21637 15515 21695 15521
rect 21726 15512 21732 15524
rect 21784 15512 21790 15564
rect 26513 15555 26571 15561
rect 26513 15521 26525 15555
rect 26559 15552 26571 15555
rect 26602 15552 26608 15564
rect 26559 15524 26608 15552
rect 26559 15521 26571 15524
rect 26513 15515 26571 15521
rect 26602 15512 26608 15524
rect 26660 15512 26666 15564
rect 30834 15512 30840 15564
rect 30892 15552 30898 15564
rect 31056 15555 31114 15561
rect 31056 15552 31068 15555
rect 30892 15524 31068 15552
rect 30892 15512 30898 15524
rect 31056 15521 31068 15524
rect 31102 15521 31114 15555
rect 34146 15552 34152 15564
rect 34107 15524 34152 15552
rect 31056 15515 31114 15521
rect 34146 15512 34152 15524
rect 34204 15512 34210 15564
rect 34606 15512 34612 15564
rect 34664 15552 34670 15564
rect 35066 15552 35072 15564
rect 34664 15524 35072 15552
rect 34664 15512 34670 15524
rect 35066 15512 35072 15524
rect 35124 15512 35130 15564
rect 36173 15555 36231 15561
rect 36173 15521 36185 15555
rect 36219 15552 36231 15555
rect 36262 15552 36268 15564
rect 36219 15524 36268 15552
rect 36219 15521 36231 15524
rect 36173 15515 36231 15521
rect 36262 15512 36268 15524
rect 36320 15512 36326 15564
rect 38194 15512 38200 15564
rect 38252 15552 38258 15564
rect 38289 15555 38347 15561
rect 38289 15552 38301 15555
rect 38252 15524 38301 15552
rect 38252 15512 38258 15524
rect 38289 15521 38301 15524
rect 38335 15521 38347 15555
rect 38746 15552 38752 15564
rect 38707 15524 38752 15552
rect 38289 15515 38347 15521
rect 38746 15512 38752 15524
rect 38804 15552 38810 15564
rect 39482 15552 39488 15564
rect 38804 15524 39488 15552
rect 38804 15512 38810 15524
rect 39482 15512 39488 15524
rect 39540 15552 39546 15564
rect 39853 15555 39911 15561
rect 39853 15552 39865 15555
rect 39540 15524 39865 15552
rect 39540 15512 39546 15524
rect 39853 15521 39865 15524
rect 39899 15521 39911 15555
rect 39853 15515 39911 15521
rect 44818 15512 44824 15564
rect 44876 15552 44882 15564
rect 44948 15555 45006 15561
rect 44948 15552 44960 15555
rect 44876 15524 44960 15552
rect 44876 15512 44882 15524
rect 44948 15521 44960 15524
rect 44994 15521 45006 15555
rect 44948 15515 45006 15521
rect 4614 15484 4620 15496
rect 4575 15456 4620 15484
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15453 9827 15487
rect 10042 15484 10048 15496
rect 10003 15456 10048 15484
rect 9769 15447 9827 15453
rect 8251 15419 8309 15425
rect 8251 15385 8263 15419
rect 8297 15416 8309 15419
rect 9784 15416 9812 15447
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 15436 15456 16129 15484
rect 15436 15444 15442 15456
rect 16117 15453 16129 15456
rect 16163 15484 16175 15487
rect 16666 15484 16672 15496
rect 16163 15456 16672 15484
rect 16163 15453 16175 15456
rect 16117 15447 16175 15453
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 22738 15484 22744 15496
rect 22699 15456 22744 15484
rect 22738 15444 22744 15456
rect 22796 15444 22802 15496
rect 23382 15484 23388 15496
rect 23343 15456 23388 15484
rect 23382 15444 23388 15456
rect 23440 15444 23446 15496
rect 24578 15484 24584 15496
rect 24539 15456 24584 15484
rect 24578 15444 24584 15456
rect 24636 15444 24642 15496
rect 29181 15487 29239 15493
rect 29181 15453 29193 15487
rect 29227 15484 29239 15487
rect 29362 15484 29368 15496
rect 29227 15456 29368 15484
rect 29227 15453 29239 15456
rect 29181 15447 29239 15453
rect 29362 15444 29368 15456
rect 29420 15444 29426 15496
rect 31938 15444 31944 15496
rect 31996 15484 32002 15496
rect 32217 15487 32275 15493
rect 32217 15484 32229 15487
rect 31996 15456 32229 15484
rect 31996 15444 32002 15456
rect 32217 15453 32229 15456
rect 32263 15484 32275 15487
rect 32950 15484 32956 15496
rect 32263 15456 32956 15484
rect 32263 15453 32275 15456
rect 32217 15447 32275 15453
rect 32950 15444 32956 15456
rect 33008 15444 33014 15496
rect 33321 15487 33379 15493
rect 33321 15453 33333 15487
rect 33367 15484 33379 15487
rect 33502 15484 33508 15496
rect 33367 15456 33508 15484
rect 33367 15453 33379 15456
rect 33321 15447 33379 15453
rect 33502 15444 33508 15456
rect 33560 15484 33566 15496
rect 38212 15484 38240 15512
rect 40954 15484 40960 15496
rect 33560 15456 38240 15484
rect 40915 15456 40960 15484
rect 33560 15444 33566 15456
rect 40954 15444 40960 15456
rect 41012 15444 41018 15496
rect 43441 15487 43499 15493
rect 43441 15453 43453 15487
rect 43487 15484 43499 15487
rect 44450 15484 44456 15496
rect 43487 15456 44456 15484
rect 43487 15453 43499 15456
rect 43441 15447 43499 15453
rect 44450 15444 44456 15456
rect 44508 15484 44514 15496
rect 45051 15487 45109 15493
rect 45051 15484 45063 15487
rect 44508 15456 45063 15484
rect 44508 15444 44514 15456
rect 45051 15453 45063 15456
rect 45097 15453 45109 15487
rect 45051 15447 45109 15453
rect 10134 15416 10140 15428
rect 8297 15388 10140 15416
rect 8297 15385 8309 15388
rect 8251 15379 8309 15385
rect 10134 15376 10140 15388
rect 10192 15376 10198 15428
rect 11514 15376 11520 15428
rect 11572 15416 11578 15428
rect 29733 15419 29791 15425
rect 11572 15388 15654 15416
rect 11572 15376 11578 15388
rect 7285 15351 7343 15357
rect 7285 15317 7297 15351
rect 7331 15348 7343 15351
rect 7558 15348 7564 15360
rect 7331 15320 7564 15348
rect 7331 15317 7343 15320
rect 7285 15311 7343 15317
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 8846 15348 8852 15360
rect 8807 15320 8852 15348
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 12066 15308 12072 15360
rect 12124 15348 12130 15360
rect 12207 15351 12265 15357
rect 12207 15348 12219 15351
rect 12124 15320 12219 15348
rect 12124 15308 12130 15320
rect 12207 15317 12219 15320
rect 12253 15317 12265 15351
rect 12526 15348 12532 15360
rect 12487 15320 12532 15348
rect 12207 15311 12265 15317
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 13998 15348 14004 15360
rect 13959 15320 14004 15348
rect 13998 15308 14004 15320
rect 14056 15308 14062 15360
rect 15626 15348 15654 15388
rect 29733 15385 29745 15419
rect 29779 15416 29791 15419
rect 32582 15416 32588 15428
rect 29779 15388 32588 15416
rect 29779 15385 29791 15388
rect 29733 15379 29791 15385
rect 32582 15376 32588 15388
rect 32640 15376 32646 15428
rect 41509 15419 41567 15425
rect 41509 15385 41521 15419
rect 41555 15416 41567 15419
rect 43714 15416 43720 15428
rect 41555 15388 43720 15416
rect 41555 15385 41567 15388
rect 41509 15379 41567 15385
rect 43714 15376 43720 15388
rect 43772 15416 43778 15428
rect 43993 15419 44051 15425
rect 43993 15416 44005 15419
rect 43772 15388 44005 15416
rect 43772 15376 43778 15388
rect 43993 15385 44005 15388
rect 44039 15385 44051 15419
rect 43993 15379 44051 15385
rect 18233 15351 18291 15357
rect 18233 15348 18245 15351
rect 15626 15320 18245 15348
rect 18233 15317 18245 15320
rect 18279 15317 18291 15351
rect 18233 15311 18291 15317
rect 21775 15351 21833 15357
rect 21775 15317 21787 15351
rect 21821 15348 21833 15351
rect 22370 15348 22376 15360
rect 21821 15320 22376 15348
rect 21821 15317 21833 15320
rect 21775 15311 21833 15317
rect 22370 15308 22376 15320
rect 22428 15308 22434 15360
rect 25222 15348 25228 15360
rect 25183 15320 25228 15348
rect 25222 15308 25228 15320
rect 25280 15308 25286 15360
rect 26878 15308 26884 15360
rect 26936 15348 26942 15360
rect 27433 15351 27491 15357
rect 27433 15348 27445 15351
rect 26936 15320 27445 15348
rect 26936 15308 26942 15320
rect 27433 15317 27445 15320
rect 27479 15317 27491 15351
rect 27433 15311 27491 15317
rect 31159 15351 31217 15357
rect 31159 15317 31171 15351
rect 31205 15348 31217 15351
rect 31754 15348 31760 15360
rect 31205 15320 31760 15348
rect 31205 15317 31217 15320
rect 31159 15311 31217 15317
rect 31754 15308 31760 15320
rect 31812 15308 31818 15360
rect 34287 15351 34345 15357
rect 34287 15317 34299 15351
rect 34333 15348 34345 15351
rect 34790 15348 34796 15360
rect 34333 15320 34796 15348
rect 34333 15317 34345 15320
rect 34287 15311 34345 15317
rect 34790 15308 34796 15320
rect 34848 15308 34854 15360
rect 34977 15351 35035 15357
rect 34977 15317 34989 15351
rect 35023 15348 35035 15351
rect 35342 15348 35348 15360
rect 35023 15320 35348 15348
rect 35023 15317 35035 15320
rect 34977 15311 35035 15317
rect 35342 15308 35348 15320
rect 35400 15308 35406 15360
rect 36311 15351 36369 15357
rect 36311 15317 36323 15351
rect 36357 15348 36369 15351
rect 36538 15348 36544 15360
rect 36357 15320 36544 15348
rect 36357 15317 36369 15320
rect 36311 15311 36369 15317
rect 36538 15308 36544 15320
rect 36596 15308 36602 15360
rect 36630 15308 36636 15360
rect 36688 15348 36694 15360
rect 40034 15348 40040 15360
rect 36688 15320 36733 15348
rect 39995 15320 40040 15348
rect 36688 15308 36694 15320
rect 40034 15308 40040 15320
rect 40092 15308 40098 15360
rect 40586 15348 40592 15360
rect 40547 15320 40592 15348
rect 40586 15308 40592 15320
rect 40644 15308 40650 15360
rect 1104 15258 48852 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 48852 15258
rect 1104 15184 48852 15206
rect 3605 15147 3663 15153
rect 3605 15113 3617 15147
rect 3651 15144 3663 15147
rect 3694 15144 3700 15156
rect 3651 15116 3700 15144
rect 3651 15113 3663 15116
rect 3605 15107 3663 15113
rect 3694 15104 3700 15116
rect 3752 15104 3758 15156
rect 3878 15144 3884 15156
rect 3839 15116 3884 15144
rect 3878 15104 3884 15116
rect 3936 15104 3942 15156
rect 6089 15147 6147 15153
rect 6089 15113 6101 15147
rect 6135 15144 6147 15147
rect 6270 15144 6276 15156
rect 6135 15116 6276 15144
rect 6135 15113 6147 15116
rect 6089 15107 6147 15113
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 8205 15147 8263 15153
rect 8205 15113 8217 15147
rect 8251 15144 8263 15147
rect 8478 15144 8484 15156
rect 8251 15116 8484 15144
rect 8251 15113 8263 15116
rect 8205 15107 8263 15113
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 10134 15144 10140 15156
rect 10095 15116 10140 15144
rect 10134 15104 10140 15116
rect 10192 15104 10198 15156
rect 11885 15147 11943 15153
rect 11885 15113 11897 15147
rect 11931 15144 11943 15147
rect 12250 15144 12256 15156
rect 11931 15116 12256 15144
rect 11931 15113 11943 15116
rect 11885 15107 11943 15113
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 13170 15104 13176 15156
rect 13228 15144 13234 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 13228 15116 13829 15144
rect 13228 15104 13234 15116
rect 13817 15113 13829 15116
rect 13863 15113 13875 15147
rect 13817 15107 13875 15113
rect 17865 15147 17923 15153
rect 17865 15113 17877 15147
rect 17911 15144 17923 15147
rect 18046 15144 18052 15156
rect 17911 15116 18052 15144
rect 17911 15113 17923 15116
rect 17865 15107 17923 15113
rect 18046 15104 18052 15116
rect 18104 15104 18110 15156
rect 18598 15144 18604 15156
rect 18559 15116 18604 15144
rect 18598 15104 18604 15116
rect 18656 15144 18662 15156
rect 19337 15147 19395 15153
rect 19337 15144 19349 15147
rect 18656 15116 19349 15144
rect 18656 15104 18662 15116
rect 19337 15113 19349 15116
rect 19383 15113 19395 15147
rect 19337 15107 19395 15113
rect 22281 15147 22339 15153
rect 22281 15113 22293 15147
rect 22327 15144 22339 15147
rect 22738 15144 22744 15156
rect 22327 15116 22744 15144
rect 22327 15113 22339 15116
rect 22281 15107 22339 15113
rect 22738 15104 22744 15116
rect 22796 15144 22802 15156
rect 23937 15147 23995 15153
rect 23937 15144 23949 15147
rect 22796 15116 23949 15144
rect 22796 15104 22802 15116
rect 23937 15113 23949 15116
rect 23983 15113 23995 15147
rect 23937 15107 23995 15113
rect 26602 15104 26608 15156
rect 26660 15144 26666 15156
rect 27709 15147 27767 15153
rect 27709 15144 27721 15147
rect 26660 15116 27721 15144
rect 26660 15104 26666 15116
rect 27709 15113 27721 15116
rect 27755 15113 27767 15147
rect 27709 15107 27767 15113
rect 28353 15147 28411 15153
rect 28353 15113 28365 15147
rect 28399 15144 28411 15147
rect 29362 15144 29368 15156
rect 28399 15116 29368 15144
rect 28399 15113 28411 15116
rect 28353 15107 28411 15113
rect 29362 15104 29368 15116
rect 29420 15104 29426 15156
rect 30834 15104 30840 15156
rect 30892 15144 30898 15156
rect 31021 15147 31079 15153
rect 31021 15144 31033 15147
rect 30892 15116 31033 15144
rect 30892 15104 30898 15116
rect 31021 15113 31033 15116
rect 31067 15113 31079 15147
rect 31021 15107 31079 15113
rect 7098 15036 7104 15088
rect 7156 15076 7162 15088
rect 9677 15079 9735 15085
rect 9677 15076 9689 15079
rect 7156 15048 9689 15076
rect 7156 15036 7162 15048
rect 9677 15045 9689 15048
rect 9723 15076 9735 15079
rect 9858 15076 9864 15088
rect 9723 15048 9864 15076
rect 9723 15045 9735 15048
rect 9677 15039 9735 15045
rect 9858 15036 9864 15048
rect 9916 15036 9922 15088
rect 12434 15036 12440 15088
rect 12492 15076 12498 15088
rect 12492 15048 12848 15076
rect 12492 15036 12498 15048
rect 4433 15011 4491 15017
rect 4433 14977 4445 15011
rect 4479 15008 4491 15011
rect 4614 15008 4620 15020
rect 4479 14980 4620 15008
rect 4479 14977 4491 14980
rect 4433 14971 4491 14977
rect 4614 14968 4620 14980
rect 4672 15008 4678 15020
rect 5629 15011 5687 15017
rect 5629 15008 5641 15011
rect 4672 14980 5641 15008
rect 4672 14968 4678 14980
rect 5629 14977 5641 14980
rect 5675 14977 5687 15011
rect 6454 15008 6460 15020
rect 6415 14980 6460 15008
rect 5629 14971 5687 14977
rect 6454 14968 6460 14980
rect 6512 14968 6518 15020
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 15008 9551 15011
rect 10042 15008 10048 15020
rect 9539 14980 10048 15008
rect 9539 14977 9551 14980
rect 9493 14971 9551 14977
rect 10042 14968 10048 14980
rect 10100 14968 10106 15020
rect 10781 15011 10839 15017
rect 10781 14977 10793 15011
rect 10827 15008 10839 15011
rect 10870 15008 10876 15020
rect 10827 14980 10876 15008
rect 10827 14977 10839 14980
rect 10781 14971 10839 14977
rect 10870 14968 10876 14980
rect 10928 14968 10934 15020
rect 11146 15008 11152 15020
rect 11107 14980 11152 15008
rect 11146 14968 11152 14980
rect 11204 14968 11210 15020
rect 12526 15008 12532 15020
rect 12487 14980 12532 15008
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 12820 15017 12848 15048
rect 16942 15036 16948 15088
rect 17000 15076 17006 15088
rect 18233 15079 18291 15085
rect 18233 15076 18245 15079
rect 17000 15048 18245 15076
rect 17000 15036 17006 15048
rect 18233 15045 18245 15048
rect 18279 15045 18291 15079
rect 18233 15039 18291 15045
rect 22511 15079 22569 15085
rect 22511 15045 22523 15079
rect 22557 15076 22569 15079
rect 23750 15076 23756 15088
rect 22557 15048 23756 15076
rect 22557 15045 22569 15048
rect 22511 15039 22569 15045
rect 23750 15036 23756 15048
rect 23808 15036 23814 15088
rect 23842 15036 23848 15088
rect 23900 15076 23906 15088
rect 26237 15079 26295 15085
rect 26237 15076 26249 15079
rect 23900 15048 26249 15076
rect 23900 15036 23906 15048
rect 26237 15045 26249 15048
rect 26283 15076 26295 15079
rect 26878 15076 26884 15088
rect 26283 15048 26884 15076
rect 26283 15045 26295 15048
rect 26237 15039 26295 15045
rect 26878 15036 26884 15048
rect 26936 15036 26942 15088
rect 28721 15079 28779 15085
rect 28721 15045 28733 15079
rect 28767 15076 28779 15079
rect 29270 15076 29276 15088
rect 28767 15048 29276 15076
rect 28767 15045 28779 15048
rect 28721 15039 28779 15045
rect 29270 15036 29276 15048
rect 29328 15036 29334 15088
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 14977 12863 15011
rect 15102 15008 15108 15020
rect 15063 14980 15108 15008
rect 12805 14971 12863 14977
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 15470 14968 15476 15020
rect 15528 15008 15534 15020
rect 16390 15008 16396 15020
rect 15528 14980 16396 15008
rect 15528 14968 15534 14980
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 16666 15008 16672 15020
rect 16627 14980 16672 15008
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 15008 19119 15011
rect 19334 15008 19340 15020
rect 19107 14980 19340 15008
rect 19107 14977 19119 14980
rect 19061 14971 19119 14977
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 23290 15008 23296 15020
rect 23251 14980 23296 15008
rect 23290 14968 23296 14980
rect 23348 14968 23354 15020
rect 23385 15011 23443 15017
rect 23385 14977 23397 15011
rect 23431 15008 23443 15011
rect 24026 15008 24032 15020
rect 23431 14980 24032 15008
rect 23431 14977 23443 14980
rect 23385 14971 23443 14977
rect 24026 14968 24032 14980
rect 24084 14968 24090 15020
rect 25222 15008 25228 15020
rect 25183 14980 25228 15008
rect 25222 14968 25228 14980
rect 25280 14968 25286 15020
rect 25866 15008 25872 15020
rect 25779 14980 25872 15008
rect 25866 14968 25872 14980
rect 25924 15008 25930 15020
rect 27065 15011 27123 15017
rect 27065 15008 27077 15011
rect 25924 14980 27077 15008
rect 25924 14968 25930 14980
rect 27065 14977 27077 14980
rect 27111 14977 27123 15011
rect 31036 15008 31064 15107
rect 31662 15104 31668 15156
rect 31720 15144 31726 15156
rect 31849 15147 31907 15153
rect 31849 15144 31861 15147
rect 31720 15116 31861 15144
rect 31720 15104 31726 15116
rect 31849 15113 31861 15116
rect 31895 15113 31907 15147
rect 31849 15107 31907 15113
rect 32030 15104 32036 15156
rect 32088 15144 32094 15156
rect 32217 15147 32275 15153
rect 32217 15144 32229 15147
rect 32088 15116 32229 15144
rect 32088 15104 32094 15116
rect 32217 15113 32229 15116
rect 32263 15113 32275 15147
rect 32217 15107 32275 15113
rect 33134 15104 33140 15156
rect 33192 15144 33198 15156
rect 33229 15147 33287 15153
rect 33229 15144 33241 15147
rect 33192 15116 33241 15144
rect 33192 15104 33198 15116
rect 33229 15113 33241 15116
rect 33275 15113 33287 15147
rect 33229 15107 33287 15113
rect 31036 14980 31800 15008
rect 27065 14971 27123 14977
rect 5810 14900 5816 14952
rect 5868 14940 5874 14952
rect 6860 14943 6918 14949
rect 6860 14940 6872 14943
rect 5868 14912 6872 14940
rect 5868 14900 5874 14912
rect 6860 14909 6872 14912
rect 6906 14940 6918 14943
rect 7285 14943 7343 14949
rect 7285 14940 7297 14943
rect 6906 14912 7297 14940
rect 6906 14909 6918 14912
rect 6860 14903 6918 14909
rect 7285 14909 7297 14912
rect 7331 14909 7343 14943
rect 7285 14903 7343 14909
rect 13354 14900 13360 14952
rect 13412 14940 13418 14952
rect 18049 14943 18107 14949
rect 13412 14912 14688 14940
rect 13412 14900 13418 14912
rect 4341 14875 4399 14881
rect 4341 14841 4353 14875
rect 4387 14872 4399 14875
rect 4795 14875 4853 14881
rect 4795 14872 4807 14875
rect 4387 14844 4807 14872
rect 4387 14841 4399 14844
rect 4341 14835 4399 14841
rect 4795 14841 4807 14844
rect 4841 14872 4853 14875
rect 4982 14872 4988 14884
rect 4841 14844 4988 14872
rect 4841 14841 4853 14844
rect 4795 14835 4853 14841
rect 4982 14832 4988 14844
rect 5040 14832 5046 14884
rect 8846 14872 8852 14884
rect 8807 14844 8852 14872
rect 8846 14832 8852 14844
rect 8904 14832 8910 14884
rect 8941 14875 8999 14881
rect 8941 14841 8953 14875
rect 8987 14872 8999 14875
rect 10594 14872 10600 14884
rect 8987 14844 10600 14872
rect 8987 14841 8999 14844
rect 8941 14835 8999 14841
rect 5350 14804 5356 14816
rect 5311 14776 5356 14804
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 6914 14764 6920 14816
rect 6972 14804 6978 14816
rect 7101 14807 7159 14813
rect 7101 14804 7113 14807
rect 6972 14776 7113 14804
rect 6972 14764 6978 14776
rect 7101 14773 7113 14776
rect 7147 14773 7159 14807
rect 7101 14767 7159 14773
rect 8478 14764 8484 14816
rect 8536 14804 8542 14816
rect 8573 14807 8631 14813
rect 8573 14804 8585 14807
rect 8536 14776 8585 14804
rect 8536 14764 8542 14776
rect 8573 14773 8585 14776
rect 8619 14804 8631 14807
rect 8956 14804 8984 14835
rect 10594 14832 10600 14844
rect 10652 14832 10658 14884
rect 10873 14875 10931 14881
rect 10873 14841 10885 14875
rect 10919 14872 10931 14875
rect 12253 14875 12311 14881
rect 12253 14872 12265 14875
rect 10919 14844 12265 14872
rect 10919 14841 10931 14844
rect 10873 14835 10931 14841
rect 12253 14841 12265 14844
rect 12299 14872 12311 14875
rect 12621 14875 12679 14881
rect 12621 14872 12633 14875
rect 12299 14844 12633 14872
rect 12299 14841 12311 14844
rect 12253 14835 12311 14841
rect 12621 14841 12633 14844
rect 12667 14872 12679 14875
rect 13814 14872 13820 14884
rect 12667 14844 13820 14872
rect 12667 14841 12679 14844
rect 12621 14835 12679 14841
rect 8619 14776 8984 14804
rect 9677 14807 9735 14813
rect 8619 14773 8631 14776
rect 8573 14767 8631 14773
rect 9677 14773 9689 14807
rect 9723 14804 9735 14807
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9723 14776 9873 14804
rect 9723 14773 9735 14776
rect 9677 14767 9735 14773
rect 9861 14773 9873 14776
rect 9907 14804 9919 14807
rect 10505 14807 10563 14813
rect 10505 14804 10517 14807
rect 9907 14776 10517 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10505 14773 10517 14776
rect 10551 14804 10563 14807
rect 10888 14804 10916 14835
rect 13814 14832 13820 14844
rect 13872 14832 13878 14884
rect 13538 14804 13544 14816
rect 10551 14776 10916 14804
rect 13499 14776 13544 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 14660 14813 14688 14912
rect 18049 14909 18061 14943
rect 18095 14940 18107 14943
rect 18322 14940 18328 14952
rect 18095 14912 18328 14940
rect 18095 14909 18107 14912
rect 18049 14903 18107 14909
rect 18322 14900 18328 14912
rect 18380 14900 18386 14952
rect 19886 14940 19892 14952
rect 19847 14912 19892 14940
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 22440 14943 22498 14949
rect 22440 14909 22452 14943
rect 22486 14940 22498 14943
rect 22922 14940 22928 14952
rect 22486 14912 22928 14940
rect 22486 14909 22498 14912
rect 22440 14903 22498 14909
rect 22922 14900 22928 14912
rect 22980 14900 22986 14952
rect 23198 14900 23204 14952
rect 23256 14940 23262 14952
rect 23728 14943 23786 14949
rect 23728 14940 23740 14943
rect 23256 14912 23740 14940
rect 23256 14900 23262 14912
rect 23728 14909 23740 14912
rect 23774 14940 23786 14943
rect 24121 14943 24179 14949
rect 24121 14940 24133 14943
rect 23774 14912 24133 14940
rect 23774 14909 23786 14912
rect 23728 14903 23786 14909
rect 24121 14909 24133 14912
rect 24167 14909 24179 14943
rect 24121 14903 24179 14909
rect 28258 14900 28264 14952
rect 28316 14940 28322 14952
rect 29273 14943 29331 14949
rect 29273 14940 29285 14943
rect 28316 14912 29285 14940
rect 28316 14900 28322 14912
rect 29273 14909 29285 14912
rect 29319 14940 29331 14943
rect 30469 14943 30527 14949
rect 30469 14940 30481 14943
rect 29319 14912 30481 14940
rect 29319 14909 29331 14912
rect 29273 14903 29331 14909
rect 30469 14909 30481 14912
rect 30515 14909 30527 14943
rect 30469 14903 30527 14909
rect 30558 14900 30564 14952
rect 30616 14940 30622 14952
rect 31440 14943 31498 14949
rect 31440 14940 31452 14943
rect 30616 14912 31452 14940
rect 30616 14900 30622 14912
rect 31440 14909 31452 14912
rect 31486 14940 31498 14943
rect 31662 14940 31668 14952
rect 31486 14912 31668 14940
rect 31486 14909 31498 14912
rect 31440 14903 31498 14909
rect 31662 14900 31668 14912
rect 31720 14900 31726 14952
rect 31772 14940 31800 14980
rect 32436 14943 32494 14949
rect 32436 14940 32448 14943
rect 31772 14912 32448 14940
rect 32436 14909 32448 14912
rect 32482 14940 32494 14943
rect 32861 14943 32919 14949
rect 32861 14940 32873 14943
rect 32482 14912 32873 14940
rect 32482 14909 32494 14912
rect 32436 14903 32494 14909
rect 32861 14909 32873 14912
rect 32907 14940 32919 14943
rect 32950 14940 32956 14952
rect 32907 14912 32956 14940
rect 32907 14909 32919 14912
rect 32861 14903 32919 14909
rect 32950 14900 32956 14912
rect 33008 14900 33014 14952
rect 33244 14940 33272 15107
rect 33870 15104 33876 15156
rect 33928 15144 33934 15156
rect 37921 15147 37979 15153
rect 33928 15116 37596 15144
rect 33928 15104 33934 15116
rect 34606 15076 34612 15088
rect 34567 15048 34612 15076
rect 34606 15036 34612 15048
rect 34664 15036 34670 15088
rect 36262 15076 36268 15088
rect 36223 15048 36268 15076
rect 36262 15036 36268 15048
rect 36320 15036 36326 15088
rect 37461 15079 37519 15085
rect 37461 15076 37473 15079
rect 36556 15048 37473 15076
rect 36556 15020 36584 15048
rect 37461 15045 37473 15048
rect 37507 15045 37519 15079
rect 37461 15039 37519 15045
rect 35250 15008 35256 15020
rect 35211 14980 35256 15008
rect 35250 14968 35256 14980
rect 35308 14968 35314 15020
rect 36538 15008 36544 15020
rect 36499 14980 36544 15008
rect 36538 14968 36544 14980
rect 36596 14968 36602 15020
rect 36814 15008 36820 15020
rect 36775 14980 36820 15008
rect 36814 14968 36820 14980
rect 36872 14968 36878 15020
rect 37568 15008 37596 15116
rect 37921 15113 37933 15147
rect 37967 15144 37979 15147
rect 38746 15144 38752 15156
rect 37967 15116 38752 15144
rect 37967 15113 37979 15116
rect 37921 15107 37979 15113
rect 38746 15104 38752 15116
rect 38804 15144 38810 15156
rect 39853 15147 39911 15153
rect 39853 15144 39865 15147
rect 38804 15116 39865 15144
rect 38804 15104 38810 15116
rect 39853 15113 39865 15116
rect 39899 15113 39911 15147
rect 40310 15144 40316 15156
rect 40271 15116 40316 15144
rect 39853 15107 39911 15113
rect 40310 15104 40316 15116
rect 40368 15104 40374 15156
rect 42981 15147 43039 15153
rect 42981 15113 42993 15147
rect 43027 15144 43039 15147
rect 43257 15147 43315 15153
rect 43257 15144 43269 15147
rect 43027 15116 43269 15144
rect 43027 15113 43039 15116
rect 42981 15107 43039 15113
rect 43257 15113 43269 15116
rect 43303 15144 43315 15147
rect 43622 15144 43628 15156
rect 43303 15116 43628 15144
rect 43303 15113 43315 15116
rect 43257 15107 43315 15113
rect 43622 15104 43628 15116
rect 43680 15104 43686 15156
rect 44450 15144 44456 15156
rect 44411 15116 44456 15144
rect 44450 15104 44456 15116
rect 44508 15104 44514 15156
rect 38194 15076 38200 15088
rect 38155 15048 38200 15076
rect 38194 15036 38200 15048
rect 38252 15036 38258 15088
rect 38565 15011 38623 15017
rect 38565 15008 38577 15011
rect 37568 14980 38577 15008
rect 38565 14977 38577 14980
rect 38611 15008 38623 15011
rect 40586 15008 40592 15020
rect 38611 14980 38792 15008
rect 40499 14980 40592 15008
rect 38611 14977 38623 14980
rect 38565 14971 38623 14977
rect 38764 14949 38792 14980
rect 40586 14968 40592 14980
rect 40644 15008 40650 15020
rect 42199 15011 42257 15017
rect 42199 15008 42211 15011
rect 40644 14980 42211 15008
rect 40644 14968 40650 14980
rect 42199 14977 42211 14980
rect 42245 14977 42257 15011
rect 42199 14971 42257 14977
rect 44726 14968 44732 15020
rect 44784 15008 44790 15020
rect 44784 14980 45115 15008
rect 44784 14968 44790 14980
rect 33413 14943 33471 14949
rect 33413 14940 33425 14943
rect 33244 14912 33425 14940
rect 33413 14909 33425 14912
rect 33459 14909 33471 14943
rect 33413 14903 33471 14909
rect 38749 14943 38807 14949
rect 38749 14909 38761 14943
rect 38795 14909 38807 14943
rect 38749 14903 38807 14909
rect 39114 14900 39120 14952
rect 39172 14940 39178 14952
rect 39301 14943 39359 14949
rect 39301 14940 39313 14943
rect 39172 14912 39313 14940
rect 39172 14900 39178 14912
rect 39301 14909 39313 14912
rect 39347 14940 39359 14943
rect 40034 14940 40040 14952
rect 39347 14912 40040 14940
rect 39347 14909 39359 14912
rect 39301 14903 39359 14909
rect 40034 14900 40040 14912
rect 40092 14900 40098 14952
rect 42112 14943 42170 14949
rect 42112 14909 42124 14943
rect 42158 14940 42170 14943
rect 42518 14940 42524 14952
rect 42158 14912 42524 14940
rect 42158 14909 42170 14912
rect 42112 14903 42170 14909
rect 42518 14900 42524 14912
rect 42576 14900 42582 14952
rect 45087 14949 45115 14980
rect 45072 14943 45130 14949
rect 45072 14909 45084 14943
rect 45118 14940 45130 14943
rect 45465 14943 45523 14949
rect 45465 14940 45477 14943
rect 45118 14912 45477 14940
rect 45118 14909 45130 14912
rect 45072 14903 45130 14909
rect 45465 14909 45477 14912
rect 45511 14909 45523 14943
rect 45465 14903 45523 14909
rect 14826 14872 14832 14884
rect 14787 14844 14832 14872
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 14921 14875 14979 14881
rect 14921 14841 14933 14875
rect 14967 14841 14979 14875
rect 14921 14835 14979 14841
rect 16209 14875 16267 14881
rect 16209 14841 16221 14875
rect 16255 14872 16267 14875
rect 16485 14875 16543 14881
rect 16485 14872 16497 14875
rect 16255 14844 16497 14872
rect 16255 14841 16267 14844
rect 16209 14835 16267 14841
rect 16485 14841 16497 14844
rect 16531 14872 16543 14875
rect 16850 14872 16856 14884
rect 16531 14844 16856 14872
rect 16531 14841 16543 14844
rect 16485 14835 16543 14841
rect 14645 14807 14703 14813
rect 14645 14773 14657 14807
rect 14691 14804 14703 14807
rect 14936 14804 14964 14835
rect 16850 14832 16856 14844
rect 16908 14832 16914 14884
rect 19797 14875 19855 14881
rect 19797 14841 19809 14875
rect 19843 14872 19855 14875
rect 20070 14872 20076 14884
rect 19843 14844 20076 14872
rect 19843 14841 19855 14844
rect 19797 14835 19855 14841
rect 20070 14832 20076 14844
rect 20128 14872 20134 14884
rect 20210 14875 20268 14881
rect 20210 14872 20222 14875
rect 20128 14844 20222 14872
rect 20128 14832 20134 14844
rect 20210 14841 20222 14844
rect 20256 14841 20268 14875
rect 20210 14835 20268 14841
rect 23290 14832 23296 14884
rect 23348 14872 23354 14884
rect 24581 14875 24639 14881
rect 24581 14872 24593 14875
rect 23348 14844 24593 14872
rect 23348 14832 23354 14844
rect 24581 14841 24593 14844
rect 24627 14872 24639 14875
rect 25041 14875 25099 14881
rect 25041 14872 25053 14875
rect 24627 14844 25053 14872
rect 24627 14841 24639 14844
rect 24581 14835 24639 14841
rect 25041 14841 25053 14844
rect 25087 14872 25099 14875
rect 25314 14872 25320 14884
rect 25087 14844 25320 14872
rect 25087 14841 25099 14844
rect 25041 14835 25099 14841
rect 25314 14832 25320 14844
rect 25372 14832 25378 14884
rect 26786 14872 26792 14884
rect 26747 14844 26792 14872
rect 26786 14832 26792 14844
rect 26844 14832 26850 14884
rect 26878 14832 26884 14884
rect 26936 14872 26942 14884
rect 29594 14875 29652 14881
rect 26936 14844 26981 14872
rect 26936 14832 26942 14844
rect 29594 14841 29606 14875
rect 29640 14872 29652 14875
rect 30282 14872 30288 14884
rect 29640 14844 30288 14872
rect 29640 14841 29652 14844
rect 29594 14835 29652 14841
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 14691 14776 15853 14804
rect 14691 14773 14703 14776
rect 14645 14767 14703 14773
rect 15841 14773 15853 14776
rect 15887 14804 15899 14807
rect 15930 14804 15936 14816
rect 15887 14776 15936 14804
rect 15887 14773 15899 14776
rect 15841 14767 15899 14773
rect 15930 14764 15936 14776
rect 15988 14764 15994 14816
rect 20806 14804 20812 14816
rect 20767 14776 20812 14804
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 21726 14804 21732 14816
rect 21639 14776 21732 14804
rect 21726 14764 21732 14776
rect 21784 14804 21790 14816
rect 23385 14807 23443 14813
rect 23385 14804 23397 14807
rect 21784 14776 23397 14804
rect 21784 14764 21790 14776
rect 23385 14773 23397 14776
rect 23431 14773 23443 14807
rect 23385 14767 23443 14773
rect 26326 14764 26332 14816
rect 26384 14804 26390 14816
rect 26513 14807 26571 14813
rect 26513 14804 26525 14807
rect 26384 14776 26525 14804
rect 26384 14764 26390 14776
rect 26513 14773 26525 14776
rect 26559 14804 26571 14807
rect 28997 14807 29055 14813
rect 28997 14804 29009 14807
rect 26559 14776 29009 14804
rect 26559 14773 26571 14776
rect 26513 14767 26571 14773
rect 28997 14773 29009 14776
rect 29043 14804 29055 14807
rect 29609 14804 29637 14835
rect 30282 14832 30288 14844
rect 30340 14832 30346 14884
rect 31527 14875 31585 14881
rect 31527 14841 31539 14875
rect 31573 14872 31585 14875
rect 34974 14872 34980 14884
rect 31573 14844 34980 14872
rect 31573 14841 31585 14844
rect 31527 14835 31585 14841
rect 34974 14832 34980 14844
rect 35032 14832 35038 14884
rect 35069 14875 35127 14881
rect 35069 14841 35081 14875
rect 35115 14872 35127 14875
rect 35342 14872 35348 14884
rect 35115 14844 35348 14872
rect 35115 14841 35127 14844
rect 35069 14835 35127 14841
rect 35342 14832 35348 14844
rect 35400 14872 35406 14884
rect 36630 14872 36636 14884
rect 35400 14844 36636 14872
rect 35400 14832 35406 14844
rect 36630 14832 36636 14844
rect 36688 14832 36694 14884
rect 39485 14875 39543 14881
rect 39485 14841 39497 14875
rect 39531 14872 39543 14875
rect 39574 14872 39580 14884
rect 39531 14844 39580 14872
rect 39531 14841 39543 14844
rect 39485 14835 39543 14841
rect 39574 14832 39580 14844
rect 39632 14832 39638 14884
rect 40310 14832 40316 14884
rect 40368 14872 40374 14884
rect 40681 14875 40739 14881
rect 40681 14872 40693 14875
rect 40368 14844 40693 14872
rect 40368 14832 40374 14844
rect 40681 14841 40693 14844
rect 40727 14841 40739 14875
rect 40681 14835 40739 14841
rect 41233 14875 41291 14881
rect 41233 14841 41245 14875
rect 41279 14872 41291 14875
rect 41690 14872 41696 14884
rect 41279 14844 41696 14872
rect 41279 14841 41291 14844
rect 41233 14835 41291 14841
rect 30190 14804 30196 14816
rect 29043 14776 29637 14804
rect 30151 14776 30196 14804
rect 29043 14773 29055 14776
rect 28997 14767 29055 14773
rect 30190 14764 30196 14776
rect 30248 14764 30254 14816
rect 32539 14807 32597 14813
rect 32539 14773 32551 14807
rect 32585 14804 32597 14807
rect 32674 14804 32680 14816
rect 32585 14776 32680 14804
rect 32585 14773 32597 14776
rect 32539 14767 32597 14773
rect 32674 14764 32680 14776
rect 32732 14764 32738 14816
rect 33597 14807 33655 14813
rect 33597 14773 33609 14807
rect 33643 14804 33655 14807
rect 33962 14804 33968 14816
rect 33643 14776 33968 14804
rect 33643 14773 33655 14776
rect 33597 14767 33655 14773
rect 33962 14764 33968 14776
rect 34020 14764 34026 14816
rect 34146 14804 34152 14816
rect 34107 14776 34152 14804
rect 34146 14764 34152 14776
rect 34204 14764 34210 14816
rect 40696 14804 40724 14835
rect 41690 14832 41696 14844
rect 41748 14832 41754 14884
rect 43530 14872 43536 14884
rect 43491 14844 43536 14872
rect 43530 14832 43536 14844
rect 43588 14832 43594 14884
rect 43622 14832 43628 14884
rect 43680 14872 43686 14884
rect 44174 14872 44180 14884
rect 43680 14844 43725 14872
rect 44135 14844 44180 14872
rect 43680 14832 43686 14844
rect 44174 14832 44180 14844
rect 44232 14832 44238 14884
rect 44818 14872 44824 14884
rect 44731 14844 44824 14872
rect 44818 14832 44824 14844
rect 44876 14872 44882 14884
rect 46934 14872 46940 14884
rect 44876 14844 46940 14872
rect 44876 14832 44882 14844
rect 46934 14832 46940 14844
rect 46992 14832 46998 14884
rect 41509 14807 41567 14813
rect 41509 14804 41521 14807
rect 40696 14776 41521 14804
rect 41509 14773 41521 14776
rect 41555 14773 41567 14807
rect 41509 14767 41567 14773
rect 44910 14764 44916 14816
rect 44968 14804 44974 14816
rect 45143 14807 45201 14813
rect 45143 14804 45155 14807
rect 44968 14776 45155 14804
rect 44968 14764 44974 14776
rect 45143 14773 45155 14776
rect 45189 14773 45201 14807
rect 45143 14767 45201 14773
rect 1104 14714 48852 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 48852 14714
rect 1104 14640 48852 14662
rect 6822 14560 6828 14612
rect 6880 14600 6886 14612
rect 6880 14572 7052 14600
rect 6880 14560 6886 14572
rect 4795 14535 4853 14541
rect 4795 14501 4807 14535
rect 4841 14532 4853 14535
rect 4982 14532 4988 14544
rect 4841 14504 4988 14532
rect 4841 14501 4853 14504
rect 4795 14495 4853 14501
rect 4982 14492 4988 14504
rect 5040 14492 5046 14544
rect 7024 14541 7052 14572
rect 12066 14560 12072 14612
rect 12124 14600 12130 14612
rect 14826 14600 14832 14612
rect 12124 14572 12204 14600
rect 14787 14572 14832 14600
rect 12124 14560 12130 14572
rect 7009 14535 7067 14541
rect 7009 14501 7021 14535
rect 7055 14501 7067 14535
rect 10502 14532 10508 14544
rect 10463 14504 10508 14532
rect 7009 14495 7067 14501
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 10594 14492 10600 14544
rect 10652 14532 10658 14544
rect 11146 14532 11152 14544
rect 10652 14504 10697 14532
rect 11107 14504 11152 14532
rect 10652 14492 10658 14504
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 12176 14541 12204 14572
rect 14826 14560 14832 14572
rect 14884 14600 14890 14612
rect 15427 14603 15485 14609
rect 15427 14600 15439 14603
rect 14884 14572 15439 14600
rect 14884 14560 14890 14572
rect 15427 14569 15439 14572
rect 15473 14569 15485 14603
rect 15838 14600 15844 14612
rect 15799 14572 15844 14600
rect 15427 14563 15485 14569
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 16390 14600 16396 14612
rect 16351 14572 16396 14600
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 18141 14603 18199 14609
rect 18141 14569 18153 14603
rect 18187 14600 18199 14603
rect 18322 14600 18328 14612
rect 18187 14572 18328 14600
rect 18187 14569 18199 14572
rect 18141 14563 18199 14569
rect 18322 14560 18328 14572
rect 18380 14560 18386 14612
rect 23014 14560 23020 14612
rect 23072 14600 23078 14612
rect 23290 14600 23296 14612
rect 23072 14572 23296 14600
rect 23072 14560 23078 14572
rect 23290 14560 23296 14572
rect 23348 14560 23354 14612
rect 24210 14600 24216 14612
rect 24171 14572 24216 14600
rect 24210 14560 24216 14572
rect 24268 14560 24274 14612
rect 24995 14603 25053 14609
rect 24995 14569 25007 14603
rect 25041 14600 25053 14603
rect 25222 14600 25228 14612
rect 25041 14572 25228 14600
rect 25041 14569 25053 14572
rect 24995 14563 25053 14569
rect 25222 14560 25228 14572
rect 25280 14560 25286 14612
rect 27338 14560 27344 14612
rect 27396 14600 27402 14612
rect 31159 14603 31217 14609
rect 27396 14572 27568 14600
rect 27396 14560 27402 14572
rect 12161 14535 12219 14541
rect 12161 14501 12173 14535
rect 12207 14501 12219 14535
rect 12161 14495 12219 14501
rect 12250 14492 12256 14544
rect 12308 14532 12314 14544
rect 13354 14532 13360 14544
rect 12308 14504 13360 14532
rect 12308 14492 12314 14504
rect 13354 14492 13360 14504
rect 13412 14492 13418 14544
rect 13814 14532 13820 14544
rect 13775 14504 13820 14532
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 14369 14535 14427 14541
rect 14369 14501 14381 14535
rect 14415 14532 14427 14535
rect 15102 14532 15108 14544
rect 14415 14504 15108 14532
rect 14415 14501 14427 14504
rect 14369 14495 14427 14501
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 16850 14532 16856 14544
rect 16811 14504 16856 14532
rect 16850 14492 16856 14504
rect 16908 14492 16914 14544
rect 19797 14535 19855 14541
rect 19797 14501 19809 14535
rect 19843 14532 19855 14535
rect 19886 14532 19892 14544
rect 19843 14504 19892 14532
rect 19843 14501 19855 14504
rect 19797 14495 19855 14501
rect 19886 14492 19892 14504
rect 19944 14532 19950 14544
rect 20073 14535 20131 14541
rect 20073 14532 20085 14535
rect 19944 14504 20085 14532
rect 19944 14492 19950 14504
rect 20073 14501 20085 14504
rect 20119 14501 20131 14535
rect 20073 14495 20131 14501
rect 20806 14492 20812 14544
rect 20864 14532 20870 14544
rect 21085 14535 21143 14541
rect 21085 14532 21097 14535
rect 20864 14504 21097 14532
rect 20864 14492 20870 14504
rect 21085 14501 21097 14504
rect 21131 14501 21143 14535
rect 21085 14495 21143 14501
rect 22370 14492 22376 14544
rect 22428 14532 22434 14544
rect 22741 14535 22799 14541
rect 22741 14532 22753 14535
rect 22428 14504 22753 14532
rect 22428 14492 22434 14504
rect 22741 14501 22753 14504
rect 22787 14501 22799 14535
rect 22741 14495 22799 14501
rect 22830 14492 22836 14544
rect 22888 14532 22894 14544
rect 23382 14532 23388 14544
rect 22888 14504 22933 14532
rect 23343 14504 23388 14532
rect 22888 14492 22894 14504
rect 23382 14492 23388 14504
rect 23440 14492 23446 14544
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 4126 14436 4445 14464
rect 3694 14356 3700 14408
rect 3752 14396 3758 14408
rect 4126 14396 4154 14436
rect 4433 14433 4445 14436
rect 4479 14464 4491 14467
rect 4890 14464 4896 14476
rect 4479 14436 4896 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 8424 14467 8482 14473
rect 8424 14464 8436 14467
rect 7616 14436 8436 14464
rect 7616 14424 7622 14436
rect 8424 14433 8436 14436
rect 8470 14464 8482 14467
rect 8849 14467 8907 14473
rect 8849 14464 8861 14467
rect 8470 14436 8861 14464
rect 8470 14433 8482 14436
rect 8424 14427 8482 14433
rect 8849 14433 8861 14436
rect 8895 14433 8907 14467
rect 8849 14427 8907 14433
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15324 14467 15382 14473
rect 15324 14464 15336 14467
rect 15252 14436 15336 14464
rect 15252 14424 15258 14436
rect 15324 14433 15336 14436
rect 15370 14433 15382 14467
rect 15324 14427 15382 14433
rect 6914 14396 6920 14408
rect 3752 14368 4154 14396
rect 6875 14368 6920 14396
rect 3752 14356 3758 14368
rect 6914 14356 6920 14368
rect 6972 14356 6978 14408
rect 12434 14396 12440 14408
rect 12395 14368 12440 14396
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 13722 14396 13728 14408
rect 13683 14368 13728 14396
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 16868 14396 16896 14492
rect 17218 14464 17224 14476
rect 17179 14436 17224 14464
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 18782 14424 18788 14476
rect 18840 14464 18846 14476
rect 19061 14467 19119 14473
rect 19061 14464 19073 14467
rect 18840 14436 19073 14464
rect 18840 14424 18846 14436
rect 19061 14433 19073 14436
rect 19107 14433 19119 14467
rect 19061 14427 19119 14433
rect 19613 14467 19671 14473
rect 19613 14433 19625 14467
rect 19659 14464 19671 14467
rect 20162 14464 20168 14476
rect 19659 14436 20168 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 24946 14473 24952 14476
rect 24924 14467 24952 14473
rect 24924 14464 24936 14467
rect 24859 14436 24936 14464
rect 24924 14433 24936 14436
rect 25004 14464 25010 14476
rect 26418 14464 26424 14476
rect 25004 14436 25544 14464
rect 26379 14436 26424 14464
rect 24924 14427 24952 14433
rect 24946 14424 24952 14427
rect 25004 14424 25010 14436
rect 13872 14368 16896 14396
rect 13872 14356 13878 14368
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20993 14399 21051 14405
rect 20993 14396 21005 14399
rect 20404 14368 21005 14396
rect 20404 14356 20410 14368
rect 20993 14365 21005 14368
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 7466 14328 7472 14340
rect 7427 14300 7472 14328
rect 7466 14288 7472 14300
rect 7524 14328 7530 14340
rect 10045 14331 10103 14337
rect 10045 14328 10057 14331
rect 7524 14300 10057 14328
rect 7524 14288 7530 14300
rect 10045 14297 10057 14300
rect 10091 14328 10103 14331
rect 10134 14328 10140 14340
rect 10091 14300 10140 14328
rect 10091 14297 10103 14300
rect 10045 14291 10103 14297
rect 10134 14288 10140 14300
rect 10192 14288 10198 14340
rect 21542 14328 21548 14340
rect 21503 14300 21548 14328
rect 21542 14288 21548 14300
rect 21600 14288 21606 14340
rect 25516 14328 25544 14436
rect 26418 14424 26424 14436
rect 26476 14424 26482 14476
rect 26651 14467 26709 14473
rect 26651 14433 26663 14467
rect 26697 14464 26709 14467
rect 26786 14464 26792 14476
rect 26697 14436 26792 14464
rect 26697 14433 26709 14436
rect 26651 14427 26709 14433
rect 26786 14424 26792 14436
rect 26844 14464 26850 14476
rect 27540 14473 27568 14572
rect 31159 14569 31171 14603
rect 31205 14600 31217 14603
rect 34057 14603 34115 14609
rect 34057 14600 34069 14603
rect 31205 14572 34069 14600
rect 31205 14569 31217 14572
rect 31159 14563 31217 14569
rect 34057 14569 34069 14572
rect 34103 14600 34115 14603
rect 39114 14600 39120 14612
rect 34103 14572 34376 14600
rect 39075 14572 39120 14600
rect 34103 14569 34115 14572
rect 34057 14563 34115 14569
rect 28258 14532 28264 14544
rect 28219 14504 28264 14532
rect 28258 14492 28264 14504
rect 28316 14492 28322 14544
rect 29270 14532 29276 14544
rect 29183 14504 29276 14532
rect 29270 14492 29276 14504
rect 29328 14532 29334 14544
rect 30190 14532 30196 14544
rect 29328 14504 30196 14532
rect 29328 14492 29334 14504
rect 30190 14492 30196 14504
rect 30248 14492 30254 14544
rect 31478 14532 31484 14544
rect 31439 14504 31484 14532
rect 31478 14492 31484 14504
rect 31536 14492 31542 14544
rect 31754 14492 31760 14544
rect 31812 14532 31818 14544
rect 32217 14535 32275 14541
rect 32217 14532 32229 14535
rect 31812 14504 32229 14532
rect 31812 14492 31818 14504
rect 32217 14501 32229 14504
rect 32263 14501 32275 14535
rect 32217 14495 32275 14501
rect 32309 14535 32367 14541
rect 32309 14501 32321 14535
rect 32355 14532 32367 14535
rect 32398 14532 32404 14544
rect 32355 14504 32404 14532
rect 32355 14501 32367 14504
rect 32309 14495 32367 14501
rect 32398 14492 32404 14504
rect 32456 14492 32462 14544
rect 34348 14541 34376 14572
rect 39114 14560 39120 14572
rect 39172 14560 39178 14612
rect 42610 14600 42616 14612
rect 39954 14572 42616 14600
rect 34333 14535 34391 14541
rect 34333 14501 34345 14535
rect 34379 14501 34391 14535
rect 34333 14495 34391 14501
rect 34422 14492 34428 14544
rect 34480 14532 34486 14544
rect 34977 14535 35035 14541
rect 34480 14504 34525 14532
rect 34480 14492 34486 14504
rect 34977 14501 34989 14535
rect 35023 14532 35035 14535
rect 35250 14532 35256 14544
rect 35023 14504 35256 14532
rect 35023 14501 35035 14504
rect 34977 14495 35035 14501
rect 35250 14492 35256 14504
rect 35308 14492 35314 14544
rect 36262 14532 36268 14544
rect 36223 14504 36268 14532
rect 36262 14492 36268 14504
rect 36320 14492 36326 14544
rect 36814 14532 36820 14544
rect 36775 14504 36820 14532
rect 36814 14492 36820 14504
rect 36872 14492 36878 14544
rect 39666 14492 39672 14544
rect 39724 14532 39730 14544
rect 39954 14541 39982 14572
rect 42610 14560 42616 14572
rect 42668 14560 42674 14612
rect 43530 14560 43536 14612
rect 43588 14600 43594 14612
rect 43901 14603 43959 14609
rect 43901 14600 43913 14603
rect 43588 14572 43913 14600
rect 43588 14560 43594 14572
rect 43901 14569 43913 14572
rect 43947 14600 43959 14603
rect 44910 14600 44916 14612
rect 43947 14572 44916 14600
rect 43947 14569 43959 14572
rect 43901 14563 43959 14569
rect 44910 14560 44916 14572
rect 44968 14560 44974 14612
rect 39939 14535 39997 14541
rect 39939 14532 39951 14535
rect 39724 14504 39951 14532
rect 39724 14492 39730 14504
rect 39939 14501 39951 14504
rect 39985 14501 39997 14535
rect 39939 14495 39997 14501
rect 41414 14492 41420 14544
rect 41472 14532 41478 14544
rect 41693 14535 41751 14541
rect 41693 14532 41705 14535
rect 41472 14504 41705 14532
rect 41472 14492 41478 14504
rect 41693 14501 41705 14504
rect 41739 14501 41751 14535
rect 42242 14532 42248 14544
rect 42203 14504 42248 14532
rect 41693 14495 41751 14501
rect 42242 14492 42248 14504
rect 42300 14492 42306 14544
rect 27341 14467 27399 14473
rect 27341 14464 27353 14467
rect 26844 14436 27353 14464
rect 26844 14424 26850 14436
rect 27341 14433 27353 14436
rect 27387 14433 27399 14467
rect 27341 14427 27399 14433
rect 27525 14467 27583 14473
rect 27525 14433 27537 14467
rect 27571 14433 27583 14467
rect 28074 14464 28080 14476
rect 27987 14436 28080 14464
rect 27525 14427 27583 14433
rect 28074 14424 28080 14436
rect 28132 14464 28138 14476
rect 28994 14464 29000 14476
rect 28132 14436 29000 14464
rect 28132 14424 28138 14436
rect 28994 14424 29000 14436
rect 29052 14424 29058 14476
rect 31088 14467 31146 14473
rect 31088 14433 31100 14467
rect 31134 14464 31146 14467
rect 31294 14464 31300 14476
rect 31134 14436 31300 14464
rect 31134 14433 31146 14436
rect 31088 14427 31146 14433
rect 31294 14424 31300 14436
rect 31352 14424 31358 14476
rect 31938 14464 31944 14476
rect 31899 14436 31944 14464
rect 31938 14424 31944 14436
rect 31996 14424 32002 14476
rect 38703 14467 38761 14473
rect 38703 14433 38715 14467
rect 38749 14464 38761 14467
rect 40865 14467 40923 14473
rect 40865 14464 40877 14467
rect 38749 14436 40877 14464
rect 38749 14433 38761 14436
rect 38703 14427 38761 14433
rect 40865 14433 40877 14436
rect 40911 14464 40923 14467
rect 40954 14464 40960 14476
rect 40911 14436 40960 14464
rect 40911 14433 40923 14436
rect 40865 14427 40923 14433
rect 40954 14424 40960 14436
rect 41012 14424 41018 14476
rect 43416 14467 43474 14473
rect 43416 14433 43428 14467
rect 43462 14464 43474 14467
rect 43530 14464 43536 14476
rect 43462 14436 43536 14464
rect 43462 14433 43474 14436
rect 43416 14427 43474 14433
rect 43530 14424 43536 14436
rect 43588 14424 43594 14476
rect 29178 14396 29184 14408
rect 29139 14368 29184 14396
rect 29178 14356 29184 14368
rect 29236 14356 29242 14408
rect 29825 14399 29883 14405
rect 29825 14365 29837 14399
rect 29871 14396 29883 14399
rect 31846 14396 31852 14408
rect 29871 14368 31852 14396
rect 29871 14365 29883 14368
rect 29825 14359 29883 14365
rect 31846 14356 31852 14368
rect 31904 14396 31910 14408
rect 32490 14396 32496 14408
rect 31904 14368 32496 14396
rect 31904 14356 31910 14368
rect 32490 14356 32496 14368
rect 32548 14356 32554 14408
rect 32674 14356 32680 14408
rect 32732 14396 32738 14408
rect 32732 14368 33134 14396
rect 32732 14356 32738 14368
rect 30834 14328 30840 14340
rect 25516 14300 30840 14328
rect 30834 14288 30840 14300
rect 30892 14288 30898 14340
rect 33106 14328 33134 14368
rect 34974 14356 34980 14408
rect 35032 14396 35038 14408
rect 35253 14399 35311 14405
rect 35253 14396 35265 14399
rect 35032 14368 35265 14396
rect 35032 14356 35038 14368
rect 35253 14365 35265 14368
rect 35299 14365 35311 14399
rect 35253 14359 35311 14365
rect 36173 14399 36231 14405
rect 36173 14365 36185 14399
rect 36219 14365 36231 14399
rect 39574 14396 39580 14408
rect 39535 14368 39580 14396
rect 36173 14359 36231 14365
rect 36188 14328 36216 14359
rect 39574 14356 39580 14368
rect 39632 14356 39638 14408
rect 41601 14399 41659 14405
rect 41601 14396 41613 14399
rect 41340 14368 41613 14396
rect 37642 14328 37648 14340
rect 33106 14300 37648 14328
rect 37642 14288 37648 14300
rect 37700 14288 37706 14340
rect 41340 14272 41368 14368
rect 41601 14365 41613 14368
rect 41647 14365 41659 14399
rect 41601 14359 41659 14365
rect 5353 14263 5411 14269
rect 5353 14229 5365 14263
rect 5399 14260 5411 14263
rect 5534 14260 5540 14272
rect 5399 14232 5540 14260
rect 5399 14229 5411 14232
rect 5353 14223 5411 14229
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 8527 14263 8585 14269
rect 8527 14229 8539 14263
rect 8573 14260 8585 14263
rect 8662 14260 8668 14272
rect 8573 14232 8668 14260
rect 8573 14229 8585 14232
rect 8527 14223 8585 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 25314 14260 25320 14272
rect 25275 14232 25320 14260
rect 25314 14220 25320 14232
rect 25372 14220 25378 14272
rect 26970 14260 26976 14272
rect 26931 14232 26976 14260
rect 26970 14220 26976 14232
rect 27028 14220 27034 14272
rect 31294 14220 31300 14272
rect 31352 14260 31358 14272
rect 32858 14260 32864 14272
rect 31352 14232 32864 14260
rect 31352 14220 31358 14232
rect 32858 14220 32864 14232
rect 32916 14260 32922 14272
rect 38473 14263 38531 14269
rect 38473 14260 38485 14263
rect 32916 14232 38485 14260
rect 32916 14220 32922 14232
rect 38473 14229 38485 14232
rect 38519 14260 38531 14263
rect 39206 14260 39212 14272
rect 38519 14232 39212 14260
rect 38519 14229 38531 14232
rect 38473 14223 38531 14229
rect 39206 14220 39212 14232
rect 39264 14220 39270 14272
rect 40494 14260 40500 14272
rect 40455 14232 40500 14260
rect 40494 14220 40500 14232
rect 40552 14220 40558 14272
rect 41322 14260 41328 14272
rect 41283 14232 41328 14260
rect 41322 14220 41328 14232
rect 41380 14220 41386 14272
rect 42978 14220 42984 14272
rect 43036 14260 43042 14272
rect 43487 14263 43545 14269
rect 43487 14260 43499 14263
rect 43036 14232 43499 14260
rect 43036 14220 43042 14232
rect 43487 14229 43499 14232
rect 43533 14229 43545 14263
rect 43487 14223 43545 14229
rect 1104 14170 48852 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 48852 14170
rect 1104 14096 48852 14118
rect 3694 14056 3700 14068
rect 3655 14028 3700 14056
rect 3694 14016 3700 14028
rect 3752 14016 3758 14068
rect 4062 14056 4068 14068
rect 3975 14028 4068 14056
rect 4062 14016 4068 14028
rect 4120 14056 4126 14068
rect 4120 14028 4568 14056
rect 4120 14016 4126 14028
rect 4540 13929 4568 14028
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 6972 14028 7849 14056
rect 6972 14016 6978 14028
rect 7837 14025 7849 14028
rect 7883 14025 7895 14059
rect 7837 14019 7895 14025
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 11149 14059 11207 14065
rect 11149 14056 11161 14059
rect 10652 14028 11161 14056
rect 10652 14016 10658 14028
rect 11149 14025 11161 14028
rect 11195 14056 11207 14059
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11195 14028 12173 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 12161 14025 12173 14028
rect 12207 14056 12219 14059
rect 12250 14056 12256 14068
rect 12207 14028 12256 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12713 14059 12771 14065
rect 12713 14056 12725 14059
rect 12584 14028 12725 14056
rect 12584 14016 12590 14028
rect 12713 14025 12725 14028
rect 12759 14025 12771 14059
rect 12713 14019 12771 14025
rect 13357 14059 13415 14065
rect 13357 14025 13369 14059
rect 13403 14056 13415 14059
rect 13587 14059 13645 14065
rect 13587 14056 13599 14059
rect 13403 14028 13599 14056
rect 13403 14025 13415 14028
rect 13357 14019 13415 14025
rect 13587 14025 13599 14028
rect 13633 14056 13645 14059
rect 13722 14056 13728 14068
rect 13633 14028 13728 14056
rect 13633 14025 13645 14028
rect 13587 14019 13645 14025
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 13909 14059 13967 14065
rect 13909 14056 13921 14059
rect 13872 14028 13921 14056
rect 13872 14016 13878 14028
rect 13909 14025 13921 14028
rect 13955 14025 13967 14059
rect 13909 14019 13967 14025
rect 13998 14016 14004 14068
rect 14056 14056 14062 14068
rect 14277 14059 14335 14065
rect 14277 14056 14289 14059
rect 14056 14028 14289 14056
rect 14056 14016 14062 14028
rect 14277 14025 14289 14028
rect 14323 14025 14335 14059
rect 14277 14019 14335 14025
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 15841 14059 15899 14065
rect 15841 14056 15853 14059
rect 15252 14028 15853 14056
rect 15252 14016 15258 14028
rect 15841 14025 15853 14028
rect 15887 14025 15899 14059
rect 15841 14019 15899 14025
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14056 20131 14059
rect 20162 14056 20168 14068
rect 20119 14028 20168 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 6822 13948 6828 14000
rect 6880 13988 6886 14000
rect 7466 13988 7472 14000
rect 6880 13960 7328 13988
rect 7427 13960 7472 13988
rect 6880 13948 6886 13960
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13889 4583 13923
rect 4525 13883 4583 13889
rect 6273 13923 6331 13929
rect 6273 13889 6285 13923
rect 6319 13920 6331 13923
rect 7098 13920 7104 13932
rect 6319 13892 7104 13920
rect 6319 13889 6331 13892
rect 6273 13883 6331 13889
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 7300 13920 7328 13960
rect 7466 13948 7472 13960
rect 7524 13948 7530 14000
rect 12066 13948 12072 14000
rect 12124 13988 12130 14000
rect 12897 13991 12955 13997
rect 12897 13988 12909 13991
rect 12124 13960 12909 13988
rect 12124 13948 12130 13960
rect 12897 13957 12909 13960
rect 12943 13957 12955 13991
rect 14016 13988 14044 14016
rect 12897 13951 12955 13957
rect 13786 13960 14044 13988
rect 8205 13923 8263 13929
rect 8205 13920 8217 13923
rect 7300 13892 8217 13920
rect 8205 13889 8217 13892
rect 8251 13889 8263 13923
rect 8205 13883 8263 13889
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13920 8539 13923
rect 8662 13920 8668 13932
rect 8527 13892 8668 13920
rect 8527 13889 8539 13892
rect 8481 13883 8539 13889
rect 4433 13855 4491 13861
rect 4433 13821 4445 13855
rect 4479 13852 4491 13855
rect 4614 13852 4620 13864
rect 4479 13824 4620 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 4614 13812 4620 13824
rect 4672 13852 4678 13864
rect 4982 13852 4988 13864
rect 4672 13824 4988 13852
rect 4672 13812 4678 13824
rect 4908 13793 4936 13824
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 4887 13787 4945 13793
rect 4887 13753 4899 13787
rect 4933 13753 4945 13787
rect 4887 13747 4945 13753
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 6917 13787 6975 13793
rect 6917 13784 6929 13787
rect 6788 13756 6929 13784
rect 6788 13744 6794 13756
rect 6917 13753 6929 13756
rect 6963 13753 6975 13787
rect 6917 13747 6975 13753
rect 7006 13744 7012 13796
rect 7064 13784 7070 13796
rect 8220 13784 8248 13883
rect 8662 13880 8668 13892
rect 8720 13920 8726 13932
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 8720 13892 9413 13920
rect 8720 13880 8726 13892
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 10134 13920 10140 13932
rect 10095 13892 10140 13920
rect 9401 13883 9459 13889
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 12504 13855 12562 13861
rect 12504 13821 12516 13855
rect 12550 13852 12562 13855
rect 12710 13852 12716 13864
rect 12550 13824 12716 13852
rect 12550 13821 12562 13824
rect 12504 13815 12562 13821
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 13500 13855 13558 13861
rect 13500 13821 13512 13855
rect 13546 13852 13558 13855
rect 13786 13852 13814 13960
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13920 14979 13923
rect 15102 13920 15108 13932
rect 14967 13892 15108 13920
rect 14967 13889 14979 13892
rect 14921 13883 14979 13889
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13920 16359 13923
rect 18509 13923 18567 13929
rect 16347 13892 17080 13920
rect 16347 13889 16359 13892
rect 16301 13883 16359 13889
rect 13546 13824 13814 13852
rect 13546 13821 13558 13824
rect 13500 13815 13558 13821
rect 15930 13812 15936 13864
rect 15988 13852 15994 13864
rect 17052 13861 17080 13892
rect 18509 13889 18521 13923
rect 18555 13920 18567 13923
rect 18555 13892 19472 13920
rect 18555 13889 18567 13892
rect 18509 13883 18567 13889
rect 19444 13864 19472 13892
rect 16393 13855 16451 13861
rect 16393 13852 16405 13855
rect 15988 13824 16405 13852
rect 15988 13812 15994 13824
rect 16393 13821 16405 13824
rect 16439 13821 16451 13855
rect 16393 13815 16451 13821
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13852 17095 13855
rect 17494 13852 17500 13864
rect 17083 13824 17500 13852
rect 17083 13821 17095 13824
rect 17037 13815 17095 13821
rect 17494 13812 17500 13824
rect 17552 13812 17558 13864
rect 18969 13855 19027 13861
rect 18969 13852 18981 13855
rect 18800 13824 18981 13852
rect 8478 13784 8484 13796
rect 7064 13756 7109 13784
rect 8220 13756 8484 13784
rect 7064 13744 7070 13756
rect 8478 13744 8484 13756
rect 8536 13784 8542 13796
rect 8573 13787 8631 13793
rect 8573 13784 8585 13787
rect 8536 13756 8585 13784
rect 8536 13744 8542 13756
rect 8573 13753 8585 13756
rect 8619 13753 8631 13787
rect 9122 13784 9128 13796
rect 9083 13756 9128 13784
rect 8573 13747 8631 13753
rect 9122 13744 9128 13756
rect 9180 13744 9186 13796
rect 10229 13787 10287 13793
rect 10229 13753 10241 13787
rect 10275 13753 10287 13787
rect 10229 13747 10287 13753
rect 10781 13787 10839 13793
rect 10781 13753 10793 13787
rect 10827 13784 10839 13787
rect 12986 13784 12992 13796
rect 10827 13756 12992 13784
rect 10827 13753 10839 13756
rect 10781 13747 10839 13753
rect 5442 13716 5448 13728
rect 5403 13688 5448 13716
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 6641 13719 6699 13725
rect 6641 13685 6653 13719
rect 6687 13716 6699 13719
rect 6822 13716 6828 13728
rect 6687 13688 6828 13716
rect 6687 13685 6699 13688
rect 6641 13679 6699 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 9950 13716 9956 13728
rect 9911 13688 9956 13716
rect 9950 13676 9956 13688
rect 10008 13716 10014 13728
rect 10244 13716 10272 13747
rect 12986 13744 12992 13756
rect 13044 13744 13050 13796
rect 14737 13787 14795 13793
rect 14737 13753 14749 13787
rect 14783 13784 14795 13787
rect 15013 13787 15071 13793
rect 15013 13784 15025 13787
rect 14783 13756 15025 13784
rect 14783 13753 14795 13756
rect 14737 13747 14795 13753
rect 15013 13753 15025 13756
rect 15059 13784 15071 13787
rect 15286 13784 15292 13796
rect 15059 13756 15292 13784
rect 15059 13753 15071 13756
rect 15013 13747 15071 13753
rect 15286 13744 15292 13756
rect 15344 13744 15350 13796
rect 15562 13784 15568 13796
rect 15523 13756 15568 13784
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 18690 13744 18696 13796
rect 18748 13784 18754 13796
rect 18800 13793 18828 13824
rect 18969 13821 18981 13824
rect 19015 13821 19027 13855
rect 18969 13815 19027 13821
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19484 13824 19533 13852
rect 19484 13812 19490 13824
rect 19521 13821 19533 13824
rect 19567 13852 19579 13855
rect 20088 13852 20116 14019
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 21361 14059 21419 14065
rect 21361 14056 21373 14059
rect 20864 14028 21373 14056
rect 20864 14016 20870 14028
rect 21361 14025 21373 14028
rect 21407 14025 21419 14059
rect 22370 14056 22376 14068
rect 22331 14028 22376 14056
rect 21361 14019 21419 14025
rect 22370 14016 22376 14028
rect 22428 14016 22434 14068
rect 23106 14056 23112 14068
rect 23067 14028 23112 14056
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 23477 14059 23535 14065
rect 23477 14056 23489 14059
rect 23216 14028 23489 14056
rect 20671 13991 20729 13997
rect 20671 13957 20683 13991
rect 20717 13988 20729 13991
rect 20898 13988 20904 14000
rect 20717 13960 20904 13988
rect 20717 13957 20729 13960
rect 20671 13951 20729 13957
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 21082 13988 21088 14000
rect 21043 13960 21088 13988
rect 21082 13948 21088 13960
rect 21140 13948 21146 14000
rect 22830 13948 22836 14000
rect 22888 13988 22894 14000
rect 23216 13988 23244 14028
rect 23477 14025 23489 14028
rect 23523 14056 23535 14059
rect 23842 14056 23848 14068
rect 23523 14028 23848 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 23842 14016 23848 14028
rect 23900 14016 23906 14068
rect 24946 14056 24952 14068
rect 24907 14028 24952 14056
rect 24946 14016 24952 14028
rect 25004 14016 25010 14068
rect 26418 14056 26424 14068
rect 26379 14028 26424 14056
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 27338 14016 27344 14068
rect 27396 14056 27402 14068
rect 27617 14059 27675 14065
rect 27617 14056 27629 14059
rect 27396 14028 27629 14056
rect 27396 14016 27402 14028
rect 27617 14025 27629 14028
rect 27663 14025 27675 14059
rect 28074 14056 28080 14068
rect 28035 14028 28080 14056
rect 27617 14019 27675 14025
rect 28074 14016 28080 14028
rect 28132 14016 28138 14068
rect 29178 14016 29184 14068
rect 29236 14056 29242 14068
rect 30653 14059 30711 14065
rect 30653 14056 30665 14059
rect 29236 14028 30665 14056
rect 29236 14016 29242 14028
rect 30653 14025 30665 14028
rect 30699 14025 30711 14059
rect 32306 14056 32312 14068
rect 30653 14019 30711 14025
rect 30852 14028 32312 14056
rect 29086 13988 29092 14000
rect 22888 13960 23244 13988
rect 23446 13960 28258 13988
rect 28999 13960 29092 13988
rect 22888 13948 22894 13960
rect 21100 13920 21128 13948
rect 20615 13892 21128 13920
rect 22097 13923 22155 13929
rect 20615 13861 20643 13892
rect 22097 13889 22109 13923
rect 22143 13920 22155 13923
rect 23446 13920 23474 13960
rect 22143 13892 23474 13920
rect 25133 13923 25191 13929
rect 22143 13889 22155 13892
rect 22097 13883 22155 13889
rect 25133 13889 25145 13923
rect 25179 13920 25191 13923
rect 25314 13920 25320 13932
rect 25179 13892 25320 13920
rect 25179 13889 25191 13892
rect 25133 13883 25191 13889
rect 19567 13824 20116 13852
rect 20584 13855 20643 13861
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 20584 13821 20596 13855
rect 20630 13824 20643 13855
rect 20630 13821 20642 13824
rect 20584 13815 20642 13821
rect 21450 13812 21456 13864
rect 21508 13852 21514 13864
rect 21612 13855 21670 13861
rect 21612 13852 21624 13855
rect 21508 13824 21624 13852
rect 21508 13812 21514 13824
rect 21612 13821 21624 13824
rect 21658 13852 21670 13855
rect 22112 13852 22140 13883
rect 25314 13880 25320 13892
rect 25372 13880 25378 13932
rect 25777 13923 25835 13929
rect 25777 13889 25789 13923
rect 25823 13920 25835 13923
rect 25866 13920 25872 13932
rect 25823 13892 25872 13920
rect 25823 13889 25835 13892
rect 25777 13883 25835 13889
rect 25866 13880 25872 13892
rect 25924 13880 25930 13932
rect 26145 13923 26203 13929
rect 26145 13889 26157 13923
rect 26191 13920 26203 13923
rect 27338 13920 27344 13932
rect 26191 13892 27344 13920
rect 26191 13889 26203 13892
rect 26145 13883 26203 13889
rect 21658 13824 22140 13852
rect 22624 13855 22682 13861
rect 21658 13821 21670 13824
rect 21612 13815 21670 13821
rect 22624 13821 22636 13855
rect 22670 13852 22682 13855
rect 23106 13852 23112 13864
rect 22670 13824 23112 13852
rect 22670 13821 22682 13824
rect 22624 13815 22682 13821
rect 23106 13812 23112 13824
rect 23164 13812 23170 13864
rect 26896 13861 26924 13892
rect 27338 13880 27344 13892
rect 27396 13880 27402 13932
rect 24096 13855 24154 13861
rect 24096 13821 24108 13855
rect 24142 13852 24154 13855
rect 26881 13855 26939 13861
rect 24142 13824 24624 13852
rect 24142 13821 24154 13824
rect 24096 13815 24154 13821
rect 18785 13787 18843 13793
rect 18785 13784 18797 13787
rect 18748 13756 18797 13784
rect 18748 13744 18754 13756
rect 18785 13753 18797 13756
rect 18831 13753 18843 13787
rect 18785 13747 18843 13753
rect 19705 13787 19763 13793
rect 19705 13753 19717 13787
rect 19751 13784 19763 13787
rect 20254 13784 20260 13796
rect 19751 13756 20260 13784
rect 19751 13753 19763 13756
rect 19705 13747 19763 13753
rect 20254 13744 20260 13756
rect 20312 13744 20318 13796
rect 24596 13793 24624 13824
rect 26881 13821 26893 13855
rect 26927 13821 26939 13855
rect 26881 13815 26939 13821
rect 26970 13812 26976 13864
rect 27028 13852 27034 13864
rect 28230 13861 28258 13960
rect 29086 13948 29092 13960
rect 29144 13988 29150 14000
rect 29270 13988 29276 14000
rect 29144 13960 29276 13988
rect 29144 13948 29150 13960
rect 29270 13948 29276 13960
rect 29328 13948 29334 14000
rect 29822 13948 29828 14000
rect 29880 13988 29886 14000
rect 29917 13991 29975 13997
rect 29917 13988 29929 13991
rect 29880 13960 29929 13988
rect 29880 13948 29886 13960
rect 29917 13957 29929 13960
rect 29963 13988 29975 13991
rect 30852 13988 30880 14028
rect 32306 14016 32312 14028
rect 32364 14016 32370 14068
rect 32398 14016 32404 14068
rect 32456 14056 32462 14068
rect 32493 14059 32551 14065
rect 32493 14056 32505 14059
rect 32456 14028 32505 14056
rect 32456 14016 32462 14028
rect 32493 14025 32505 14028
rect 32539 14056 32551 14059
rect 32861 14059 32919 14065
rect 32861 14056 32873 14059
rect 32539 14028 32873 14056
rect 32539 14025 32551 14028
rect 32493 14019 32551 14025
rect 32861 14025 32873 14028
rect 32907 14056 32919 14059
rect 33318 14056 33324 14068
rect 32907 14028 33324 14056
rect 32907 14025 32919 14028
rect 32861 14019 32919 14025
rect 33318 14016 33324 14028
rect 33376 14016 33382 14068
rect 34333 14059 34391 14065
rect 34333 14025 34345 14059
rect 34379 14056 34391 14059
rect 34422 14056 34428 14068
rect 34379 14028 34428 14056
rect 34379 14025 34391 14028
rect 34333 14019 34391 14025
rect 34422 14016 34428 14028
rect 34480 14056 34486 14068
rect 36081 14059 36139 14065
rect 36081 14056 36093 14059
rect 34480 14028 36093 14056
rect 34480 14016 34486 14028
rect 36081 14025 36093 14028
rect 36127 14056 36139 14059
rect 36262 14056 36268 14068
rect 36127 14028 36268 14056
rect 36127 14025 36139 14028
rect 36081 14019 36139 14025
rect 36262 14016 36268 14028
rect 36320 14016 36326 14068
rect 37642 14056 37648 14068
rect 37603 14028 37648 14056
rect 37642 14016 37648 14028
rect 37700 14016 37706 14068
rect 38105 14059 38163 14065
rect 38105 14025 38117 14059
rect 38151 14056 38163 14059
rect 38378 14056 38384 14068
rect 38151 14028 38384 14056
rect 38151 14025 38163 14028
rect 38105 14019 38163 14025
rect 29963 13960 30880 13988
rect 31113 13991 31171 13997
rect 29963 13957 29975 13960
rect 29917 13951 29975 13957
rect 31113 13957 31125 13991
rect 31159 13988 31171 13991
rect 31294 13988 31300 14000
rect 31159 13960 31300 13988
rect 31159 13957 31171 13960
rect 31113 13951 31171 13957
rect 31294 13948 31300 13960
rect 31352 13948 31358 14000
rect 31478 13948 31484 14000
rect 31536 13988 31542 14000
rect 31536 13960 31616 13988
rect 31536 13948 31542 13960
rect 31588 13929 31616 13960
rect 34514 13948 34520 14000
rect 34572 13988 34578 14000
rect 34609 13991 34667 13997
rect 34609 13988 34621 13991
rect 34572 13960 34621 13988
rect 34572 13948 34578 13960
rect 34609 13957 34621 13960
rect 34655 13957 34667 13991
rect 38120 13988 38148 14019
rect 38378 14016 38384 14028
rect 38436 14016 38442 14068
rect 39206 14056 39212 14068
rect 39167 14028 39212 14056
rect 39206 14016 39212 14028
rect 39264 14016 39270 14068
rect 39574 14016 39580 14068
rect 39632 14056 39638 14068
rect 39945 14059 40003 14065
rect 39945 14056 39957 14059
rect 39632 14028 39957 14056
rect 39632 14016 39638 14028
rect 39945 14025 39957 14028
rect 39991 14025 40003 14059
rect 39945 14019 40003 14025
rect 40635 14059 40693 14065
rect 40635 14025 40647 14059
rect 40681 14056 40693 14059
rect 41322 14056 41328 14068
rect 40681 14028 41328 14056
rect 40681 14025 40693 14028
rect 40635 14019 40693 14025
rect 41322 14016 41328 14028
rect 41380 14016 41386 14068
rect 42978 14056 42984 14068
rect 42766 14028 42984 14056
rect 34609 13951 34667 13957
rect 37384 13960 38148 13988
rect 28307 13923 28365 13929
rect 28307 13889 28319 13923
rect 28353 13920 28365 13923
rect 29365 13923 29423 13929
rect 29365 13920 29377 13923
rect 28353 13892 29377 13920
rect 28353 13889 28365 13892
rect 28307 13883 28365 13889
rect 29365 13889 29377 13892
rect 29411 13920 29423 13923
rect 30285 13923 30343 13929
rect 30285 13920 30297 13923
rect 29411 13892 30297 13920
rect 29411 13889 29423 13892
rect 29365 13883 29423 13889
rect 30285 13889 30297 13892
rect 30331 13889 30343 13923
rect 30285 13883 30343 13889
rect 31573 13923 31631 13929
rect 31573 13889 31585 13923
rect 31619 13889 31631 13923
rect 31846 13920 31852 13932
rect 31807 13892 31852 13920
rect 31573 13883 31631 13889
rect 31846 13880 31852 13892
rect 31904 13880 31910 13932
rect 32950 13880 32956 13932
rect 33008 13920 33014 13932
rect 33413 13923 33471 13929
rect 33413 13920 33425 13923
rect 33008 13892 33425 13920
rect 33008 13880 33014 13892
rect 33413 13889 33425 13892
rect 33459 13889 33471 13923
rect 33413 13883 33471 13889
rect 34146 13880 34152 13932
rect 34204 13920 34210 13932
rect 35894 13920 35900 13932
rect 34204 13892 35900 13920
rect 34204 13880 34210 13892
rect 35894 13880 35900 13892
rect 35952 13880 35958 13932
rect 36814 13880 36820 13932
rect 36872 13920 36878 13932
rect 37182 13920 37188 13932
rect 36872 13892 37188 13920
rect 36872 13880 36878 13892
rect 37182 13880 37188 13892
rect 37240 13880 37246 13932
rect 27065 13855 27123 13861
rect 27065 13852 27077 13855
rect 27028 13824 27077 13852
rect 27028 13812 27034 13824
rect 27065 13821 27077 13824
rect 27111 13821 27123 13855
rect 27065 13815 27123 13821
rect 28220 13855 28278 13861
rect 28220 13821 28232 13855
rect 28266 13852 28278 13855
rect 28721 13855 28779 13861
rect 28721 13852 28733 13855
rect 28266 13824 28733 13852
rect 28266 13821 28278 13824
rect 28220 13815 28278 13821
rect 28721 13821 28733 13824
rect 28767 13852 28779 13855
rect 28810 13852 28816 13864
rect 28767 13824 28816 13852
rect 28767 13821 28779 13824
rect 28721 13815 28779 13821
rect 28810 13812 28816 13824
rect 28868 13812 28874 13864
rect 34882 13852 34888 13864
rect 34843 13824 34888 13852
rect 34882 13812 34888 13824
rect 34940 13812 34946 13864
rect 24581 13787 24639 13793
rect 24581 13784 24593 13787
rect 24559 13756 24593 13784
rect 24581 13753 24593 13756
rect 24627 13784 24639 13787
rect 24946 13784 24952 13796
rect 24627 13756 24952 13784
rect 24627 13753 24639 13756
rect 24581 13747 24639 13753
rect 24946 13744 24952 13756
rect 25004 13744 25010 13796
rect 25222 13784 25228 13796
rect 25183 13756 25228 13784
rect 25222 13744 25228 13756
rect 25280 13744 25286 13796
rect 29086 13744 29092 13796
rect 29144 13784 29150 13796
rect 29454 13784 29460 13796
rect 29144 13756 29460 13784
rect 29144 13744 29150 13756
rect 29454 13744 29460 13756
rect 29512 13744 29518 13796
rect 31570 13744 31576 13796
rect 31628 13784 31634 13796
rect 31665 13787 31723 13793
rect 31665 13784 31677 13787
rect 31628 13756 31677 13784
rect 31628 13744 31634 13756
rect 31665 13753 31677 13756
rect 31711 13784 31723 13787
rect 32030 13784 32036 13796
rect 31711 13756 32036 13784
rect 31711 13753 31723 13756
rect 31665 13747 31723 13753
rect 32030 13744 32036 13756
rect 32088 13744 32094 13796
rect 32398 13744 32404 13796
rect 32456 13784 32462 13796
rect 33126 13787 33184 13793
rect 33126 13784 33138 13787
rect 32456 13756 33138 13784
rect 32456 13744 32462 13756
rect 33126 13753 33138 13756
rect 33172 13753 33184 13787
rect 33126 13747 33184 13753
rect 33222 13787 33280 13793
rect 33222 13753 33234 13787
rect 33268 13784 33280 13787
rect 33318 13784 33324 13796
rect 33268 13756 33324 13784
rect 33268 13753 33280 13756
rect 33222 13747 33280 13753
rect 33318 13744 33324 13756
rect 33376 13744 33382 13796
rect 34514 13744 34520 13796
rect 34572 13784 34578 13796
rect 35206 13787 35264 13793
rect 35206 13784 35218 13787
rect 34572 13756 35218 13784
rect 34572 13744 34578 13756
rect 35206 13753 35218 13756
rect 35252 13753 35264 13787
rect 36722 13784 36728 13796
rect 36683 13756 36728 13784
rect 35206 13747 35264 13753
rect 36722 13744 36728 13756
rect 36780 13744 36786 13796
rect 36817 13787 36875 13793
rect 36817 13753 36829 13787
rect 36863 13784 36875 13787
rect 37384 13784 37412 13960
rect 38194 13948 38200 14000
rect 38252 13988 38258 14000
rect 39666 13988 39672 14000
rect 38252 13960 38332 13988
rect 39627 13960 39672 13988
rect 38252 13948 38258 13960
rect 38304 13929 38332 13960
rect 39666 13948 39672 13960
rect 39724 13948 39730 14000
rect 40494 13948 40500 14000
rect 40552 13988 40558 14000
rect 41414 13988 41420 14000
rect 40552 13960 41420 13988
rect 40552 13948 40558 13960
rect 38289 13923 38347 13929
rect 38289 13889 38301 13923
rect 38335 13889 38347 13923
rect 38289 13883 38347 13889
rect 38470 13880 38476 13932
rect 38528 13920 38534 13932
rect 38565 13923 38623 13929
rect 38565 13920 38577 13923
rect 38528 13892 38577 13920
rect 38528 13880 38534 13892
rect 38565 13889 38577 13892
rect 38611 13889 38623 13923
rect 40954 13920 40960 13932
rect 38565 13883 38623 13889
rect 40547 13892 40960 13920
rect 40547 13861 40575 13892
rect 40954 13880 40960 13892
rect 41012 13880 41018 13932
rect 40532 13855 40590 13861
rect 40532 13821 40544 13855
rect 40578 13821 40590 13855
rect 40532 13815 40590 13821
rect 36863 13756 37412 13784
rect 36863 13753 36875 13756
rect 36817 13747 36875 13753
rect 10008 13688 10272 13716
rect 10008 13676 10014 13688
rect 17218 13676 17224 13728
rect 17276 13716 17282 13728
rect 17405 13719 17463 13725
rect 17405 13716 17417 13719
rect 17276 13688 17417 13716
rect 17276 13676 17282 13688
rect 17405 13685 17417 13688
rect 17451 13685 17463 13719
rect 20346 13716 20352 13728
rect 20307 13688 20352 13716
rect 17405 13679 17463 13685
rect 20346 13676 20352 13688
rect 20404 13676 20410 13728
rect 21683 13719 21741 13725
rect 21683 13685 21695 13719
rect 21729 13716 21741 13719
rect 22370 13716 22376 13728
rect 21729 13688 22376 13716
rect 21729 13685 21741 13688
rect 21683 13679 21741 13685
rect 22370 13676 22376 13688
rect 22428 13676 22434 13728
rect 22695 13719 22753 13725
rect 22695 13685 22707 13719
rect 22741 13716 22753 13719
rect 23106 13716 23112 13728
rect 22741 13688 23112 13716
rect 22741 13685 22753 13688
rect 22695 13679 22753 13685
rect 23106 13676 23112 13688
rect 23164 13676 23170 13728
rect 24167 13719 24225 13725
rect 24167 13685 24179 13719
rect 24213 13716 24225 13719
rect 24394 13716 24400 13728
rect 24213 13688 24400 13716
rect 24213 13685 24225 13688
rect 24167 13679 24225 13685
rect 24394 13676 24400 13688
rect 24452 13676 24458 13728
rect 26694 13716 26700 13728
rect 26655 13688 26700 13716
rect 26694 13676 26700 13688
rect 26752 13676 26758 13728
rect 32766 13676 32772 13728
rect 32824 13716 32830 13728
rect 32950 13716 32956 13728
rect 32824 13688 32956 13716
rect 32824 13676 32830 13688
rect 32950 13676 32956 13688
rect 33008 13676 33014 13728
rect 35805 13719 35863 13725
rect 35805 13685 35817 13719
rect 35851 13716 35863 13719
rect 36262 13716 36268 13728
rect 35851 13688 36268 13716
rect 35851 13685 35863 13688
rect 35805 13679 35863 13685
rect 36262 13676 36268 13688
rect 36320 13716 36326 13728
rect 36541 13719 36599 13725
rect 36541 13716 36553 13719
rect 36320 13688 36553 13716
rect 36320 13676 36326 13688
rect 36541 13685 36553 13688
rect 36587 13716 36599 13719
rect 36832 13716 36860 13747
rect 38378 13744 38384 13796
rect 38436 13784 38442 13796
rect 41340 13784 41368 13960
rect 41414 13948 41420 13960
rect 41472 13948 41478 14000
rect 42150 13988 42156 14000
rect 42111 13960 42156 13988
rect 42150 13948 42156 13960
rect 42208 13948 42214 14000
rect 41601 13923 41659 13929
rect 41601 13889 41613 13923
rect 41647 13920 41659 13923
rect 42766 13920 42794 14028
rect 42978 14016 42984 14028
rect 43036 14016 43042 14068
rect 43898 13920 43904 13932
rect 41647 13892 42794 13920
rect 43088 13892 43904 13920
rect 41647 13889 41659 13892
rect 41601 13883 41659 13889
rect 43088 13861 43116 13892
rect 43898 13880 43904 13892
rect 43956 13880 43962 13932
rect 43088 13855 43166 13861
rect 43088 13824 43120 13855
rect 43108 13821 43120 13824
rect 43154 13821 43166 13855
rect 43108 13815 43166 13821
rect 41598 13784 41604 13796
rect 38436 13756 38481 13784
rect 41340 13756 41604 13784
rect 38436 13744 38442 13756
rect 41598 13744 41604 13756
rect 41656 13784 41662 13796
rect 41693 13787 41751 13793
rect 41693 13784 41705 13787
rect 41656 13756 41705 13784
rect 41656 13744 41662 13756
rect 41693 13753 41705 13756
rect 41739 13753 41751 13787
rect 41693 13747 41751 13753
rect 36587 13688 36860 13716
rect 41708 13716 41736 13747
rect 42521 13719 42579 13725
rect 42521 13716 42533 13719
rect 41708 13688 42533 13716
rect 36587 13685 36599 13688
rect 36541 13679 36599 13685
rect 42521 13685 42533 13688
rect 42567 13685 42579 13719
rect 42521 13679 42579 13685
rect 42610 13676 42616 13728
rect 42668 13716 42674 13728
rect 43211 13719 43269 13725
rect 43211 13716 43223 13719
rect 42668 13688 43223 13716
rect 42668 13676 42674 13688
rect 43211 13685 43223 13688
rect 43257 13685 43269 13719
rect 43530 13716 43536 13728
rect 43491 13688 43536 13716
rect 43211 13679 43269 13685
rect 43530 13676 43536 13688
rect 43588 13676 43594 13728
rect 1104 13626 48852 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 48852 13626
rect 1104 13552 48852 13574
rect 4614 13512 4620 13524
rect 4575 13484 4620 13512
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 5629 13515 5687 13521
rect 5629 13481 5641 13515
rect 5675 13512 5687 13515
rect 10502 13512 10508 13524
rect 5675 13484 8559 13512
rect 10463 13484 10508 13512
rect 5675 13481 5687 13484
rect 5629 13475 5687 13481
rect 4632 13444 4660 13472
rect 5030 13447 5088 13453
rect 5030 13444 5042 13447
rect 4632 13416 5042 13444
rect 5030 13413 5042 13416
rect 5076 13413 5088 13447
rect 7098 13444 7104 13456
rect 7059 13416 7104 13444
rect 5030 13407 5088 13413
rect 7098 13404 7104 13416
rect 7156 13404 7162 13456
rect 4706 13376 4712 13388
rect 4667 13348 4712 13376
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 8531 13385 8559 13484
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 12529 13515 12587 13521
rect 12529 13481 12541 13515
rect 12575 13512 12587 13515
rect 12710 13512 12716 13524
rect 12575 13484 12716 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 14921 13515 14979 13521
rect 14921 13481 14933 13515
rect 14967 13512 14979 13515
rect 15102 13512 15108 13524
rect 14967 13484 15108 13512
rect 14967 13481 14979 13484
rect 14921 13475 14979 13481
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 16758 13472 16764 13524
rect 16816 13512 16822 13524
rect 18322 13512 18328 13524
rect 16816 13484 18328 13512
rect 16816 13472 16822 13484
rect 18322 13472 18328 13484
rect 18380 13512 18386 13524
rect 21450 13512 21456 13524
rect 18380 13484 21456 13512
rect 18380 13472 18386 13484
rect 21450 13472 21456 13484
rect 21508 13472 21514 13524
rect 23106 13472 23112 13524
rect 23164 13512 23170 13524
rect 23750 13512 23756 13524
rect 23164 13484 23756 13512
rect 23164 13472 23170 13484
rect 23750 13472 23756 13484
rect 23808 13472 23814 13524
rect 24903 13515 24961 13521
rect 24903 13481 24915 13515
rect 24949 13512 24961 13515
rect 25314 13512 25320 13524
rect 24949 13484 25320 13512
rect 24949 13481 24961 13484
rect 24903 13475 24961 13481
rect 25314 13472 25320 13484
rect 25372 13472 25378 13524
rect 28859 13515 28917 13521
rect 28859 13481 28871 13515
rect 28905 13512 28917 13515
rect 29178 13512 29184 13524
rect 28905 13484 29184 13512
rect 28905 13481 28917 13484
rect 28859 13475 28917 13481
rect 29178 13472 29184 13484
rect 29236 13472 29242 13524
rect 29273 13515 29331 13521
rect 29273 13481 29285 13515
rect 29319 13512 29331 13515
rect 29454 13512 29460 13524
rect 29319 13484 29460 13512
rect 29319 13481 29331 13484
rect 29273 13475 29331 13481
rect 29454 13472 29460 13484
rect 29512 13472 29518 13524
rect 31570 13512 31576 13524
rect 31531 13484 31576 13512
rect 31570 13472 31576 13484
rect 31628 13472 31634 13524
rect 31754 13472 31760 13524
rect 31812 13512 31818 13524
rect 31849 13515 31907 13521
rect 31849 13512 31861 13515
rect 31812 13484 31861 13512
rect 31812 13472 31818 13484
rect 31849 13481 31861 13484
rect 31895 13481 31907 13515
rect 31849 13475 31907 13481
rect 36722 13472 36728 13524
rect 36780 13512 36786 13524
rect 37093 13515 37151 13521
rect 37093 13512 37105 13515
rect 36780 13484 37105 13512
rect 36780 13472 36786 13484
rect 37093 13481 37105 13484
rect 37139 13512 37151 13515
rect 37875 13515 37933 13521
rect 37875 13512 37887 13515
rect 37139 13484 37887 13512
rect 37139 13481 37151 13484
rect 37093 13475 37151 13481
rect 37875 13481 37887 13484
rect 37921 13481 37933 13515
rect 37875 13475 37933 13481
rect 11238 13444 11244 13456
rect 11199 13416 11244 13444
rect 11238 13404 11244 13416
rect 11296 13444 11302 13456
rect 12805 13447 12863 13453
rect 12805 13444 12817 13447
rect 11296 13416 12817 13444
rect 11296 13404 11302 13416
rect 12805 13413 12817 13416
rect 12851 13444 12863 13447
rect 15473 13447 15531 13453
rect 15473 13444 15485 13447
rect 12851 13416 15485 13444
rect 12851 13413 12863 13416
rect 12805 13407 12863 13413
rect 15473 13413 15485 13416
rect 15519 13444 15531 13447
rect 15838 13444 15844 13456
rect 15519 13416 15844 13444
rect 15519 13413 15531 13416
rect 15473 13407 15531 13413
rect 15838 13404 15844 13416
rect 15896 13404 15902 13456
rect 18782 13404 18788 13456
rect 18840 13444 18846 13456
rect 19061 13447 19119 13453
rect 19061 13444 19073 13447
rect 18840 13416 19073 13444
rect 18840 13404 18846 13416
rect 19061 13413 19073 13416
rect 19107 13413 19119 13447
rect 21174 13444 21180 13456
rect 21135 13416 21180 13444
rect 19061 13407 19119 13413
rect 21174 13404 21180 13416
rect 21232 13404 21238 13456
rect 23385 13447 23443 13453
rect 23385 13413 23397 13447
rect 23431 13444 23443 13447
rect 23474 13444 23480 13456
rect 23431 13416 23480 13444
rect 23431 13413 23443 13416
rect 23385 13407 23443 13413
rect 23474 13404 23480 13416
rect 23532 13444 23538 13456
rect 25222 13444 25228 13456
rect 23532 13416 25228 13444
rect 23532 13404 23538 13416
rect 25222 13404 25228 13416
rect 25280 13404 25286 13456
rect 26326 13404 26332 13456
rect 26384 13444 26390 13456
rect 26834 13447 26892 13453
rect 26834 13444 26846 13447
rect 26384 13416 26846 13444
rect 26384 13404 26390 13416
rect 26834 13413 26846 13416
rect 26880 13413 26892 13447
rect 31588 13444 31616 13472
rect 32309 13447 32367 13453
rect 32309 13444 32321 13447
rect 31588 13416 32321 13444
rect 26834 13407 26892 13413
rect 32309 13413 32321 13416
rect 32355 13444 32367 13447
rect 32490 13444 32496 13456
rect 32355 13416 32496 13444
rect 32355 13413 32367 13416
rect 32309 13407 32367 13413
rect 32490 13404 32496 13416
rect 32548 13404 32554 13456
rect 32858 13444 32864 13456
rect 32819 13416 32864 13444
rect 32858 13404 32864 13416
rect 32916 13404 32922 13456
rect 34609 13447 34667 13453
rect 34609 13413 34621 13447
rect 34655 13444 34667 13447
rect 34882 13444 34888 13456
rect 34655 13416 34888 13444
rect 34655 13413 34667 13416
rect 34609 13407 34667 13413
rect 34882 13404 34888 13416
rect 34940 13444 34946 13456
rect 35253 13447 35311 13453
rect 35253 13444 35265 13447
rect 34940 13416 35265 13444
rect 34940 13404 34946 13416
rect 35253 13413 35265 13416
rect 35299 13413 35311 13447
rect 36262 13444 36268 13456
rect 36223 13416 36268 13444
rect 35253 13407 35311 13413
rect 36262 13404 36268 13416
rect 36320 13404 36326 13456
rect 39666 13404 39672 13456
rect 39724 13444 39730 13456
rect 39898 13447 39956 13453
rect 39898 13444 39910 13447
rect 39724 13416 39910 13444
rect 39724 13404 39730 13416
rect 39898 13413 39910 13416
rect 39944 13413 39956 13447
rect 41598 13444 41604 13456
rect 41559 13416 41604 13444
rect 39898 13407 39956 13413
rect 41598 13404 41604 13416
rect 41656 13404 41662 13456
rect 8516 13379 8574 13385
rect 8516 13345 8528 13379
rect 8562 13376 8574 13379
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8562 13348 8953 13376
rect 8562 13345 8574 13348
rect 8516 13339 8574 13345
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 9214 13336 9220 13388
rect 9272 13376 9278 13388
rect 9677 13379 9735 13385
rect 9677 13376 9689 13379
rect 9272 13348 9689 13376
rect 9272 13336 9278 13348
rect 9677 13345 9689 13348
rect 9723 13345 9735 13379
rect 14182 13376 14188 13388
rect 14143 13348 14188 13376
rect 9677 13339 9735 13345
rect 14182 13336 14188 13348
rect 14240 13336 14246 13388
rect 18116 13379 18174 13385
rect 18116 13345 18128 13379
rect 18162 13376 18174 13379
rect 18598 13376 18604 13388
rect 18162 13348 18604 13376
rect 18162 13345 18174 13348
rect 18116 13339 18174 13345
rect 18598 13336 18604 13348
rect 18656 13336 18662 13388
rect 19242 13376 19248 13388
rect 19203 13348 19248 13376
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 19705 13379 19763 13385
rect 19705 13376 19717 13379
rect 19484 13348 19717 13376
rect 19484 13336 19490 13348
rect 19705 13345 19717 13348
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 24765 13379 24823 13385
rect 24765 13345 24777 13379
rect 24811 13376 24823 13379
rect 24854 13376 24860 13388
rect 24811 13348 24860 13376
rect 24811 13345 24823 13348
rect 24765 13339 24823 13345
rect 24854 13336 24860 13348
rect 24912 13336 24918 13388
rect 26513 13379 26571 13385
rect 26513 13345 26525 13379
rect 26559 13376 26571 13379
rect 26694 13376 26700 13388
rect 26559 13348 26700 13376
rect 26559 13345 26571 13348
rect 26513 13339 26571 13345
rect 26694 13336 26700 13348
rect 26752 13336 26758 13388
rect 28629 13379 28687 13385
rect 28629 13345 28641 13379
rect 28675 13376 28687 13379
rect 28810 13376 28816 13388
rect 28675 13348 28816 13376
rect 28675 13345 28687 13348
rect 28629 13339 28687 13345
rect 28810 13336 28816 13348
rect 28868 13336 28874 13388
rect 30044 13379 30102 13385
rect 30044 13376 30056 13379
rect 29885 13348 30056 13376
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13277 7067 13311
rect 7650 13308 7656 13320
rect 7611 13280 7656 13308
rect 7009 13271 7067 13277
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 7024 13240 7052 13271
rect 7650 13268 7656 13280
rect 7708 13268 7714 13320
rect 11146 13308 11152 13320
rect 11059 13280 11152 13308
rect 11146 13268 11152 13280
rect 11204 13308 11210 13320
rect 11422 13308 11428 13320
rect 11204 13280 11428 13308
rect 11204 13268 11210 13280
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 11606 13308 11612 13320
rect 11567 13280 11612 13308
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 12434 13308 12440 13320
rect 11940 13280 12440 13308
rect 11940 13268 11946 13280
rect 12434 13268 12440 13280
rect 12492 13308 12498 13320
rect 12713 13311 12771 13317
rect 12713 13308 12725 13311
rect 12492 13280 12725 13308
rect 12492 13268 12498 13280
rect 12713 13277 12725 13280
rect 12759 13277 12771 13311
rect 12986 13308 12992 13320
rect 12947 13280 12992 13308
rect 12713 13271 12771 13277
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 15102 13268 15108 13320
rect 15160 13308 15166 13320
rect 15378 13308 15384 13320
rect 15160 13280 15384 13308
rect 15160 13268 15166 13280
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13277 15715 13311
rect 17034 13308 17040 13320
rect 16995 13280 17040 13308
rect 15657 13271 15715 13277
rect 8619 13243 8677 13249
rect 8619 13240 8631 13243
rect 6880 13212 8631 13240
rect 6880 13200 6886 13212
rect 8619 13209 8631 13212
rect 8665 13209 8677 13243
rect 8619 13203 8677 13209
rect 13998 13200 14004 13252
rect 14056 13240 14062 13252
rect 15562 13240 15568 13252
rect 14056 13212 15568 13240
rect 14056 13200 14062 13212
rect 15562 13200 15568 13212
rect 15620 13240 15626 13252
rect 15672 13240 15700 13271
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 19981 13311 20039 13317
rect 19981 13277 19993 13311
rect 20027 13308 20039 13311
rect 20162 13308 20168 13320
rect 20027 13280 20168 13308
rect 20027 13277 20039 13280
rect 19981 13271 20039 13277
rect 20162 13268 20168 13280
rect 20220 13308 20226 13320
rect 20257 13311 20315 13317
rect 20257 13308 20269 13311
rect 20220 13280 20269 13308
rect 20220 13268 20226 13280
rect 20257 13277 20269 13280
rect 20303 13277 20315 13311
rect 20257 13271 20315 13277
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13308 21143 13311
rect 21358 13308 21364 13320
rect 21131 13280 21364 13308
rect 21131 13277 21143 13280
rect 21085 13271 21143 13277
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 21542 13308 21548 13320
rect 21503 13280 21548 13308
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 22370 13268 22376 13320
rect 22428 13308 22434 13320
rect 23293 13311 23351 13317
rect 23293 13308 23305 13311
rect 22428 13280 23305 13308
rect 22428 13268 22434 13280
rect 23293 13277 23305 13280
rect 23339 13277 23351 13311
rect 23566 13308 23572 13320
rect 23527 13280 23572 13308
rect 23293 13271 23351 13277
rect 23566 13268 23572 13280
rect 23624 13268 23630 13320
rect 24118 13268 24124 13320
rect 24176 13308 24182 13320
rect 29885 13308 29913 13348
rect 30044 13345 30056 13348
rect 30090 13376 30102 13379
rect 30558 13376 30564 13388
rect 30090 13348 30564 13376
rect 30090 13345 30102 13348
rect 30044 13339 30102 13345
rect 30558 13336 30564 13348
rect 30616 13336 30622 13388
rect 31072 13379 31130 13385
rect 31072 13345 31084 13379
rect 31118 13376 31130 13379
rect 31294 13376 31300 13388
rect 31118 13348 31300 13376
rect 31118 13345 31130 13348
rect 31072 13339 31130 13345
rect 31294 13336 31300 13348
rect 31352 13336 31358 13388
rect 33870 13376 33876 13388
rect 33831 13348 33876 13376
rect 33870 13336 33876 13348
rect 33928 13336 33934 13388
rect 33962 13336 33968 13388
rect 34020 13376 34026 13388
rect 34333 13379 34391 13385
rect 34333 13376 34345 13379
rect 34020 13348 34345 13376
rect 34020 13336 34026 13348
rect 34333 13345 34345 13348
rect 34379 13376 34391 13379
rect 34514 13376 34520 13388
rect 34379 13348 34520 13376
rect 34379 13345 34391 13348
rect 34333 13339 34391 13345
rect 34514 13336 34520 13348
rect 34572 13376 34578 13388
rect 34977 13379 35035 13385
rect 34977 13376 34989 13379
rect 34572 13348 34989 13376
rect 34572 13336 34578 13348
rect 34977 13345 34989 13348
rect 35023 13345 35035 13379
rect 34977 13339 35035 13345
rect 37645 13379 37703 13385
rect 37645 13345 37657 13379
rect 37691 13376 37703 13379
rect 37826 13376 37832 13388
rect 37691 13348 37832 13376
rect 37691 13345 37703 13348
rect 37645 13339 37703 13345
rect 37826 13336 37832 13348
rect 37884 13336 37890 13388
rect 43254 13376 43260 13388
rect 43215 13348 43260 13376
rect 43254 13336 43260 13348
rect 43312 13336 43318 13388
rect 24176 13280 29913 13308
rect 30147 13311 30205 13317
rect 24176 13268 24182 13280
rect 30147 13277 30159 13311
rect 30193 13308 30205 13311
rect 32217 13311 32275 13317
rect 32217 13308 32229 13311
rect 30193 13280 32229 13308
rect 30193 13277 30205 13280
rect 30147 13271 30205 13277
rect 32217 13277 32229 13280
rect 32263 13308 32275 13311
rect 32858 13308 32864 13320
rect 32263 13280 32864 13308
rect 32263 13277 32275 13280
rect 32217 13271 32275 13277
rect 32858 13268 32864 13280
rect 32916 13268 32922 13320
rect 34790 13268 34796 13320
rect 34848 13308 34854 13320
rect 36170 13308 36176 13320
rect 34848 13280 36176 13308
rect 34848 13268 34854 13280
rect 36170 13268 36176 13280
rect 36228 13268 36234 13320
rect 36630 13268 36636 13320
rect 36688 13308 36694 13320
rect 36817 13311 36875 13317
rect 36817 13308 36829 13311
rect 36688 13280 36829 13308
rect 36688 13268 36694 13280
rect 36817 13277 36829 13280
rect 36863 13308 36875 13311
rect 37182 13308 37188 13320
rect 36863 13280 37188 13308
rect 36863 13277 36875 13280
rect 36817 13271 36875 13277
rect 37182 13268 37188 13280
rect 37240 13268 37246 13320
rect 39574 13308 39580 13320
rect 39535 13280 39580 13308
rect 39574 13268 39580 13280
rect 39632 13268 39638 13320
rect 41509 13311 41567 13317
rect 41509 13277 41521 13311
rect 41555 13308 41567 13311
rect 42610 13308 42616 13320
rect 41555 13280 42616 13308
rect 41555 13277 41567 13280
rect 41509 13271 41567 13277
rect 42610 13268 42616 13280
rect 42668 13268 42674 13320
rect 15620 13212 15700 13240
rect 15620 13200 15626 13212
rect 26878 13200 26884 13252
rect 26936 13240 26942 13252
rect 31386 13240 31392 13252
rect 26936 13212 31392 13240
rect 26936 13200 26942 13212
rect 31386 13200 31392 13212
rect 31444 13200 31450 13252
rect 34330 13200 34336 13252
rect 34388 13240 34394 13252
rect 38286 13240 38292 13252
rect 34388 13212 38292 13240
rect 34388 13200 34394 13212
rect 38286 13200 38292 13212
rect 38344 13200 38350 13252
rect 40862 13200 40868 13252
rect 40920 13240 40926 13252
rect 41690 13240 41696 13252
rect 40920 13212 41696 13240
rect 40920 13200 40926 13212
rect 41690 13200 41696 13212
rect 41748 13240 41754 13252
rect 42061 13243 42119 13249
rect 42061 13240 42073 13243
rect 41748 13212 42073 13240
rect 41748 13200 41754 13212
rect 42061 13209 42073 13212
rect 42107 13240 42119 13243
rect 44174 13240 44180 13252
rect 42107 13212 44180 13240
rect 42107 13209 42119 13212
rect 42061 13203 42119 13209
rect 44174 13200 44180 13212
rect 44232 13200 44238 13252
rect 6730 13172 6736 13184
rect 6691 13144 6736 13172
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 9861 13175 9919 13181
rect 9861 13141 9873 13175
rect 9907 13172 9919 13175
rect 10042 13172 10048 13184
rect 9907 13144 10048 13172
rect 9907 13141 9919 13144
rect 9861 13135 9919 13141
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 14366 13172 14372 13184
rect 14327 13144 14372 13172
rect 14366 13132 14372 13144
rect 14424 13132 14430 13184
rect 18046 13132 18052 13184
rect 18104 13172 18110 13184
rect 18187 13175 18245 13181
rect 18187 13172 18199 13175
rect 18104 13144 18199 13172
rect 18104 13132 18110 13144
rect 18187 13141 18199 13144
rect 18233 13141 18245 13175
rect 18598 13172 18604 13184
rect 18559 13144 18604 13172
rect 18187 13135 18245 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 23750 13132 23756 13184
rect 23808 13172 23814 13184
rect 24213 13175 24271 13181
rect 24213 13172 24225 13175
rect 23808 13144 24225 13172
rect 23808 13132 23814 13144
rect 24213 13141 24225 13144
rect 24259 13141 24271 13175
rect 24213 13135 24271 13141
rect 25222 13132 25228 13184
rect 25280 13172 25286 13184
rect 25317 13175 25375 13181
rect 25317 13172 25329 13175
rect 25280 13144 25329 13172
rect 25280 13132 25286 13144
rect 25317 13141 25329 13144
rect 25363 13172 25375 13175
rect 27433 13175 27491 13181
rect 27433 13172 27445 13175
rect 25363 13144 27445 13172
rect 25363 13141 25375 13144
rect 25317 13135 25375 13141
rect 27433 13141 27445 13144
rect 27479 13141 27491 13175
rect 27433 13135 27491 13141
rect 29641 13175 29699 13181
rect 29641 13141 29653 13175
rect 29687 13172 29699 13175
rect 29730 13172 29736 13184
rect 29687 13144 29736 13172
rect 29687 13141 29699 13144
rect 29641 13135 29699 13141
rect 29730 13132 29736 13144
rect 29788 13132 29794 13184
rect 31159 13175 31217 13181
rect 31159 13141 31171 13175
rect 31205 13172 31217 13175
rect 32398 13172 32404 13184
rect 31205 13144 32404 13172
rect 31205 13141 31217 13144
rect 31159 13135 31217 13141
rect 32398 13132 32404 13144
rect 32456 13172 32462 13184
rect 33137 13175 33195 13181
rect 33137 13172 33149 13175
rect 32456 13144 33149 13172
rect 32456 13132 32462 13144
rect 33137 13141 33149 13144
rect 33183 13141 33195 13175
rect 38194 13172 38200 13184
rect 38155 13144 38200 13172
rect 33137 13135 33195 13141
rect 38194 13132 38200 13144
rect 38252 13132 38258 13184
rect 40497 13175 40555 13181
rect 40497 13141 40509 13175
rect 40543 13172 40555 13175
rect 40773 13175 40831 13181
rect 40773 13172 40785 13175
rect 40543 13144 40785 13172
rect 40543 13141 40555 13144
rect 40497 13135 40555 13141
rect 40773 13141 40785 13144
rect 40819 13172 40831 13175
rect 40954 13172 40960 13184
rect 40819 13144 40960 13172
rect 40819 13141 40831 13144
rect 40773 13135 40831 13141
rect 40954 13132 40960 13144
rect 41012 13132 41018 13184
rect 43162 13132 43168 13184
rect 43220 13172 43226 13184
rect 43487 13175 43545 13181
rect 43487 13172 43499 13175
rect 43220 13144 43499 13172
rect 43220 13132 43226 13144
rect 43487 13141 43499 13144
rect 43533 13141 43545 13175
rect 43487 13135 43545 13141
rect 1104 13082 48852 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 48852 13082
rect 1104 13008 48852 13030
rect 4433 12971 4491 12977
rect 4433 12937 4445 12971
rect 4479 12968 4491 12971
rect 4706 12968 4712 12980
rect 4479 12940 4712 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5350 12968 5356 12980
rect 5311 12940 5356 12968
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 5675 12971 5733 12977
rect 5675 12937 5687 12971
rect 5721 12968 5733 12971
rect 6730 12968 6736 12980
rect 5721 12940 6736 12968
rect 5721 12937 5733 12940
rect 5675 12931 5733 12937
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9493 12971 9551 12977
rect 9493 12968 9505 12971
rect 9272 12940 9505 12968
rect 9272 12928 9278 12940
rect 9493 12937 9505 12940
rect 9539 12937 9551 12971
rect 11422 12968 11428 12980
rect 11383 12940 11428 12968
rect 9493 12931 9551 12937
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 11882 12968 11888 12980
rect 11843 12940 11888 12968
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 15286 12968 15292 12980
rect 13786 12940 15292 12968
rect 7561 12903 7619 12909
rect 7561 12869 7573 12903
rect 7607 12900 7619 12903
rect 9122 12900 9128 12912
rect 7607 12872 9128 12900
rect 7607 12869 7619 12872
rect 7561 12863 7619 12869
rect 9122 12860 9128 12872
rect 9180 12860 9186 12912
rect 9858 12860 9864 12912
rect 9916 12900 9922 12912
rect 11057 12903 11115 12909
rect 11057 12900 11069 12903
rect 9916 12872 11069 12900
rect 9916 12860 9922 12872
rect 11057 12869 11069 12872
rect 11103 12900 11115 12903
rect 11238 12900 11244 12912
rect 11103 12872 11244 12900
rect 11103 12869 11115 12872
rect 11057 12863 11115 12869
rect 11238 12860 11244 12872
rect 11296 12860 11302 12912
rect 13786 12900 13814 12940
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 15838 12968 15844 12980
rect 15799 12940 15844 12968
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 19613 12971 19671 12977
rect 19613 12968 19625 12971
rect 19484 12940 19625 12968
rect 19484 12928 19490 12940
rect 19613 12937 19625 12940
rect 19659 12937 19671 12971
rect 20070 12968 20076 12980
rect 20031 12940 20076 12968
rect 19613 12931 19671 12937
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 21358 12968 21364 12980
rect 21319 12940 21364 12968
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 22370 12968 22376 12980
rect 22331 12940 22376 12968
rect 22370 12928 22376 12940
rect 22428 12928 22434 12980
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 27525 12971 27583 12977
rect 23532 12940 23577 12968
rect 23532 12928 23538 12940
rect 27525 12937 27537 12971
rect 27571 12968 27583 12971
rect 27614 12968 27620 12980
rect 27571 12940 27620 12968
rect 27571 12937 27583 12940
rect 27525 12931 27583 12937
rect 27614 12928 27620 12940
rect 27672 12928 27678 12980
rect 30558 12968 30564 12980
rect 30519 12940 30564 12968
rect 30558 12928 30564 12940
rect 30616 12928 30622 12980
rect 31113 12971 31171 12977
rect 31113 12937 31125 12971
rect 31159 12968 31171 12971
rect 31294 12968 31300 12980
rect 31159 12940 31300 12968
rect 31159 12937 31171 12940
rect 31113 12931 31171 12937
rect 31294 12928 31300 12940
rect 31352 12928 31358 12980
rect 32490 12968 32496 12980
rect 32451 12940 32496 12968
rect 32490 12928 32496 12940
rect 32548 12928 32554 12980
rect 32858 12968 32864 12980
rect 32819 12940 32864 12968
rect 32858 12928 32864 12940
rect 32916 12928 32922 12980
rect 33689 12971 33747 12977
rect 33689 12937 33701 12971
rect 33735 12968 33747 12971
rect 33870 12968 33876 12980
rect 33735 12940 33876 12968
rect 33735 12937 33747 12940
rect 33689 12931 33747 12937
rect 33870 12928 33876 12940
rect 33928 12928 33934 12980
rect 34330 12968 34336 12980
rect 34291 12940 34336 12968
rect 34330 12928 34336 12940
rect 34388 12928 34394 12980
rect 34514 12928 34520 12980
rect 34572 12968 34578 12980
rect 34609 12971 34667 12977
rect 34609 12968 34621 12971
rect 34572 12940 34621 12968
rect 34572 12928 34578 12940
rect 34609 12937 34621 12940
rect 34655 12968 34667 12971
rect 35342 12968 35348 12980
rect 34655 12940 35348 12968
rect 34655 12937 34667 12940
rect 34609 12931 34667 12937
rect 35342 12928 35348 12940
rect 35400 12928 35406 12980
rect 36173 12971 36231 12977
rect 36173 12937 36185 12971
rect 36219 12968 36231 12971
rect 36262 12968 36268 12980
rect 36219 12940 36268 12968
rect 36219 12937 36231 12940
rect 36173 12931 36231 12937
rect 36262 12928 36268 12940
rect 36320 12928 36326 12980
rect 37826 12968 37832 12980
rect 37787 12940 37832 12968
rect 37826 12928 37832 12940
rect 37884 12928 37890 12980
rect 39666 12928 39672 12980
rect 39724 12968 39730 12980
rect 39853 12971 39911 12977
rect 39853 12968 39865 12971
rect 39724 12940 39865 12968
rect 39724 12928 39730 12940
rect 39853 12937 39865 12940
rect 39899 12937 39911 12971
rect 39853 12931 39911 12937
rect 41598 12928 41604 12980
rect 41656 12968 41662 12980
rect 41785 12971 41843 12977
rect 41785 12968 41797 12971
rect 41656 12940 41797 12968
rect 41656 12928 41662 12940
rect 41785 12937 41797 12940
rect 41831 12937 41843 12971
rect 41785 12931 41843 12937
rect 42245 12971 42303 12977
rect 42245 12937 42257 12971
rect 42291 12968 42303 12971
rect 42610 12968 42616 12980
rect 42291 12940 42616 12968
rect 42291 12937 42303 12940
rect 42245 12931 42303 12937
rect 42610 12928 42616 12940
rect 42668 12928 42674 12980
rect 43254 12928 43260 12980
rect 43312 12968 43318 12980
rect 44085 12971 44143 12977
rect 44085 12968 44097 12971
rect 43312 12940 44097 12968
rect 43312 12928 43318 12940
rect 44085 12937 44097 12940
rect 44131 12937 44143 12971
rect 44085 12931 44143 12937
rect 11716 12872 13814 12900
rect 21085 12903 21143 12909
rect 4614 12792 4620 12844
rect 4672 12832 4678 12844
rect 4709 12835 4767 12841
rect 4709 12832 4721 12835
rect 4672 12804 4721 12832
rect 4672 12792 4678 12804
rect 4709 12801 4721 12804
rect 4755 12801 4767 12835
rect 7006 12832 7012 12844
rect 6919 12804 7012 12832
rect 4709 12795 4767 12801
rect 7006 12792 7012 12804
rect 7064 12832 7070 12844
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 7064 12804 7941 12832
rect 7064 12792 7070 12804
rect 7929 12801 7941 12804
rect 7975 12801 7987 12835
rect 7929 12795 7987 12801
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12832 10839 12835
rect 11606 12832 11612 12844
rect 10827 12804 11612 12832
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 5350 12724 5356 12776
rect 5408 12764 5414 12776
rect 5572 12767 5630 12773
rect 5572 12764 5584 12767
rect 5408 12736 5584 12764
rect 5408 12724 5414 12736
rect 5572 12733 5584 12736
rect 5618 12733 5630 12767
rect 5572 12727 5630 12733
rect 6273 12699 6331 12705
rect 6273 12665 6285 12699
rect 6319 12696 6331 12699
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 6319 12668 6653 12696
rect 6319 12665 6331 12668
rect 6273 12659 6331 12665
rect 6641 12665 6653 12668
rect 6687 12696 6699 12699
rect 7098 12696 7104 12708
rect 6687 12668 7104 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 7742 12656 7748 12708
rect 7800 12696 7806 12708
rect 8573 12699 8631 12705
rect 8573 12696 8585 12699
rect 7800 12668 8585 12696
rect 7800 12656 7806 12668
rect 8573 12665 8585 12668
rect 8619 12665 8631 12699
rect 8573 12659 8631 12665
rect 8665 12699 8723 12705
rect 8665 12665 8677 12699
rect 8711 12665 8723 12699
rect 9214 12696 9220 12708
rect 9175 12668 9220 12696
rect 8665 12659 8723 12665
rect 8389 12631 8447 12637
rect 8389 12597 8401 12631
rect 8435 12628 8447 12631
rect 8680 12628 8708 12659
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 10134 12696 10140 12708
rect 10095 12668 10140 12696
rect 10134 12656 10140 12668
rect 10192 12656 10198 12708
rect 10229 12699 10287 12705
rect 10229 12665 10241 12699
rect 10275 12696 10287 12699
rect 11716 12696 11744 12872
rect 21085 12869 21097 12903
rect 21131 12900 21143 12903
rect 21174 12900 21180 12912
rect 21131 12872 21180 12900
rect 21131 12869 21143 12872
rect 21085 12863 21143 12869
rect 21174 12860 21180 12872
rect 21232 12900 21238 12912
rect 21729 12903 21787 12909
rect 21729 12900 21741 12903
rect 21232 12872 21741 12900
rect 21232 12860 21238 12872
rect 21729 12869 21741 12872
rect 21775 12869 21787 12903
rect 21729 12863 21787 12869
rect 30466 12860 30472 12912
rect 30524 12900 30530 12912
rect 32125 12903 32183 12909
rect 32125 12900 32137 12903
rect 30524 12872 32137 12900
rect 30524 12860 30530 12872
rect 32125 12869 32137 12872
rect 32171 12900 32183 12903
rect 32674 12900 32680 12912
rect 32171 12872 32680 12900
rect 32171 12869 32183 12872
rect 32125 12863 32183 12869
rect 32674 12860 32680 12872
rect 32732 12860 32738 12912
rect 34698 12860 34704 12912
rect 34756 12900 34762 12912
rect 38657 12903 38715 12909
rect 38657 12900 38669 12903
rect 34756 12872 38669 12900
rect 34756 12860 34762 12872
rect 38657 12869 38669 12872
rect 38703 12869 38715 12903
rect 38657 12863 38715 12869
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12832 12955 12835
rect 12986 12832 12992 12844
rect 12943 12804 12992 12832
rect 12943 12801 12955 12804
rect 12897 12795 12955 12801
rect 12986 12792 12992 12804
rect 13044 12832 13050 12844
rect 13817 12835 13875 12841
rect 13817 12832 13829 12835
rect 13044 12804 13829 12832
rect 13044 12792 13050 12804
rect 13817 12801 13829 12804
rect 13863 12801 13875 12835
rect 13817 12795 13875 12801
rect 17681 12835 17739 12841
rect 17681 12801 17693 12835
rect 17727 12832 17739 12835
rect 18414 12832 18420 12844
rect 17727 12804 18420 12832
rect 17727 12801 17739 12804
rect 17681 12795 17739 12801
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 20162 12832 20168 12844
rect 20123 12804 20168 12832
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 23750 12832 23756 12844
rect 23711 12804 23756 12832
rect 23750 12792 23756 12804
rect 23808 12792 23814 12844
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12832 24455 12835
rect 24578 12832 24584 12844
rect 24443 12804 24584 12832
rect 24443 12801 24455 12804
rect 24397 12795 24455 12801
rect 24578 12792 24584 12804
rect 24636 12792 24642 12844
rect 24854 12832 24860 12844
rect 24767 12804 24860 12832
rect 24854 12792 24860 12804
rect 24912 12832 24918 12844
rect 28810 12832 28816 12844
rect 24912 12804 28816 12832
rect 24912 12792 24918 12804
rect 28810 12792 28816 12804
rect 28868 12792 28874 12844
rect 29641 12835 29699 12841
rect 29641 12801 29653 12835
rect 29687 12832 29699 12835
rect 29914 12832 29920 12844
rect 29687 12804 29920 12832
rect 29687 12801 29699 12804
rect 29641 12795 29699 12801
rect 29914 12792 29920 12804
rect 29972 12832 29978 12844
rect 32582 12832 32588 12844
rect 29972 12804 32588 12832
rect 29972 12792 29978 12804
rect 32582 12792 32588 12804
rect 32640 12792 32646 12844
rect 34422 12792 34428 12844
rect 34480 12832 34486 12844
rect 36633 12835 36691 12841
rect 36633 12832 36645 12835
rect 34480 12804 36645 12832
rect 34480 12792 34486 12804
rect 36633 12801 36645 12804
rect 36679 12801 36691 12835
rect 36633 12795 36691 12801
rect 36909 12835 36967 12841
rect 36909 12801 36921 12835
rect 36955 12832 36967 12835
rect 37090 12832 37096 12844
rect 36955 12804 37096 12832
rect 36955 12801 36967 12804
rect 36909 12795 36967 12801
rect 14737 12767 14795 12773
rect 14737 12733 14749 12767
rect 14783 12764 14795 12767
rect 15473 12767 15531 12773
rect 15473 12764 15485 12767
rect 14783 12736 15485 12764
rect 14783 12733 14795 12736
rect 14737 12727 14795 12733
rect 15473 12733 15485 12736
rect 15519 12764 15531 12767
rect 15746 12764 15752 12776
rect 15519 12736 15752 12764
rect 15519 12733 15531 12736
rect 15473 12727 15531 12733
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 16393 12767 16451 12773
rect 16393 12733 16405 12767
rect 16439 12733 16451 12767
rect 16942 12764 16948 12776
rect 16903 12736 16948 12764
rect 16393 12727 16451 12733
rect 10275 12668 11744 12696
rect 12253 12699 12311 12705
rect 10275 12665 10287 12668
rect 10229 12659 10287 12665
rect 12253 12665 12265 12699
rect 12299 12696 12311 12699
rect 12989 12699 13047 12705
rect 12989 12696 13001 12699
rect 12299 12668 13001 12696
rect 12299 12665 12311 12668
rect 12253 12659 12311 12665
rect 12989 12665 13001 12668
rect 13035 12696 13047 12699
rect 13170 12696 13176 12708
rect 13035 12668 13176 12696
rect 13035 12665 13047 12668
rect 12989 12659 13047 12665
rect 9950 12628 9956 12640
rect 8435 12600 9956 12628
rect 8435 12597 8447 12600
rect 8389 12591 8447 12597
rect 9950 12588 9956 12600
rect 10008 12628 10014 12640
rect 10244 12628 10272 12659
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 13541 12699 13599 12705
rect 13541 12665 13553 12699
rect 13587 12696 13599 12699
rect 13630 12696 13636 12708
rect 13587 12668 13636 12696
rect 13587 12665 13599 12668
rect 13541 12659 13599 12665
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 13814 12656 13820 12708
rect 13872 12696 13878 12708
rect 16209 12699 16267 12705
rect 16209 12696 16221 12699
rect 13872 12668 16221 12696
rect 13872 12656 13878 12668
rect 16209 12665 16221 12668
rect 16255 12696 16267 12699
rect 16408 12696 16436 12727
rect 16942 12724 16948 12736
rect 17000 12724 17006 12776
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12764 17187 12767
rect 17497 12767 17555 12773
rect 17497 12764 17509 12767
rect 17175 12736 17509 12764
rect 17175 12733 17187 12736
rect 17129 12727 17187 12733
rect 17497 12733 17509 12736
rect 17543 12764 17555 12767
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17543 12736 18061 12764
rect 17543 12733 17555 12736
rect 17497 12727 17555 12733
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 19242 12764 19248 12776
rect 18049 12727 18107 12733
rect 18248 12736 19248 12764
rect 18248 12708 18276 12736
rect 19242 12724 19248 12736
rect 19300 12724 19306 12776
rect 22624 12767 22682 12773
rect 22624 12733 22636 12767
rect 22670 12764 22682 12767
rect 25774 12764 25780 12776
rect 22670 12736 23152 12764
rect 25735 12736 25780 12764
rect 22670 12733 22682 12736
rect 22624 12727 22682 12733
rect 18230 12696 18236 12708
rect 16255 12668 18236 12696
rect 16255 12665 16267 12668
rect 16209 12659 16267 12665
rect 18230 12656 18236 12668
rect 18288 12656 18294 12708
rect 20070 12696 20076 12708
rect 18432 12668 20076 12696
rect 18432 12640 18460 12668
rect 20070 12656 20076 12668
rect 20128 12696 20134 12708
rect 20486 12699 20544 12705
rect 20486 12696 20498 12699
rect 20128 12668 20498 12696
rect 20128 12656 20134 12668
rect 20486 12665 20498 12668
rect 20532 12665 20544 12699
rect 20486 12659 20544 12665
rect 23124 12640 23152 12736
rect 25774 12724 25780 12736
rect 25832 12724 25838 12776
rect 27614 12764 27620 12776
rect 27575 12736 27620 12764
rect 27614 12724 27620 12736
rect 27672 12724 27678 12776
rect 28074 12764 28080 12776
rect 28035 12736 28080 12764
rect 28074 12724 28080 12736
rect 28132 12724 28138 12776
rect 33778 12764 33784 12776
rect 33742 12736 33784 12764
rect 33778 12724 33784 12736
rect 33836 12773 33842 12776
rect 33836 12767 33890 12773
rect 33836 12733 33844 12767
rect 33878 12764 33890 12767
rect 34330 12764 34336 12776
rect 33878 12736 34336 12764
rect 33878 12733 33890 12736
rect 33836 12727 33890 12733
rect 33836 12724 33842 12727
rect 34330 12724 34336 12736
rect 34388 12724 34394 12776
rect 34698 12724 34704 12776
rect 34756 12764 34762 12776
rect 34885 12767 34943 12773
rect 34885 12764 34897 12767
rect 34756 12736 34897 12764
rect 34756 12724 34762 12736
rect 34885 12733 34897 12736
rect 34931 12733 34943 12767
rect 35342 12764 35348 12776
rect 35303 12736 35348 12764
rect 34885 12727 34943 12733
rect 35342 12724 35348 12736
rect 35400 12724 35406 12776
rect 23474 12656 23480 12708
rect 23532 12696 23538 12708
rect 23845 12699 23903 12705
rect 23845 12696 23857 12699
rect 23532 12668 23857 12696
rect 23532 12656 23538 12668
rect 23845 12665 23857 12668
rect 23891 12696 23903 12699
rect 23934 12696 23940 12708
rect 23891 12668 23940 12696
rect 23891 12665 23903 12668
rect 23845 12659 23903 12665
rect 23934 12656 23940 12668
rect 23992 12656 23998 12708
rect 26098 12699 26156 12705
rect 26098 12696 26110 12699
rect 25608 12668 26110 12696
rect 10008 12600 10272 12628
rect 10008 12588 10014 12600
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 11296 12600 12633 12628
rect 11296 12588 11302 12600
rect 12621 12597 12633 12600
rect 12667 12597 12679 12631
rect 14182 12628 14188 12640
rect 14143 12600 14188 12628
rect 12621 12591 12679 12597
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 16758 12588 16764 12640
rect 16816 12628 16822 12640
rect 17681 12631 17739 12637
rect 17681 12628 17693 12631
rect 16816 12600 17693 12628
rect 16816 12588 16822 12600
rect 17681 12597 17693 12600
rect 17727 12628 17739 12631
rect 17773 12631 17831 12637
rect 17773 12628 17785 12631
rect 17727 12600 17785 12628
rect 17727 12597 17739 12600
rect 17681 12591 17739 12597
rect 17773 12597 17785 12600
rect 17819 12597 17831 12631
rect 18414 12628 18420 12640
rect 18375 12600 18420 12628
rect 17773 12591 17831 12597
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 18966 12628 18972 12640
rect 18927 12600 18972 12628
rect 18966 12588 18972 12600
rect 19024 12588 19030 12640
rect 22695 12631 22753 12637
rect 22695 12597 22707 12631
rect 22741 12628 22753 12631
rect 22830 12628 22836 12640
rect 22741 12600 22836 12628
rect 22741 12597 22753 12600
rect 22695 12591 22753 12597
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 23106 12628 23112 12640
rect 23067 12600 23112 12628
rect 23106 12588 23112 12600
rect 23164 12588 23170 12640
rect 25406 12588 25412 12640
rect 25464 12628 25470 12640
rect 25608 12637 25636 12668
rect 26098 12665 26110 12668
rect 26144 12696 26156 12699
rect 26326 12696 26332 12708
rect 26144 12668 26332 12696
rect 26144 12665 26156 12668
rect 26098 12659 26156 12665
rect 26326 12656 26332 12668
rect 26384 12696 26390 12708
rect 26973 12699 27031 12705
rect 26973 12696 26985 12699
rect 26384 12668 26985 12696
rect 26384 12656 26390 12668
rect 26973 12665 26985 12668
rect 27019 12665 27031 12699
rect 26973 12659 27031 12665
rect 28353 12699 28411 12705
rect 28353 12665 28365 12699
rect 28399 12696 28411 12699
rect 28626 12696 28632 12708
rect 28399 12668 28632 12696
rect 28399 12665 28411 12668
rect 28353 12659 28411 12665
rect 28626 12656 28632 12668
rect 28684 12656 28690 12708
rect 29730 12656 29736 12708
rect 29788 12696 29794 12708
rect 30285 12699 30343 12705
rect 29788 12668 29833 12696
rect 29788 12656 29794 12668
rect 30285 12665 30297 12699
rect 30331 12696 30343 12699
rect 31294 12696 31300 12708
rect 30331 12668 31300 12696
rect 30331 12665 30343 12668
rect 30285 12659 30343 12665
rect 31294 12656 31300 12668
rect 31352 12656 31358 12708
rect 31570 12696 31576 12708
rect 31531 12668 31576 12696
rect 31570 12656 31576 12668
rect 31628 12656 31634 12708
rect 31662 12656 31668 12708
rect 31720 12696 31726 12708
rect 33919 12699 33977 12705
rect 31720 12668 31765 12696
rect 31720 12656 31726 12668
rect 33919 12665 33931 12699
rect 33965 12696 33977 12699
rect 36538 12696 36544 12708
rect 33965 12668 36544 12696
rect 33965 12665 33977 12668
rect 33919 12659 33977 12665
rect 36538 12656 36544 12668
rect 36596 12656 36602 12708
rect 36648 12696 36676 12795
rect 37090 12792 37096 12804
rect 37148 12792 37154 12844
rect 37182 12792 37188 12844
rect 37240 12832 37246 12844
rect 37240 12804 37285 12832
rect 37240 12792 37246 12804
rect 38672 12764 38700 12863
rect 41506 12860 41512 12912
rect 41564 12900 41570 12912
rect 41564 12872 43484 12900
rect 41564 12860 41570 12872
rect 42260 12844 42288 12872
rect 39574 12832 39580 12844
rect 39487 12804 39580 12832
rect 39574 12792 39580 12804
rect 39632 12832 39638 12844
rect 40221 12835 40279 12841
rect 40221 12832 40233 12835
rect 39632 12804 40233 12832
rect 39632 12792 39638 12804
rect 40221 12801 40233 12804
rect 40267 12801 40279 12835
rect 40221 12795 40279 12801
rect 42242 12792 42248 12844
rect 42300 12792 42306 12844
rect 43162 12832 43168 12844
rect 43123 12804 43168 12832
rect 43162 12792 43168 12804
rect 43220 12792 43226 12844
rect 43456 12841 43484 12872
rect 43441 12835 43499 12841
rect 43441 12801 43453 12835
rect 43487 12801 43499 12835
rect 43441 12795 43499 12801
rect 38841 12767 38899 12773
rect 38841 12764 38853 12767
rect 38672 12736 38853 12764
rect 38841 12733 38853 12736
rect 38887 12733 38899 12767
rect 38841 12727 38899 12733
rect 39114 12724 39120 12776
rect 39172 12764 39178 12776
rect 39301 12767 39359 12773
rect 39301 12764 39313 12767
rect 39172 12736 39313 12764
rect 39172 12724 39178 12736
rect 39301 12733 39313 12736
rect 39347 12733 39359 12767
rect 39301 12727 39359 12733
rect 43990 12724 43996 12776
rect 44048 12764 44054 12776
rect 44672 12767 44730 12773
rect 44672 12764 44684 12767
rect 44048 12736 44684 12764
rect 44048 12724 44054 12736
rect 44672 12733 44684 12736
rect 44718 12764 44730 12767
rect 45097 12767 45155 12773
rect 45097 12764 45109 12767
rect 44718 12736 45109 12764
rect 44718 12733 44730 12736
rect 44672 12727 44730 12733
rect 45097 12733 45109 12736
rect 45143 12733 45155 12767
rect 45097 12727 45155 12733
rect 36998 12696 37004 12708
rect 36648 12668 37004 12696
rect 36998 12656 37004 12668
rect 37056 12656 37062 12708
rect 40862 12696 40868 12708
rect 40823 12668 40868 12696
rect 40862 12656 40868 12668
rect 40920 12656 40926 12708
rect 40954 12656 40960 12708
rect 41012 12696 41018 12708
rect 41509 12699 41567 12705
rect 41012 12668 41057 12696
rect 41012 12656 41018 12668
rect 41509 12665 41521 12699
rect 41555 12696 41567 12699
rect 41874 12696 41880 12708
rect 41555 12668 41880 12696
rect 41555 12665 41567 12668
rect 41509 12659 41567 12665
rect 41874 12656 41880 12668
rect 41932 12656 41938 12708
rect 43257 12699 43315 12705
rect 43257 12665 43269 12699
rect 43303 12665 43315 12699
rect 43257 12659 43315 12665
rect 25593 12631 25651 12637
rect 25593 12628 25605 12631
rect 25464 12600 25605 12628
rect 25464 12588 25470 12600
rect 25593 12597 25605 12600
rect 25639 12597 25651 12631
rect 25593 12591 25651 12597
rect 25682 12588 25688 12640
rect 25740 12628 25746 12640
rect 26697 12631 26755 12637
rect 26697 12628 26709 12631
rect 25740 12600 26709 12628
rect 25740 12588 25746 12600
rect 26697 12597 26709 12600
rect 26743 12597 26755 12631
rect 26697 12591 26755 12597
rect 35161 12631 35219 12637
rect 35161 12597 35173 12631
rect 35207 12628 35219 12631
rect 35250 12628 35256 12640
rect 35207 12600 35256 12628
rect 35207 12597 35219 12600
rect 35161 12591 35219 12597
rect 35250 12588 35256 12600
rect 35308 12588 35314 12640
rect 42981 12631 43039 12637
rect 42981 12597 42993 12631
rect 43027 12628 43039 12631
rect 43272 12628 43300 12659
rect 43530 12628 43536 12640
rect 43027 12600 43536 12628
rect 43027 12597 43039 12600
rect 42981 12591 43039 12597
rect 43530 12588 43536 12600
rect 43588 12588 43594 12640
rect 44450 12588 44456 12640
rect 44508 12628 44514 12640
rect 44775 12631 44833 12637
rect 44775 12628 44787 12631
rect 44508 12600 44787 12628
rect 44508 12588 44514 12600
rect 44775 12597 44787 12600
rect 44821 12597 44833 12631
rect 44775 12591 44833 12597
rect 1104 12538 48852 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 48852 12538
rect 1104 12464 48852 12486
rect 5951 12427 6009 12433
rect 5951 12393 5963 12427
rect 5997 12424 6009 12427
rect 7006 12424 7012 12436
rect 5997 12396 7012 12424
rect 5997 12393 6009 12396
rect 5951 12387 6009 12393
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 8711 12427 8769 12433
rect 8711 12393 8723 12427
rect 8757 12424 8769 12427
rect 8846 12424 8852 12436
rect 8757 12396 8852 12424
rect 8757 12393 8769 12396
rect 8711 12387 8769 12393
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 10192 12396 10701 12424
rect 10192 12384 10198 12396
rect 10689 12393 10701 12396
rect 10735 12393 10747 12427
rect 15102 12424 15108 12436
rect 15063 12396 15108 12424
rect 10689 12387 10747 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15838 12424 15844 12436
rect 15799 12396 15844 12424
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 15930 12384 15936 12436
rect 15988 12424 15994 12436
rect 16485 12427 16543 12433
rect 16485 12424 16497 12427
rect 15988 12396 16497 12424
rect 15988 12384 15994 12396
rect 16485 12393 16497 12396
rect 16531 12424 16543 12427
rect 16942 12424 16948 12436
rect 16531 12396 16948 12424
rect 16531 12393 16543 12396
rect 16485 12387 16543 12393
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 19935 12427 19993 12433
rect 19935 12393 19947 12427
rect 19981 12424 19993 12427
rect 20346 12424 20352 12436
rect 19981 12396 20352 12424
rect 19981 12393 19993 12396
rect 19935 12387 19993 12393
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 22922 12384 22928 12436
rect 22980 12424 22986 12436
rect 24026 12424 24032 12436
rect 22980 12396 23152 12424
rect 22980 12384 22986 12396
rect 6822 12356 6828 12368
rect 6783 12328 6828 12356
rect 6822 12316 6828 12328
rect 6880 12316 6886 12368
rect 7098 12356 7104 12368
rect 7059 12328 7104 12356
rect 7098 12316 7104 12328
rect 7156 12316 7162 12368
rect 7650 12356 7656 12368
rect 7611 12328 7656 12356
rect 7650 12316 7656 12328
rect 7708 12356 7714 12368
rect 9033 12359 9091 12365
rect 9033 12356 9045 12359
rect 7708 12328 9045 12356
rect 7708 12316 7714 12328
rect 9033 12325 9045 12328
rect 9079 12325 9091 12359
rect 9033 12319 9091 12325
rect 9122 12316 9128 12368
rect 9180 12356 9186 12368
rect 9766 12356 9772 12368
rect 9180 12328 9772 12356
rect 9180 12316 9186 12328
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 9858 12316 9864 12368
rect 9916 12356 9922 12368
rect 9916 12328 9961 12356
rect 9916 12316 9922 12328
rect 11606 12316 11612 12368
rect 11664 12356 11670 12368
rect 12802 12356 12808 12368
rect 11664 12328 12808 12356
rect 11664 12316 11670 12328
rect 12802 12316 12808 12328
rect 12860 12316 12866 12368
rect 12897 12359 12955 12365
rect 12897 12325 12909 12359
rect 12943 12356 12955 12359
rect 13170 12356 13176 12368
rect 12943 12328 13176 12356
rect 12943 12325 12955 12328
rect 12897 12319 12955 12325
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 17034 12316 17040 12368
rect 17092 12356 17098 12368
rect 17862 12356 17868 12368
rect 17092 12328 17868 12356
rect 17092 12316 17098 12328
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 17954 12316 17960 12368
rect 18012 12356 18018 12368
rect 18966 12356 18972 12368
rect 18012 12328 18972 12356
rect 18012 12316 18018 12328
rect 18966 12316 18972 12328
rect 19024 12316 19030 12368
rect 20254 12356 20260 12368
rect 20215 12328 20260 12356
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 21082 12356 21088 12368
rect 21043 12328 21088 12356
rect 21082 12316 21088 12328
rect 21140 12316 21146 12368
rect 22830 12316 22836 12368
rect 22888 12356 22894 12368
rect 23124 12365 23152 12396
rect 23676 12396 24032 12424
rect 23676 12365 23704 12396
rect 24026 12384 24032 12396
rect 24084 12424 24090 12436
rect 24305 12427 24363 12433
rect 24305 12424 24317 12427
rect 24084 12396 24317 12424
rect 24084 12384 24090 12396
rect 24305 12393 24317 12396
rect 24351 12424 24363 12427
rect 24578 12424 24584 12436
rect 24351 12396 24584 12424
rect 24351 12393 24363 12396
rect 24305 12387 24363 12393
rect 24578 12384 24584 12396
rect 24636 12384 24642 12436
rect 26329 12427 26387 12433
rect 26329 12393 26341 12427
rect 26375 12424 26387 12427
rect 26694 12424 26700 12436
rect 26375 12396 26700 12424
rect 26375 12393 26387 12396
rect 26329 12387 26387 12393
rect 26694 12384 26700 12396
rect 26752 12384 26758 12436
rect 27709 12427 27767 12433
rect 27709 12393 27721 12427
rect 27755 12424 27767 12427
rect 28074 12424 28080 12436
rect 27755 12396 28080 12424
rect 27755 12393 27767 12396
rect 27709 12387 27767 12393
rect 28074 12384 28080 12396
rect 28132 12384 28138 12436
rect 28902 12384 28908 12436
rect 28960 12424 28966 12436
rect 28997 12427 29055 12433
rect 28997 12424 29009 12427
rect 28960 12396 29009 12424
rect 28960 12384 28966 12396
rect 28997 12393 29009 12396
rect 29043 12393 29055 12427
rect 28997 12387 29055 12393
rect 29549 12427 29607 12433
rect 29549 12393 29561 12427
rect 29595 12424 29607 12427
rect 29730 12424 29736 12436
rect 29595 12396 29736 12424
rect 29595 12393 29607 12396
rect 29549 12387 29607 12393
rect 29730 12384 29736 12396
rect 29788 12384 29794 12436
rect 29914 12424 29920 12436
rect 29875 12396 29920 12424
rect 29914 12384 29920 12396
rect 29972 12384 29978 12436
rect 31573 12427 31631 12433
rect 31573 12393 31585 12427
rect 31619 12424 31631 12427
rect 31662 12424 31668 12436
rect 31619 12396 31668 12424
rect 31619 12393 31631 12396
rect 31573 12387 31631 12393
rect 31662 12384 31668 12396
rect 31720 12384 31726 12436
rect 34698 12384 34704 12436
rect 34756 12424 34762 12436
rect 35253 12427 35311 12433
rect 35253 12424 35265 12427
rect 34756 12396 35265 12424
rect 34756 12384 34762 12396
rect 35253 12393 35265 12396
rect 35299 12393 35311 12427
rect 36170 12424 36176 12436
rect 36131 12396 36176 12424
rect 35253 12387 35311 12393
rect 36170 12384 36176 12396
rect 36228 12384 36234 12436
rect 37875 12427 37933 12433
rect 37875 12393 37887 12427
rect 37921 12424 37933 12427
rect 38194 12424 38200 12436
rect 37921 12396 38200 12424
rect 37921 12393 37933 12396
rect 37875 12387 37933 12393
rect 38194 12384 38200 12396
rect 38252 12384 38258 12436
rect 38933 12427 38991 12433
rect 38933 12393 38945 12427
rect 38979 12424 38991 12427
rect 39114 12424 39120 12436
rect 38979 12396 39120 12424
rect 38979 12393 38991 12396
rect 38933 12387 38991 12393
rect 39114 12384 39120 12396
rect 39172 12384 39178 12436
rect 40589 12427 40647 12433
rect 40589 12393 40601 12427
rect 40635 12424 40647 12427
rect 43162 12424 43168 12436
rect 40635 12396 41644 12424
rect 43123 12396 43168 12424
rect 40635 12393 40647 12396
rect 40589 12387 40647 12393
rect 23017 12359 23075 12365
rect 23017 12356 23029 12359
rect 22888 12328 23029 12356
rect 22888 12316 22894 12328
rect 23017 12325 23029 12328
rect 23063 12325 23075 12359
rect 23017 12319 23075 12325
rect 23109 12359 23167 12365
rect 23109 12325 23121 12359
rect 23155 12325 23167 12359
rect 23109 12319 23167 12325
rect 23661 12359 23719 12365
rect 23661 12325 23673 12359
rect 23707 12325 23719 12359
rect 23934 12356 23940 12368
rect 23895 12328 23940 12356
rect 23661 12319 23719 12325
rect 23934 12316 23940 12328
rect 23992 12316 23998 12368
rect 24394 12316 24400 12368
rect 24452 12356 24458 12368
rect 24765 12359 24823 12365
rect 24765 12356 24777 12359
rect 24452 12328 24777 12356
rect 24452 12316 24458 12328
rect 24765 12325 24777 12328
rect 24811 12325 24823 12359
rect 24765 12319 24823 12325
rect 24857 12359 24915 12365
rect 24857 12325 24869 12359
rect 24903 12356 24915 12359
rect 25222 12356 25228 12368
rect 24903 12328 25228 12356
rect 24903 12325 24915 12328
rect 24857 12319 24915 12325
rect 25222 12316 25228 12328
rect 25280 12316 25286 12368
rect 25409 12359 25467 12365
rect 25409 12325 25421 12359
rect 25455 12356 25467 12359
rect 25866 12356 25872 12368
rect 25455 12328 25872 12356
rect 25455 12325 25467 12328
rect 25409 12319 25467 12325
rect 25866 12316 25872 12328
rect 25924 12316 25930 12368
rect 27614 12356 27620 12368
rect 26804 12328 27620 12356
rect 5442 12248 5448 12300
rect 5500 12288 5506 12300
rect 5848 12291 5906 12297
rect 5848 12288 5860 12291
rect 5500 12260 5860 12288
rect 5500 12248 5506 12260
rect 5848 12257 5860 12260
rect 5894 12288 5906 12291
rect 6086 12288 6092 12300
rect 5894 12260 6092 12288
rect 5894 12257 5906 12260
rect 5848 12251 5906 12257
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 8481 12291 8539 12297
rect 8481 12257 8493 12291
rect 8527 12288 8539 12291
rect 8570 12288 8576 12300
rect 8527 12260 8576 12288
rect 8527 12257 8539 12260
rect 8481 12251 8539 12257
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 15378 12248 15384 12300
rect 15436 12288 15442 12300
rect 15473 12291 15531 12297
rect 15473 12288 15485 12291
rect 15436 12260 15485 12288
rect 15436 12248 15442 12260
rect 15473 12257 15485 12260
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 18874 12248 18880 12300
rect 18932 12288 18938 12300
rect 19150 12288 19156 12300
rect 18932 12260 19156 12288
rect 18932 12248 18938 12260
rect 19150 12248 19156 12260
rect 19208 12288 19214 12300
rect 19832 12291 19890 12297
rect 19832 12288 19844 12291
rect 19208 12260 19844 12288
rect 19208 12248 19214 12260
rect 19832 12257 19844 12260
rect 19878 12257 19890 12291
rect 19832 12251 19890 12257
rect 26602 12248 26608 12300
rect 26660 12288 26666 12300
rect 26804 12297 26832 12328
rect 27614 12316 27620 12328
rect 27672 12316 27678 12368
rect 30558 12356 30564 12368
rect 30519 12328 30564 12356
rect 30558 12316 30564 12328
rect 30616 12316 30622 12368
rect 31680 12356 31708 12384
rect 32030 12356 32036 12368
rect 31680 12328 32036 12356
rect 32030 12316 32036 12328
rect 32088 12356 32094 12368
rect 32309 12359 32367 12365
rect 32309 12356 32321 12359
rect 32088 12328 32321 12356
rect 32088 12316 32094 12328
rect 32309 12325 32321 12328
rect 32355 12325 32367 12359
rect 34422 12356 34428 12368
rect 34383 12328 34428 12356
rect 32309 12319 32367 12325
rect 34422 12316 34428 12328
rect 34480 12316 34486 12368
rect 34790 12316 34796 12368
rect 34848 12356 34854 12368
rect 34977 12359 35035 12365
rect 34977 12356 34989 12359
rect 34848 12328 34989 12356
rect 34848 12316 34854 12328
rect 34977 12325 34989 12328
rect 35023 12356 35035 12359
rect 35158 12356 35164 12368
rect 35023 12328 35164 12356
rect 35023 12325 35035 12328
rect 34977 12319 35035 12325
rect 35158 12316 35164 12328
rect 35216 12316 35222 12368
rect 39666 12316 39672 12368
rect 39724 12356 39730 12368
rect 39942 12356 39948 12368
rect 39724 12328 39948 12356
rect 39724 12316 39730 12328
rect 39942 12316 39948 12328
rect 40000 12365 40006 12368
rect 40000 12359 40048 12365
rect 40000 12325 40002 12359
rect 40036 12325 40048 12359
rect 40862 12356 40868 12368
rect 40823 12328 40868 12356
rect 40000 12319 40048 12325
rect 40000 12316 40006 12319
rect 40862 12316 40868 12328
rect 40920 12316 40926 12368
rect 41616 12365 41644 12396
rect 43162 12384 43168 12396
rect 43220 12384 43226 12436
rect 41601 12359 41659 12365
rect 41601 12325 41613 12359
rect 41647 12356 41659 12359
rect 42242 12356 42248 12368
rect 41647 12328 42248 12356
rect 41647 12325 41659 12328
rect 41601 12319 41659 12325
rect 42242 12316 42248 12328
rect 42300 12316 42306 12368
rect 43530 12356 43536 12368
rect 43491 12328 43536 12356
rect 43530 12316 43536 12328
rect 43588 12316 43594 12368
rect 44085 12359 44143 12365
rect 44085 12325 44097 12359
rect 44131 12356 44143 12359
rect 44174 12356 44180 12368
rect 44131 12328 44180 12356
rect 44131 12325 44143 12328
rect 44085 12319 44143 12325
rect 44174 12316 44180 12328
rect 44232 12316 44238 12368
rect 26789 12291 26847 12297
rect 26789 12288 26801 12291
rect 26660 12260 26801 12288
rect 26660 12248 26666 12260
rect 26789 12257 26801 12260
rect 26835 12257 26847 12291
rect 26970 12288 26976 12300
rect 26931 12260 26976 12288
rect 26789 12251 26847 12257
rect 26970 12248 26976 12260
rect 27028 12248 27034 12300
rect 31113 12291 31171 12297
rect 31113 12257 31125 12291
rect 31159 12288 31171 12291
rect 31294 12288 31300 12300
rect 31159 12260 31300 12288
rect 31159 12257 31171 12260
rect 31113 12251 31171 12257
rect 31294 12248 31300 12260
rect 31352 12248 31358 12300
rect 36078 12248 36084 12300
rect 36136 12288 36142 12300
rect 36633 12291 36691 12297
rect 36633 12288 36645 12291
rect 36136 12260 36645 12288
rect 36136 12248 36142 12260
rect 36633 12257 36645 12260
rect 36679 12288 36691 12291
rect 36722 12288 36728 12300
rect 36679 12260 36728 12288
rect 36679 12257 36691 12260
rect 36633 12251 36691 12257
rect 36722 12248 36728 12260
rect 36780 12248 36786 12300
rect 37804 12291 37862 12297
rect 37804 12257 37816 12291
rect 37850 12288 37862 12291
rect 38010 12288 38016 12300
rect 37850 12260 38016 12288
rect 37850 12257 37862 12260
rect 37804 12251 37862 12257
rect 38010 12248 38016 12260
rect 38068 12248 38074 12300
rect 7006 12220 7012 12232
rect 6967 12192 7012 12220
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 10045 12223 10103 12229
rect 10045 12220 10057 12223
rect 9272 12192 10057 12220
rect 9272 12180 9278 12192
rect 10045 12189 10057 12192
rect 10091 12220 10103 12223
rect 12158 12220 12164 12232
rect 10091 12192 12164 12220
rect 10091 12189 10103 12192
rect 10045 12183 10103 12189
rect 12158 12180 12164 12192
rect 12216 12180 12222 12232
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 14274 12220 14280 12232
rect 13495 12192 14280 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 20990 12220 20996 12232
rect 20951 12192 20996 12220
rect 20990 12180 20996 12192
rect 21048 12180 21054 12232
rect 25774 12180 25780 12232
rect 25832 12220 25838 12232
rect 25869 12223 25927 12229
rect 25869 12220 25881 12223
rect 25832 12192 25881 12220
rect 25832 12180 25838 12192
rect 25869 12189 25881 12192
rect 25915 12220 25927 12223
rect 27065 12223 27123 12229
rect 27065 12220 27077 12223
rect 25915 12192 27077 12220
rect 25915 12189 25927 12192
rect 25869 12183 25927 12189
rect 27065 12189 27077 12192
rect 27111 12189 27123 12223
rect 28626 12220 28632 12232
rect 28587 12192 28632 12220
rect 27065 12183 27123 12189
rect 28626 12180 28632 12192
rect 28684 12180 28690 12232
rect 30466 12220 30472 12232
rect 30427 12192 30472 12220
rect 30466 12180 30472 12192
rect 30524 12180 30530 12232
rect 32214 12220 32220 12232
rect 32175 12192 32220 12220
rect 32214 12180 32220 12192
rect 32272 12180 32278 12232
rect 32582 12220 32588 12232
rect 32543 12192 32588 12220
rect 32582 12180 32588 12192
rect 32640 12180 32646 12232
rect 34333 12223 34391 12229
rect 34333 12189 34345 12223
rect 34379 12189 34391 12223
rect 39666 12220 39672 12232
rect 39627 12192 39672 12220
rect 34333 12183 34391 12189
rect 18414 12152 18420 12164
rect 18375 12124 18420 12152
rect 18414 12112 18420 12124
rect 18472 12112 18478 12164
rect 21542 12152 21548 12164
rect 21503 12124 21548 12152
rect 21542 12112 21548 12124
rect 21600 12112 21606 12164
rect 34238 12112 34244 12164
rect 34296 12152 34302 12164
rect 34348 12152 34376 12183
rect 39666 12180 39672 12192
rect 39724 12180 39730 12232
rect 40770 12180 40776 12232
rect 40828 12220 40834 12232
rect 41506 12220 41512 12232
rect 40828 12192 41512 12220
rect 40828 12180 40834 12192
rect 41506 12180 41512 12192
rect 41564 12180 41570 12232
rect 41874 12220 41880 12232
rect 41835 12192 41880 12220
rect 41874 12180 41880 12192
rect 41932 12180 41938 12232
rect 43441 12223 43499 12229
rect 43441 12189 43453 12223
rect 43487 12220 43499 12223
rect 44450 12220 44456 12232
rect 43487 12192 44456 12220
rect 43487 12189 43499 12192
rect 43441 12183 43499 12189
rect 44450 12180 44456 12192
rect 44508 12180 44514 12232
rect 41322 12152 41328 12164
rect 34296 12124 34376 12152
rect 41235 12124 41328 12152
rect 34296 12112 34302 12124
rect 41322 12112 41328 12124
rect 41380 12152 41386 12164
rect 42150 12152 42156 12164
rect 41380 12124 42156 12152
rect 41380 12112 41386 12124
rect 42150 12112 42156 12124
rect 42208 12152 42214 12164
rect 43346 12152 43352 12164
rect 42208 12124 43352 12152
rect 42208 12112 42214 12124
rect 43346 12112 43352 12124
rect 43404 12112 43410 12164
rect 11606 12084 11612 12096
rect 11567 12056 11612 12084
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 11839 12087 11897 12093
rect 11839 12053 11851 12087
rect 11885 12084 11897 12087
rect 13262 12084 13268 12096
rect 11885 12056 13268 12084
rect 11885 12053 11897 12056
rect 11839 12047 11897 12053
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 23198 12084 23204 12096
rect 14148 12056 23204 12084
rect 14148 12044 14154 12056
rect 23198 12044 23204 12056
rect 23256 12044 23262 12096
rect 31570 12044 31576 12096
rect 31628 12084 31634 12096
rect 31941 12087 31999 12093
rect 31941 12084 31953 12087
rect 31628 12056 31953 12084
rect 31628 12044 31634 12056
rect 31941 12053 31953 12056
rect 31987 12084 31999 12087
rect 33778 12084 33784 12096
rect 31987 12056 33784 12084
rect 31987 12053 31999 12056
rect 31941 12047 31999 12053
rect 33778 12044 33784 12056
rect 33836 12044 33842 12096
rect 36771 12087 36829 12093
rect 36771 12053 36783 12087
rect 36817 12084 36829 12087
rect 36906 12084 36912 12096
rect 36817 12056 36912 12084
rect 36817 12053 36829 12056
rect 36771 12047 36829 12053
rect 36906 12044 36912 12056
rect 36964 12044 36970 12096
rect 37090 12084 37096 12096
rect 37051 12056 37096 12084
rect 37090 12044 37096 12056
rect 37148 12044 37154 12096
rect 1104 11994 48852 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 48852 11994
rect 1104 11920 48852 11942
rect 5767 11883 5825 11889
rect 5767 11849 5779 11883
rect 5813 11880 5825 11883
rect 7006 11880 7012 11892
rect 5813 11852 7012 11880
rect 5813 11849 5825 11852
rect 5767 11843 5825 11849
rect 7006 11840 7012 11852
rect 7064 11880 7070 11892
rect 7377 11883 7435 11889
rect 7377 11880 7389 11883
rect 7064 11852 7389 11880
rect 7064 11840 7070 11852
rect 7377 11849 7389 11852
rect 7423 11849 7435 11883
rect 8570 11880 8576 11892
rect 8531 11852 8576 11880
rect 7377 11843 7435 11849
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 10045 11883 10103 11889
rect 10045 11880 10057 11883
rect 9824 11852 10057 11880
rect 9824 11840 9830 11852
rect 10045 11849 10057 11852
rect 10091 11849 10103 11883
rect 10045 11843 10103 11849
rect 11425 11883 11483 11889
rect 11425 11849 11437 11883
rect 11471 11880 11483 11883
rect 11514 11880 11520 11892
rect 11471 11852 11520 11880
rect 11471 11849 11483 11852
rect 11425 11843 11483 11849
rect 6086 11812 6092 11824
rect 6047 11784 6092 11812
rect 6086 11772 6092 11784
rect 6144 11772 6150 11824
rect 7098 11812 7104 11824
rect 7059 11784 7104 11812
rect 7098 11772 7104 11784
rect 7156 11772 7162 11824
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11744 9827 11747
rect 9858 11744 9864 11756
rect 9815 11716 9864 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 5664 11679 5722 11685
rect 5664 11676 5676 11679
rect 5592 11648 5676 11676
rect 5592 11636 5598 11648
rect 5664 11645 5676 11648
rect 5710 11676 5722 11679
rect 6457 11679 6515 11685
rect 6457 11676 6469 11679
rect 5710 11648 6469 11676
rect 5710 11645 5722 11648
rect 5664 11639 5722 11645
rect 6457 11645 6469 11648
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 10873 11679 10931 11685
rect 10873 11645 10885 11679
rect 10919 11676 10931 11679
rect 11440 11676 11468 11843
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 13265 11883 13323 11889
rect 13265 11880 13277 11883
rect 12860 11852 13277 11880
rect 12860 11840 12866 11852
rect 13265 11849 13277 11852
rect 13311 11849 13323 11883
rect 13265 11843 13323 11849
rect 14182 11840 14188 11892
rect 14240 11840 14246 11892
rect 14366 11840 14372 11892
rect 14424 11880 14430 11892
rect 14921 11883 14979 11889
rect 14921 11880 14933 11883
rect 14424 11852 14933 11880
rect 14424 11840 14430 11852
rect 14921 11849 14933 11852
rect 14967 11849 14979 11883
rect 17862 11880 17868 11892
rect 17823 11852 17868 11880
rect 14921 11843 14979 11849
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 11793 11815 11851 11821
rect 11793 11812 11805 11815
rect 11664 11784 11805 11812
rect 11664 11772 11670 11784
rect 11793 11781 11805 11784
rect 11839 11812 11851 11815
rect 14200 11812 14228 11840
rect 14826 11812 14832 11824
rect 11839 11784 14832 11812
rect 11839 11781 11851 11784
rect 11793 11775 11851 11781
rect 14826 11772 14832 11784
rect 14884 11772 14890 11824
rect 12575 11747 12633 11753
rect 12575 11713 12587 11747
rect 12621 11744 12633 11747
rect 14090 11744 14096 11756
rect 12621 11716 14096 11744
rect 12621 11713 12633 11716
rect 12575 11707 12633 11713
rect 14090 11704 14096 11716
rect 14148 11704 14154 11756
rect 14274 11744 14280 11756
rect 14235 11716 14280 11744
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 12472 11679 12530 11685
rect 12472 11676 12484 11679
rect 10919 11648 11468 11676
rect 12268 11648 12484 11676
rect 10919 11645 10931 11648
rect 10873 11639 10931 11645
rect 12268 11552 12296 11648
rect 12472 11645 12484 11648
rect 12518 11645 12530 11679
rect 14936 11676 14964 11843
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 18322 11840 18328 11892
rect 18380 11880 18386 11892
rect 18463 11883 18521 11889
rect 18463 11880 18475 11883
rect 18380 11852 18475 11880
rect 18380 11840 18386 11852
rect 18463 11849 18475 11852
rect 18509 11849 18521 11883
rect 18463 11843 18521 11849
rect 19334 11840 19340 11892
rect 19392 11880 19398 11892
rect 19613 11883 19671 11889
rect 19613 11880 19625 11883
rect 19392 11852 19625 11880
rect 19392 11840 19398 11852
rect 19613 11849 19625 11852
rect 19659 11880 19671 11883
rect 20070 11880 20076 11892
rect 19659 11852 20076 11880
rect 19659 11849 19671 11852
rect 19613 11843 19671 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 20625 11883 20683 11889
rect 20625 11849 20637 11883
rect 20671 11880 20683 11883
rect 20993 11883 21051 11889
rect 20993 11880 21005 11883
rect 20671 11852 21005 11880
rect 20671 11849 20683 11852
rect 20625 11843 20683 11849
rect 20993 11849 21005 11852
rect 21039 11880 21051 11883
rect 21082 11880 21088 11892
rect 21039 11852 21088 11880
rect 21039 11849 21051 11852
rect 20993 11843 21051 11849
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 22603 11883 22661 11889
rect 22603 11849 22615 11883
rect 22649 11880 22661 11883
rect 24118 11880 24124 11892
rect 22649 11852 24124 11880
rect 22649 11849 22661 11852
rect 22603 11843 22661 11849
rect 24118 11840 24124 11852
rect 24176 11840 24182 11892
rect 26602 11880 26608 11892
rect 26563 11852 26608 11880
rect 26602 11840 26608 11852
rect 26660 11840 26666 11892
rect 30193 11883 30251 11889
rect 30193 11849 30205 11883
rect 30239 11880 30251 11883
rect 30558 11880 30564 11892
rect 30239 11852 30564 11880
rect 30239 11849 30251 11852
rect 30193 11843 30251 11849
rect 30558 11840 30564 11852
rect 30616 11840 30622 11892
rect 32030 11840 32036 11892
rect 32088 11880 32094 11892
rect 32125 11883 32183 11889
rect 32125 11880 32137 11883
rect 32088 11852 32137 11880
rect 32088 11840 32094 11852
rect 32125 11849 32137 11852
rect 32171 11849 32183 11883
rect 32125 11843 32183 11849
rect 34422 11840 34428 11892
rect 34480 11880 34486 11892
rect 34609 11883 34667 11889
rect 34609 11880 34621 11883
rect 34480 11852 34621 11880
rect 34480 11840 34486 11852
rect 34609 11849 34621 11852
rect 34655 11849 34667 11883
rect 38010 11880 38016 11892
rect 37971 11852 38016 11880
rect 34609 11843 34667 11849
rect 38010 11840 38016 11852
rect 38068 11840 38074 11892
rect 38654 11880 38660 11892
rect 38615 11852 38660 11880
rect 38654 11840 38660 11852
rect 38712 11840 38718 11892
rect 39942 11880 39948 11892
rect 39903 11852 39948 11880
rect 39942 11840 39948 11852
rect 40000 11840 40006 11892
rect 40770 11880 40776 11892
rect 40731 11852 40776 11880
rect 40770 11840 40776 11852
rect 40828 11840 40834 11892
rect 42242 11880 42248 11892
rect 42203 11852 42248 11880
rect 42242 11840 42248 11852
rect 42300 11840 42306 11892
rect 43070 11840 43076 11892
rect 43128 11880 43134 11892
rect 44450 11880 44456 11892
rect 43128 11852 44220 11880
rect 44411 11852 44456 11880
rect 43128 11840 43134 11852
rect 17497 11815 17555 11821
rect 17497 11781 17509 11815
rect 17543 11812 17555 11815
rect 17954 11812 17960 11824
rect 17543 11784 17960 11812
rect 17543 11781 17555 11784
rect 17497 11775 17555 11781
rect 17954 11772 17960 11784
rect 18012 11772 18018 11824
rect 23566 11772 23572 11824
rect 23624 11812 23630 11824
rect 25498 11812 25504 11824
rect 23624 11784 25504 11812
rect 23624 11772 23630 11784
rect 19705 11747 19763 11753
rect 19705 11713 19717 11747
rect 19751 11744 19763 11747
rect 20254 11744 20260 11756
rect 19751 11716 20260 11744
rect 19751 11713 19763 11716
rect 19705 11707 19763 11713
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 21358 11704 21364 11756
rect 21416 11744 21422 11756
rect 21453 11747 21511 11753
rect 21453 11744 21465 11747
rect 21416 11716 21465 11744
rect 21416 11704 21422 11716
rect 21453 11713 21465 11716
rect 21499 11713 21511 11747
rect 24026 11744 24032 11756
rect 23987 11716 24032 11744
rect 21453 11707 21511 11713
rect 24026 11704 24032 11716
rect 24084 11704 24090 11756
rect 24320 11753 24348 11784
rect 25498 11772 25504 11784
rect 25556 11812 25562 11824
rect 26145 11815 26203 11821
rect 26145 11812 26157 11815
rect 25556 11784 26157 11812
rect 25556 11772 25562 11784
rect 26145 11781 26157 11784
rect 26191 11781 26203 11815
rect 26145 11775 26203 11781
rect 30466 11772 30472 11824
rect 30524 11812 30530 11824
rect 30837 11815 30895 11821
rect 30837 11812 30849 11815
rect 30524 11784 30849 11812
rect 30524 11772 30530 11784
rect 30837 11781 30849 11784
rect 30883 11781 30895 11815
rect 36722 11812 36728 11824
rect 36635 11784 36728 11812
rect 30837 11775 30895 11781
rect 36722 11772 36728 11784
rect 36780 11812 36786 11824
rect 41874 11812 41880 11824
rect 36780 11784 41736 11812
rect 41835 11784 41880 11812
rect 36780 11772 36786 11784
rect 41708 11756 41736 11784
rect 41874 11772 41880 11784
rect 41932 11772 41938 11824
rect 44192 11812 44220 11852
rect 44450 11840 44456 11852
rect 44508 11840 44514 11892
rect 44683 11815 44741 11821
rect 44683 11812 44695 11815
rect 42766 11784 44128 11812
rect 44192 11784 44695 11812
rect 24305 11747 24363 11753
rect 24305 11713 24317 11747
rect 24351 11713 24363 11747
rect 24305 11707 24363 11713
rect 25593 11747 25651 11753
rect 25593 11713 25605 11747
rect 25639 11744 25651 11747
rect 25866 11744 25872 11756
rect 25639 11716 25872 11744
rect 25639 11713 25651 11716
rect 25593 11707 25651 11713
rect 25866 11704 25872 11716
rect 25924 11704 25930 11756
rect 31435 11747 31493 11753
rect 31435 11713 31447 11747
rect 31481 11744 31493 11747
rect 32214 11744 32220 11756
rect 31481 11716 32220 11744
rect 31481 11713 31493 11716
rect 31435 11707 31493 11713
rect 32214 11704 32220 11716
rect 32272 11744 32278 11756
rect 32493 11747 32551 11753
rect 32493 11744 32505 11747
rect 32272 11716 32505 11744
rect 32272 11704 32278 11716
rect 32493 11713 32505 11716
rect 32539 11713 32551 11747
rect 35250 11744 35256 11756
rect 35211 11716 35256 11744
rect 32493 11707 32551 11713
rect 35250 11704 35256 11716
rect 35308 11704 35314 11756
rect 36538 11704 36544 11756
rect 36596 11744 36602 11756
rect 37093 11747 37151 11753
rect 37093 11744 37105 11747
rect 36596 11716 37105 11744
rect 36596 11704 36602 11716
rect 37093 11713 37105 11716
rect 37139 11744 37151 11747
rect 37458 11744 37464 11756
rect 37139 11716 37464 11744
rect 37139 11713 37151 11716
rect 37093 11707 37151 11713
rect 37458 11704 37464 11716
rect 37516 11704 37522 11756
rect 37737 11747 37795 11753
rect 37737 11713 37749 11747
rect 37783 11744 37795 11747
rect 37918 11744 37924 11756
rect 37783 11716 37924 11744
rect 37783 11713 37795 11716
rect 37737 11707 37795 11713
rect 37918 11704 37924 11716
rect 37976 11744 37982 11756
rect 38470 11744 38476 11756
rect 37976 11716 38476 11744
rect 37976 11704 37982 11716
rect 38470 11704 38476 11716
rect 38528 11704 38534 11756
rect 39577 11747 39635 11753
rect 39577 11713 39589 11747
rect 39623 11744 39635 11747
rect 39666 11744 39672 11756
rect 39623 11716 39672 11744
rect 39623 11713 39635 11716
rect 39577 11707 39635 11713
rect 39666 11704 39672 11716
rect 39724 11744 39730 11756
rect 40221 11747 40279 11753
rect 40221 11744 40233 11747
rect 39724 11716 40233 11744
rect 39724 11704 39730 11716
rect 40221 11713 40233 11716
rect 40267 11713 40279 11747
rect 41322 11744 41328 11756
rect 41283 11716 41328 11744
rect 40221 11707 40279 11713
rect 41322 11704 41328 11716
rect 41380 11704 41386 11756
rect 41690 11704 41696 11756
rect 41748 11744 41754 11756
rect 42766 11744 42794 11784
rect 43070 11744 43076 11756
rect 41748 11716 42794 11744
rect 43031 11716 43076 11744
rect 41748 11704 41754 11716
rect 43070 11704 43076 11716
rect 43128 11704 43134 11756
rect 43346 11744 43352 11756
rect 43307 11716 43352 11744
rect 43346 11704 43352 11716
rect 43404 11704 43410 11756
rect 15565 11679 15623 11685
rect 15565 11676 15577 11679
rect 14936 11648 15577 11676
rect 12472 11639 12530 11645
rect 15565 11645 15577 11648
rect 15611 11645 15623 11679
rect 15565 11639 15623 11645
rect 17678 11636 17684 11688
rect 17736 11676 17742 11688
rect 18414 11685 18420 11688
rect 18360 11679 18420 11685
rect 18360 11676 18372 11679
rect 17736 11648 18372 11676
rect 17736 11636 17742 11648
rect 18360 11645 18372 11648
rect 18406 11645 18420 11679
rect 18360 11639 18420 11645
rect 18414 11636 18420 11639
rect 18472 11676 18478 11688
rect 18785 11679 18843 11685
rect 18785 11676 18797 11679
rect 18472 11648 18797 11676
rect 18472 11636 18478 11648
rect 18785 11645 18797 11648
rect 18831 11645 18843 11679
rect 18785 11639 18843 11645
rect 21542 11636 21548 11688
rect 21600 11676 21606 11688
rect 22500 11679 22558 11685
rect 22500 11676 22512 11679
rect 21600 11648 22512 11676
rect 21600 11636 21606 11648
rect 22500 11645 22512 11648
rect 22546 11676 22558 11679
rect 22925 11679 22983 11685
rect 22925 11676 22937 11679
rect 22546 11648 22937 11676
rect 22546 11645 22558 11648
rect 22500 11639 22558 11645
rect 22925 11645 22937 11648
rect 22971 11645 22983 11679
rect 27522 11676 27528 11688
rect 27435 11648 27528 11676
rect 22925 11639 22983 11645
rect 27522 11636 27528 11648
rect 27580 11676 27586 11688
rect 27798 11676 27804 11688
rect 27580 11648 27804 11676
rect 27580 11636 27586 11648
rect 27798 11636 27804 11648
rect 27856 11636 27862 11688
rect 28074 11676 28080 11688
rect 28035 11648 28080 11676
rect 28074 11636 28080 11648
rect 28132 11636 28138 11688
rect 28353 11679 28411 11685
rect 28353 11645 28365 11679
rect 28399 11676 28411 11679
rect 29270 11676 29276 11688
rect 28399 11648 29276 11676
rect 28399 11645 28411 11648
rect 28353 11639 28411 11645
rect 29270 11636 29276 11648
rect 29328 11636 29334 11688
rect 31202 11636 31208 11688
rect 31260 11676 31266 11688
rect 31332 11679 31390 11685
rect 31332 11676 31344 11679
rect 31260 11648 31344 11676
rect 31260 11636 31266 11648
rect 31332 11645 31344 11648
rect 31378 11676 31390 11679
rect 31754 11676 31760 11688
rect 31378 11648 31760 11676
rect 31378 11645 31390 11648
rect 31332 11639 31390 11645
rect 31754 11636 31760 11648
rect 31812 11636 31818 11688
rect 33226 11676 33232 11688
rect 33187 11648 33232 11676
rect 33226 11636 33232 11648
rect 33284 11636 33290 11688
rect 33781 11679 33839 11685
rect 33781 11645 33793 11679
rect 33827 11676 33839 11679
rect 33962 11676 33968 11688
rect 33827 11648 33968 11676
rect 33827 11645 33839 11648
rect 33781 11639 33839 11645
rect 13998 11608 14004 11620
rect 13959 11580 14004 11608
rect 13998 11568 14004 11580
rect 14056 11568 14062 11620
rect 14093 11611 14151 11617
rect 14093 11577 14105 11611
rect 14139 11577 14151 11611
rect 15473 11611 15531 11617
rect 15473 11608 15485 11611
rect 14093 11571 14151 11577
rect 14752 11580 15485 11608
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 10284 11512 11069 11540
rect 10284 11500 10290 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 12250 11540 12256 11552
rect 12211 11512 12256 11540
rect 11057 11503 11115 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 12989 11543 13047 11549
rect 12989 11509 13001 11543
rect 13035 11540 13047 11543
rect 13170 11540 13176 11552
rect 13035 11512 13176 11540
rect 13035 11509 13047 11512
rect 12989 11503 13047 11509
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13354 11500 13360 11552
rect 13412 11540 13418 11552
rect 13817 11543 13875 11549
rect 13817 11540 13829 11543
rect 13412 11512 13829 11540
rect 13412 11500 13418 11512
rect 13817 11509 13829 11512
rect 13863 11540 13875 11543
rect 14108 11540 14136 11571
rect 14752 11540 14780 11580
rect 15473 11577 15485 11580
rect 15519 11577 15531 11611
rect 24118 11608 24124 11620
rect 24079 11580 24124 11608
rect 15473 11571 15531 11577
rect 24118 11568 24124 11580
rect 24176 11568 24182 11620
rect 25682 11568 25688 11620
rect 25740 11608 25746 11620
rect 27157 11611 27215 11617
rect 25740 11580 25785 11608
rect 25740 11568 25746 11580
rect 27157 11577 27169 11611
rect 27203 11608 27215 11611
rect 28092 11608 28120 11636
rect 29594 11611 29652 11617
rect 29594 11608 29606 11611
rect 27203 11580 28120 11608
rect 29012 11580 29606 11608
rect 27203 11577 27215 11580
rect 27157 11571 27215 11577
rect 15378 11540 15384 11552
rect 13863 11512 14780 11540
rect 15339 11512 15384 11540
rect 13863 11509 13875 11512
rect 13817 11503 13875 11509
rect 15378 11500 15384 11512
rect 15436 11500 15442 11552
rect 18874 11500 18880 11552
rect 18932 11540 18938 11552
rect 19153 11543 19211 11549
rect 19153 11540 19165 11543
rect 18932 11512 19165 11540
rect 18932 11500 18938 11512
rect 19153 11509 19165 11512
rect 19199 11509 19211 11543
rect 20070 11540 20076 11552
rect 20031 11512 20076 11540
rect 19153 11503 19211 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20438 11500 20444 11552
rect 20496 11540 20502 11552
rect 20990 11540 20996 11552
rect 20496 11512 20996 11540
rect 20496 11500 20502 11512
rect 20990 11500 20996 11512
rect 21048 11540 21054 11552
rect 21269 11543 21327 11549
rect 21269 11540 21281 11543
rect 21048 11512 21281 11540
rect 21048 11500 21054 11512
rect 21269 11509 21281 11512
rect 21315 11509 21327 11543
rect 21269 11503 21327 11509
rect 22922 11500 22928 11552
rect 22980 11540 22986 11552
rect 23385 11543 23443 11549
rect 23385 11540 23397 11543
rect 22980 11512 23397 11540
rect 22980 11500 22986 11512
rect 23385 11509 23397 11512
rect 23431 11540 23443 11543
rect 25041 11543 25099 11549
rect 25041 11540 25053 11543
rect 23431 11512 25053 11540
rect 23431 11509 23443 11512
rect 23385 11503 23443 11509
rect 25041 11509 25053 11512
rect 25087 11540 25099 11543
rect 25222 11540 25228 11552
rect 25087 11512 25228 11540
rect 25087 11509 25099 11512
rect 25041 11503 25099 11509
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 25409 11543 25467 11549
rect 25409 11509 25421 11543
rect 25455 11540 25467 11543
rect 25700 11540 25728 11568
rect 25455 11512 25728 11540
rect 25455 11509 25467 11512
rect 25409 11503 25467 11509
rect 26694 11500 26700 11552
rect 26752 11540 26758 11552
rect 28629 11543 28687 11549
rect 28629 11540 28641 11543
rect 26752 11512 28641 11540
rect 26752 11500 26758 11512
rect 28629 11509 28641 11512
rect 28675 11540 28687 11543
rect 28902 11540 28908 11552
rect 28675 11512 28908 11540
rect 28675 11509 28687 11512
rect 28629 11503 28687 11509
rect 28902 11500 28908 11512
rect 28960 11540 28966 11552
rect 29012 11549 29040 11580
rect 29594 11577 29606 11580
rect 29640 11577 29652 11611
rect 29594 11571 29652 11577
rect 33137 11611 33195 11617
rect 33137 11577 33149 11611
rect 33183 11608 33195 11611
rect 33796 11608 33824 11639
rect 33962 11636 33968 11648
rect 34020 11636 34026 11688
rect 38654 11636 38660 11688
rect 38712 11676 38718 11688
rect 38841 11679 38899 11685
rect 38841 11676 38853 11679
rect 38712 11648 38853 11676
rect 38712 11636 38718 11648
rect 38841 11645 38853 11648
rect 38887 11645 38899 11679
rect 38841 11639 38899 11645
rect 39114 11636 39120 11688
rect 39172 11676 39178 11688
rect 39301 11679 39359 11685
rect 39301 11676 39313 11679
rect 39172 11648 39313 11676
rect 39172 11636 39178 11648
rect 39301 11645 39313 11648
rect 39347 11645 39359 11679
rect 44100 11676 44128 11784
rect 44683 11781 44695 11784
rect 44729 11781 44741 11815
rect 44683 11775 44741 11781
rect 44580 11679 44638 11685
rect 44580 11676 44592 11679
rect 44100 11648 44592 11676
rect 39301 11639 39359 11645
rect 44580 11645 44592 11648
rect 44626 11676 44638 11679
rect 45005 11679 45063 11685
rect 45005 11676 45017 11679
rect 44626 11648 45017 11676
rect 44626 11645 44638 11648
rect 44580 11639 44638 11645
rect 45005 11645 45017 11648
rect 45051 11645 45063 11679
rect 45005 11639 45063 11645
rect 35574 11611 35632 11617
rect 35574 11608 35586 11611
rect 33183 11580 33824 11608
rect 35084 11580 35586 11608
rect 33183 11577 33195 11580
rect 33137 11571 33195 11577
rect 35084 11552 35112 11580
rect 35574 11577 35586 11580
rect 35620 11577 35632 11611
rect 35574 11571 35632 11577
rect 37185 11611 37243 11617
rect 37185 11577 37197 11611
rect 37231 11577 37243 11611
rect 37185 11571 37243 11577
rect 41417 11611 41475 11617
rect 41417 11577 41429 11611
rect 41463 11608 41475 11611
rect 41506 11608 41512 11620
rect 41463 11580 41512 11608
rect 41463 11577 41475 11580
rect 41417 11571 41475 11577
rect 28997 11543 29055 11549
rect 28997 11540 29009 11543
rect 28960 11512 29009 11540
rect 28960 11500 28966 11512
rect 28997 11509 29009 11512
rect 29043 11509 29055 11543
rect 33502 11540 33508 11552
rect 33463 11512 33508 11540
rect 28997 11503 29055 11509
rect 33502 11500 33508 11512
rect 33560 11500 33566 11552
rect 34238 11540 34244 11552
rect 34199 11512 34244 11540
rect 34238 11500 34244 11512
rect 34296 11500 34302 11552
rect 35066 11540 35072 11552
rect 35027 11512 35072 11540
rect 35066 11500 35072 11512
rect 35124 11500 35130 11552
rect 36170 11540 36176 11552
rect 36131 11512 36176 11540
rect 36170 11500 36176 11512
rect 36228 11500 36234 11552
rect 36998 11500 37004 11552
rect 37056 11540 37062 11552
rect 37200 11540 37228 11571
rect 37734 11540 37740 11552
rect 37056 11512 37740 11540
rect 37056 11500 37062 11512
rect 37734 11500 37740 11512
rect 37792 11500 37798 11552
rect 41141 11543 41199 11549
rect 41141 11509 41153 11543
rect 41187 11540 41199 11543
rect 41432 11540 41460 11571
rect 41506 11568 41512 11580
rect 41564 11568 41570 11620
rect 43165 11611 43223 11617
rect 43165 11577 43177 11611
rect 43211 11577 43223 11611
rect 43165 11571 43223 11577
rect 42886 11540 42892 11552
rect 41187 11512 41460 11540
rect 42799 11512 42892 11540
rect 41187 11509 41199 11512
rect 41141 11503 41199 11509
rect 42886 11500 42892 11512
rect 42944 11540 42950 11552
rect 43180 11540 43208 11571
rect 43530 11540 43536 11552
rect 42944 11512 43536 11540
rect 42944 11500 42950 11512
rect 43530 11500 43536 11512
rect 43588 11540 43594 11552
rect 44085 11543 44143 11549
rect 44085 11540 44097 11543
rect 43588 11512 44097 11540
rect 43588 11500 43594 11512
rect 44085 11509 44097 11512
rect 44131 11540 44143 11543
rect 44174 11540 44180 11552
rect 44131 11512 44180 11540
rect 44131 11509 44143 11512
rect 44085 11503 44143 11509
rect 44174 11500 44180 11512
rect 44232 11500 44238 11552
rect 1104 11450 48852 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 48852 11450
rect 1104 11376 48852 11398
rect 10042 11336 10048 11348
rect 9955 11308 10048 11336
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 9968 11209 9996 11308
rect 10042 11296 10048 11308
rect 10100 11336 10106 11348
rect 13814 11336 13820 11348
rect 10100 11308 13820 11336
rect 10100 11296 10106 11308
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 13998 11336 14004 11348
rect 13959 11308 14004 11336
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 19058 11336 19064 11348
rect 19019 11308 19064 11336
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 22830 11296 22836 11348
rect 22888 11336 22894 11348
rect 22925 11339 22983 11345
rect 22925 11336 22937 11339
rect 22888 11308 22937 11336
rect 22888 11296 22894 11308
rect 22925 11305 22937 11308
rect 22971 11305 22983 11339
rect 22925 11299 22983 11305
rect 24394 11296 24400 11348
rect 24452 11336 24458 11348
rect 24673 11339 24731 11345
rect 24673 11336 24685 11339
rect 24452 11308 24685 11336
rect 24452 11296 24458 11308
rect 24673 11305 24685 11308
rect 24719 11305 24731 11339
rect 24673 11299 24731 11305
rect 25593 11339 25651 11345
rect 25593 11305 25605 11339
rect 25639 11305 25651 11339
rect 25866 11336 25872 11348
rect 25827 11308 25872 11336
rect 25593 11299 25651 11305
rect 11422 11268 11428 11280
rect 11383 11240 11428 11268
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 12158 11228 12164 11280
rect 12216 11268 12222 11280
rect 12989 11271 13047 11277
rect 12989 11268 13001 11271
rect 12216 11240 13001 11268
rect 12216 11228 12222 11240
rect 12989 11237 13001 11240
rect 13035 11237 13047 11271
rect 12989 11231 13047 11237
rect 13081 11271 13139 11277
rect 13081 11237 13093 11271
rect 13127 11268 13139 11271
rect 13354 11268 13360 11280
rect 13127 11240 13360 11268
rect 13127 11237 13139 11240
rect 13081 11231 13139 11237
rect 13354 11228 13360 11240
rect 13412 11228 13418 11280
rect 13630 11268 13636 11280
rect 13591 11240 13636 11268
rect 13630 11228 13636 11240
rect 13688 11228 13694 11280
rect 17126 11268 17132 11280
rect 17087 11240 17132 11268
rect 17126 11228 17132 11240
rect 17184 11228 17190 11280
rect 19150 11228 19156 11280
rect 19208 11268 19214 11280
rect 23382 11268 23388 11280
rect 19208 11240 20944 11268
rect 23343 11240 23388 11268
rect 19208 11228 19214 11240
rect 9953 11203 10011 11209
rect 9953 11200 9965 11203
rect 9916 11172 9965 11200
rect 9916 11160 9922 11172
rect 9953 11169 9965 11172
rect 9999 11169 10011 11203
rect 10226 11200 10232 11212
rect 10187 11172 10232 11200
rect 9953 11163 10011 11169
rect 10226 11160 10232 11172
rect 10284 11160 10290 11212
rect 15654 11200 15660 11212
rect 15615 11172 15660 11200
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 15930 11200 15936 11212
rect 15891 11172 15936 11200
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 18782 11160 18788 11212
rect 18840 11200 18846 11212
rect 18969 11203 19027 11209
rect 18969 11200 18981 11203
rect 18840 11172 18981 11200
rect 18840 11160 18846 11172
rect 18969 11169 18981 11172
rect 19015 11169 19027 11203
rect 19426 11200 19432 11212
rect 19387 11172 19432 11200
rect 18969 11163 19027 11169
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 20916 11209 20944 11240
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 23477 11271 23535 11277
rect 23477 11237 23489 11271
rect 23523 11268 23535 11271
rect 23566 11268 23572 11280
rect 23523 11240 23572 11268
rect 23523 11237 23535 11240
rect 23477 11231 23535 11237
rect 23566 11228 23572 11240
rect 23624 11228 23630 11280
rect 25608 11268 25636 11299
rect 25866 11296 25872 11308
rect 25924 11296 25930 11348
rect 26329 11339 26387 11345
rect 26329 11305 26341 11339
rect 26375 11336 26387 11339
rect 26970 11336 26976 11348
rect 26375 11308 26976 11336
rect 26375 11305 26387 11308
rect 26329 11299 26387 11305
rect 26344 11268 26372 11299
rect 26970 11296 26976 11308
rect 27028 11296 27034 11348
rect 28626 11296 28632 11348
rect 28684 11336 28690 11348
rect 29181 11339 29239 11345
rect 29181 11336 29193 11339
rect 28684 11308 29193 11336
rect 28684 11296 28690 11308
rect 29181 11305 29193 11308
rect 29227 11305 29239 11339
rect 29181 11299 29239 11305
rect 29270 11296 29276 11348
rect 29328 11336 29334 11348
rect 29549 11339 29607 11345
rect 29549 11336 29561 11339
rect 29328 11308 29561 11336
rect 29328 11296 29334 11308
rect 29549 11305 29561 11308
rect 29595 11305 29607 11339
rect 29549 11299 29607 11305
rect 30742 11296 30748 11348
rect 30800 11336 30806 11348
rect 30837 11339 30895 11345
rect 30837 11336 30849 11339
rect 30800 11308 30849 11336
rect 30800 11296 30806 11308
rect 30837 11305 30849 11308
rect 30883 11336 30895 11339
rect 32766 11336 32772 11348
rect 30883 11308 32772 11336
rect 30883 11305 30895 11308
rect 30837 11299 30895 11305
rect 32766 11296 32772 11308
rect 32824 11296 32830 11348
rect 34422 11296 34428 11348
rect 34480 11336 34486 11348
rect 34609 11339 34667 11345
rect 34609 11336 34621 11339
rect 34480 11308 34621 11336
rect 34480 11296 34486 11308
rect 34609 11305 34621 11308
rect 34655 11305 34667 11339
rect 35250 11336 35256 11348
rect 35211 11308 35256 11336
rect 34609 11299 34667 11305
rect 35250 11296 35256 11308
rect 35308 11296 35314 11348
rect 36998 11296 37004 11348
rect 37056 11336 37062 11348
rect 37093 11339 37151 11345
rect 37093 11336 37105 11339
rect 37056 11308 37105 11336
rect 37056 11296 37062 11308
rect 37093 11305 37105 11308
rect 37139 11305 37151 11339
rect 37458 11336 37464 11348
rect 37419 11308 37464 11336
rect 37093 11299 37151 11305
rect 37458 11296 37464 11308
rect 37516 11296 37522 11348
rect 37734 11296 37740 11348
rect 37792 11336 37798 11348
rect 38933 11339 38991 11345
rect 37792 11308 37964 11336
rect 37792 11296 37798 11308
rect 25608 11240 26372 11268
rect 26694 11228 26700 11280
rect 26752 11268 26758 11280
rect 26834 11271 26892 11277
rect 26834 11268 26846 11271
rect 26752 11240 26846 11268
rect 26752 11228 26758 11240
rect 26834 11237 26846 11240
rect 26880 11237 26892 11271
rect 29914 11268 29920 11280
rect 29875 11240 29920 11268
rect 26834 11231 26892 11237
rect 29914 11228 29920 11240
rect 29972 11228 29978 11280
rect 32030 11228 32036 11280
rect 32088 11268 32094 11280
rect 32309 11271 32367 11277
rect 32309 11268 32321 11271
rect 32088 11240 32321 11268
rect 32088 11228 32094 11240
rect 32309 11237 32321 11240
rect 32355 11237 32367 11271
rect 32309 11231 32367 11237
rect 33594 11228 33600 11280
rect 33652 11268 33658 11280
rect 34010 11271 34068 11277
rect 34010 11268 34022 11271
rect 33652 11240 34022 11268
rect 33652 11228 33658 11240
rect 34010 11237 34022 11240
rect 34056 11268 34068 11271
rect 35066 11268 35072 11280
rect 34056 11240 35072 11268
rect 34056 11237 34068 11240
rect 34010 11231 34068 11237
rect 35066 11228 35072 11240
rect 35124 11228 35130 11280
rect 36170 11228 36176 11280
rect 36228 11268 36234 11280
rect 36265 11271 36323 11277
rect 36265 11268 36277 11271
rect 36228 11240 36277 11268
rect 36228 11228 36234 11240
rect 36265 11237 36277 11240
rect 36311 11237 36323 11271
rect 36265 11231 36323 11237
rect 36906 11228 36912 11280
rect 36964 11268 36970 11280
rect 37826 11268 37832 11280
rect 36964 11240 37832 11268
rect 36964 11228 36970 11240
rect 37826 11228 37832 11240
rect 37884 11228 37890 11280
rect 37936 11277 37964 11308
rect 38933 11305 38945 11339
rect 38979 11336 38991 11339
rect 39114 11336 39120 11348
rect 38979 11308 39120 11336
rect 38979 11305 38991 11308
rect 38933 11299 38991 11305
rect 39114 11296 39120 11308
rect 39172 11296 39178 11348
rect 43070 11336 43076 11348
rect 43031 11308 43076 11336
rect 43070 11296 43076 11308
rect 43128 11296 43134 11348
rect 37921 11271 37979 11277
rect 37921 11237 37933 11271
rect 37967 11237 37979 11271
rect 39132 11268 39160 11296
rect 41414 11268 41420 11280
rect 39132 11240 39804 11268
rect 41375 11240 41420 11268
rect 37921 11231 37979 11237
rect 20901 11203 20959 11209
rect 20901 11169 20913 11203
rect 20947 11200 20959 11203
rect 21450 11200 21456 11212
rect 20947 11172 21456 11200
rect 20947 11169 20959 11172
rect 20901 11163 20959 11169
rect 21450 11160 21456 11172
rect 21508 11160 21514 11212
rect 22097 11203 22155 11209
rect 22097 11169 22109 11203
rect 22143 11200 22155 11203
rect 22922 11200 22928 11212
rect 22143 11172 22928 11200
rect 22143 11169 22155 11172
rect 22097 11163 22155 11169
rect 22922 11160 22928 11172
rect 22980 11160 22986 11212
rect 25409 11203 25467 11209
rect 25409 11169 25421 11203
rect 25455 11200 25467 11203
rect 27154 11200 27160 11212
rect 25455 11172 27160 11200
rect 25455 11169 25467 11172
rect 25409 11163 25467 11169
rect 27154 11160 27160 11172
rect 27212 11160 27218 11212
rect 28629 11203 28687 11209
rect 28629 11169 28641 11203
rect 28675 11200 28687 11203
rect 28718 11200 28724 11212
rect 28675 11172 28724 11200
rect 28675 11169 28687 11172
rect 28629 11163 28687 11169
rect 28718 11160 28724 11172
rect 28776 11160 28782 11212
rect 33502 11160 33508 11212
rect 33560 11200 33566 11212
rect 33689 11203 33747 11209
rect 33689 11200 33701 11203
rect 33560 11172 33701 11200
rect 33560 11160 33566 11172
rect 33689 11169 33701 11172
rect 33735 11169 33747 11203
rect 39298 11200 39304 11212
rect 39259 11172 39304 11200
rect 33689 11163 33747 11169
rect 39298 11160 39304 11172
rect 39356 11160 39362 11212
rect 39776 11209 39804 11240
rect 41414 11228 41420 11240
rect 41472 11228 41478 11280
rect 43533 11271 43591 11277
rect 43533 11237 43545 11271
rect 43579 11268 43591 11271
rect 44174 11268 44180 11280
rect 43579 11240 44180 11268
rect 43579 11237 43591 11240
rect 43533 11231 43591 11237
rect 44174 11228 44180 11240
rect 44232 11228 44238 11280
rect 39761 11203 39819 11209
rect 39761 11169 39773 11203
rect 39807 11169 39819 11203
rect 39761 11163 39819 11169
rect 10318 11092 10324 11144
rect 10376 11132 10382 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 10376 11104 10425 11132
rect 10376 11092 10382 11104
rect 10413 11101 10425 11104
rect 10459 11132 10471 11135
rect 10689 11135 10747 11141
rect 10689 11132 10701 11135
rect 10459 11104 10701 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 10689 11101 10701 11104
rect 10735 11101 10747 11135
rect 11330 11132 11336 11144
rect 11291 11104 11336 11132
rect 10689 11095 10747 11101
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 15672 11132 15700 11160
rect 16114 11132 16120 11144
rect 11440 11104 15700 11132
rect 16075 11104 16120 11132
rect 10134 11024 10140 11076
rect 10192 11064 10198 11076
rect 11440 11064 11468 11104
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 17037 11135 17095 11141
rect 17037 11132 17049 11135
rect 16724 11104 17049 11132
rect 16724 11092 16730 11104
rect 17037 11101 17049 11104
rect 17083 11101 17095 11135
rect 17678 11132 17684 11144
rect 17639 11104 17684 11132
rect 17037 11095 17095 11101
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 22278 11132 22284 11144
rect 22239 11104 22284 11132
rect 22278 11092 22284 11104
rect 22336 11092 22342 11144
rect 23474 11092 23480 11144
rect 23532 11132 23538 11144
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 23532 11104 23673 11132
rect 23532 11092 23538 11104
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 26510 11132 26516 11144
rect 26471 11104 26516 11132
rect 23661 11095 23719 11101
rect 26510 11092 26516 11104
rect 26568 11092 26574 11144
rect 29822 11132 29828 11144
rect 29783 11104 29828 11132
rect 29822 11092 29828 11104
rect 29880 11092 29886 11144
rect 30101 11135 30159 11141
rect 30101 11101 30113 11135
rect 30147 11101 30159 11135
rect 30101 11095 30159 11101
rect 10192 11036 11468 11064
rect 11885 11067 11943 11073
rect 10192 11024 10198 11036
rect 11885 11033 11897 11067
rect 11931 11064 11943 11067
rect 12250 11064 12256 11076
rect 11931 11036 12256 11064
rect 11931 11033 11943 11036
rect 11885 11027 11943 11033
rect 12250 11024 12256 11036
rect 12308 11064 12314 11076
rect 13078 11064 13084 11076
rect 12308 11036 13084 11064
rect 12308 11024 12314 11036
rect 13078 11024 13084 11036
rect 13136 11024 13142 11076
rect 24118 11024 24124 11076
rect 24176 11064 24182 11076
rect 24397 11067 24455 11073
rect 24397 11064 24409 11067
rect 24176 11036 24409 11064
rect 24176 11024 24182 11036
rect 24397 11033 24409 11036
rect 24443 11064 24455 11067
rect 27433 11067 27491 11073
rect 27433 11064 27445 11067
rect 24443 11036 27445 11064
rect 24443 11033 24455 11036
rect 24397 11027 24455 11033
rect 27433 11033 27445 11036
rect 27479 11033 27491 11067
rect 27433 11027 27491 11033
rect 28718 11024 28724 11076
rect 28776 11064 28782 11076
rect 30116 11064 30144 11095
rect 31938 11092 31944 11144
rect 31996 11132 32002 11144
rect 32217 11135 32275 11141
rect 32217 11132 32229 11135
rect 31996 11104 32229 11132
rect 31996 11092 32002 11104
rect 32217 11101 32229 11104
rect 32263 11101 32275 11135
rect 32217 11095 32275 11101
rect 32306 11092 32312 11144
rect 32364 11132 32370 11144
rect 32493 11135 32551 11141
rect 32493 11132 32505 11135
rect 32364 11104 32505 11132
rect 32364 11092 32370 11104
rect 32493 11101 32505 11104
rect 32539 11101 32551 11135
rect 32493 11095 32551 11101
rect 36173 11135 36231 11141
rect 36173 11101 36185 11135
rect 36219 11132 36231 11135
rect 36906 11132 36912 11144
rect 36219 11104 36912 11132
rect 36219 11101 36231 11104
rect 36173 11095 36231 11101
rect 36906 11092 36912 11104
rect 36964 11132 36970 11144
rect 37182 11132 37188 11144
rect 36964 11104 37188 11132
rect 36964 11092 36970 11104
rect 37182 11092 37188 11104
rect 37240 11092 37246 11144
rect 38105 11135 38163 11141
rect 38105 11101 38117 11135
rect 38151 11101 38163 11135
rect 40034 11132 40040 11144
rect 39995 11104 40040 11132
rect 38105 11095 38163 11101
rect 31294 11064 31300 11076
rect 28776 11036 31300 11064
rect 28776 11024 28782 11036
rect 31294 11024 31300 11036
rect 31352 11024 31358 11076
rect 36722 11064 36728 11076
rect 36683 11036 36728 11064
rect 36722 11024 36728 11036
rect 36780 11024 36786 11076
rect 36814 11024 36820 11076
rect 36872 11064 36878 11076
rect 38120 11064 38148 11095
rect 40034 11092 40040 11104
rect 40092 11092 40098 11144
rect 41322 11132 41328 11144
rect 41235 11104 41328 11132
rect 41322 11092 41328 11104
rect 41380 11132 41386 11144
rect 43438 11132 43444 11144
rect 41380 11104 42794 11132
rect 43399 11104 43444 11132
rect 41380 11092 41386 11104
rect 41874 11064 41880 11076
rect 36872 11036 38148 11064
rect 41835 11036 41880 11064
rect 36872 11024 36878 11036
rect 41874 11024 41880 11036
rect 41932 11024 41938 11076
rect 42766 11064 42794 11104
rect 43438 11092 43444 11104
rect 43496 11092 43502 11144
rect 43714 11132 43720 11144
rect 43675 11104 43720 11132
rect 43714 11092 43720 11104
rect 43772 11092 43778 11144
rect 43732 11064 43760 11092
rect 42766 11036 43760 11064
rect 19978 10996 19984 11008
rect 19939 10968 19984 10996
rect 19978 10956 19984 10968
rect 20036 10996 20042 11008
rect 21085 10999 21143 11005
rect 21085 10996 21097 10999
rect 20036 10968 21097 10996
rect 20036 10956 20042 10968
rect 21085 10965 21097 10968
rect 21131 10965 21143 10999
rect 25130 10996 25136 11008
rect 25091 10968 25136 10996
rect 21085 10959 21143 10965
rect 25130 10956 25136 10968
rect 25188 10956 25194 11008
rect 26326 10956 26332 11008
rect 26384 10996 26390 11008
rect 28859 10999 28917 11005
rect 28859 10996 28871 10999
rect 26384 10968 28871 10996
rect 26384 10956 26390 10968
rect 28859 10965 28871 10968
rect 28905 10965 28917 10999
rect 33226 10996 33232 11008
rect 33187 10968 33232 10996
rect 28859 10959 28917 10965
rect 33226 10956 33232 10968
rect 33284 10956 33290 11008
rect 38654 10956 38660 11008
rect 38712 10996 38718 11008
rect 39022 10996 39028 11008
rect 38712 10968 39028 10996
rect 38712 10956 38718 10968
rect 39022 10956 39028 10968
rect 39080 10956 39086 11008
rect 1104 10906 48852 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 48852 10906
rect 1104 10832 48852 10854
rect 9858 10792 9864 10804
rect 9819 10764 9864 10792
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 11241 10795 11299 10801
rect 11241 10761 11253 10795
rect 11287 10792 11299 10795
rect 11422 10792 11428 10804
rect 11287 10764 11428 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 12158 10792 12164 10804
rect 12119 10764 12164 10792
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12989 10795 13047 10801
rect 12989 10761 13001 10795
rect 13035 10792 13047 10795
rect 13354 10792 13360 10804
rect 13035 10764 13360 10792
rect 13035 10761 13047 10764
rect 12989 10755 13047 10761
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 14737 10795 14795 10801
rect 14737 10761 14749 10795
rect 14783 10792 14795 10795
rect 15010 10792 15016 10804
rect 14783 10764 15016 10792
rect 14783 10761 14795 10764
rect 14737 10755 14795 10761
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 15335 10795 15393 10801
rect 15335 10761 15347 10795
rect 15381 10792 15393 10795
rect 16666 10792 16672 10804
rect 15381 10764 16672 10792
rect 15381 10761 15393 10764
rect 15335 10755 15393 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 17126 10792 17132 10804
rect 17087 10764 17132 10792
rect 17126 10752 17132 10764
rect 17184 10792 17190 10804
rect 17405 10795 17463 10801
rect 17405 10792 17417 10795
rect 17184 10764 17417 10792
rect 17184 10752 17190 10764
rect 17405 10761 17417 10764
rect 17451 10761 17463 10795
rect 17405 10755 17463 10761
rect 17494 10752 17500 10804
rect 17552 10792 17558 10804
rect 18187 10795 18245 10801
rect 18187 10792 18199 10795
rect 17552 10764 18199 10792
rect 17552 10752 17558 10764
rect 18187 10761 18199 10764
rect 18233 10761 18245 10795
rect 18187 10755 18245 10761
rect 18782 10752 18788 10804
rect 18840 10792 18846 10804
rect 18969 10795 19027 10801
rect 18969 10792 18981 10795
rect 18840 10764 18981 10792
rect 18840 10752 18846 10764
rect 18969 10761 18981 10764
rect 19015 10761 19027 10795
rect 21450 10792 21456 10804
rect 21411 10764 21456 10792
rect 18969 10755 19027 10761
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 25222 10752 25228 10804
rect 25280 10792 25286 10804
rect 25961 10795 26019 10801
rect 25961 10792 25973 10795
rect 25280 10764 25973 10792
rect 25280 10752 25286 10764
rect 25961 10761 25973 10764
rect 26007 10761 26019 10795
rect 25961 10755 26019 10761
rect 26510 10752 26516 10804
rect 26568 10792 26574 10804
rect 27614 10792 27620 10804
rect 26568 10764 27620 10792
rect 26568 10752 26574 10764
rect 27614 10752 27620 10764
rect 27672 10792 27678 10804
rect 28169 10795 28227 10801
rect 28169 10792 28181 10795
rect 27672 10764 28181 10792
rect 27672 10752 27678 10764
rect 28169 10761 28181 10764
rect 28215 10761 28227 10795
rect 28718 10792 28724 10804
rect 28679 10764 28724 10792
rect 28169 10755 28227 10761
rect 28718 10752 28724 10764
rect 28776 10752 28782 10804
rect 29549 10795 29607 10801
rect 29549 10761 29561 10795
rect 29595 10792 29607 10795
rect 29822 10792 29828 10804
rect 29595 10764 29828 10792
rect 29595 10761 29607 10764
rect 29549 10755 29607 10761
rect 29822 10752 29828 10764
rect 29880 10752 29886 10804
rect 29914 10752 29920 10804
rect 29972 10792 29978 10804
rect 30469 10795 30527 10801
rect 30469 10792 30481 10795
rect 29972 10764 30481 10792
rect 29972 10752 29978 10764
rect 30469 10761 30481 10764
rect 30515 10761 30527 10795
rect 30469 10755 30527 10761
rect 31757 10795 31815 10801
rect 31757 10761 31769 10795
rect 31803 10792 31815 10795
rect 32030 10792 32036 10804
rect 31803 10764 32036 10792
rect 31803 10761 31815 10764
rect 31757 10755 31815 10761
rect 32030 10752 32036 10764
rect 32088 10752 32094 10804
rect 33321 10795 33379 10801
rect 33321 10761 33333 10795
rect 33367 10792 33379 10795
rect 33502 10792 33508 10804
rect 33367 10764 33508 10792
rect 33367 10761 33379 10764
rect 33321 10755 33379 10761
rect 33502 10752 33508 10764
rect 33560 10752 33566 10804
rect 33778 10752 33784 10804
rect 33836 10792 33842 10804
rect 33919 10795 33977 10801
rect 33919 10792 33931 10795
rect 33836 10764 33931 10792
rect 33836 10752 33842 10764
rect 33919 10761 33931 10764
rect 33965 10761 33977 10795
rect 34330 10792 34336 10804
rect 34291 10764 34336 10792
rect 33919 10755 33977 10761
rect 34330 10752 34336 10764
rect 34388 10752 34394 10804
rect 36170 10792 36176 10804
rect 36131 10764 36176 10792
rect 36170 10752 36176 10764
rect 36228 10752 36234 10804
rect 37734 10792 37740 10804
rect 37695 10764 37740 10792
rect 37734 10752 37740 10764
rect 37792 10752 37798 10804
rect 37826 10752 37832 10804
rect 37884 10792 37890 10804
rect 38105 10795 38163 10801
rect 38105 10792 38117 10795
rect 37884 10764 38117 10792
rect 37884 10752 37890 10764
rect 38105 10761 38117 10764
rect 38151 10761 38163 10795
rect 38654 10792 38660 10804
rect 38615 10764 38660 10792
rect 38105 10755 38163 10761
rect 38654 10752 38660 10764
rect 38712 10752 38718 10804
rect 39298 10752 39304 10804
rect 39356 10792 39362 10804
rect 39853 10795 39911 10801
rect 39853 10792 39865 10795
rect 39356 10764 39865 10792
rect 39356 10752 39362 10764
rect 39853 10761 39865 10764
rect 39899 10761 39911 10795
rect 39853 10755 39911 10761
rect 41325 10795 41383 10801
rect 41325 10761 41337 10795
rect 41371 10792 41383 10795
rect 41414 10792 41420 10804
rect 41371 10764 41420 10792
rect 41371 10761 41383 10764
rect 41325 10755 41383 10761
rect 41414 10752 41420 10764
rect 41472 10752 41478 10804
rect 42886 10792 42892 10804
rect 42847 10764 42892 10792
rect 42886 10752 42892 10764
rect 42944 10752 42950 10804
rect 43438 10792 43444 10804
rect 43399 10764 43444 10792
rect 43438 10752 43444 10764
rect 43496 10792 43502 10804
rect 44174 10792 44180 10804
rect 43496 10764 43760 10792
rect 44135 10764 44180 10792
rect 43496 10752 43502 10764
rect 15105 10727 15163 10733
rect 15105 10693 15117 10727
rect 15151 10724 15163 10727
rect 15930 10724 15936 10736
rect 15151 10696 15936 10724
rect 15151 10693 15163 10696
rect 15105 10687 15163 10693
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 16684 10724 16712 10752
rect 17773 10727 17831 10733
rect 17773 10724 17785 10727
rect 16684 10696 17785 10724
rect 17773 10693 17785 10696
rect 17819 10693 17831 10727
rect 18800 10724 18828 10752
rect 17773 10687 17831 10693
rect 17880 10696 18828 10724
rect 22649 10727 22707 10733
rect 10318 10656 10324 10668
rect 10279 10628 10324 10656
rect 10318 10616 10324 10628
rect 10376 10616 10382 10668
rect 13170 10656 13176 10668
rect 13131 10628 13176 10656
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 16114 10616 16120 10668
rect 16172 10656 16178 10668
rect 16209 10659 16267 10665
rect 16209 10656 16221 10659
rect 16172 10628 16221 10656
rect 16172 10616 16178 10628
rect 16209 10625 16221 10628
rect 16255 10625 16267 10659
rect 16209 10619 16267 10625
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 11330 10588 11336 10600
rect 9355 10560 11336 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 11330 10548 11336 10560
rect 11388 10588 11394 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 11388 10560 11529 10588
rect 11388 10548 11394 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 13262 10588 13268 10600
rect 13223 10560 13268 10588
rect 11517 10551 11575 10557
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 15010 10548 15016 10600
rect 15068 10588 15074 10600
rect 15232 10591 15290 10597
rect 15232 10588 15244 10591
rect 15068 10560 15244 10588
rect 15068 10548 15074 10560
rect 15232 10557 15244 10560
rect 15278 10557 15290 10591
rect 15232 10551 15290 10557
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 15749 10591 15807 10597
rect 15749 10588 15761 10591
rect 15712 10560 15761 10588
rect 15712 10548 15718 10560
rect 15749 10557 15761 10560
rect 15795 10588 15807 10591
rect 17880 10588 17908 10696
rect 22649 10693 22661 10727
rect 22695 10724 22707 10727
rect 23382 10724 23388 10736
rect 22695 10696 23388 10724
rect 22695 10693 22707 10696
rect 22649 10687 22707 10693
rect 23382 10684 23388 10696
rect 23440 10724 23446 10736
rect 24489 10727 24547 10733
rect 24489 10724 24501 10727
rect 23440 10696 24501 10724
rect 23440 10684 23446 10696
rect 24489 10693 24501 10696
rect 24535 10693 24547 10727
rect 31294 10724 31300 10736
rect 31255 10696 31300 10724
rect 24489 10687 24547 10693
rect 31294 10684 31300 10696
rect 31352 10684 31358 10736
rect 33686 10684 33692 10736
rect 33744 10724 33750 10736
rect 36722 10724 36728 10736
rect 33744 10696 36728 10724
rect 33744 10684 33750 10696
rect 18230 10616 18236 10668
rect 18288 10656 18294 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18288 10628 18613 10656
rect 18288 10616 18294 10628
rect 18601 10625 18613 10628
rect 18647 10656 18659 10659
rect 21913 10659 21971 10665
rect 18647 10628 19380 10656
rect 18647 10625 18659 10628
rect 18601 10619 18659 10625
rect 15795 10560 17908 10588
rect 17957 10591 18015 10597
rect 15795 10557 15807 10560
rect 15749 10551 15807 10557
rect 17957 10557 17969 10591
rect 18003 10588 18015 10591
rect 18046 10588 18052 10600
rect 18003 10560 18052 10588
rect 18003 10557 18015 10560
rect 17957 10551 18015 10557
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 19352 10597 19380 10628
rect 21913 10625 21925 10659
rect 21959 10656 21971 10659
rect 22097 10659 22155 10665
rect 22097 10656 22109 10659
rect 21959 10628 22109 10656
rect 21959 10625 21971 10628
rect 21913 10619 21971 10625
rect 22097 10625 22109 10628
rect 22143 10656 22155 10659
rect 22278 10656 22284 10668
rect 22143 10628 22284 10656
rect 22143 10625 22155 10628
rect 22097 10619 22155 10625
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 24213 10659 24271 10665
rect 24213 10625 24225 10659
rect 24259 10656 24271 10659
rect 29779 10659 29837 10665
rect 24259 10628 27384 10656
rect 24259 10625 24271 10628
rect 24213 10619 24271 10625
rect 19337 10591 19395 10597
rect 19337 10557 19349 10591
rect 19383 10557 19395 10591
rect 19337 10551 19395 10557
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 19797 10591 19855 10597
rect 19797 10588 19809 10591
rect 19484 10560 19809 10588
rect 19484 10548 19490 10560
rect 19797 10557 19809 10560
rect 19843 10588 19855 10591
rect 19978 10588 19984 10600
rect 19843 10560 19984 10588
rect 19843 10557 19855 10560
rect 19797 10551 19855 10557
rect 19978 10548 19984 10560
rect 20036 10588 20042 10600
rect 20349 10591 20407 10597
rect 20349 10588 20361 10591
rect 20036 10560 20361 10588
rect 20036 10548 20042 10560
rect 20349 10557 20361 10560
rect 20395 10557 20407 10591
rect 20349 10551 20407 10557
rect 23385 10591 23443 10597
rect 23385 10557 23397 10591
rect 23431 10588 23443 10591
rect 23566 10588 23572 10600
rect 23431 10560 23572 10588
rect 23431 10557 23443 10560
rect 23385 10551 23443 10557
rect 23566 10548 23572 10560
rect 23624 10548 23630 10600
rect 23750 10597 23756 10600
rect 23728 10591 23756 10597
rect 23728 10588 23740 10591
rect 23663 10560 23740 10588
rect 23728 10557 23740 10560
rect 23808 10588 23814 10600
rect 24228 10588 24256 10619
rect 23808 10560 24256 10588
rect 25041 10591 25099 10597
rect 23728 10551 23756 10557
rect 23750 10548 23756 10551
rect 23808 10548 23814 10560
rect 25041 10557 25053 10591
rect 25087 10588 25099 10591
rect 25130 10588 25136 10600
rect 25087 10560 25136 10588
rect 25087 10557 25099 10560
rect 25041 10551 25099 10557
rect 25130 10548 25136 10560
rect 25188 10588 25194 10600
rect 26142 10588 26148 10600
rect 25188 10560 26148 10588
rect 25188 10548 25194 10560
rect 26142 10548 26148 10560
rect 26200 10548 26206 10600
rect 26878 10588 26884 10600
rect 26839 10560 26884 10588
rect 26878 10548 26884 10560
rect 26936 10548 26942 10600
rect 26970 10548 26976 10600
rect 27028 10588 27034 10600
rect 27246 10588 27252 10600
rect 27028 10560 27252 10588
rect 27028 10548 27034 10560
rect 27246 10548 27252 10560
rect 27304 10548 27310 10600
rect 27356 10588 27384 10628
rect 29779 10625 29791 10659
rect 29825 10656 29837 10659
rect 31938 10656 31944 10668
rect 29825 10628 31944 10656
rect 29825 10625 29837 10628
rect 29779 10619 29837 10625
rect 31938 10616 31944 10628
rect 31996 10616 32002 10668
rect 32766 10656 32772 10668
rect 32727 10628 32772 10656
rect 32766 10616 32772 10628
rect 32824 10616 32830 10668
rect 34790 10616 34796 10668
rect 34848 10656 34854 10668
rect 35268 10665 35296 10696
rect 36722 10684 36728 10696
rect 36780 10724 36786 10736
rect 36780 10696 37136 10724
rect 36780 10684 36786 10696
rect 34977 10659 35035 10665
rect 34977 10656 34989 10659
rect 34848 10628 34989 10656
rect 34848 10616 34854 10628
rect 34977 10625 34989 10628
rect 35023 10625 35035 10659
rect 34977 10619 35035 10625
rect 35253 10659 35311 10665
rect 35253 10625 35265 10659
rect 35299 10625 35311 10659
rect 36814 10656 36820 10668
rect 36775 10628 36820 10656
rect 35253 10619 35311 10625
rect 36814 10616 36820 10628
rect 36872 10616 36878 10668
rect 37108 10665 37136 10696
rect 39942 10684 39948 10736
rect 40000 10724 40006 10736
rect 41785 10727 41843 10733
rect 41785 10724 41797 10727
rect 40000 10696 41797 10724
rect 40000 10684 40006 10696
rect 41785 10693 41797 10696
rect 41831 10724 41843 10727
rect 41831 10696 42104 10724
rect 41831 10693 41843 10696
rect 41785 10687 41843 10693
rect 37093 10659 37151 10665
rect 37093 10625 37105 10659
rect 37139 10656 37151 10659
rect 38102 10656 38108 10668
rect 37139 10628 38108 10656
rect 37139 10625 37151 10628
rect 37093 10619 37151 10625
rect 38102 10616 38108 10628
rect 38160 10616 38166 10668
rect 40034 10616 40040 10668
rect 40092 10656 40098 10668
rect 41966 10656 41972 10668
rect 40092 10628 41972 10656
rect 40092 10616 40098 10628
rect 41966 10616 41972 10628
rect 42024 10616 42030 10668
rect 29692 10591 29750 10597
rect 29692 10588 29704 10591
rect 27356 10560 29704 10588
rect 29692 10557 29704 10560
rect 29738 10588 29750 10591
rect 30190 10588 30196 10600
rect 29738 10560 30196 10588
rect 29738 10557 29750 10560
rect 29692 10551 29750 10557
rect 30190 10548 30196 10560
rect 30248 10548 30254 10600
rect 33848 10591 33906 10597
rect 33848 10557 33860 10591
rect 33894 10588 33906 10591
rect 34330 10588 34336 10600
rect 33894 10560 34336 10588
rect 33894 10557 33906 10560
rect 33848 10551 33906 10557
rect 34330 10548 34336 10560
rect 34388 10548 34394 10600
rect 38654 10548 38660 10600
rect 38712 10588 38718 10600
rect 38841 10591 38899 10597
rect 38841 10588 38853 10591
rect 38712 10560 38853 10588
rect 38712 10548 38718 10560
rect 38841 10557 38853 10560
rect 38887 10557 38899 10591
rect 38841 10551 38899 10557
rect 39114 10548 39120 10600
rect 39172 10588 39178 10600
rect 39301 10591 39359 10597
rect 39301 10588 39313 10591
rect 39172 10560 39313 10588
rect 39172 10548 39178 10560
rect 39301 10557 39313 10560
rect 39347 10557 39359 10591
rect 39301 10551 39359 10557
rect 40313 10591 40371 10597
rect 40313 10557 40325 10591
rect 40359 10588 40371 10591
rect 40532 10591 40590 10597
rect 40532 10588 40544 10591
rect 40359 10560 40544 10588
rect 40359 10557 40371 10560
rect 40313 10551 40371 10557
rect 40532 10557 40544 10560
rect 40578 10588 40590 10591
rect 41874 10588 41880 10600
rect 40578 10560 41880 10588
rect 40578 10557 40590 10560
rect 40532 10551 40590 10557
rect 41874 10548 41880 10560
rect 41932 10548 41938 10600
rect 9217 10523 9275 10529
rect 9217 10489 9229 10523
rect 9263 10520 9275 10523
rect 10226 10520 10232 10532
rect 9263 10492 10232 10520
rect 9263 10489 9275 10492
rect 9217 10483 9275 10489
rect 10226 10480 10232 10492
rect 10284 10480 10290 10532
rect 10502 10480 10508 10532
rect 10560 10520 10566 10532
rect 10642 10523 10700 10529
rect 10642 10520 10654 10523
rect 10560 10492 10654 10520
rect 10560 10480 10566 10492
rect 10642 10489 10654 10492
rect 10688 10520 10700 10523
rect 13538 10520 13544 10532
rect 10688 10492 13544 10520
rect 10688 10489 10700 10492
rect 10642 10483 10700 10489
rect 13538 10480 13544 10492
rect 13596 10520 13602 10532
rect 16025 10523 16083 10529
rect 16025 10520 16037 10523
rect 13596 10492 16037 10520
rect 13596 10480 13602 10492
rect 16025 10489 16037 10492
rect 16071 10520 16083 10523
rect 16530 10523 16588 10529
rect 16530 10520 16542 10523
rect 16071 10492 16542 10520
rect 16071 10489 16083 10492
rect 16025 10483 16083 10489
rect 16530 10489 16542 10492
rect 16576 10520 16588 10523
rect 16666 10520 16672 10532
rect 16576 10492 16672 10520
rect 16576 10489 16588 10492
rect 16530 10483 16588 10489
rect 16666 10480 16672 10492
rect 16724 10480 16730 10532
rect 20070 10520 20076 10532
rect 20031 10492 20076 10520
rect 20070 10480 20076 10492
rect 20128 10480 20134 10532
rect 22189 10523 22247 10529
rect 22189 10489 22201 10523
rect 22235 10520 22247 10523
rect 22922 10520 22928 10532
rect 22235 10492 22928 10520
rect 22235 10489 22247 10492
rect 22189 10483 22247 10489
rect 22922 10480 22928 10492
rect 22980 10520 22986 10532
rect 23474 10520 23480 10532
rect 22980 10492 23480 10520
rect 22980 10480 22986 10492
rect 23474 10480 23480 10492
rect 23532 10480 23538 10532
rect 27264 10520 27292 10548
rect 27801 10523 27859 10529
rect 27801 10520 27813 10523
rect 27264 10492 27813 10520
rect 27801 10489 27813 10492
rect 27847 10489 27859 10523
rect 30742 10520 30748 10532
rect 30703 10492 30748 10520
rect 27801 10483 27859 10489
rect 30742 10480 30748 10492
rect 30800 10480 30806 10532
rect 30834 10480 30840 10532
rect 30892 10520 30898 10532
rect 32122 10520 32128 10532
rect 30892 10492 30937 10520
rect 32035 10492 32128 10520
rect 30892 10480 30898 10492
rect 32122 10480 32128 10492
rect 32180 10520 32186 10532
rect 32309 10523 32367 10529
rect 32309 10520 32321 10523
rect 32180 10492 32321 10520
rect 32180 10480 32186 10492
rect 32309 10489 32321 10492
rect 32355 10489 32367 10523
rect 32309 10483 32367 10489
rect 32401 10523 32459 10529
rect 32401 10489 32413 10523
rect 32447 10489 32459 10523
rect 32401 10483 32459 10489
rect 35069 10523 35127 10529
rect 35069 10489 35081 10523
rect 35115 10489 35127 10523
rect 35069 10483 35127 10489
rect 36909 10523 36967 10529
rect 36909 10489 36921 10523
rect 36955 10489 36967 10523
rect 39574 10520 39580 10532
rect 39535 10492 39580 10520
rect 36909 10483 36967 10489
rect 10137 10455 10195 10461
rect 10137 10421 10149 10455
rect 10183 10452 10195 10455
rect 10520 10452 10548 10480
rect 20990 10452 20996 10464
rect 10183 10424 10548 10452
rect 20951 10424 20996 10452
rect 10183 10421 10195 10424
rect 10137 10415 10195 10421
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 23382 10412 23388 10464
rect 23440 10452 23446 10464
rect 23799 10455 23857 10461
rect 23799 10452 23811 10455
rect 23440 10424 23811 10452
rect 23440 10412 23446 10424
rect 23799 10421 23811 10424
rect 23845 10421 23857 10455
rect 23799 10415 23857 10421
rect 24670 10412 24676 10464
rect 24728 10452 24734 10464
rect 24857 10455 24915 10461
rect 24857 10452 24869 10455
rect 24728 10424 24869 10452
rect 24728 10412 24734 10424
rect 24857 10421 24869 10424
rect 24903 10421 24915 10455
rect 25406 10452 25412 10464
rect 25367 10424 25412 10452
rect 24857 10415 24915 10421
rect 25406 10412 25412 10424
rect 25464 10452 25470 10464
rect 26513 10455 26571 10461
rect 26513 10452 26525 10455
rect 25464 10424 26525 10452
rect 25464 10412 25470 10424
rect 26513 10421 26525 10424
rect 26559 10452 26571 10455
rect 26694 10452 26700 10464
rect 26559 10424 26700 10452
rect 26559 10421 26571 10424
rect 26513 10415 26571 10421
rect 26694 10412 26700 10424
rect 26752 10412 26758 10464
rect 26878 10452 26884 10464
rect 26839 10424 26884 10452
rect 26878 10412 26884 10424
rect 26936 10412 26942 10464
rect 32030 10412 32036 10464
rect 32088 10452 32094 10464
rect 32416 10452 32444 10483
rect 32582 10452 32588 10464
rect 32088 10424 32588 10452
rect 32088 10412 32094 10424
rect 32582 10412 32588 10424
rect 32640 10412 32646 10464
rect 33134 10412 33140 10464
rect 33192 10452 33198 10464
rect 33594 10452 33600 10464
rect 33192 10424 33600 10452
rect 33192 10412 33198 10424
rect 33594 10412 33600 10424
rect 33652 10412 33658 10464
rect 34606 10452 34612 10464
rect 34567 10424 34612 10452
rect 34606 10412 34612 10424
rect 34664 10452 34670 10464
rect 35084 10452 35112 10483
rect 34664 10424 35112 10452
rect 36633 10455 36691 10461
rect 34664 10412 34670 10424
rect 36633 10421 36645 10455
rect 36679 10452 36691 10455
rect 36722 10452 36728 10464
rect 36679 10424 36728 10452
rect 36679 10421 36691 10424
rect 36633 10415 36691 10421
rect 36722 10412 36728 10424
rect 36780 10452 36786 10464
rect 36924 10452 36952 10483
rect 39574 10480 39580 10492
rect 39632 10480 39638 10532
rect 42076 10520 42104 10696
rect 43732 10665 43760 10764
rect 44174 10752 44180 10764
rect 44232 10752 44238 10804
rect 43717 10659 43775 10665
rect 43717 10625 43729 10659
rect 43763 10625 43775 10659
rect 43717 10619 43775 10625
rect 42290 10523 42348 10529
rect 42290 10520 42302 10523
rect 42076 10492 42302 10520
rect 42290 10489 42302 10492
rect 42336 10489 42348 10523
rect 42290 10483 42348 10489
rect 36780 10424 36952 10452
rect 36780 10412 36786 10424
rect 40494 10412 40500 10464
rect 40552 10452 40558 10464
rect 40635 10455 40693 10461
rect 40635 10452 40647 10455
rect 40552 10424 40647 10452
rect 40552 10412 40558 10424
rect 40635 10421 40647 10424
rect 40681 10421 40693 10455
rect 40635 10415 40693 10421
rect 1104 10362 48852 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 48852 10362
rect 1104 10288 48852 10310
rect 11333 10251 11391 10257
rect 11333 10217 11345 10251
rect 11379 10248 11391 10251
rect 11422 10248 11428 10260
rect 11379 10220 11428 10248
rect 11379 10217 11391 10220
rect 11333 10211 11391 10217
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 11790 10248 11796 10260
rect 11751 10220 11796 10248
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 13262 10248 13268 10260
rect 13223 10220 13268 10248
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13688 10220 13768 10248
rect 13688 10208 13694 10220
rect 13740 10189 13768 10220
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 15795 10251 15853 10257
rect 15795 10248 15807 10251
rect 15436 10220 15807 10248
rect 15436 10208 15442 10220
rect 15795 10217 15807 10220
rect 15841 10217 15853 10251
rect 15795 10211 15853 10217
rect 16114 10208 16120 10260
rect 16172 10248 16178 10260
rect 16209 10251 16267 10257
rect 16209 10248 16221 10251
rect 16172 10220 16221 10248
rect 16172 10208 16178 10220
rect 16209 10217 16221 10220
rect 16255 10217 16267 10251
rect 18046 10248 18052 10260
rect 18007 10220 18052 10248
rect 16209 10211 16267 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18969 10251 19027 10257
rect 18969 10217 18981 10251
rect 19015 10248 19027 10251
rect 19058 10248 19064 10260
rect 19015 10220 19064 10248
rect 19015 10217 19027 10220
rect 18969 10211 19027 10217
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 23566 10208 23572 10260
rect 23624 10248 23630 10260
rect 23937 10251 23995 10257
rect 23937 10248 23949 10251
rect 23624 10220 23949 10248
rect 23624 10208 23630 10220
rect 23937 10217 23949 10220
rect 23983 10217 23995 10251
rect 23937 10211 23995 10217
rect 25869 10251 25927 10257
rect 25869 10217 25881 10251
rect 25915 10248 25927 10251
rect 27154 10248 27160 10260
rect 25915 10220 27160 10248
rect 25915 10217 25927 10220
rect 25869 10211 25927 10217
rect 27154 10208 27160 10220
rect 27212 10208 27218 10260
rect 27246 10208 27252 10260
rect 27304 10248 27310 10260
rect 27433 10251 27491 10257
rect 27433 10248 27445 10251
rect 27304 10220 27445 10248
rect 27304 10208 27310 10220
rect 27433 10217 27445 10220
rect 27479 10217 27491 10251
rect 27433 10211 27491 10217
rect 28902 10208 28908 10260
rect 28960 10248 28966 10260
rect 29273 10251 29331 10257
rect 29273 10248 29285 10251
rect 28960 10220 29285 10248
rect 28960 10208 28966 10220
rect 29273 10217 29285 10220
rect 29319 10248 29331 10251
rect 30469 10251 30527 10257
rect 29319 10220 29913 10248
rect 29319 10217 29331 10220
rect 29273 10211 29331 10217
rect 12897 10183 12955 10189
rect 10612 10152 12204 10180
rect 10134 10112 10140 10124
rect 10095 10084 10140 10112
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10612 10121 10640 10152
rect 12176 10124 12204 10152
rect 12897 10149 12909 10183
rect 12943 10180 12955 10183
rect 13725 10183 13783 10189
rect 13725 10180 13737 10183
rect 12943 10152 13737 10180
rect 12943 10149 12955 10152
rect 12897 10143 12955 10149
rect 13725 10149 13737 10152
rect 13771 10149 13783 10183
rect 13725 10143 13783 10149
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 13872 10152 13917 10180
rect 13872 10140 13878 10152
rect 16666 10140 16672 10192
rect 16724 10180 16730 10192
rect 16990 10183 17048 10189
rect 16990 10180 17002 10183
rect 16724 10152 17002 10180
rect 16724 10140 16730 10152
rect 16990 10149 17002 10152
rect 17036 10149 17048 10183
rect 16990 10143 17048 10149
rect 10597 10115 10655 10121
rect 10597 10112 10609 10115
rect 10284 10084 10609 10112
rect 10284 10072 10290 10084
rect 10597 10081 10609 10084
rect 10643 10081 10655 10115
rect 11698 10112 11704 10124
rect 11659 10084 11704 10112
rect 10597 10075 10655 10081
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 12158 10112 12164 10124
rect 12119 10084 12164 10112
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 19076 10121 19104 10208
rect 19150 10140 19156 10192
rect 19208 10180 19214 10192
rect 19334 10180 19340 10192
rect 19208 10152 19340 10180
rect 19208 10140 19214 10152
rect 19334 10140 19340 10152
rect 19392 10189 19398 10192
rect 19392 10183 19440 10189
rect 19392 10149 19394 10183
rect 19428 10180 19440 10183
rect 19978 10180 19984 10192
rect 19428 10152 19984 10180
rect 19428 10149 19440 10152
rect 19392 10143 19440 10149
rect 19392 10140 19398 10143
rect 19978 10140 19984 10152
rect 20036 10180 20042 10192
rect 21222 10183 21280 10189
rect 21222 10180 21234 10183
rect 20036 10152 21234 10180
rect 20036 10140 20042 10152
rect 21222 10149 21234 10152
rect 21268 10180 21280 10183
rect 22922 10180 22928 10192
rect 21268 10152 22928 10180
rect 21268 10149 21280 10152
rect 21222 10143 21280 10149
rect 22922 10140 22928 10152
rect 22980 10180 22986 10192
rect 23338 10183 23396 10189
rect 23338 10180 23350 10183
rect 22980 10152 23350 10180
rect 22980 10140 22986 10152
rect 23338 10149 23350 10152
rect 23384 10180 23396 10183
rect 24670 10180 24676 10192
rect 23384 10152 24676 10180
rect 23384 10149 23396 10152
rect 23338 10143 23396 10149
rect 24670 10140 24676 10152
rect 24728 10140 24734 10192
rect 24946 10180 24952 10192
rect 24907 10152 24952 10180
rect 24946 10140 24952 10152
rect 25004 10140 25010 10192
rect 25498 10180 25504 10192
rect 25459 10152 25504 10180
rect 25498 10140 25504 10152
rect 25556 10140 25562 10192
rect 26786 10180 26792 10192
rect 26747 10152 26792 10180
rect 26786 10140 26792 10152
rect 26844 10140 26850 10192
rect 29885 10189 29913 10220
rect 30469 10217 30481 10251
rect 30515 10248 30527 10251
rect 30834 10248 30840 10260
rect 30515 10220 30840 10248
rect 30515 10217 30527 10220
rect 30469 10211 30527 10217
rect 30834 10208 30840 10220
rect 30892 10208 30898 10260
rect 32122 10248 32128 10260
rect 32083 10220 32128 10248
rect 32122 10208 32128 10220
rect 32180 10208 32186 10260
rect 32582 10248 32588 10260
rect 32543 10220 32588 10248
rect 32582 10208 32588 10220
rect 32640 10208 32646 10260
rect 34425 10251 34483 10257
rect 34425 10217 34437 10251
rect 34471 10248 34483 10251
rect 34606 10248 34612 10260
rect 34471 10220 34612 10248
rect 34471 10217 34483 10220
rect 34425 10211 34483 10217
rect 34606 10208 34612 10220
rect 34664 10208 34670 10260
rect 34790 10208 34796 10260
rect 34848 10248 34854 10260
rect 34885 10251 34943 10257
rect 34885 10248 34897 10251
rect 34848 10220 34897 10248
rect 34848 10208 34854 10220
rect 34885 10217 34897 10220
rect 34931 10217 34943 10251
rect 36078 10248 36084 10260
rect 36039 10220 36084 10248
rect 34885 10211 34943 10217
rect 36078 10208 36084 10220
rect 36136 10208 36142 10260
rect 36633 10251 36691 10257
rect 36633 10217 36645 10251
rect 36679 10248 36691 10251
rect 37734 10248 37740 10260
rect 36679 10220 37740 10248
rect 36679 10217 36691 10220
rect 36633 10211 36691 10217
rect 37734 10208 37740 10220
rect 37792 10248 37798 10260
rect 38933 10251 38991 10257
rect 37792 10220 37964 10248
rect 37792 10208 37798 10220
rect 29870 10183 29928 10189
rect 29870 10149 29882 10183
rect 29916 10149 29928 10183
rect 29870 10143 29928 10149
rect 31938 10140 31944 10192
rect 31996 10180 32002 10192
rect 32953 10183 33011 10189
rect 32953 10180 32965 10183
rect 31996 10152 32965 10180
rect 31996 10140 32002 10152
rect 32953 10149 32965 10152
rect 32999 10149 33011 10183
rect 32953 10143 33011 10149
rect 33134 10140 33140 10192
rect 33192 10180 33198 10192
rect 33826 10183 33884 10189
rect 33826 10180 33838 10183
rect 33192 10152 33838 10180
rect 33192 10140 33198 10152
rect 33826 10149 33838 10152
rect 33872 10149 33884 10183
rect 36906 10180 36912 10192
rect 36867 10152 36912 10180
rect 33826 10143 33884 10149
rect 36906 10140 36912 10152
rect 36964 10140 36970 10192
rect 37936 10189 37964 10220
rect 38933 10217 38945 10251
rect 38979 10248 38991 10251
rect 39114 10248 39120 10260
rect 38979 10220 39120 10248
rect 38979 10217 38991 10220
rect 38933 10211 38991 10217
rect 39114 10208 39120 10220
rect 39172 10248 39178 10260
rect 39301 10251 39359 10257
rect 39301 10248 39313 10251
rect 39172 10220 39313 10248
rect 39172 10208 39178 10220
rect 39301 10217 39313 10220
rect 39347 10217 39359 10251
rect 39301 10211 39359 10217
rect 41049 10251 41107 10257
rect 41049 10217 41061 10251
rect 41095 10248 41107 10251
rect 41414 10248 41420 10260
rect 41095 10220 41420 10248
rect 41095 10217 41107 10220
rect 41049 10211 41107 10217
rect 41414 10208 41420 10220
rect 41472 10208 41478 10260
rect 41966 10248 41972 10260
rect 41927 10220 41972 10248
rect 41966 10208 41972 10220
rect 42024 10208 42030 10260
rect 37921 10183 37979 10189
rect 37921 10149 37933 10183
rect 37967 10149 37979 10183
rect 37921 10143 37979 10149
rect 39942 10140 39948 10192
rect 40000 10180 40006 10192
rect 40450 10183 40508 10189
rect 40450 10180 40462 10183
rect 40000 10152 40462 10180
rect 40000 10140 40006 10152
rect 40450 10149 40462 10152
rect 40496 10149 40508 10183
rect 41322 10180 41328 10192
rect 41283 10152 41328 10180
rect 40450 10143 40508 10149
rect 41322 10140 41328 10152
rect 41380 10140 41386 10192
rect 15724 10115 15782 10121
rect 15724 10081 15736 10115
rect 15770 10081 15782 10115
rect 15724 10075 15782 10081
rect 19061 10115 19119 10121
rect 19061 10081 19073 10115
rect 19107 10081 19119 10115
rect 19061 10075 19119 10081
rect 26973 10115 27031 10121
rect 26973 10081 26985 10115
rect 27019 10112 27031 10115
rect 27062 10112 27068 10124
rect 27019 10084 27068 10112
rect 27019 10081 27031 10084
rect 26973 10075 27031 10081
rect 10686 10044 10692 10056
rect 10647 10016 10692 10044
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 15739 10044 15767 10075
rect 27062 10072 27068 10084
rect 27120 10072 27126 10124
rect 27985 10115 28043 10121
rect 27985 10081 27997 10115
rect 28031 10081 28043 10115
rect 27985 10075 28043 10081
rect 15838 10044 15844 10056
rect 15739 10016 15844 10044
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 16669 10047 16727 10053
rect 16669 10044 16681 10047
rect 16540 10016 16681 10044
rect 16540 10004 16546 10016
rect 16669 10013 16681 10016
rect 16715 10013 16727 10047
rect 16669 10007 16727 10013
rect 20070 10004 20076 10056
rect 20128 10044 20134 10056
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20128 10016 20913 10044
rect 20128 10004 20134 10016
rect 20901 10013 20913 10016
rect 20947 10044 20959 10047
rect 22462 10044 22468 10056
rect 20947 10016 22468 10044
rect 20947 10013 20959 10016
rect 20901 10007 20959 10013
rect 22462 10004 22468 10016
rect 22520 10004 22526 10056
rect 23014 10044 23020 10056
rect 22975 10016 23020 10044
rect 23014 10004 23020 10016
rect 23072 10004 23078 10056
rect 23658 10004 23664 10056
rect 23716 10044 23722 10056
rect 24854 10044 24860 10056
rect 23716 10016 24860 10044
rect 23716 10004 23722 10016
rect 24854 10004 24860 10016
rect 24912 10004 24918 10056
rect 11698 9936 11704 9988
rect 11756 9976 11762 9988
rect 13906 9976 13912 9988
rect 11756 9948 13912 9976
rect 11756 9936 11762 9948
rect 13906 9936 13912 9948
rect 13964 9936 13970 9988
rect 14274 9976 14280 9988
rect 14235 9948 14280 9976
rect 14274 9936 14280 9948
rect 14332 9936 14338 9988
rect 26878 9976 26884 9988
rect 25694 9948 26884 9976
rect 17586 9908 17592 9920
rect 17547 9880 17592 9908
rect 17586 9868 17592 9880
rect 17644 9868 17650 9920
rect 19981 9911 20039 9917
rect 19981 9877 19993 9911
rect 20027 9908 20039 9911
rect 21266 9908 21272 9920
rect 20027 9880 21272 9908
rect 20027 9877 20039 9880
rect 19981 9871 20039 9877
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 21358 9868 21364 9920
rect 21416 9908 21422 9920
rect 21821 9911 21879 9917
rect 21821 9908 21833 9911
rect 21416 9880 21833 9908
rect 21416 9868 21422 9880
rect 21821 9877 21833 9880
rect 21867 9877 21879 9911
rect 21821 9871 21879 9877
rect 23014 9868 23020 9920
rect 23072 9908 23078 9920
rect 25694 9908 25722 9948
rect 26878 9936 26884 9948
rect 26936 9936 26942 9988
rect 28000 9976 28028 10075
rect 28074 10072 28080 10124
rect 28132 10112 28138 10124
rect 28442 10112 28448 10124
rect 28132 10084 28448 10112
rect 28132 10072 28138 10084
rect 28442 10072 28448 10084
rect 28500 10072 28506 10124
rect 31754 10072 31760 10124
rect 31812 10112 31818 10124
rect 36538 10112 36544 10124
rect 31812 10084 36544 10112
rect 31812 10072 31818 10084
rect 36538 10072 36544 10084
rect 36596 10072 36602 10124
rect 36814 10072 36820 10124
rect 36872 10112 36878 10124
rect 37277 10115 37335 10121
rect 37277 10112 37289 10115
rect 36872 10084 37289 10112
rect 36872 10072 36878 10084
rect 37277 10081 37289 10084
rect 37323 10081 37335 10115
rect 37277 10075 37335 10081
rect 39574 10072 39580 10124
rect 39632 10112 39638 10124
rect 40126 10112 40132 10124
rect 39632 10084 40132 10112
rect 39632 10072 39638 10084
rect 40126 10072 40132 10084
rect 40184 10072 40190 10124
rect 28718 10044 28724 10056
rect 28679 10016 28724 10044
rect 28718 10004 28724 10016
rect 28776 10004 28782 10056
rect 29546 10044 29552 10056
rect 29507 10016 29552 10044
rect 29546 10004 29552 10016
rect 29604 10004 29610 10056
rect 33505 10047 33563 10053
rect 33505 10013 33517 10047
rect 33551 10044 33563 10047
rect 33778 10044 33784 10056
rect 33551 10016 33784 10044
rect 33551 10013 33563 10016
rect 33505 10007 33563 10013
rect 33778 10004 33784 10016
rect 33836 10004 33842 10056
rect 35710 10044 35716 10056
rect 35671 10016 35716 10044
rect 35710 10004 35716 10016
rect 35768 10004 35774 10056
rect 37829 10047 37887 10053
rect 37829 10013 37841 10047
rect 37875 10044 37887 10047
rect 37918 10044 37924 10056
rect 37875 10016 37924 10044
rect 37875 10013 37887 10016
rect 37829 10007 37887 10013
rect 37918 10004 37924 10016
rect 37976 10004 37982 10056
rect 38102 10044 38108 10056
rect 38063 10016 38108 10044
rect 38102 10004 38108 10016
rect 38160 10004 38166 10056
rect 28166 9976 28172 9988
rect 28000 9948 28172 9976
rect 28166 9936 28172 9948
rect 28224 9976 28230 9988
rect 32950 9976 32956 9988
rect 28224 9948 32956 9976
rect 28224 9936 28230 9948
rect 32950 9936 32956 9948
rect 33008 9976 33014 9988
rect 34698 9976 34704 9988
rect 33008 9948 34704 9976
rect 33008 9936 33014 9948
rect 34698 9936 34704 9948
rect 34756 9936 34762 9988
rect 23072 9880 25722 9908
rect 23072 9868 23078 9880
rect 1104 9818 48852 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 48852 9818
rect 1104 9744 48852 9766
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 10226 9704 10232 9716
rect 9815 9676 10232 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 10502 9704 10508 9716
rect 10463 9676 10508 9704
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11756 9676 11805 9704
rect 11756 9664 11762 9676
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 12158 9704 12164 9716
rect 12119 9676 12164 9704
rect 11793 9667 11851 9673
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 13906 9704 13912 9716
rect 13819 9676 13912 9704
rect 13906 9664 13912 9676
rect 13964 9704 13970 9716
rect 15289 9707 15347 9713
rect 13964 9676 15056 9704
rect 13964 9664 13970 9676
rect 10134 9636 10140 9648
rect 10095 9608 10140 9636
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 14182 9636 14188 9648
rect 13924 9608 14188 9636
rect 10597 9571 10655 9577
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 10686 9568 10692 9580
rect 10643 9540 10692 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 13924 9577 13952 9608
rect 14182 9596 14188 9608
rect 14240 9596 14246 9648
rect 15028 9636 15056 9676
rect 15289 9673 15301 9707
rect 15335 9704 15347 9707
rect 15838 9704 15844 9716
rect 15335 9676 15844 9704
rect 15335 9673 15347 9676
rect 15289 9667 15347 9673
rect 15838 9664 15844 9676
rect 15896 9664 15902 9716
rect 16666 9704 16672 9716
rect 16627 9676 16672 9704
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 18506 9704 18512 9716
rect 18467 9676 18512 9704
rect 18506 9664 18512 9676
rect 18564 9664 18570 9716
rect 19150 9704 19156 9716
rect 19111 9676 19156 9704
rect 19150 9664 19156 9676
rect 19208 9704 19214 9716
rect 19521 9707 19579 9713
rect 19521 9704 19533 9707
rect 19208 9676 19533 9704
rect 19208 9664 19214 9676
rect 19521 9673 19533 9676
rect 19567 9673 19579 9707
rect 21266 9704 21272 9716
rect 21227 9676 21272 9704
rect 19521 9667 19579 9673
rect 21266 9664 21272 9676
rect 21324 9664 21330 9716
rect 22462 9704 22468 9716
rect 22423 9676 22468 9704
rect 22462 9664 22468 9676
rect 22520 9664 22526 9716
rect 22922 9664 22928 9716
rect 22980 9704 22986 9716
rect 23017 9707 23075 9713
rect 23017 9704 23029 9707
rect 22980 9676 23029 9704
rect 22980 9664 22986 9676
rect 23017 9673 23029 9676
rect 23063 9673 23075 9707
rect 23017 9667 23075 9673
rect 24670 9664 24676 9716
rect 24728 9704 24734 9716
rect 25041 9707 25099 9713
rect 25041 9704 25053 9707
rect 24728 9676 25053 9704
rect 24728 9664 24734 9676
rect 25041 9673 25053 9676
rect 25087 9704 25099 9707
rect 25133 9707 25191 9713
rect 25133 9704 25145 9707
rect 25087 9676 25145 9704
rect 25087 9673 25099 9676
rect 25041 9667 25099 9673
rect 25133 9673 25145 9676
rect 25179 9704 25191 9707
rect 25406 9704 25412 9716
rect 25179 9676 25412 9704
rect 25179 9673 25191 9676
rect 25133 9667 25191 9673
rect 25406 9664 25412 9676
rect 25464 9664 25470 9716
rect 26605 9707 26663 9713
rect 26605 9673 26617 9707
rect 26651 9704 26663 9707
rect 27062 9704 27068 9716
rect 26651 9676 27068 9704
rect 26651 9673 26663 9676
rect 26605 9667 26663 9673
rect 27062 9664 27068 9676
rect 27120 9664 27126 9716
rect 28166 9704 28172 9716
rect 28127 9676 28172 9704
rect 28166 9664 28172 9676
rect 28224 9664 28230 9716
rect 28442 9704 28448 9716
rect 28403 9676 28448 9704
rect 28442 9664 28448 9676
rect 28500 9664 28506 9716
rect 28902 9664 28908 9716
rect 28960 9704 28966 9716
rect 28997 9707 29055 9713
rect 28997 9704 29009 9707
rect 28960 9676 29009 9704
rect 28960 9664 28966 9676
rect 28997 9673 29009 9676
rect 29043 9673 29055 9707
rect 28997 9667 29055 9673
rect 29914 9664 29920 9716
rect 29972 9704 29978 9716
rect 30193 9707 30251 9713
rect 30193 9704 30205 9707
rect 29972 9676 30205 9704
rect 29972 9664 29978 9676
rect 30193 9673 30205 9676
rect 30239 9673 30251 9707
rect 30193 9667 30251 9673
rect 31941 9707 31999 9713
rect 31941 9673 31953 9707
rect 31987 9704 31999 9707
rect 32030 9704 32036 9716
rect 31987 9676 32036 9704
rect 31987 9673 31999 9676
rect 31941 9667 31999 9673
rect 32030 9664 32036 9676
rect 32088 9664 32094 9716
rect 36722 9704 36728 9716
rect 36683 9676 36728 9704
rect 36722 9664 36728 9676
rect 36780 9664 36786 9716
rect 37734 9704 37740 9716
rect 37695 9676 37740 9704
rect 37734 9664 37740 9676
rect 37792 9664 37798 9716
rect 37918 9664 37924 9716
rect 37976 9704 37982 9716
rect 38105 9707 38163 9713
rect 38105 9704 38117 9707
rect 37976 9676 38117 9704
rect 37976 9664 37982 9676
rect 38105 9673 38117 9676
rect 38151 9673 38163 9707
rect 38105 9667 38163 9673
rect 39942 9664 39948 9716
rect 40000 9704 40006 9716
rect 40129 9707 40187 9713
rect 40129 9704 40141 9707
rect 40000 9676 40141 9704
rect 40000 9664 40006 9676
rect 40129 9673 40141 9676
rect 40175 9673 40187 9707
rect 40129 9667 40187 9673
rect 41417 9707 41475 9713
rect 41417 9673 41429 9707
rect 41463 9704 41475 9707
rect 41506 9704 41512 9716
rect 41463 9676 41512 9704
rect 41463 9673 41475 9676
rect 41417 9667 41475 9673
rect 41506 9664 41512 9676
rect 41564 9664 41570 9716
rect 16574 9636 16580 9648
rect 15028 9608 16580 9636
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 23658 9596 23664 9648
rect 23716 9636 23722 9648
rect 24857 9639 24915 9645
rect 23716 9608 24072 9636
rect 23716 9596 23722 9608
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9537 13967 9571
rect 14274 9568 14280 9580
rect 14235 9540 14280 9568
rect 13909 9531 13967 9537
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 17083 9571 17141 9577
rect 17083 9537 17095 9571
rect 17129 9568 17141 9571
rect 21542 9568 21548 9580
rect 17129 9540 21548 9568
rect 17129 9537 17141 9540
rect 17083 9531 17141 9537
rect 21542 9528 21548 9540
rect 21600 9528 21606 9580
rect 21818 9568 21824 9580
rect 21779 9540 21824 9568
rect 21818 9528 21824 9540
rect 21876 9528 21882 9580
rect 23382 9528 23388 9580
rect 23440 9568 23446 9580
rect 24044 9577 24072 9608
rect 24857 9605 24869 9639
rect 24903 9636 24915 9639
rect 24946 9636 24952 9648
rect 24903 9608 24952 9636
rect 24903 9605 24915 9608
rect 24857 9599 24915 9605
rect 24946 9596 24952 9608
rect 25004 9636 25010 9648
rect 26237 9639 26295 9645
rect 26237 9636 26249 9639
rect 25004 9608 26249 9636
rect 25004 9596 25010 9608
rect 26237 9605 26249 9608
rect 26283 9605 26295 9639
rect 26237 9599 26295 9605
rect 28810 9596 28816 9648
rect 28868 9636 28874 9648
rect 32861 9639 32919 9645
rect 32861 9636 32873 9639
rect 28868 9608 32873 9636
rect 28868 9596 28874 9608
rect 32861 9605 32873 9608
rect 32907 9605 32919 9639
rect 32861 9599 32919 9605
rect 23753 9571 23811 9577
rect 23753 9568 23765 9571
rect 23440 9540 23765 9568
rect 23440 9528 23446 9540
rect 23753 9537 23765 9540
rect 23799 9537 23811 9571
rect 23753 9531 23811 9537
rect 24029 9571 24087 9577
rect 24029 9537 24041 9571
rect 24075 9537 24087 9571
rect 27614 9568 27620 9580
rect 27575 9540 27620 9568
rect 24029 9531 24087 9537
rect 27614 9528 27620 9540
rect 27672 9528 27678 9580
rect 28718 9528 28724 9580
rect 28776 9568 28782 9580
rect 29270 9568 29276 9580
rect 28776 9540 29276 9568
rect 28776 9528 28782 9540
rect 29270 9528 29276 9540
rect 29328 9528 29334 9580
rect 29546 9528 29552 9580
rect 29604 9568 29610 9580
rect 30469 9571 30527 9577
rect 30469 9568 30481 9571
rect 29604 9540 30481 9568
rect 29604 9528 29610 9540
rect 30469 9537 30481 9540
rect 30515 9537 30527 9571
rect 30469 9531 30527 9537
rect 12504 9503 12562 9509
rect 12504 9469 12516 9503
rect 12550 9469 12562 9503
rect 14918 9500 14924 9512
rect 14831 9472 14924 9500
rect 12504 9463 12562 9469
rect 10502 9392 10508 9444
rect 10560 9432 10566 9444
rect 10918 9435 10976 9441
rect 10918 9432 10930 9435
rect 10560 9404 10930 9432
rect 10560 9392 10566 9404
rect 10918 9401 10930 9404
rect 10964 9432 10976 9435
rect 11238 9432 11244 9444
rect 10964 9404 11244 9432
rect 10964 9401 10976 9404
rect 10918 9395 10976 9401
rect 11238 9392 11244 9404
rect 11296 9392 11302 9444
rect 12519 9432 12547 9463
rect 14918 9460 14924 9472
rect 14976 9500 14982 9512
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 14976 9472 15485 9500
rect 14976 9460 14982 9472
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 16996 9503 17054 9509
rect 16996 9469 17008 9503
rect 17042 9500 17054 9503
rect 18116 9503 18174 9509
rect 17042 9472 17540 9500
rect 17042 9469 17054 9472
rect 16996 9463 17054 9469
rect 12989 9435 13047 9441
rect 12989 9432 13001 9435
rect 12519 9404 13001 9432
rect 12989 9401 13001 9404
rect 13035 9432 13047 9435
rect 13538 9432 13544 9444
rect 13035 9404 13544 9432
rect 13035 9401 13047 9404
rect 12989 9395 13047 9401
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 13725 9435 13783 9441
rect 13725 9401 13737 9435
rect 13771 9432 13783 9435
rect 14001 9435 14059 9441
rect 14001 9432 14013 9435
rect 13771 9404 14013 9432
rect 13771 9401 13783 9404
rect 13725 9395 13783 9401
rect 14001 9401 14013 9404
rect 14047 9432 14059 9435
rect 15381 9435 15439 9441
rect 15381 9432 15393 9435
rect 14047 9404 15393 9432
rect 14047 9401 14059 9404
rect 14001 9395 14059 9401
rect 15381 9401 15393 9404
rect 15427 9401 15439 9435
rect 15381 9395 15439 9401
rect 11514 9364 11520 9376
rect 11475 9336 11520 9364
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12575 9367 12633 9373
rect 12575 9364 12587 9367
rect 12492 9336 12587 9364
rect 12492 9324 12498 9336
rect 12575 9333 12587 9336
rect 12621 9333 12633 9367
rect 12575 9327 12633 9333
rect 13357 9367 13415 9373
rect 13357 9333 13369 9367
rect 13403 9364 13415 9367
rect 13630 9364 13636 9376
rect 13403 9336 13636 9364
rect 13403 9333 13415 9336
rect 13357 9327 13415 9333
rect 13630 9324 13636 9336
rect 13688 9364 13694 9376
rect 13814 9364 13820 9376
rect 13688 9336 13820 9364
rect 13688 9324 13694 9336
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 17512 9373 17540 9472
rect 18116 9469 18128 9503
rect 18162 9500 18174 9503
rect 18506 9500 18512 9512
rect 18162 9472 18512 9500
rect 18162 9469 18174 9472
rect 18116 9463 18174 9469
rect 18506 9460 18512 9472
rect 18564 9460 18570 9512
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 19886 9500 19892 9512
rect 19751 9472 19892 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 19886 9460 19892 9472
rect 19944 9460 19950 9512
rect 23477 9503 23535 9509
rect 23477 9469 23489 9503
rect 23523 9500 23535 9503
rect 23566 9500 23572 9512
rect 23523 9472 23572 9500
rect 23523 9469 23535 9472
rect 23477 9463 23535 9469
rect 23566 9460 23572 9472
rect 23624 9460 23630 9512
rect 25314 9500 25320 9512
rect 25275 9472 25320 9500
rect 25314 9460 25320 9472
rect 25372 9460 25378 9512
rect 26973 9503 27031 9509
rect 26973 9469 26985 9503
rect 27019 9500 27031 9503
rect 27157 9503 27215 9509
rect 27157 9500 27169 9503
rect 27019 9472 27169 9500
rect 27019 9469 27031 9472
rect 26973 9463 27031 9469
rect 27157 9469 27169 9472
rect 27203 9469 27215 9503
rect 27157 9463 27215 9469
rect 20901 9435 20959 9441
rect 20901 9432 20913 9435
rect 20088 9404 20913 9432
rect 17497 9367 17555 9373
rect 17497 9333 17509 9367
rect 17543 9364 17555 9367
rect 18187 9367 18245 9373
rect 18187 9364 18199 9367
rect 17543 9336 18199 9364
rect 17543 9333 17555 9336
rect 17497 9327 17555 9333
rect 18187 9333 18199 9336
rect 18233 9364 18245 9367
rect 18506 9364 18512 9376
rect 18233 9336 18512 9364
rect 18233 9333 18245 9336
rect 18187 9327 18245 9333
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 19978 9324 19984 9376
rect 20036 9364 20042 9376
rect 20088 9373 20116 9404
rect 20901 9401 20913 9404
rect 20947 9401 20959 9435
rect 20901 9395 20959 9401
rect 21637 9435 21695 9441
rect 21637 9401 21649 9435
rect 21683 9401 21695 9435
rect 23584 9432 23612 9460
rect 23845 9435 23903 9441
rect 23845 9432 23857 9435
rect 23584 9404 23857 9432
rect 21637 9395 21695 9401
rect 23845 9401 23857 9404
rect 23891 9401 23903 9435
rect 23845 9395 23903 9401
rect 25041 9435 25099 9441
rect 25041 9401 25053 9435
rect 25087 9432 25099 9435
rect 25638 9435 25696 9441
rect 25638 9432 25650 9435
rect 25087 9404 25650 9432
rect 25087 9401 25099 9404
rect 25041 9395 25099 9401
rect 25638 9401 25650 9404
rect 25684 9401 25696 9435
rect 27172 9432 27200 9463
rect 27246 9460 27252 9512
rect 27304 9500 27310 9512
rect 27525 9503 27583 9509
rect 27525 9500 27537 9503
rect 27304 9472 27537 9500
rect 27304 9460 27310 9472
rect 27525 9469 27537 9472
rect 27571 9469 27583 9503
rect 31018 9500 31024 9512
rect 30979 9472 31024 9500
rect 27525 9463 27583 9469
rect 31018 9460 31024 9472
rect 31076 9460 31082 9512
rect 32876 9500 32904 9599
rect 34514 9596 34520 9648
rect 34572 9636 34578 9648
rect 38562 9636 38568 9648
rect 34572 9608 38568 9636
rect 34572 9596 34578 9608
rect 38562 9596 38568 9608
rect 38620 9596 38626 9648
rect 33778 9568 33784 9580
rect 33691 9540 33784 9568
rect 33778 9528 33784 9540
rect 33836 9568 33842 9580
rect 34425 9571 34483 9577
rect 34425 9568 34437 9571
rect 33836 9540 34437 9568
rect 33836 9528 33842 9540
rect 34425 9537 34437 9540
rect 34471 9537 34483 9571
rect 34425 9531 34483 9537
rect 34698 9528 34704 9580
rect 34756 9568 34762 9580
rect 38657 9571 38715 9577
rect 38657 9568 38669 9571
rect 34756 9540 38669 9568
rect 34756 9528 34762 9540
rect 38657 9537 38669 9540
rect 38703 9537 38715 9571
rect 38657 9531 38715 9537
rect 33045 9503 33103 9509
rect 33045 9500 33057 9503
rect 32876 9472 33057 9500
rect 33045 9469 33057 9472
rect 33091 9469 33103 9503
rect 33045 9463 33103 9469
rect 33597 9503 33655 9509
rect 33597 9469 33609 9503
rect 33643 9500 33655 9503
rect 33962 9500 33968 9512
rect 33643 9472 33968 9500
rect 33643 9469 33655 9472
rect 33597 9463 33655 9469
rect 33962 9460 33968 9472
rect 34020 9460 34026 9512
rect 35802 9500 35808 9512
rect 35763 9472 35808 9500
rect 35802 9460 35808 9472
rect 35860 9460 35866 9512
rect 38672 9500 38700 9531
rect 38841 9503 38899 9509
rect 38841 9500 38853 9503
rect 38672 9472 38853 9500
rect 38841 9469 38853 9472
rect 38887 9469 38899 9503
rect 38841 9463 38899 9469
rect 39114 9460 39120 9512
rect 39172 9500 39178 9512
rect 39301 9503 39359 9509
rect 39301 9500 39313 9503
rect 39172 9472 39313 9500
rect 39172 9460 39178 9472
rect 39301 9469 39313 9472
rect 39347 9469 39359 9503
rect 39301 9463 39359 9469
rect 39577 9503 39635 9509
rect 39577 9469 39589 9503
rect 39623 9500 39635 9503
rect 40494 9500 40500 9512
rect 39623 9472 40500 9500
rect 39623 9469 39635 9472
rect 39577 9463 39635 9469
rect 40494 9460 40500 9472
rect 40552 9460 40558 9512
rect 27798 9432 27804 9444
rect 27172 9404 27804 9432
rect 25638 9395 25696 9401
rect 20073 9367 20131 9373
rect 20073 9364 20085 9367
rect 20036 9336 20085 9364
rect 20036 9324 20042 9336
rect 20073 9333 20085 9336
rect 20119 9333 20131 9367
rect 20622 9364 20628 9376
rect 20583 9336 20628 9364
rect 20073 9327 20131 9333
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 21266 9324 21272 9376
rect 21324 9364 21330 9376
rect 21652 9364 21680 9395
rect 27798 9392 27804 9404
rect 27856 9392 27862 9444
rect 28902 9392 28908 9444
rect 28960 9432 28966 9444
rect 29594 9435 29652 9441
rect 29594 9432 29606 9435
rect 28960 9404 29606 9432
rect 28960 9392 28966 9404
rect 29594 9401 29606 9404
rect 29640 9432 29652 9435
rect 30837 9435 30895 9441
rect 30837 9432 30849 9435
rect 29640 9404 30849 9432
rect 29640 9401 29652 9404
rect 29594 9395 29652 9401
rect 30837 9401 30849 9404
rect 30883 9432 30895 9435
rect 31342 9435 31400 9441
rect 31342 9432 31354 9435
rect 30883 9404 31354 9432
rect 30883 9401 30895 9404
rect 30837 9395 30895 9401
rect 31342 9401 31354 9404
rect 31388 9432 31400 9435
rect 33134 9432 33140 9444
rect 31388 9404 33140 9432
rect 31388 9401 31400 9404
rect 31342 9395 31400 9401
rect 33134 9392 33140 9404
rect 33192 9432 33198 9444
rect 34057 9435 34115 9441
rect 34057 9432 34069 9435
rect 33192 9404 34069 9432
rect 33192 9392 33198 9404
rect 34057 9401 34069 9404
rect 34103 9432 34115 9435
rect 35253 9435 35311 9441
rect 35253 9432 35265 9435
rect 34103 9404 35265 9432
rect 34103 9401 34115 9404
rect 34057 9395 34115 9401
rect 35253 9401 35265 9404
rect 35299 9432 35311 9435
rect 35621 9435 35679 9441
rect 35621 9432 35633 9435
rect 35299 9404 35633 9432
rect 35299 9401 35311 9404
rect 35253 9395 35311 9401
rect 35621 9401 35633 9404
rect 35667 9432 35679 9435
rect 36078 9432 36084 9444
rect 35667 9404 36084 9432
rect 35667 9401 35679 9404
rect 35621 9395 35679 9401
rect 36078 9392 36084 9404
rect 36136 9441 36142 9444
rect 36136 9435 36184 9441
rect 36136 9401 36138 9435
rect 36172 9401 36184 9435
rect 36136 9395 36184 9401
rect 36136 9392 36142 9395
rect 39942 9392 39948 9444
rect 40000 9432 40006 9444
rect 40818 9435 40876 9441
rect 40818 9432 40830 9435
rect 40000 9404 40830 9432
rect 40000 9392 40006 9404
rect 40818 9401 40830 9404
rect 40864 9401 40876 9435
rect 40818 9395 40876 9401
rect 21324 9336 21680 9364
rect 21324 9324 21330 9336
rect 1104 9274 48852 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 48852 9274
rect 1104 9200 48852 9222
rect 10686 9160 10692 9172
rect 10647 9132 10692 9160
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11238 9160 11244 9172
rect 11199 9132 11244 9160
rect 11238 9120 11244 9132
rect 11296 9120 11302 9172
rect 12434 9160 12440 9172
rect 12395 9132 12440 9160
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 13909 9163 13967 9169
rect 13909 9129 13921 9163
rect 13955 9160 13967 9163
rect 14182 9160 14188 9172
rect 13955 9132 14188 9160
rect 13955 9129 13967 9132
rect 13909 9123 13967 9129
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 21542 9120 21548 9172
rect 21600 9160 21606 9172
rect 21913 9163 21971 9169
rect 21913 9160 21925 9163
rect 21600 9132 21925 9160
rect 21600 9120 21606 9132
rect 21913 9129 21925 9132
rect 21959 9129 21971 9163
rect 21913 9123 21971 9129
rect 22603 9163 22661 9169
rect 22603 9129 22615 9163
rect 22649 9160 22661 9163
rect 23198 9160 23204 9172
rect 22649 9132 23204 9160
rect 22649 9129 22661 9132
rect 22603 9123 22661 9129
rect 23198 9120 23204 9132
rect 23256 9120 23262 9172
rect 23382 9120 23388 9172
rect 23440 9160 23446 9172
rect 23661 9163 23719 9169
rect 23661 9160 23673 9163
rect 23440 9132 23673 9160
rect 23440 9120 23446 9132
rect 23661 9129 23673 9132
rect 23707 9129 23719 9163
rect 24854 9160 24860 9172
rect 24815 9132 24860 9160
rect 23661 9123 23719 9129
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 25314 9120 25320 9172
rect 25372 9160 25378 9172
rect 25409 9163 25467 9169
rect 25409 9160 25421 9163
rect 25372 9132 25421 9160
rect 25372 9120 25378 9132
rect 25409 9129 25421 9132
rect 25455 9160 25467 9163
rect 26605 9163 26663 9169
rect 26605 9160 26617 9163
rect 25455 9132 26617 9160
rect 25455 9129 25467 9132
rect 25409 9123 25467 9129
rect 26605 9129 26617 9132
rect 26651 9129 26663 9163
rect 26605 9123 26663 9129
rect 29270 9120 29276 9172
rect 29328 9160 29334 9172
rect 29733 9163 29791 9169
rect 29733 9160 29745 9163
rect 29328 9132 29745 9160
rect 29328 9120 29334 9132
rect 29733 9129 29745 9132
rect 29779 9129 29791 9163
rect 29733 9123 29791 9129
rect 33137 9163 33195 9169
rect 33137 9129 33149 9163
rect 33183 9160 33195 9163
rect 33962 9160 33968 9172
rect 33183 9132 33968 9160
rect 33183 9129 33195 9132
rect 33137 9123 33195 9129
rect 33962 9120 33968 9132
rect 34020 9120 34026 9172
rect 35710 9160 35716 9172
rect 35671 9132 35716 9160
rect 35710 9120 35716 9132
rect 35768 9120 35774 9172
rect 36679 9163 36737 9169
rect 36679 9129 36691 9163
rect 36725 9160 36737 9163
rect 37090 9160 37096 9172
rect 36725 9132 37096 9160
rect 36725 9129 36737 9132
rect 36679 9123 36737 9129
rect 37090 9120 37096 9132
rect 37148 9120 37154 9172
rect 38933 9163 38991 9169
rect 38933 9129 38945 9163
rect 38979 9160 38991 9163
rect 39114 9160 39120 9172
rect 38979 9132 39120 9160
rect 38979 9129 38991 9132
rect 38933 9123 38991 9129
rect 39114 9120 39120 9132
rect 39172 9120 39178 9172
rect 40126 9160 40132 9172
rect 40087 9132 40132 9160
rect 40126 9120 40132 9132
rect 40184 9120 40190 9172
rect 40494 9120 40500 9172
rect 40552 9160 40558 9172
rect 40865 9163 40923 9169
rect 40865 9160 40877 9163
rect 40552 9132 40877 9160
rect 40552 9120 40558 9132
rect 40865 9129 40877 9132
rect 40911 9129 40923 9163
rect 40865 9123 40923 9129
rect 12805 9095 12863 9101
rect 12805 9092 12817 9095
rect 12487 9064 12817 9092
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 9024 10931 9027
rect 11698 9024 11704 9036
rect 10919 8996 11704 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 9024 11851 9027
rect 12487 9024 12515 9064
rect 12805 9061 12817 9064
rect 12851 9092 12863 9095
rect 13446 9092 13452 9104
rect 12851 9064 13452 9092
rect 12851 9061 12863 9064
rect 12805 9055 12863 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 13538 9052 13544 9104
rect 13596 9092 13602 9104
rect 15427 9095 15485 9101
rect 15427 9092 15439 9095
rect 13596 9064 15439 9092
rect 13596 9052 13602 9064
rect 15427 9061 15439 9064
rect 15473 9061 15485 9095
rect 15427 9055 15485 9061
rect 17313 9095 17371 9101
rect 17313 9061 17325 9095
rect 17359 9092 17371 9095
rect 17586 9092 17592 9104
rect 17359 9064 17592 9092
rect 17359 9061 17371 9064
rect 17313 9055 17371 9061
rect 17586 9052 17592 9064
rect 17644 9052 17650 9104
rect 19705 9095 19763 9101
rect 19705 9061 19717 9095
rect 19751 9092 19763 9095
rect 19886 9092 19892 9104
rect 19751 9064 19892 9092
rect 19751 9061 19763 9064
rect 19705 9055 19763 9061
rect 19886 9052 19892 9064
rect 19944 9092 19950 9104
rect 19981 9095 20039 9101
rect 19981 9092 19993 9095
rect 19944 9064 19993 9092
rect 19944 9052 19950 9064
rect 19981 9061 19993 9064
rect 20027 9061 20039 9095
rect 19981 9055 20039 9061
rect 20622 9052 20628 9104
rect 20680 9092 20686 9104
rect 21085 9095 21143 9101
rect 21085 9092 21097 9095
rect 20680 9064 21097 9092
rect 20680 9052 20686 9064
rect 21085 9061 21097 9064
rect 21131 9061 21143 9095
rect 21085 9055 21143 9061
rect 21637 9095 21695 9101
rect 21637 9061 21649 9095
rect 21683 9092 21695 9095
rect 21818 9092 21824 9104
rect 21683 9064 21824 9092
rect 21683 9061 21695 9064
rect 21637 9055 21695 9061
rect 21818 9052 21824 9064
rect 21876 9092 21882 9104
rect 23014 9092 23020 9104
rect 21876 9064 22600 9092
rect 22975 9064 23020 9092
rect 21876 9052 21882 9064
rect 14182 9024 14188 9036
rect 11839 8996 12515 9024
rect 14143 8996 14188 9024
rect 11839 8993 11851 8996
rect 11793 8987 11851 8993
rect 14182 8984 14188 8996
rect 14240 8984 14246 9036
rect 14274 8984 14280 9036
rect 14332 9024 14338 9036
rect 15324 9027 15382 9033
rect 15324 9024 15336 9027
rect 14332 8996 15336 9024
rect 14332 8984 14338 8996
rect 15324 8993 15336 8996
rect 15370 9024 15382 9027
rect 15749 9027 15807 9033
rect 15749 9024 15761 9027
rect 15370 8996 15761 9024
rect 15370 8993 15382 8996
rect 15324 8987 15382 8993
rect 15749 8993 15761 8996
rect 15795 8993 15807 9027
rect 15749 8987 15807 8993
rect 18690 8984 18696 9036
rect 18748 9024 18754 9036
rect 18969 9027 19027 9033
rect 18969 9024 18981 9027
rect 18748 8996 18981 9024
rect 18748 8984 18754 8996
rect 18969 8993 18981 8996
rect 19015 8993 19027 9027
rect 19426 9024 19432 9036
rect 19387 8996 19432 9024
rect 18969 8987 19027 8993
rect 19426 8984 19432 8996
rect 19484 8984 19490 9036
rect 22572 9033 22600 9064
rect 23014 9052 23020 9064
rect 23072 9052 23078 9104
rect 26786 9052 26792 9104
rect 26844 9092 26850 9104
rect 26844 9064 28247 9092
rect 26844 9052 26850 9064
rect 22532 9027 22600 9033
rect 22532 8993 22544 9027
rect 22578 8996 22600 9027
rect 26697 9027 26755 9033
rect 22578 8993 22590 8996
rect 22532 8987 22590 8993
rect 26697 8993 26709 9027
rect 26743 8993 26755 9027
rect 26697 8987 26755 8993
rect 27065 9027 27123 9033
rect 27065 8993 27077 9027
rect 27111 9024 27123 9027
rect 27246 9024 27252 9036
rect 27111 8996 27252 9024
rect 27111 8993 27123 8996
rect 27065 8987 27123 8993
rect 12710 8956 12716 8968
rect 12671 8928 12716 8956
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 13078 8956 13084 8968
rect 13039 8928 13084 8956
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 17221 8959 17279 8965
rect 17221 8925 17233 8959
rect 17267 8956 17279 8959
rect 17494 8956 17500 8968
rect 17267 8928 17500 8956
rect 17267 8925 17279 8928
rect 17221 8919 17279 8925
rect 17494 8916 17500 8928
rect 17552 8916 17558 8968
rect 17678 8956 17684 8968
rect 17639 8928 17684 8956
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 20993 8959 21051 8965
rect 20993 8925 21005 8959
rect 21039 8956 21051 8959
rect 21174 8956 21180 8968
rect 21039 8928 21180 8956
rect 21039 8925 21051 8928
rect 20993 8919 21051 8925
rect 21174 8916 21180 8928
rect 21232 8916 21238 8968
rect 26712 8956 26740 8987
rect 27246 8984 27252 8996
rect 27304 8984 27310 9036
rect 28219 9024 28247 9064
rect 28442 9052 28448 9104
rect 28500 9092 28506 9104
rect 29457 9095 29515 9101
rect 28500 9064 29224 9092
rect 28500 9052 28506 9064
rect 28718 9024 28724 9036
rect 28219 8996 28724 9024
rect 28718 8984 28724 8996
rect 28776 8984 28782 9036
rect 29196 9033 29224 9064
rect 29457 9061 29469 9095
rect 29503 9092 29515 9095
rect 29546 9092 29552 9104
rect 29503 9064 29552 9092
rect 29503 9061 29515 9064
rect 29457 9055 29515 9061
rect 29546 9052 29552 9064
rect 29604 9052 29610 9104
rect 33980 9092 34008 9120
rect 35437 9095 35495 9101
rect 33980 9064 35204 9092
rect 29181 9027 29239 9033
rect 29181 8993 29193 9027
rect 29227 9024 29239 9027
rect 29730 9024 29736 9036
rect 29227 8996 29736 9024
rect 29227 8993 29239 8996
rect 29181 8987 29239 8993
rect 29730 8984 29736 8996
rect 29788 8984 29794 9036
rect 33594 9024 33600 9036
rect 33555 8996 33600 9024
rect 33594 8984 33600 8996
rect 33652 8984 33658 9036
rect 34698 9024 34704 9036
rect 34659 8996 34704 9024
rect 34698 8984 34704 8996
rect 34756 8984 34762 9036
rect 35176 9033 35204 9064
rect 35437 9061 35449 9095
rect 35483 9092 35495 9095
rect 35802 9092 35808 9104
rect 35483 9064 35808 9092
rect 35483 9061 35495 9064
rect 35437 9055 35495 9061
rect 35802 9052 35808 9064
rect 35860 9092 35866 9104
rect 36081 9095 36139 9101
rect 36081 9092 36093 9095
rect 35860 9064 36093 9092
rect 35860 9052 35866 9064
rect 36081 9061 36093 9064
rect 36127 9061 36139 9095
rect 36081 9055 36139 9061
rect 35161 9027 35219 9033
rect 35161 8993 35173 9027
rect 35207 8993 35219 9027
rect 36538 9024 36544 9036
rect 36499 8996 36544 9024
rect 35161 8987 35219 8993
rect 36538 8984 36544 8996
rect 36596 8984 36602 9036
rect 39942 8984 39948 9036
rect 40000 9024 40006 9036
rect 40497 9027 40555 9033
rect 40497 9024 40509 9027
rect 40000 8996 40509 9024
rect 40000 8984 40006 8996
rect 40497 8993 40509 8996
rect 40543 8993 40555 9027
rect 40497 8987 40555 8993
rect 27154 8956 27160 8968
rect 26712 8928 27160 8956
rect 27154 8916 27160 8928
rect 27212 8956 27218 8968
rect 28166 8956 28172 8968
rect 27212 8928 28172 8956
rect 27212 8916 27218 8928
rect 28166 8916 28172 8928
rect 28224 8916 28230 8968
rect 14366 8820 14372 8832
rect 14327 8792 14372 8820
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 16482 8780 16488 8832
rect 16540 8820 16546 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 16540 8792 16681 8820
rect 16540 8780 16546 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16669 8783 16727 8789
rect 30006 8780 30012 8832
rect 30064 8820 30070 8832
rect 31018 8820 31024 8832
rect 30064 8792 31024 8820
rect 30064 8780 30070 8792
rect 31018 8780 31024 8792
rect 31076 8780 31082 8832
rect 33410 8780 33416 8832
rect 33468 8820 33474 8832
rect 33735 8823 33793 8829
rect 33735 8820 33747 8823
rect 33468 8792 33747 8820
rect 33468 8780 33474 8792
rect 33735 8789 33747 8792
rect 33781 8789 33793 8823
rect 33735 8783 33793 8789
rect 1104 8730 48852 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 48852 8730
rect 1104 8656 48852 8678
rect 10965 8619 11023 8625
rect 10965 8585 10977 8619
rect 11011 8616 11023 8619
rect 11238 8616 11244 8628
rect 11011 8588 11244 8616
rect 11011 8585 11023 8588
rect 10965 8579 11023 8585
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11572 8588 12173 8616
rect 11572 8576 11578 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 12161 8579 12219 8585
rect 11333 8551 11391 8557
rect 11333 8517 11345 8551
rect 11379 8548 11391 8551
rect 11790 8548 11796 8560
rect 11379 8520 11796 8548
rect 11379 8517 11391 8520
rect 11333 8511 11391 8517
rect 11790 8508 11796 8520
rect 11848 8508 11854 8560
rect 12176 8344 12204 8579
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 17586 8576 17592 8628
rect 17644 8616 17650 8628
rect 17681 8619 17739 8625
rect 17681 8616 17693 8619
rect 17644 8588 17693 8616
rect 17644 8576 17650 8588
rect 17681 8585 17693 8588
rect 17727 8585 17739 8619
rect 17681 8579 17739 8585
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 18969 8619 19027 8625
rect 18969 8616 18981 8619
rect 18748 8588 18981 8616
rect 18748 8576 18754 8588
rect 18969 8585 18981 8588
rect 19015 8585 19027 8619
rect 19426 8616 19432 8628
rect 19387 8588 19432 8616
rect 18969 8579 19027 8585
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 20027 8619 20085 8625
rect 20027 8585 20039 8619
rect 20073 8616 20085 8619
rect 20438 8616 20444 8628
rect 20073 8588 20444 8616
rect 20073 8585 20085 8588
rect 20027 8579 20085 8585
rect 20438 8576 20444 8588
rect 20496 8576 20502 8628
rect 20622 8616 20628 8628
rect 20583 8588 20628 8616
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 20990 8616 20996 8628
rect 20951 8588 20996 8616
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 27154 8616 27160 8628
rect 27115 8588 27160 8616
rect 27154 8576 27160 8588
rect 27212 8576 27218 8628
rect 28442 8616 28448 8628
rect 28403 8588 28448 8616
rect 28442 8576 28448 8588
rect 28500 8576 28506 8628
rect 28718 8616 28724 8628
rect 28679 8588 28724 8616
rect 28718 8576 28724 8588
rect 28776 8576 28782 8628
rect 33594 8616 33600 8628
rect 33555 8588 33600 8616
rect 33594 8576 33600 8588
rect 33652 8576 33658 8628
rect 33962 8576 33968 8628
rect 34020 8616 34026 8628
rect 34241 8619 34299 8625
rect 34241 8616 34253 8619
rect 34020 8588 34253 8616
rect 34020 8576 34026 8588
rect 34241 8585 34253 8588
rect 34287 8616 34299 8619
rect 34609 8619 34667 8625
rect 34609 8616 34621 8619
rect 34287 8588 34621 8616
rect 34287 8585 34299 8588
rect 34241 8579 34299 8585
rect 34609 8585 34621 8588
rect 34655 8585 34667 8619
rect 36538 8616 36544 8628
rect 36499 8588 36544 8616
rect 34609 8579 34667 8585
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 13078 8548 13084 8560
rect 12492 8520 12572 8548
rect 13039 8520 13084 8548
rect 12492 8508 12498 8520
rect 12544 8489 12572 8520
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 16574 8508 16580 8560
rect 16632 8548 16638 8560
rect 18708 8548 18736 8576
rect 16632 8520 18736 8548
rect 16632 8508 16638 8520
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 13688 8452 14013 8480
rect 13688 8440 13694 8452
rect 14001 8449 14013 8452
rect 14047 8449 14059 8483
rect 21008 8480 21036 8576
rect 21818 8508 21824 8560
rect 21876 8548 21882 8560
rect 22557 8551 22615 8557
rect 22557 8548 22569 8551
rect 21876 8520 22569 8548
rect 21876 8508 21882 8520
rect 21928 8489 21956 8520
rect 22557 8517 22569 8520
rect 22603 8517 22615 8551
rect 22557 8511 22615 8517
rect 21269 8483 21327 8489
rect 21269 8480 21281 8483
rect 21008 8452 21281 8480
rect 14001 8443 14059 8449
rect 21269 8449 21281 8452
rect 21315 8449 21327 8483
rect 21913 8483 21971 8489
rect 21913 8480 21925 8483
rect 21891 8452 21925 8480
rect 21269 8443 21327 8449
rect 21913 8449 21925 8452
rect 21959 8449 21971 8483
rect 30006 8480 30012 8492
rect 29967 8452 30012 8480
rect 21913 8443 21971 8449
rect 30006 8440 30012 8452
rect 30064 8440 30070 8492
rect 33781 8483 33839 8489
rect 33781 8449 33793 8483
rect 33827 8480 33839 8483
rect 34238 8480 34244 8492
rect 33827 8452 34244 8480
rect 33827 8449 33839 8452
rect 33781 8443 33839 8449
rect 34238 8440 34244 8452
rect 34296 8440 34302 8492
rect 34624 8480 34652 8579
rect 36538 8576 36544 8588
rect 36596 8576 36602 8628
rect 35621 8483 35679 8489
rect 34624 8452 35388 8480
rect 13909 8415 13967 8421
rect 13909 8381 13921 8415
rect 13955 8412 13967 8415
rect 14366 8412 14372 8424
rect 13955 8384 14372 8412
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 17405 8415 17463 8421
rect 17405 8381 17417 8415
rect 17451 8412 17463 8415
rect 17770 8412 17776 8424
rect 17451 8384 17776 8412
rect 17451 8381 17463 8384
rect 17405 8375 17463 8381
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 17862 8372 17868 8424
rect 17920 8412 17926 8424
rect 18084 8415 18142 8421
rect 18084 8412 18096 8415
rect 17920 8384 18096 8412
rect 17920 8372 17926 8384
rect 18084 8381 18096 8384
rect 18130 8412 18142 8415
rect 18509 8415 18567 8421
rect 18509 8412 18521 8415
rect 18130 8384 18521 8412
rect 18130 8381 18142 8384
rect 18084 8375 18142 8381
rect 18509 8381 18521 8384
rect 18555 8381 18567 8415
rect 18509 8375 18567 8381
rect 19797 8415 19855 8421
rect 19797 8381 19809 8415
rect 19843 8412 19855 8415
rect 19956 8415 20014 8421
rect 19956 8412 19968 8415
rect 19843 8384 19968 8412
rect 19843 8381 19855 8384
rect 19797 8375 19855 8381
rect 19956 8381 19968 8384
rect 20002 8412 20014 8415
rect 20346 8412 20352 8424
rect 20002 8384 20352 8412
rect 20002 8381 20014 8384
rect 19956 8375 20014 8381
rect 20346 8372 20352 8384
rect 20404 8372 20410 8424
rect 26329 8415 26387 8421
rect 26329 8381 26341 8415
rect 26375 8381 26387 8415
rect 26329 8375 26387 8381
rect 12621 8347 12679 8353
rect 12621 8344 12633 8347
rect 12176 8316 12633 8344
rect 12621 8313 12633 8316
rect 12667 8313 12679 8347
rect 12621 8307 12679 8313
rect 14090 8304 14096 8356
rect 14148 8344 14154 8356
rect 15473 8347 15531 8353
rect 15473 8344 15485 8347
rect 14148 8316 15485 8344
rect 14148 8304 14154 8316
rect 15473 8313 15485 8316
rect 15519 8344 15531 8347
rect 15657 8347 15715 8353
rect 15657 8344 15669 8347
rect 15519 8316 15669 8344
rect 15519 8313 15531 8316
rect 15473 8307 15531 8313
rect 15657 8313 15669 8316
rect 15703 8313 15715 8347
rect 15657 8307 15715 8313
rect 17494 8304 17500 8356
rect 17552 8344 17558 8356
rect 18187 8347 18245 8353
rect 18187 8344 18199 8347
rect 17552 8316 18199 8344
rect 17552 8304 17558 8316
rect 18187 8313 18199 8316
rect 18233 8313 18245 8347
rect 18187 8307 18245 8313
rect 21358 8304 21364 8356
rect 21416 8344 21422 8356
rect 25961 8347 26019 8353
rect 21416 8316 21461 8344
rect 21416 8304 21422 8316
rect 25961 8313 25973 8347
rect 26007 8344 26019 8347
rect 26344 8344 26372 8375
rect 26418 8372 26424 8424
rect 26476 8412 26482 8424
rect 26605 8415 26663 8421
rect 26605 8412 26617 8415
rect 26476 8384 26617 8412
rect 26476 8372 26482 8384
rect 26605 8381 26617 8384
rect 26651 8412 26663 8415
rect 27246 8412 27252 8424
rect 26651 8384 27252 8412
rect 26651 8381 26663 8384
rect 26605 8375 26663 8381
rect 27246 8372 27252 8384
rect 27304 8372 27310 8424
rect 29549 8415 29607 8421
rect 29549 8381 29561 8415
rect 29595 8381 29607 8415
rect 29730 8412 29736 8424
rect 29691 8384 29736 8412
rect 29549 8375 29607 8381
rect 29362 8344 29368 8356
rect 26007 8316 29368 8344
rect 26007 8313 26019 8316
rect 25961 8307 26019 8313
rect 29362 8304 29368 8316
rect 29420 8344 29426 8356
rect 29564 8344 29592 8375
rect 29730 8372 29736 8384
rect 29788 8372 29794 8424
rect 34514 8372 34520 8424
rect 34572 8412 34578 8424
rect 34885 8415 34943 8421
rect 34885 8412 34897 8415
rect 34572 8384 34897 8412
rect 34572 8372 34578 8384
rect 34885 8381 34897 8384
rect 34931 8412 34943 8415
rect 35066 8412 35072 8424
rect 34931 8384 35072 8412
rect 34931 8381 34943 8384
rect 34885 8375 34943 8381
rect 35066 8372 35072 8384
rect 35124 8372 35130 8424
rect 35360 8421 35388 8452
rect 35621 8449 35633 8483
rect 35667 8480 35679 8483
rect 35710 8480 35716 8492
rect 35667 8452 35716 8480
rect 35667 8449 35679 8452
rect 35621 8443 35679 8449
rect 35710 8440 35716 8452
rect 35768 8440 35774 8492
rect 35345 8415 35403 8421
rect 35345 8381 35357 8415
rect 35391 8381 35403 8415
rect 35345 8375 35403 8381
rect 33226 8344 33232 8356
rect 29420 8316 33232 8344
rect 29420 8304 29426 8316
rect 33226 8304 33232 8316
rect 33284 8304 33290 8356
rect 15102 8276 15108 8288
rect 15063 8248 15108 8276
rect 15102 8236 15108 8248
rect 15160 8236 15166 8288
rect 21174 8236 21180 8288
rect 21232 8276 21238 8288
rect 22189 8279 22247 8285
rect 22189 8276 22201 8279
rect 21232 8248 22201 8276
rect 21232 8236 21238 8248
rect 22189 8245 22201 8248
rect 22235 8245 22247 8279
rect 26142 8276 26148 8288
rect 26103 8248 26148 8276
rect 22189 8239 22247 8245
rect 26142 8236 26148 8248
rect 26200 8236 26206 8288
rect 1104 8186 48852 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 48852 8186
rect 1104 8112 48852 8134
rect 12710 8072 12716 8084
rect 12671 8044 12716 8072
rect 12710 8032 12716 8044
rect 12768 8072 12774 8084
rect 13219 8075 13277 8081
rect 13219 8072 13231 8075
rect 12768 8044 13231 8072
rect 12768 8032 12774 8044
rect 13219 8041 13231 8044
rect 13265 8041 13277 8075
rect 13219 8035 13277 8041
rect 14323 8075 14381 8081
rect 14323 8041 14335 8075
rect 14369 8072 14381 8075
rect 14918 8072 14924 8084
rect 14369 8044 14924 8072
rect 14369 8041 14381 8044
rect 14323 8035 14381 8041
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 15746 8072 15752 8084
rect 15707 8044 15752 8072
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 15838 8032 15844 8084
rect 15896 8072 15902 8084
rect 16025 8075 16083 8081
rect 16025 8072 16037 8075
rect 15896 8044 16037 8072
rect 15896 8032 15902 8044
rect 16025 8041 16037 8044
rect 16071 8041 16083 8075
rect 16482 8072 16488 8084
rect 16443 8044 16488 8072
rect 16025 8035 16083 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 17218 8072 17224 8084
rect 17179 8044 17224 8072
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 17494 8072 17500 8084
rect 17455 8044 17500 8072
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 19981 8075 20039 8081
rect 19981 8041 19993 8075
rect 20027 8072 20039 8075
rect 21174 8072 21180 8084
rect 20027 8044 20944 8072
rect 21135 8044 21180 8072
rect 20027 8041 20039 8044
rect 19981 8035 20039 8041
rect 14093 8007 14151 8013
rect 14093 7973 14105 8007
rect 14139 8004 14151 8007
rect 14182 8004 14188 8016
rect 14139 7976 14188 8004
rect 14139 7973 14151 7976
rect 14093 7967 14151 7973
rect 14182 7964 14188 7976
rect 14240 8004 14246 8016
rect 15102 8004 15108 8016
rect 14240 7976 15108 8004
rect 14240 7964 14246 7976
rect 15102 7964 15108 7976
rect 15160 7964 15166 8016
rect 13078 7936 13084 7948
rect 13039 7908 13084 7936
rect 13078 7896 13084 7908
rect 13136 7896 13142 7948
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7936 15623 7939
rect 15856 7936 15884 8032
rect 15930 7964 15936 8016
rect 15988 8004 15994 8016
rect 15988 7976 16712 8004
rect 15988 7964 15994 7976
rect 15611 7908 15884 7936
rect 16485 7939 16543 7945
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 16485 7905 16497 7939
rect 16531 7936 16543 7939
rect 16574 7936 16580 7948
rect 16531 7908 16580 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 16684 7945 16712 7976
rect 18782 7964 18788 8016
rect 18840 7964 18846 8016
rect 20916 7948 20944 8044
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 21358 8072 21364 8084
rect 21319 8044 21364 8072
rect 21358 8032 21364 8044
rect 21416 8032 21422 8084
rect 26145 8075 26203 8081
rect 26145 8041 26157 8075
rect 26191 8072 26203 8075
rect 26418 8072 26424 8084
rect 26191 8044 26424 8072
rect 26191 8041 26203 8044
rect 26145 8035 26203 8041
rect 26418 8032 26424 8044
rect 26476 8072 26482 8084
rect 26697 8075 26755 8081
rect 26697 8072 26709 8075
rect 26476 8044 26709 8072
rect 26476 8032 26482 8044
rect 26697 8041 26709 8044
rect 26743 8041 26755 8075
rect 29362 8072 29368 8084
rect 29323 8044 29368 8072
rect 26697 8035 26755 8041
rect 29362 8032 29368 8044
rect 29420 8032 29426 8084
rect 29730 8072 29736 8084
rect 29691 8044 29736 8072
rect 29730 8032 29736 8044
rect 29788 8032 29794 8084
rect 34698 8072 34704 8084
rect 34659 8044 34704 8072
rect 34698 8032 34704 8044
rect 34756 8032 34762 8084
rect 35066 8072 35072 8084
rect 35027 8044 35072 8072
rect 35066 8032 35072 8044
rect 35124 8032 35130 8084
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7905 16727 7939
rect 16669 7899 16727 7905
rect 17037 7939 17095 7945
rect 17037 7905 17049 7939
rect 17083 7936 17095 7939
rect 17126 7936 17132 7948
rect 17083 7908 17132 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 17126 7896 17132 7908
rect 17184 7936 17190 7948
rect 17954 7936 17960 7948
rect 17184 7908 17960 7936
rect 17184 7896 17190 7908
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 19521 7939 19579 7945
rect 19521 7905 19533 7939
rect 19567 7936 19579 7939
rect 19610 7936 19616 7948
rect 19567 7908 19616 7936
rect 19567 7905 19579 7908
rect 19521 7899 19579 7905
rect 19610 7896 19616 7908
rect 19668 7896 19674 7948
rect 20898 7936 20904 7948
rect 20956 7945 20962 7948
rect 20956 7939 20994 7945
rect 20811 7908 20904 7936
rect 20898 7896 20904 7908
rect 20982 7905 20994 7939
rect 20956 7899 20994 7905
rect 20956 7896 20962 7899
rect 17678 7868 17684 7880
rect 17639 7840 17684 7868
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7868 18107 7871
rect 18506 7868 18512 7880
rect 18095 7840 18512 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 13170 7692 13176 7744
rect 13228 7732 13234 7744
rect 13541 7735 13599 7741
rect 13541 7732 13553 7735
rect 13228 7704 13553 7732
rect 13228 7692 13234 7704
rect 13541 7701 13553 7704
rect 13587 7701 13599 7735
rect 13541 7695 13599 7701
rect 1104 7642 48852 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 48852 7642
rect 1104 7568 48852 7590
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 13078 7528 13084 7540
rect 12299 7500 13084 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 13078 7488 13084 7500
rect 13136 7528 13142 7540
rect 15473 7531 15531 7537
rect 15473 7528 15485 7531
rect 13136 7500 15485 7528
rect 13136 7488 13142 7500
rect 15473 7497 15485 7500
rect 15519 7497 15531 7531
rect 15930 7528 15936 7540
rect 15891 7500 15936 7528
rect 15473 7491 15531 7497
rect 15930 7488 15936 7500
rect 15988 7488 15994 7540
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 16574 7528 16580 7540
rect 16347 7500 16580 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 16574 7488 16580 7500
rect 16632 7488 16638 7540
rect 20346 7528 20352 7540
rect 20307 7500 20352 7528
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 20898 7528 20904 7540
rect 20859 7500 20904 7528
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 13170 7392 13176 7404
rect 13131 7364 13176 7392
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7392 18475 7395
rect 18874 7392 18880 7404
rect 18463 7364 18880 7392
rect 18463 7361 18475 7364
rect 18417 7355 18475 7361
rect 18874 7352 18880 7364
rect 18932 7352 18938 7404
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7324 12771 7327
rect 13538 7324 13544 7336
rect 12759 7296 13544 7324
rect 12759 7293 12771 7296
rect 12713 7287 12771 7293
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 15013 7327 15071 7333
rect 15013 7293 15025 7327
rect 15059 7293 15071 7327
rect 15013 7287 15071 7293
rect 8570 7216 8576 7268
rect 8628 7256 8634 7268
rect 12989 7259 13047 7265
rect 12989 7256 13001 7259
rect 8628 7228 13001 7256
rect 8628 7216 8634 7228
rect 12989 7225 13001 7228
rect 13035 7225 13047 7259
rect 12989 7219 13047 7225
rect 13004 7188 13032 7219
rect 14642 7216 14648 7268
rect 14700 7216 14706 7268
rect 15028 7188 15056 7287
rect 17770 7284 17776 7336
rect 17828 7324 17834 7336
rect 17865 7327 17923 7333
rect 17865 7324 17877 7327
rect 17828 7296 17877 7324
rect 17828 7284 17834 7296
rect 17865 7293 17877 7296
rect 17911 7293 17923 7327
rect 18046 7324 18052 7336
rect 18007 7296 18052 7324
rect 17865 7287 17923 7293
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7293 19947 7327
rect 19889 7287 19947 7293
rect 17129 7259 17187 7265
rect 17129 7256 17141 7259
rect 15580 7228 17141 7256
rect 15580 7200 15608 7228
rect 17129 7225 17141 7228
rect 17175 7256 17187 7259
rect 17402 7256 17408 7268
rect 17175 7228 17408 7256
rect 17175 7225 17187 7228
rect 17129 7219 17187 7225
rect 17402 7216 17408 7228
rect 17460 7256 17466 7268
rect 17497 7259 17555 7265
rect 17497 7256 17509 7259
rect 17460 7228 17509 7256
rect 17460 7216 17466 7228
rect 17497 7225 17509 7228
rect 17543 7256 17555 7259
rect 17543 7228 18184 7256
rect 17543 7225 17555 7228
rect 17497 7219 17555 7225
rect 15562 7188 15568 7200
rect 13004 7160 15568 7188
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 16853 7191 16911 7197
rect 16853 7157 16865 7191
rect 16899 7188 16911 7191
rect 17034 7188 17040 7200
rect 16899 7160 17040 7188
rect 16899 7157 16911 7160
rect 16853 7151 16911 7157
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 17678 7188 17684 7200
rect 17591 7160 17684 7188
rect 17678 7148 17684 7160
rect 17736 7188 17742 7200
rect 18046 7188 18052 7200
rect 17736 7160 18052 7188
rect 17736 7148 17742 7160
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18156 7188 18184 7228
rect 18782 7216 18788 7268
rect 18840 7216 18846 7268
rect 19610 7216 19616 7268
rect 19668 7216 19674 7268
rect 19628 7188 19656 7216
rect 19904 7188 19932 7287
rect 18156 7160 19932 7188
rect 1104 7098 48852 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 48852 7098
rect 1104 7024 48852 7046
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 13228 6956 13553 6984
rect 13228 6944 13234 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13541 6947 13599 6953
rect 14277 6987 14335 6993
rect 14277 6953 14289 6987
rect 14323 6984 14335 6987
rect 15102 6984 15108 6996
rect 14323 6956 15108 6984
rect 14323 6953 14335 6956
rect 14277 6947 14335 6953
rect 13556 6780 13584 6947
rect 15102 6944 15108 6956
rect 15160 6944 15166 6996
rect 17862 6984 17868 6996
rect 17823 6956 17868 6984
rect 17862 6944 17868 6956
rect 17920 6944 17926 6996
rect 18506 6984 18512 6996
rect 18467 6956 18512 6984
rect 18506 6944 18512 6956
rect 18564 6944 18570 6996
rect 18874 6984 18880 6996
rect 18835 6956 18880 6984
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 17034 6876 17040 6928
rect 17092 6916 17098 6928
rect 18233 6919 18291 6925
rect 18233 6916 18245 6919
rect 17092 6888 18245 6916
rect 17092 6876 17098 6888
rect 18233 6885 18245 6888
rect 18279 6916 18291 6919
rect 18782 6916 18788 6928
rect 18279 6888 18788 6916
rect 18279 6885 18291 6888
rect 18233 6879 18291 6885
rect 18782 6876 18788 6888
rect 18840 6876 18846 6928
rect 13722 6848 13728 6860
rect 13683 6820 13728 6848
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 15010 6808 15016 6860
rect 15068 6848 15074 6860
rect 15930 6848 15936 6860
rect 15068 6820 15936 6848
rect 15068 6808 15074 6820
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 17402 6848 17408 6860
rect 17363 6820 17408 6848
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 15194 6780 15200 6792
rect 13556 6752 15200 6780
rect 15194 6740 15200 6752
rect 15252 6780 15258 6792
rect 15565 6783 15623 6789
rect 15565 6780 15577 6783
rect 15252 6752 15577 6780
rect 15252 6740 15258 6752
rect 15565 6749 15577 6752
rect 15611 6749 15623 6783
rect 15565 6743 15623 6749
rect 14642 6712 14648 6724
rect 13188 6684 14648 6712
rect 13188 6656 13216 6684
rect 14642 6672 14648 6684
rect 14700 6672 14706 6724
rect 13170 6644 13176 6656
rect 13131 6616 13176 6644
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 1104 6554 48852 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 48852 6554
rect 1104 6480 48852 6502
rect 15194 6440 15200 6452
rect 15155 6412 15200 6440
rect 15194 6400 15200 6412
rect 15252 6400 15258 6452
rect 15562 6440 15568 6452
rect 15523 6412 15568 6440
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16301 6443 16359 6449
rect 16301 6440 16313 6443
rect 15988 6412 16313 6440
rect 15988 6400 15994 6412
rect 16301 6409 16313 6412
rect 16347 6409 16359 6443
rect 17126 6440 17132 6452
rect 17087 6412 17132 6440
rect 16301 6403 16359 6409
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 18046 6400 18052 6452
rect 18104 6440 18110 6452
rect 18325 6443 18383 6449
rect 18325 6440 18337 6443
rect 18104 6412 18337 6440
rect 18104 6400 18110 6412
rect 18325 6409 18337 6412
rect 18371 6440 18383 6443
rect 18601 6443 18659 6449
rect 18601 6440 18613 6443
rect 18371 6412 18613 6440
rect 18371 6409 18383 6412
rect 18325 6403 18383 6409
rect 18601 6409 18613 6412
rect 18647 6409 18659 6443
rect 18601 6403 18659 6409
rect 13633 6375 13691 6381
rect 13633 6341 13645 6375
rect 13679 6372 13691 6375
rect 13722 6372 13728 6384
rect 13679 6344 13728 6372
rect 13679 6341 13691 6344
rect 13633 6335 13691 6341
rect 13722 6332 13728 6344
rect 13780 6372 13786 6384
rect 17681 6375 17739 6381
rect 17681 6372 17693 6375
rect 13780 6344 17693 6372
rect 13780 6332 13786 6344
rect 17681 6341 17693 6344
rect 17727 6372 17739 6375
rect 17770 6372 17776 6384
rect 17727 6344 17776 6372
rect 17727 6341 17739 6344
rect 17681 6335 17739 6341
rect 17770 6332 17776 6344
rect 17828 6332 17834 6384
rect 14642 6264 14648 6316
rect 14700 6304 14706 6316
rect 16025 6307 16083 6313
rect 16025 6304 16037 6307
rect 14700 6276 16037 6304
rect 14700 6264 14706 6276
rect 16025 6273 16037 6276
rect 16071 6304 16083 6307
rect 17034 6304 17040 6316
rect 16071 6276 17040 6304
rect 16071 6273 16083 6276
rect 16025 6267 16083 6273
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 1104 6010 48852 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 48852 6010
rect 1104 5936 48852 5958
rect 1104 5466 48852 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 48852 5466
rect 1104 5392 48852 5414
rect 1104 4922 48852 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 48852 4922
rect 1104 4848 48852 4870
rect 1104 4378 48852 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 48852 4378
rect 1104 4304 48852 4326
rect 1104 3834 48852 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 48852 3834
rect 1104 3760 48852 3782
rect 1104 3290 48852 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 48852 3290
rect 1104 3216 48852 3238
rect 1104 2746 48852 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 48852 2746
rect 1104 2672 48852 2694
rect 1104 2202 48852 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 48852 2202
rect 1104 2128 48852 2150
rect 28534 76 28540 128
rect 28592 116 28598 128
rect 30466 116 30472 128
rect 28592 88 30472 116
rect 28592 76 28598 88
rect 30466 76 30472 88
rect 30524 76 30530 128
<< via1 >>
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 30748 44319 30800 44328
rect 30748 44285 30766 44319
rect 30766 44285 30800 44319
rect 38016 44344 38068 44396
rect 30748 44276 30800 44285
rect 31852 44276 31904 44328
rect 31024 44140 31076 44192
rect 34796 44140 34848 44192
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 31024 43936 31076 43988
rect 32588 43936 32640 43988
rect 33692 43868 33744 43920
rect 23112 43843 23164 43852
rect 23112 43809 23121 43843
rect 23121 43809 23155 43843
rect 23155 43809 23164 43843
rect 23112 43800 23164 43809
rect 25044 43800 25096 43852
rect 30840 43800 30892 43852
rect 33324 43775 33376 43784
rect 33324 43741 33333 43775
rect 33333 43741 33367 43775
rect 33367 43741 33376 43775
rect 33324 43732 33376 43741
rect 31208 43664 31260 43716
rect 33508 43664 33560 43716
rect 23572 43596 23624 43648
rect 23848 43596 23900 43648
rect 24032 43639 24084 43648
rect 24032 43605 24041 43639
rect 24041 43605 24075 43639
rect 24075 43605 24084 43639
rect 24032 43596 24084 43605
rect 25412 43596 25464 43648
rect 25596 43639 25648 43648
rect 25596 43605 25605 43639
rect 25605 43605 25639 43639
rect 25639 43605 25648 43639
rect 25596 43596 25648 43605
rect 30380 43596 30432 43648
rect 31024 43639 31076 43648
rect 31024 43605 31033 43639
rect 31033 43605 31067 43639
rect 31067 43605 31076 43639
rect 31024 43596 31076 43605
rect 31300 43639 31352 43648
rect 31300 43605 31309 43639
rect 31309 43605 31343 43639
rect 31343 43605 31352 43639
rect 31300 43596 31352 43605
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 22376 43392 22428 43444
rect 23112 43435 23164 43444
rect 23112 43401 23121 43435
rect 23121 43401 23155 43435
rect 23155 43401 23164 43435
rect 23112 43392 23164 43401
rect 25044 43435 25096 43444
rect 25044 43401 25053 43435
rect 25053 43401 25087 43435
rect 25087 43401 25096 43435
rect 25044 43392 25096 43401
rect 23204 43324 23256 43376
rect 26608 43324 26660 43376
rect 23480 43256 23532 43308
rect 24032 43256 24084 43308
rect 24216 43256 24268 43308
rect 21640 43052 21692 43104
rect 27528 43231 27580 43240
rect 27528 43197 27537 43231
rect 27537 43197 27571 43231
rect 27571 43197 27580 43231
rect 27528 43188 27580 43197
rect 27988 43231 28040 43240
rect 27988 43197 27997 43231
rect 27997 43197 28031 43231
rect 28031 43197 28040 43231
rect 27988 43188 28040 43197
rect 30472 43392 30524 43444
rect 30840 43435 30892 43444
rect 30840 43401 30849 43435
rect 30849 43401 30883 43435
rect 30883 43401 30892 43435
rect 30840 43392 30892 43401
rect 30564 43324 30616 43376
rect 33324 43392 33376 43444
rect 33876 43435 33928 43444
rect 33876 43401 33885 43435
rect 33885 43401 33919 43435
rect 33919 43401 33928 43435
rect 33876 43392 33928 43401
rect 31300 43256 31352 43308
rect 32588 43299 32640 43308
rect 32588 43265 32597 43299
rect 32597 43265 32631 43299
rect 32631 43265 32640 43299
rect 32588 43256 32640 43265
rect 37096 43324 37148 43376
rect 23848 43163 23900 43172
rect 23848 43129 23857 43163
rect 23857 43129 23891 43163
rect 23891 43129 23900 43163
rect 23848 43120 23900 43129
rect 25504 43163 25556 43172
rect 25504 43129 25513 43163
rect 25513 43129 25547 43163
rect 25547 43129 25556 43163
rect 25504 43120 25556 43129
rect 25596 43163 25648 43172
rect 25596 43129 25605 43163
rect 25605 43129 25639 43163
rect 25639 43129 25648 43163
rect 25596 43120 25648 43129
rect 31024 43120 31076 43172
rect 31668 43163 31720 43172
rect 23020 43052 23072 43104
rect 27620 43095 27672 43104
rect 27620 43061 27629 43095
rect 27629 43061 27663 43095
rect 27663 43061 27672 43095
rect 27620 43052 27672 43061
rect 31668 43129 31677 43163
rect 31677 43129 31711 43163
rect 31711 43129 31720 43163
rect 31668 43120 31720 43129
rect 33692 43052 33744 43104
rect 34244 43052 34296 43104
rect 35440 43095 35492 43104
rect 35440 43061 35449 43095
rect 35449 43061 35483 43095
rect 35483 43061 35492 43095
rect 35440 43052 35492 43061
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 27988 42848 28040 42900
rect 23572 42823 23624 42832
rect 23572 42789 23581 42823
rect 23581 42789 23615 42823
rect 23615 42789 23624 42823
rect 23572 42780 23624 42789
rect 23664 42823 23716 42832
rect 23664 42789 23673 42823
rect 23673 42789 23707 42823
rect 23707 42789 23716 42823
rect 24216 42823 24268 42832
rect 23664 42780 23716 42789
rect 24216 42789 24225 42823
rect 24225 42789 24259 42823
rect 24259 42789 24268 42823
rect 24216 42780 24268 42789
rect 25412 42780 25464 42832
rect 26240 42780 26292 42832
rect 26700 42823 26752 42832
rect 26700 42789 26709 42823
rect 26709 42789 26743 42823
rect 26743 42789 26752 42823
rect 26700 42780 26752 42789
rect 30380 42780 30432 42832
rect 31024 42780 31076 42832
rect 31208 42823 31260 42832
rect 31208 42789 31217 42823
rect 31217 42789 31251 42823
rect 31251 42789 31260 42823
rect 31208 42780 31260 42789
rect 33692 42848 33744 42900
rect 34796 42780 34848 42832
rect 35716 42780 35768 42832
rect 23112 42712 23164 42764
rect 25320 42712 25372 42764
rect 27528 42712 27580 42764
rect 29184 42755 29236 42764
rect 29184 42721 29193 42755
rect 29193 42721 29227 42755
rect 29227 42721 29236 42755
rect 29184 42712 29236 42721
rect 29552 42712 29604 42764
rect 32496 42712 32548 42764
rect 37096 42712 37148 42764
rect 38200 42712 38252 42764
rect 39856 42755 39908 42764
rect 39856 42721 39865 42755
rect 39865 42721 39899 42755
rect 39899 42721 39908 42755
rect 39856 42712 39908 42721
rect 24400 42644 24452 42696
rect 29644 42687 29696 42696
rect 29644 42653 29653 42687
rect 29653 42653 29687 42687
rect 29687 42653 29696 42687
rect 29644 42644 29696 42653
rect 34244 42644 34296 42696
rect 35532 42687 35584 42696
rect 35532 42653 35541 42687
rect 35541 42653 35575 42687
rect 35575 42653 35584 42687
rect 35532 42644 35584 42653
rect 31668 42576 31720 42628
rect 34060 42619 34112 42628
rect 34060 42585 34069 42619
rect 34069 42585 34103 42619
rect 34103 42585 34112 42619
rect 34060 42576 34112 42585
rect 35440 42576 35492 42628
rect 39764 42576 39816 42628
rect 41420 42576 41472 42628
rect 22100 42508 22152 42560
rect 23756 42508 23808 42560
rect 25596 42508 25648 42560
rect 34704 42508 34756 42560
rect 38476 42508 38528 42560
rect 38568 42551 38620 42560
rect 38568 42517 38577 42551
rect 38577 42517 38611 42551
rect 38611 42517 38620 42551
rect 38568 42508 38620 42517
rect 40316 42508 40368 42560
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 18512 42304 18564 42356
rect 19340 42304 19392 42356
rect 25320 42347 25372 42356
rect 25320 42313 25329 42347
rect 25329 42313 25363 42347
rect 25363 42313 25372 42347
rect 25320 42304 25372 42313
rect 21364 41964 21416 42016
rect 23664 42236 23716 42288
rect 26700 42236 26752 42288
rect 22100 42211 22152 42220
rect 22100 42177 22109 42211
rect 22109 42177 22143 42211
rect 22143 42177 22152 42211
rect 22100 42168 22152 42177
rect 23020 42168 23072 42220
rect 23756 42211 23808 42220
rect 23756 42177 23765 42211
rect 23765 42177 23799 42211
rect 23799 42177 23808 42211
rect 23756 42168 23808 42177
rect 24400 42211 24452 42220
rect 24400 42177 24409 42211
rect 24409 42177 24443 42211
rect 24443 42177 24452 42211
rect 24400 42168 24452 42177
rect 25596 42211 25648 42220
rect 25596 42177 25605 42211
rect 25605 42177 25639 42211
rect 25639 42177 25648 42211
rect 25596 42168 25648 42177
rect 27620 42168 27672 42220
rect 29644 42168 29696 42220
rect 29460 42100 29512 42152
rect 31024 42347 31076 42356
rect 31024 42313 31033 42347
rect 31033 42313 31067 42347
rect 31067 42313 31076 42347
rect 31024 42304 31076 42313
rect 33876 42304 33928 42356
rect 34244 42347 34296 42356
rect 34244 42313 34253 42347
rect 34253 42313 34287 42347
rect 34287 42313 34296 42347
rect 34244 42304 34296 42313
rect 34796 42304 34848 42356
rect 35716 42347 35768 42356
rect 35716 42313 35725 42347
rect 35725 42313 35759 42347
rect 35759 42313 35768 42347
rect 35716 42304 35768 42313
rect 39856 42347 39908 42356
rect 30380 42236 30432 42288
rect 30288 42168 30340 42220
rect 22744 42075 22796 42084
rect 22744 42041 22753 42075
rect 22753 42041 22787 42075
rect 22787 42041 22796 42075
rect 22744 42032 22796 42041
rect 23204 42032 23256 42084
rect 25688 42075 25740 42084
rect 22652 41964 22704 42016
rect 23112 42007 23164 42016
rect 23112 41973 23121 42007
rect 23121 41973 23155 42007
rect 23155 41973 23164 42007
rect 23112 41964 23164 41973
rect 23756 41964 23808 42016
rect 25688 42041 25697 42075
rect 25697 42041 25731 42075
rect 25731 42041 25740 42075
rect 25688 42032 25740 42041
rect 26608 42032 26660 42084
rect 26700 41964 26752 42016
rect 27252 42007 27304 42016
rect 27252 41973 27261 42007
rect 27261 41973 27295 42007
rect 27295 41973 27304 42007
rect 29184 42032 29236 42084
rect 30748 42100 30800 42152
rect 33692 42236 33744 42288
rect 35624 42236 35676 42288
rect 39856 42313 39865 42347
rect 39865 42313 39899 42347
rect 39899 42313 39908 42347
rect 39856 42304 39908 42313
rect 35900 42236 35952 42288
rect 27252 41964 27304 41973
rect 29460 41964 29512 42016
rect 32036 41964 32088 42016
rect 32496 42007 32548 42016
rect 32496 41973 32505 42007
rect 32505 41973 32539 42007
rect 32539 41973 32548 42007
rect 32496 41964 32548 41973
rect 35256 42168 35308 42220
rect 35440 42100 35492 42152
rect 35808 42100 35860 42152
rect 38476 42211 38528 42220
rect 38476 42177 38485 42211
rect 38485 42177 38519 42211
rect 38519 42177 38528 42211
rect 38476 42168 38528 42177
rect 36176 42100 36228 42152
rect 33692 42032 33744 42084
rect 38292 42032 38344 42084
rect 38568 42075 38620 42084
rect 38568 42041 38577 42075
rect 38577 42041 38611 42075
rect 38611 42041 38620 42075
rect 38568 42032 38620 42041
rect 40132 42032 40184 42084
rect 32956 41964 33008 42016
rect 33968 41964 34020 42016
rect 35440 42007 35492 42016
rect 35440 41973 35449 42007
rect 35449 41973 35483 42007
rect 35483 41973 35492 42007
rect 35440 41964 35492 41973
rect 37740 41964 37792 42016
rect 38200 42007 38252 42016
rect 38200 41973 38209 42007
rect 38209 41973 38243 42007
rect 38243 41973 38252 42007
rect 38200 41964 38252 41973
rect 40776 41964 40828 42016
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 22100 41803 22152 41812
rect 22100 41769 22109 41803
rect 22109 41769 22143 41803
rect 22143 41769 22152 41803
rect 22100 41760 22152 41769
rect 23480 41760 23532 41812
rect 23572 41760 23624 41812
rect 25504 41760 25556 41812
rect 25688 41803 25740 41812
rect 25688 41769 25697 41803
rect 25697 41769 25731 41803
rect 25731 41769 25740 41803
rect 25688 41760 25740 41769
rect 26240 41803 26292 41812
rect 26240 41769 26249 41803
rect 26249 41769 26283 41803
rect 26283 41769 26292 41803
rect 26240 41760 26292 41769
rect 29644 41760 29696 41812
rect 34704 41760 34756 41812
rect 21364 41692 21416 41744
rect 23296 41735 23348 41744
rect 23296 41701 23305 41735
rect 23305 41701 23339 41735
rect 23339 41701 23348 41735
rect 23296 41692 23348 41701
rect 23664 41692 23716 41744
rect 24400 41692 24452 41744
rect 26700 41735 26752 41744
rect 26700 41701 26709 41735
rect 26709 41701 26743 41735
rect 26743 41701 26752 41735
rect 26700 41692 26752 41701
rect 30656 41735 30708 41744
rect 30656 41701 30665 41735
rect 30665 41701 30699 41735
rect 30699 41701 30708 41735
rect 30656 41692 30708 41701
rect 33692 41735 33744 41744
rect 33692 41701 33701 41735
rect 33701 41701 33735 41735
rect 33735 41701 33744 41735
rect 33692 41692 33744 41701
rect 34612 41692 34664 41744
rect 35256 41735 35308 41744
rect 35256 41701 35265 41735
rect 35265 41701 35299 41735
rect 35299 41701 35308 41735
rect 35256 41692 35308 41701
rect 38568 41692 38620 41744
rect 40316 41735 40368 41744
rect 40316 41701 40325 41735
rect 40325 41701 40359 41735
rect 40359 41701 40368 41735
rect 40316 41692 40368 41701
rect 40408 41735 40460 41744
rect 40408 41701 40417 41735
rect 40417 41701 40451 41735
rect 40451 41701 40460 41735
rect 42248 41735 42300 41744
rect 40408 41692 40460 41701
rect 42248 41701 42257 41735
rect 42257 41701 42291 41735
rect 42291 41701 42300 41735
rect 42248 41692 42300 41701
rect 22100 41624 22152 41676
rect 24768 41624 24820 41676
rect 29276 41624 29328 41676
rect 26608 41599 26660 41608
rect 26608 41565 26617 41599
rect 26617 41565 26651 41599
rect 26651 41565 26660 41599
rect 26608 41556 26660 41565
rect 26884 41599 26936 41608
rect 26884 41565 26893 41599
rect 26893 41565 26927 41599
rect 26927 41565 26936 41599
rect 26884 41556 26936 41565
rect 29552 41624 29604 41676
rect 32312 41624 32364 41676
rect 42064 41624 42116 41676
rect 46940 41624 46992 41676
rect 30104 41556 30156 41608
rect 30564 41599 30616 41608
rect 30564 41565 30573 41599
rect 30573 41565 30607 41599
rect 30607 41565 30616 41599
rect 30564 41556 30616 41565
rect 32220 41556 32272 41608
rect 34060 41599 34112 41608
rect 34060 41565 34069 41599
rect 34069 41565 34103 41599
rect 34103 41565 34112 41599
rect 34060 41556 34112 41565
rect 35532 41599 35584 41608
rect 35532 41565 35541 41599
rect 35541 41565 35575 41599
rect 35575 41565 35584 41599
rect 35532 41556 35584 41565
rect 38568 41599 38620 41608
rect 38568 41565 38577 41599
rect 38577 41565 38611 41599
rect 38611 41565 38620 41599
rect 38568 41556 38620 41565
rect 40132 41556 40184 41608
rect 30840 41488 30892 41540
rect 38660 41488 38712 41540
rect 40868 41488 40920 41540
rect 33416 41420 33468 41472
rect 36636 41463 36688 41472
rect 36636 41429 36645 41463
rect 36645 41429 36679 41463
rect 36679 41429 36688 41463
rect 36636 41420 36688 41429
rect 42156 41420 42208 41472
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 23480 41216 23532 41268
rect 23664 41216 23716 41268
rect 23848 41216 23900 41268
rect 24768 41259 24820 41268
rect 24768 41225 24777 41259
rect 24777 41225 24811 41259
rect 24811 41225 24820 41259
rect 24768 41216 24820 41225
rect 26608 41216 26660 41268
rect 29460 41216 29512 41268
rect 19248 41148 19300 41200
rect 26700 41148 26752 41200
rect 23848 41080 23900 41132
rect 19064 41012 19116 41064
rect 22468 40944 22520 40996
rect 22100 40876 22152 40928
rect 23112 41012 23164 41064
rect 23204 41012 23256 41064
rect 23940 40944 23992 40996
rect 27344 41080 27396 41132
rect 30104 41123 30156 41132
rect 30104 41089 30113 41123
rect 30113 41089 30147 41123
rect 30147 41089 30156 41123
rect 30104 41080 30156 41089
rect 25228 41055 25280 41064
rect 25228 41021 25237 41055
rect 25237 41021 25271 41055
rect 25271 41021 25280 41055
rect 25228 41012 25280 41021
rect 30656 41216 30708 41268
rect 33692 41216 33744 41268
rect 37740 41216 37792 41268
rect 30564 41148 30616 41200
rect 31668 41080 31720 41132
rect 31944 41123 31996 41132
rect 31944 41089 31953 41123
rect 31953 41089 31987 41123
rect 31987 41089 31996 41123
rect 31944 41080 31996 41089
rect 32220 41123 32272 41132
rect 32220 41089 32229 41123
rect 32229 41089 32263 41123
rect 32263 41089 32272 41123
rect 32220 41080 32272 41089
rect 34704 41080 34756 41132
rect 35532 41148 35584 41200
rect 38568 41080 38620 41132
rect 40776 41080 40828 41132
rect 40868 41123 40920 41132
rect 40868 41089 40877 41123
rect 40877 41089 40911 41123
rect 40911 41089 40920 41123
rect 42432 41123 42484 41132
rect 40868 41080 40920 41089
rect 42432 41089 42441 41123
rect 42441 41089 42475 41123
rect 42475 41089 42484 41123
rect 42432 41080 42484 41089
rect 32772 41012 32824 41064
rect 36636 41055 36688 41064
rect 36636 41021 36645 41055
rect 36645 41021 36679 41055
rect 36679 41021 36688 41055
rect 36636 41012 36688 41021
rect 27252 40944 27304 40996
rect 30472 40944 30524 40996
rect 24584 40876 24636 40928
rect 25688 40876 25740 40928
rect 29276 40876 29328 40928
rect 29552 40919 29604 40928
rect 29552 40885 29561 40919
rect 29561 40885 29595 40919
rect 29595 40885 29604 40919
rect 29552 40876 29604 40885
rect 31668 40919 31720 40928
rect 31668 40885 31677 40919
rect 31677 40885 31711 40919
rect 31711 40885 31720 40919
rect 33692 40944 33744 40996
rect 31668 40876 31720 40885
rect 32312 40876 32364 40928
rect 33324 40876 33376 40928
rect 34612 40876 34664 40928
rect 36544 40919 36596 40928
rect 36544 40885 36553 40919
rect 36553 40885 36587 40919
rect 36587 40885 36596 40919
rect 38476 40944 38528 40996
rect 39120 40987 39172 40996
rect 39120 40953 39129 40987
rect 39129 40953 39163 40987
rect 39163 40953 39172 40987
rect 39120 40944 39172 40953
rect 39948 40919 40000 40928
rect 36544 40876 36596 40885
rect 39948 40885 39957 40919
rect 39957 40885 39991 40919
rect 39991 40885 40000 40919
rect 39948 40876 40000 40885
rect 40408 40876 40460 40928
rect 41696 40944 41748 40996
rect 42064 40876 42116 40928
rect 42248 40987 42300 40996
rect 42248 40953 42257 40987
rect 42257 40953 42291 40987
rect 42291 40953 42300 40987
rect 42248 40944 42300 40953
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 23296 40672 23348 40724
rect 25228 40672 25280 40724
rect 30564 40672 30616 40724
rect 31668 40672 31720 40724
rect 31944 40715 31996 40724
rect 31944 40681 31953 40715
rect 31953 40681 31987 40715
rect 31987 40681 31996 40715
rect 31944 40672 31996 40681
rect 32036 40672 32088 40724
rect 22928 40604 22980 40656
rect 24492 40604 24544 40656
rect 30472 40604 30524 40656
rect 33416 40647 33468 40656
rect 33416 40613 33425 40647
rect 33425 40613 33459 40647
rect 33459 40613 33468 40647
rect 33416 40604 33468 40613
rect 33692 40604 33744 40656
rect 34060 40647 34112 40656
rect 34060 40613 34069 40647
rect 34069 40613 34103 40647
rect 34103 40613 34112 40647
rect 34060 40604 34112 40613
rect 21180 40536 21232 40588
rect 27620 40579 27672 40588
rect 27620 40545 27629 40579
rect 27629 40545 27663 40579
rect 27663 40545 27672 40579
rect 27620 40536 27672 40545
rect 27988 40536 28040 40588
rect 28724 40536 28776 40588
rect 32128 40579 32180 40588
rect 22468 40511 22520 40520
rect 22468 40477 22477 40511
rect 22477 40477 22511 40511
rect 22511 40477 22520 40511
rect 22468 40468 22520 40477
rect 22744 40511 22796 40520
rect 22744 40477 22753 40511
rect 22753 40477 22787 40511
rect 22787 40477 22796 40511
rect 22744 40468 22796 40477
rect 23296 40400 23348 40452
rect 24400 40511 24452 40520
rect 24400 40477 24409 40511
rect 24409 40477 24443 40511
rect 24443 40477 24452 40511
rect 24400 40468 24452 40477
rect 32128 40545 32137 40579
rect 32137 40545 32171 40579
rect 32171 40545 32180 40579
rect 32128 40536 32180 40545
rect 34796 40536 34848 40588
rect 35256 40672 35308 40724
rect 38568 40672 38620 40724
rect 40316 40672 40368 40724
rect 40776 40715 40828 40724
rect 40776 40681 40785 40715
rect 40785 40681 40819 40715
rect 40819 40681 40828 40715
rect 40776 40672 40828 40681
rect 42156 40672 42208 40724
rect 43260 40672 43312 40724
rect 36636 40647 36688 40656
rect 36636 40613 36645 40647
rect 36645 40613 36679 40647
rect 36679 40613 36688 40647
rect 36636 40604 36688 40613
rect 41696 40604 41748 40656
rect 41788 40647 41840 40656
rect 41788 40613 41797 40647
rect 41797 40613 41831 40647
rect 41831 40613 41840 40647
rect 41788 40604 41840 40613
rect 42432 40604 42484 40656
rect 36268 40536 36320 40588
rect 30012 40511 30064 40520
rect 30012 40477 30021 40511
rect 30021 40477 30055 40511
rect 30055 40477 30064 40511
rect 30012 40468 30064 40477
rect 35716 40468 35768 40520
rect 38016 40536 38068 40588
rect 38476 40536 38528 40588
rect 39764 40536 39816 40588
rect 29276 40400 29328 40452
rect 33140 40400 33192 40452
rect 41604 40400 41656 40452
rect 27344 40332 27396 40384
rect 29552 40375 29604 40384
rect 29552 40341 29561 40375
rect 29561 40341 29595 40375
rect 29595 40341 29604 40375
rect 29552 40332 29604 40341
rect 31300 40332 31352 40384
rect 33692 40332 33744 40384
rect 38752 40332 38804 40384
rect 41696 40332 41748 40384
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 23296 40128 23348 40180
rect 24400 40128 24452 40180
rect 32128 40171 32180 40180
rect 23572 40060 23624 40112
rect 32128 40137 32137 40171
rect 32137 40137 32171 40171
rect 32171 40137 32180 40171
rect 32128 40128 32180 40137
rect 34520 40128 34572 40180
rect 34796 40128 34848 40180
rect 36268 40171 36320 40180
rect 36268 40137 36277 40171
rect 36277 40137 36311 40171
rect 36311 40137 36320 40171
rect 36268 40128 36320 40137
rect 38016 40128 38068 40180
rect 39120 40128 39172 40180
rect 42432 40128 42484 40180
rect 26792 40060 26844 40112
rect 25780 40035 25832 40044
rect 25780 40001 25789 40035
rect 25789 40001 25823 40035
rect 25823 40001 25832 40035
rect 25780 39992 25832 40001
rect 23020 39924 23072 39976
rect 29276 39992 29328 40044
rect 30012 40035 30064 40044
rect 30012 40001 30021 40035
rect 30021 40001 30055 40035
rect 30055 40001 30064 40035
rect 30012 39992 30064 40001
rect 27988 39924 28040 39976
rect 22560 39856 22612 39908
rect 12808 39788 12860 39840
rect 12992 39831 13044 39840
rect 12992 39797 13001 39831
rect 13001 39797 13035 39831
rect 13035 39797 13044 39831
rect 12992 39788 13044 39797
rect 21180 39788 21232 39840
rect 22284 39831 22336 39840
rect 22284 39797 22293 39831
rect 22293 39797 22327 39831
rect 22327 39797 22336 39831
rect 22284 39788 22336 39797
rect 22928 39788 22980 39840
rect 23664 39788 23716 39840
rect 24492 39831 24544 39840
rect 24492 39797 24501 39831
rect 24501 39797 24535 39831
rect 24535 39797 24544 39831
rect 24492 39788 24544 39797
rect 25688 39856 25740 39908
rect 27620 39856 27672 39908
rect 29552 39924 29604 39976
rect 33324 40035 33376 40044
rect 33324 40001 33333 40035
rect 33333 40001 33367 40035
rect 33367 40001 33376 40035
rect 33324 39992 33376 40001
rect 33508 39992 33560 40044
rect 35808 39992 35860 40044
rect 30840 39967 30892 39976
rect 30840 39933 30849 39967
rect 30849 39933 30883 39967
rect 30883 39933 30892 39967
rect 30840 39924 30892 39933
rect 31300 39967 31352 39976
rect 31300 39933 31309 39967
rect 31309 39933 31343 39967
rect 31343 39933 31352 39967
rect 31300 39924 31352 39933
rect 35256 39967 35308 39976
rect 35256 39933 35265 39967
rect 35265 39933 35299 39967
rect 35299 39933 35308 39967
rect 35256 39924 35308 39933
rect 35716 39967 35768 39976
rect 35716 39933 35725 39967
rect 35725 39933 35759 39967
rect 35759 39933 35768 39967
rect 35716 39924 35768 39933
rect 36912 39924 36964 39976
rect 30380 39856 30432 39908
rect 31576 39899 31628 39908
rect 31576 39865 31585 39899
rect 31585 39865 31619 39899
rect 31619 39865 31628 39899
rect 31576 39856 31628 39865
rect 33048 39856 33100 39908
rect 33600 39856 33652 39908
rect 27344 39831 27396 39840
rect 27344 39797 27353 39831
rect 27353 39797 27387 39831
rect 27387 39797 27396 39831
rect 27344 39788 27396 39797
rect 28724 39831 28776 39840
rect 28724 39797 28733 39831
rect 28733 39797 28767 39831
rect 28767 39797 28776 39831
rect 28724 39788 28776 39797
rect 29460 39788 29512 39840
rect 36544 39788 36596 39840
rect 37004 39788 37056 39840
rect 37740 39831 37792 39840
rect 37740 39797 37749 39831
rect 37749 39797 37783 39831
rect 37783 39797 37792 39831
rect 37740 39788 37792 39797
rect 39764 40060 39816 40112
rect 41328 40060 41380 40112
rect 40868 39992 40920 40044
rect 43260 40035 43312 40044
rect 43260 40001 43269 40035
rect 43269 40001 43303 40035
rect 43303 40001 43312 40035
rect 43260 39992 43312 40001
rect 38752 39899 38804 39908
rect 38752 39865 38761 39899
rect 38761 39865 38795 39899
rect 38795 39865 38804 39899
rect 39304 39899 39356 39908
rect 38752 39856 38804 39865
rect 39304 39865 39313 39899
rect 39313 39865 39347 39899
rect 39347 39865 39356 39899
rect 39304 39856 39356 39865
rect 41144 39924 41196 39976
rect 41696 39899 41748 39908
rect 41696 39865 41705 39899
rect 41705 39865 41739 39899
rect 41739 39865 41748 39899
rect 41696 39856 41748 39865
rect 41788 39899 41840 39908
rect 41788 39865 41797 39899
rect 41797 39865 41831 39899
rect 41831 39865 41840 39899
rect 43076 39899 43128 39908
rect 41788 39856 41840 39865
rect 43076 39865 43085 39899
rect 43085 39865 43119 39899
rect 43119 39865 43128 39899
rect 43076 39856 43128 39865
rect 40960 39788 41012 39840
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 22192 39627 22244 39636
rect 22192 39593 22201 39627
rect 22201 39593 22235 39627
rect 22235 39593 22244 39627
rect 22192 39584 22244 39593
rect 22468 39584 22520 39636
rect 27988 39584 28040 39636
rect 28172 39627 28224 39636
rect 28172 39593 28181 39627
rect 28181 39593 28215 39627
rect 28215 39593 28224 39627
rect 28172 39584 28224 39593
rect 30012 39627 30064 39636
rect 30012 39593 30021 39627
rect 30021 39593 30055 39627
rect 30055 39593 30064 39627
rect 30012 39584 30064 39593
rect 32404 39584 32456 39636
rect 33048 39627 33100 39636
rect 33048 39593 33057 39627
rect 33057 39593 33091 39627
rect 33091 39593 33100 39627
rect 33048 39584 33100 39593
rect 33324 39584 33376 39636
rect 36912 39627 36964 39636
rect 36912 39593 36921 39627
rect 36921 39593 36955 39627
rect 36955 39593 36964 39627
rect 36912 39584 36964 39593
rect 41604 39627 41656 39636
rect 41604 39593 41613 39627
rect 41613 39593 41647 39627
rect 41647 39593 41656 39627
rect 41604 39584 41656 39593
rect 22928 39516 22980 39568
rect 24492 39516 24544 39568
rect 26700 39559 26752 39568
rect 26700 39525 26709 39559
rect 26709 39525 26743 39559
rect 26743 39525 26752 39559
rect 26700 39516 26752 39525
rect 30656 39559 30708 39568
rect 11980 39491 12032 39500
rect 11980 39457 11989 39491
rect 11989 39457 12023 39491
rect 12023 39457 12032 39491
rect 11980 39448 12032 39457
rect 14832 39448 14884 39500
rect 16120 39448 16172 39500
rect 25136 39491 25188 39500
rect 25136 39457 25145 39491
rect 25145 39457 25179 39491
rect 25179 39457 25188 39491
rect 25136 39448 25188 39457
rect 28356 39491 28408 39500
rect 28356 39457 28365 39491
rect 28365 39457 28399 39491
rect 28399 39457 28408 39491
rect 28356 39448 28408 39457
rect 30656 39525 30665 39559
rect 30665 39525 30699 39559
rect 30699 39525 30708 39559
rect 30656 39516 30708 39525
rect 33416 39559 33468 39568
rect 33416 39525 33425 39559
rect 33425 39525 33459 39559
rect 33459 39525 33468 39559
rect 33416 39516 33468 39525
rect 33968 39559 34020 39568
rect 33968 39525 33977 39559
rect 33977 39525 34011 39559
rect 34011 39525 34020 39559
rect 33968 39516 34020 39525
rect 34612 39516 34664 39568
rect 37740 39516 37792 39568
rect 38568 39516 38620 39568
rect 40132 39516 40184 39568
rect 40960 39516 41012 39568
rect 41512 39516 41564 39568
rect 43076 39516 43128 39568
rect 31576 39448 31628 39500
rect 32680 39448 32732 39500
rect 36176 39491 36228 39500
rect 36176 39457 36185 39491
rect 36185 39457 36219 39491
rect 36219 39457 36228 39491
rect 36176 39448 36228 39457
rect 10968 39380 11020 39432
rect 12992 39380 13044 39432
rect 21456 39380 21508 39432
rect 23664 39423 23716 39432
rect 23664 39389 23673 39423
rect 23673 39389 23707 39423
rect 23707 39389 23716 39423
rect 23664 39380 23716 39389
rect 25320 39380 25372 39432
rect 26884 39423 26936 39432
rect 17316 39312 17368 39364
rect 24032 39312 24084 39364
rect 24216 39355 24268 39364
rect 24216 39321 24225 39355
rect 24225 39321 24259 39355
rect 24259 39321 24268 39355
rect 24216 39312 24268 39321
rect 26240 39312 26292 39364
rect 26884 39389 26893 39423
rect 26893 39389 26927 39423
rect 26927 39389 26936 39423
rect 26884 39380 26936 39389
rect 13636 39244 13688 39296
rect 15016 39244 15068 39296
rect 22928 39244 22980 39296
rect 24400 39244 24452 39296
rect 25780 39244 25832 39296
rect 31116 39355 31168 39364
rect 31116 39321 31125 39355
rect 31125 39321 31159 39355
rect 31159 39321 31168 39355
rect 31116 39312 31168 39321
rect 33140 39380 33192 39432
rect 35256 39423 35308 39432
rect 35256 39389 35265 39423
rect 35265 39389 35299 39423
rect 35299 39389 35308 39423
rect 35256 39380 35308 39389
rect 42432 39491 42484 39500
rect 42432 39457 42441 39491
rect 42441 39457 42475 39491
rect 42475 39457 42484 39491
rect 42432 39448 42484 39457
rect 43168 39448 43220 39500
rect 36636 39423 36688 39432
rect 33508 39312 33560 39364
rect 36636 39389 36645 39423
rect 36645 39389 36679 39423
rect 36679 39389 36688 39423
rect 36636 39380 36688 39389
rect 38660 39380 38712 39432
rect 40224 39380 40276 39432
rect 39304 39312 39356 39364
rect 29460 39244 29512 39296
rect 35716 39287 35768 39296
rect 35716 39253 35725 39287
rect 35725 39253 35759 39287
rect 35759 39253 35768 39287
rect 35716 39244 35768 39253
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 22192 39083 22244 39092
rect 22192 39049 22201 39083
rect 22201 39049 22235 39083
rect 22235 39049 22244 39083
rect 22192 39040 22244 39049
rect 23480 39083 23532 39092
rect 23480 39049 23489 39083
rect 23489 39049 23523 39083
rect 23523 39049 23532 39083
rect 23480 39040 23532 39049
rect 23664 39040 23716 39092
rect 30656 39040 30708 39092
rect 32680 39083 32732 39092
rect 32680 39049 32689 39083
rect 32689 39049 32723 39083
rect 32723 39049 32732 39083
rect 32680 39040 32732 39049
rect 38568 39083 38620 39092
rect 38568 39049 38577 39083
rect 38577 39049 38611 39083
rect 38611 39049 38620 39083
rect 38568 39040 38620 39049
rect 40224 39040 40276 39092
rect 41696 39040 41748 39092
rect 42708 39040 42760 39092
rect 43168 39083 43220 39092
rect 43168 39049 43177 39083
rect 43177 39049 43211 39083
rect 43211 39049 43220 39083
rect 43168 39040 43220 39049
rect 26700 38972 26752 39024
rect 31116 38972 31168 39024
rect 32220 38972 32272 39024
rect 38752 38972 38804 39024
rect 39304 39015 39356 39024
rect 39304 38981 39313 39015
rect 39313 38981 39347 39015
rect 39347 38981 39356 39015
rect 39304 38972 39356 38981
rect 8300 38904 8352 38956
rect 11152 38947 11204 38956
rect 11152 38913 11161 38947
rect 11161 38913 11195 38947
rect 11195 38913 11204 38947
rect 11152 38904 11204 38913
rect 21180 38947 21232 38956
rect 21180 38913 21189 38947
rect 21189 38913 21223 38947
rect 21223 38913 21232 38947
rect 21180 38904 21232 38913
rect 24216 38947 24268 38956
rect 24216 38913 24225 38947
rect 24225 38913 24259 38947
rect 24259 38913 24268 38947
rect 24216 38904 24268 38913
rect 25780 38947 25832 38956
rect 25780 38913 25789 38947
rect 25789 38913 25823 38947
rect 25823 38913 25832 38947
rect 25780 38904 25832 38913
rect 28172 38904 28224 38956
rect 11980 38836 12032 38888
rect 12808 38836 12860 38888
rect 14832 38879 14884 38888
rect 10876 38811 10928 38820
rect 10876 38777 10885 38811
rect 10885 38777 10919 38811
rect 10919 38777 10928 38811
rect 10876 38768 10928 38777
rect 10968 38811 11020 38820
rect 10968 38777 10977 38811
rect 10977 38777 11011 38811
rect 11011 38777 11020 38811
rect 13728 38811 13780 38820
rect 10968 38768 11020 38777
rect 13728 38777 13737 38811
rect 13737 38777 13771 38811
rect 13771 38777 13780 38811
rect 13728 38768 13780 38777
rect 14832 38845 14841 38879
rect 14841 38845 14875 38879
rect 14875 38845 14884 38879
rect 14832 38836 14884 38845
rect 22100 38836 22152 38888
rect 29276 38836 29328 38888
rect 23388 38768 23440 38820
rect 23572 38768 23624 38820
rect 11888 38700 11940 38752
rect 15844 38743 15896 38752
rect 15844 38709 15853 38743
rect 15853 38709 15887 38743
rect 15887 38709 15896 38743
rect 15844 38700 15896 38709
rect 16120 38743 16172 38752
rect 16120 38709 16129 38743
rect 16129 38709 16163 38743
rect 16163 38709 16172 38743
rect 16120 38700 16172 38709
rect 16304 38700 16356 38752
rect 16856 38743 16908 38752
rect 16856 38709 16865 38743
rect 16865 38709 16899 38743
rect 16899 38709 16908 38743
rect 16856 38700 16908 38709
rect 20996 38700 21048 38752
rect 21456 38743 21508 38752
rect 21456 38709 21465 38743
rect 21465 38709 21499 38743
rect 21499 38709 21508 38743
rect 21456 38700 21508 38709
rect 21548 38700 21600 38752
rect 22468 38743 22520 38752
rect 22468 38709 22477 38743
rect 22477 38709 22511 38743
rect 22511 38709 22520 38743
rect 22468 38700 22520 38709
rect 22928 38700 22980 38752
rect 23480 38700 23532 38752
rect 25320 38768 25372 38820
rect 25596 38811 25648 38820
rect 25596 38777 25605 38811
rect 25605 38777 25639 38811
rect 25639 38777 25648 38811
rect 25596 38768 25648 38777
rect 24032 38700 24084 38752
rect 25136 38700 25188 38752
rect 25688 38700 25740 38752
rect 27252 38743 27304 38752
rect 27252 38709 27261 38743
rect 27261 38709 27295 38743
rect 27295 38709 27304 38743
rect 29460 38768 29512 38820
rect 29920 38768 29972 38820
rect 27252 38700 27304 38709
rect 28356 38700 28408 38752
rect 29092 38700 29144 38752
rect 31116 38743 31168 38752
rect 31116 38709 31125 38743
rect 31125 38709 31159 38743
rect 31159 38709 31168 38743
rect 33600 38768 33652 38820
rect 34612 38904 34664 38956
rect 36636 38904 36688 38956
rect 43076 38972 43128 39024
rect 43444 38972 43496 39024
rect 35256 38879 35308 38888
rect 35256 38845 35265 38879
rect 35265 38845 35299 38879
rect 35299 38845 35308 38879
rect 35256 38836 35308 38845
rect 35716 38879 35768 38888
rect 35716 38845 35725 38879
rect 35725 38845 35759 38879
rect 35759 38845 35768 38879
rect 35716 38836 35768 38845
rect 34336 38768 34388 38820
rect 35900 38811 35952 38820
rect 35900 38777 35909 38811
rect 35909 38777 35943 38811
rect 35943 38777 35952 38811
rect 35900 38768 35952 38777
rect 38752 38811 38804 38820
rect 38752 38777 38761 38811
rect 38761 38777 38795 38811
rect 38795 38777 38804 38811
rect 38752 38768 38804 38777
rect 32312 38743 32364 38752
rect 31116 38700 31168 38709
rect 32312 38709 32321 38743
rect 32321 38709 32355 38743
rect 32355 38709 32364 38743
rect 32312 38700 32364 38709
rect 33048 38743 33100 38752
rect 33048 38709 33057 38743
rect 33057 38709 33091 38743
rect 33091 38709 33100 38743
rect 33048 38700 33100 38709
rect 36176 38700 36228 38752
rect 36360 38700 36412 38752
rect 36912 38700 36964 38752
rect 37096 38743 37148 38752
rect 37096 38709 37105 38743
rect 37105 38709 37139 38743
rect 37139 38709 37148 38743
rect 37096 38700 37148 38709
rect 38108 38743 38160 38752
rect 38108 38709 38117 38743
rect 38117 38709 38151 38743
rect 38151 38709 38160 38743
rect 41420 38768 41472 38820
rect 41880 38811 41932 38820
rect 41880 38777 41889 38811
rect 41889 38777 41923 38811
rect 41923 38777 41932 38811
rect 41880 38768 41932 38777
rect 40040 38743 40092 38752
rect 38108 38700 38160 38709
rect 40040 38709 40049 38743
rect 40049 38709 40083 38743
rect 40083 38709 40092 38743
rect 40040 38700 40092 38709
rect 41144 38743 41196 38752
rect 41144 38709 41153 38743
rect 41153 38709 41187 38743
rect 41187 38709 41196 38743
rect 41144 38700 41196 38709
rect 41604 38743 41656 38752
rect 41604 38709 41613 38743
rect 41613 38709 41647 38743
rect 41647 38709 41656 38743
rect 41604 38700 41656 38709
rect 43444 38811 43496 38820
rect 43444 38777 43453 38811
rect 43453 38777 43487 38811
rect 43487 38777 43496 38811
rect 43444 38768 43496 38777
rect 43536 38700 43588 38752
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 10232 38428 10284 38480
rect 13728 38496 13780 38548
rect 23388 38496 23440 38548
rect 24584 38496 24636 38548
rect 26240 38539 26292 38548
rect 13820 38471 13872 38480
rect 13820 38437 13829 38471
rect 13829 38437 13863 38471
rect 13863 38437 13872 38471
rect 15476 38471 15528 38480
rect 13820 38428 13872 38437
rect 15476 38437 15485 38471
rect 15485 38437 15519 38471
rect 15519 38437 15528 38471
rect 15476 38428 15528 38437
rect 20996 38471 21048 38480
rect 20996 38437 21005 38471
rect 21005 38437 21039 38471
rect 21039 38437 21048 38471
rect 20996 38428 21048 38437
rect 21088 38471 21140 38480
rect 21088 38437 21097 38471
rect 21097 38437 21131 38471
rect 21131 38437 21140 38471
rect 21088 38428 21140 38437
rect 22284 38428 22336 38480
rect 22836 38471 22888 38480
rect 22836 38437 22845 38471
rect 22845 38437 22879 38471
rect 22879 38437 22888 38471
rect 22836 38428 22888 38437
rect 22928 38471 22980 38480
rect 22928 38437 22937 38471
rect 22937 38437 22971 38471
rect 22971 38437 22980 38471
rect 22928 38428 22980 38437
rect 24400 38471 24452 38480
rect 24400 38437 24409 38471
rect 24409 38437 24443 38471
rect 24443 38437 24452 38471
rect 24400 38428 24452 38437
rect 25136 38428 25188 38480
rect 26240 38505 26249 38539
rect 26249 38505 26283 38539
rect 26283 38505 26292 38539
rect 26240 38496 26292 38505
rect 27988 38496 28040 38548
rect 29276 38539 29328 38548
rect 26608 38471 26660 38480
rect 26608 38437 26617 38471
rect 26617 38437 26651 38471
rect 26651 38437 26660 38471
rect 26608 38428 26660 38437
rect 26700 38471 26752 38480
rect 26700 38437 26709 38471
rect 26709 38437 26743 38471
rect 26743 38437 26752 38471
rect 29276 38505 29285 38539
rect 29285 38505 29319 38539
rect 29319 38505 29328 38539
rect 29276 38496 29328 38505
rect 33048 38496 33100 38548
rect 33600 38496 33652 38548
rect 33968 38496 34020 38548
rect 36636 38496 36688 38548
rect 40040 38496 40092 38548
rect 41512 38539 41564 38548
rect 41512 38505 41521 38539
rect 41521 38505 41555 38539
rect 41555 38505 41564 38539
rect 41512 38496 41564 38505
rect 41880 38496 41932 38548
rect 43536 38539 43588 38548
rect 43536 38505 43545 38539
rect 43545 38505 43579 38539
rect 43579 38505 43588 38539
rect 43536 38496 43588 38505
rect 33692 38471 33744 38480
rect 26700 38428 26752 38437
rect 33692 38437 33701 38471
rect 33701 38437 33735 38471
rect 33735 38437 33744 38471
rect 33692 38428 33744 38437
rect 33784 38471 33836 38480
rect 33784 38437 33793 38471
rect 33793 38437 33827 38471
rect 33827 38437 33836 38471
rect 33784 38428 33836 38437
rect 35716 38428 35768 38480
rect 37004 38428 37056 38480
rect 38752 38428 38804 38480
rect 39120 38428 39172 38480
rect 11888 38403 11940 38412
rect 11888 38369 11897 38403
rect 11897 38369 11931 38403
rect 11931 38369 11940 38403
rect 11888 38360 11940 38369
rect 17776 38360 17828 38412
rect 19064 38360 19116 38412
rect 29552 38403 29604 38412
rect 10048 38335 10100 38344
rect 7196 38224 7248 38276
rect 10048 38301 10057 38335
rect 10057 38301 10091 38335
rect 10091 38301 10100 38335
rect 10048 38292 10100 38301
rect 10876 38292 10928 38344
rect 11244 38335 11296 38344
rect 11244 38301 11253 38335
rect 11253 38301 11287 38335
rect 11287 38301 11296 38335
rect 11244 38292 11296 38301
rect 13176 38292 13228 38344
rect 15384 38335 15436 38344
rect 11152 38224 11204 38276
rect 15384 38301 15393 38335
rect 15393 38301 15427 38335
rect 15427 38301 15436 38335
rect 15384 38292 15436 38301
rect 16120 38292 16172 38344
rect 21916 38292 21968 38344
rect 16856 38224 16908 38276
rect 25320 38292 25372 38344
rect 29092 38292 29144 38344
rect 29552 38369 29561 38403
rect 29561 38369 29595 38403
rect 29595 38369 29604 38403
rect 29552 38360 29604 38369
rect 30564 38403 30616 38412
rect 30564 38369 30573 38403
rect 30573 38369 30607 38403
rect 30607 38369 30616 38403
rect 30564 38360 30616 38369
rect 32864 38360 32916 38412
rect 33048 38360 33100 38412
rect 36084 38403 36136 38412
rect 36084 38369 36093 38403
rect 36093 38369 36127 38403
rect 36127 38369 36136 38403
rect 36084 38360 36136 38369
rect 36544 38403 36596 38412
rect 36544 38369 36553 38403
rect 36553 38369 36587 38403
rect 36587 38369 36596 38403
rect 36544 38360 36596 38369
rect 39488 38403 39540 38412
rect 39488 38369 39497 38403
rect 39497 38369 39531 38403
rect 39531 38369 39540 38403
rect 39488 38360 39540 38369
rect 41880 38360 41932 38412
rect 43812 38360 43864 38412
rect 34336 38335 34388 38344
rect 7656 38199 7708 38208
rect 7656 38165 7665 38199
rect 7665 38165 7699 38199
rect 7699 38165 7708 38199
rect 7656 38156 7708 38165
rect 19340 38156 19392 38208
rect 19616 38199 19668 38208
rect 19616 38165 19625 38199
rect 19625 38165 19659 38199
rect 19659 38165 19668 38199
rect 19616 38156 19668 38165
rect 21088 38156 21140 38208
rect 21732 38156 21784 38208
rect 25504 38199 25556 38208
rect 25504 38165 25513 38199
rect 25513 38165 25547 38199
rect 25547 38165 25556 38199
rect 25504 38156 25556 38165
rect 30196 38199 30248 38208
rect 30196 38165 30205 38199
rect 30205 38165 30239 38199
rect 30239 38165 30248 38199
rect 30196 38156 30248 38165
rect 34336 38301 34345 38335
rect 34345 38301 34379 38335
rect 34379 38301 34388 38335
rect 34336 38292 34388 38301
rect 35900 38292 35952 38344
rect 37924 38292 37976 38344
rect 38660 38292 38712 38344
rect 41696 38335 41748 38344
rect 41696 38301 41705 38335
rect 41705 38301 41739 38335
rect 41739 38301 41748 38335
rect 41696 38292 41748 38301
rect 41420 38224 41472 38276
rect 35256 38199 35308 38208
rect 35256 38165 35265 38199
rect 35265 38165 35299 38199
rect 35299 38165 35308 38199
rect 35256 38156 35308 38165
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 11888 37995 11940 38004
rect 11888 37961 11897 37995
rect 11897 37961 11931 37995
rect 11931 37961 11940 37995
rect 11888 37952 11940 37961
rect 11980 37952 12032 38004
rect 12808 37952 12860 38004
rect 13820 37952 13872 38004
rect 15476 37952 15528 38004
rect 17776 37995 17828 38004
rect 17776 37961 17785 37995
rect 17785 37961 17819 37995
rect 17819 37961 17828 37995
rect 17776 37952 17828 37961
rect 19064 37995 19116 38004
rect 19064 37961 19073 37995
rect 19073 37961 19107 37995
rect 19107 37961 19116 37995
rect 19064 37952 19116 37961
rect 20996 37952 21048 38004
rect 22836 37995 22888 38004
rect 22836 37961 22845 37995
rect 22845 37961 22879 37995
rect 22879 37961 22888 37995
rect 22836 37952 22888 37961
rect 23756 37952 23808 38004
rect 25136 37995 25188 38004
rect 25136 37961 25145 37995
rect 25145 37961 25179 37995
rect 25179 37961 25188 37995
rect 25136 37952 25188 37961
rect 25504 37952 25556 38004
rect 29092 37995 29144 38004
rect 29092 37961 29101 37995
rect 29101 37961 29135 37995
rect 29135 37961 29144 37995
rect 29092 37952 29144 37961
rect 29920 37995 29972 38004
rect 29920 37961 29929 37995
rect 29929 37961 29963 37995
rect 29963 37961 29972 37995
rect 29920 37952 29972 37961
rect 31116 37952 31168 38004
rect 33692 37952 33744 38004
rect 37004 37995 37056 38004
rect 37004 37961 37013 37995
rect 37013 37961 37047 37995
rect 37047 37961 37056 37995
rect 37004 37952 37056 37961
rect 38108 37995 38160 38004
rect 38108 37961 38117 37995
rect 38117 37961 38151 37995
rect 38151 37961 38160 37995
rect 38108 37952 38160 37961
rect 10232 37927 10284 37936
rect 10232 37893 10241 37927
rect 10241 37893 10275 37927
rect 10275 37893 10284 37927
rect 10232 37884 10284 37893
rect 8300 37859 8352 37868
rect 8300 37825 8309 37859
rect 8309 37825 8343 37859
rect 8343 37825 8352 37859
rect 8300 37816 8352 37825
rect 7656 37723 7708 37732
rect 7656 37689 7665 37723
rect 7665 37689 7699 37723
rect 7699 37689 7708 37723
rect 7656 37680 7708 37689
rect 9496 37816 9548 37868
rect 10048 37816 10100 37868
rect 14004 37884 14056 37936
rect 13912 37816 13964 37868
rect 12808 37748 12860 37800
rect 13636 37748 13688 37800
rect 16856 37791 16908 37800
rect 9036 37723 9088 37732
rect 9036 37689 9045 37723
rect 9045 37689 9079 37723
rect 9079 37689 9088 37723
rect 9036 37680 9088 37689
rect 9220 37723 9272 37732
rect 9220 37689 9229 37723
rect 9229 37689 9263 37723
rect 9263 37689 9272 37723
rect 9220 37680 9272 37689
rect 9496 37680 9548 37732
rect 10876 37723 10928 37732
rect 10876 37689 10885 37723
rect 10885 37689 10919 37723
rect 10919 37689 10928 37723
rect 10876 37680 10928 37689
rect 11244 37680 11296 37732
rect 13176 37680 13228 37732
rect 16856 37757 16865 37791
rect 16865 37757 16899 37791
rect 16899 37757 16908 37791
rect 16856 37748 16908 37757
rect 26608 37884 26660 37936
rect 30840 37884 30892 37936
rect 19340 37816 19392 37868
rect 21088 37816 21140 37868
rect 21732 37816 21784 37868
rect 21916 37859 21968 37868
rect 21916 37825 21925 37859
rect 21925 37825 21959 37859
rect 21959 37825 21968 37859
rect 21916 37816 21968 37825
rect 29736 37816 29788 37868
rect 30564 37816 30616 37868
rect 33784 37927 33836 37936
rect 33784 37893 33793 37927
rect 33793 37893 33827 37927
rect 33827 37893 33836 37927
rect 33784 37884 33836 37893
rect 36084 37884 36136 37936
rect 34336 37816 34388 37868
rect 37556 37816 37608 37868
rect 37832 37816 37884 37868
rect 19248 37748 19300 37800
rect 26516 37791 26568 37800
rect 19616 37723 19668 37732
rect 19616 37689 19625 37723
rect 19625 37689 19659 37723
rect 19659 37689 19668 37723
rect 19616 37680 19668 37689
rect 20168 37723 20220 37732
rect 20168 37689 20177 37723
rect 20177 37689 20211 37723
rect 20211 37689 20220 37723
rect 20168 37680 20220 37689
rect 18328 37612 18380 37664
rect 21824 37612 21876 37664
rect 23848 37612 23900 37664
rect 26516 37757 26525 37791
rect 26525 37757 26559 37791
rect 26559 37757 26568 37791
rect 26516 37748 26568 37757
rect 29552 37791 29604 37800
rect 29552 37757 29561 37791
rect 29561 37757 29595 37791
rect 29595 37757 29604 37791
rect 29552 37748 29604 37757
rect 29920 37748 29972 37800
rect 30196 37748 30248 37800
rect 32404 37748 32456 37800
rect 37004 37748 37056 37800
rect 26700 37680 26752 37732
rect 30012 37680 30064 37732
rect 32312 37723 32364 37732
rect 32312 37689 32321 37723
rect 32321 37689 32355 37723
rect 32355 37689 32364 37723
rect 32312 37680 32364 37689
rect 34796 37680 34848 37732
rect 36544 37723 36596 37732
rect 25688 37612 25740 37664
rect 25964 37655 26016 37664
rect 25964 37621 25973 37655
rect 25973 37621 26007 37655
rect 26007 37621 26016 37655
rect 25964 37612 26016 37621
rect 27252 37612 27304 37664
rect 34612 37655 34664 37664
rect 34612 37621 34621 37655
rect 34621 37621 34655 37655
rect 34655 37621 34664 37655
rect 36544 37689 36553 37723
rect 36553 37689 36587 37723
rect 36587 37689 36596 37723
rect 36544 37680 36596 37689
rect 37096 37680 37148 37732
rect 39304 37952 39356 38004
rect 39488 37952 39540 38004
rect 41420 37952 41472 38004
rect 41696 37995 41748 38004
rect 41696 37961 41705 37995
rect 41705 37961 41739 37995
rect 41739 37961 41748 37995
rect 41696 37952 41748 37961
rect 41788 37884 41840 37936
rect 40408 37748 40460 37800
rect 43628 37748 43680 37800
rect 39120 37680 39172 37732
rect 41880 37680 41932 37732
rect 36084 37655 36136 37664
rect 34612 37612 34664 37621
rect 36084 37621 36093 37655
rect 36093 37621 36127 37655
rect 36127 37621 36136 37655
rect 36084 37612 36136 37621
rect 42432 37612 42484 37664
rect 43812 37655 43864 37664
rect 43812 37621 43821 37655
rect 43821 37621 43855 37655
rect 43855 37621 43864 37655
rect 43812 37612 43864 37621
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 9220 37451 9272 37460
rect 9220 37417 9229 37451
rect 9229 37417 9263 37451
rect 9263 37417 9272 37451
rect 9220 37408 9272 37417
rect 10876 37451 10928 37460
rect 10876 37417 10885 37451
rect 10885 37417 10919 37451
rect 10919 37417 10928 37451
rect 10876 37408 10928 37417
rect 13636 37408 13688 37460
rect 15384 37408 15436 37460
rect 19340 37408 19392 37460
rect 21732 37408 21784 37460
rect 23480 37408 23532 37460
rect 25964 37408 26016 37460
rect 26516 37408 26568 37460
rect 34612 37408 34664 37460
rect 37924 37451 37976 37460
rect 37924 37417 37933 37451
rect 37933 37417 37967 37451
rect 37967 37417 37976 37451
rect 37924 37408 37976 37417
rect 39948 37408 40000 37460
rect 40684 37408 40736 37460
rect 41604 37408 41656 37460
rect 41880 37408 41932 37460
rect 42432 37451 42484 37460
rect 42432 37417 42441 37451
rect 42441 37417 42475 37451
rect 42475 37417 42484 37451
rect 42432 37408 42484 37417
rect 7104 37340 7156 37392
rect 10232 37340 10284 37392
rect 11428 37383 11480 37392
rect 11428 37349 11437 37383
rect 11437 37349 11471 37383
rect 11471 37349 11480 37383
rect 11428 37340 11480 37349
rect 12992 37383 13044 37392
rect 12992 37349 13001 37383
rect 13001 37349 13035 37383
rect 13035 37349 13044 37383
rect 12992 37340 13044 37349
rect 18420 37340 18472 37392
rect 21548 37383 21600 37392
rect 21548 37349 21557 37383
rect 21557 37349 21591 37383
rect 21591 37349 21600 37383
rect 21548 37340 21600 37349
rect 21824 37340 21876 37392
rect 22928 37340 22980 37392
rect 23848 37340 23900 37392
rect 30196 37383 30248 37392
rect 16304 37315 16356 37324
rect 16304 37281 16313 37315
rect 16313 37281 16347 37315
rect 16347 37281 16356 37315
rect 16304 37272 16356 37281
rect 17868 37272 17920 37324
rect 18512 37272 18564 37324
rect 22652 37272 22704 37324
rect 26608 37272 26660 37324
rect 30196 37349 30205 37383
rect 30205 37349 30239 37383
rect 30239 37349 30248 37383
rect 30196 37340 30248 37349
rect 32312 37340 32364 37392
rect 33232 37383 33284 37392
rect 33232 37349 33235 37383
rect 33235 37349 33269 37383
rect 33269 37349 33284 37383
rect 33232 37340 33284 37349
rect 39120 37340 39172 37392
rect 41512 37340 41564 37392
rect 27988 37272 28040 37324
rect 28356 37315 28408 37324
rect 28356 37281 28365 37315
rect 28365 37281 28399 37315
rect 28399 37281 28408 37315
rect 28356 37272 28408 37281
rect 29460 37315 29512 37324
rect 29460 37281 29469 37315
rect 29469 37281 29503 37315
rect 29503 37281 29512 37315
rect 29460 37272 29512 37281
rect 29920 37315 29972 37324
rect 29920 37281 29929 37315
rect 29929 37281 29963 37315
rect 29963 37281 29972 37315
rect 29920 37272 29972 37281
rect 31116 37315 31168 37324
rect 31116 37281 31134 37315
rect 31134 37281 31168 37315
rect 31116 37272 31168 37281
rect 6920 37247 6972 37256
rect 6920 37213 6929 37247
rect 6929 37213 6963 37247
rect 6963 37213 6972 37247
rect 6920 37204 6972 37213
rect 7196 37247 7248 37256
rect 7196 37213 7205 37247
rect 7205 37213 7239 37247
rect 7239 37213 7248 37247
rect 7196 37204 7248 37213
rect 8944 37204 8996 37256
rect 11336 37247 11388 37256
rect 11336 37213 11345 37247
rect 11345 37213 11379 37247
rect 11379 37213 11388 37247
rect 11336 37204 11388 37213
rect 7656 37136 7708 37188
rect 12900 37247 12952 37256
rect 12900 37213 12909 37247
rect 12909 37213 12943 37247
rect 12943 37213 12952 37247
rect 12900 37204 12952 37213
rect 13176 37247 13228 37256
rect 13176 37213 13185 37247
rect 13185 37213 13219 37247
rect 13219 37213 13228 37247
rect 13176 37204 13228 37213
rect 15752 37247 15804 37256
rect 15752 37213 15761 37247
rect 15761 37213 15795 37247
rect 15795 37213 15804 37247
rect 15752 37204 15804 37213
rect 18972 37247 19024 37256
rect 18972 37213 18981 37247
rect 18981 37213 19015 37247
rect 19015 37213 19024 37247
rect 18972 37204 19024 37213
rect 19340 37247 19392 37256
rect 19340 37213 19349 37247
rect 19349 37213 19383 37247
rect 19383 37213 19392 37247
rect 19340 37204 19392 37213
rect 20168 37204 20220 37256
rect 24032 37204 24084 37256
rect 29368 37204 29420 37256
rect 32864 37247 32916 37256
rect 32864 37213 32873 37247
rect 32873 37213 32907 37247
rect 32907 37213 32916 37247
rect 32864 37204 32916 37213
rect 35808 37272 35860 37324
rect 35992 37315 36044 37324
rect 35992 37281 36001 37315
rect 36001 37281 36035 37315
rect 36035 37281 36044 37315
rect 35992 37272 36044 37281
rect 43352 37272 43404 37324
rect 35440 37204 35492 37256
rect 35900 37204 35952 37256
rect 36176 37247 36228 37256
rect 36176 37213 36185 37247
rect 36185 37213 36219 37247
rect 36219 37213 36228 37247
rect 36176 37204 36228 37213
rect 38660 37247 38712 37256
rect 38660 37213 38669 37247
rect 38669 37213 38703 37247
rect 38703 37213 38712 37247
rect 38660 37204 38712 37213
rect 40776 37247 40828 37256
rect 40776 37213 40785 37247
rect 40785 37213 40819 37247
rect 40819 37213 40828 37247
rect 40776 37204 40828 37213
rect 40592 37136 40644 37188
rect 18420 37111 18472 37120
rect 18420 37077 18429 37111
rect 18429 37077 18463 37111
rect 18463 37077 18472 37111
rect 18420 37068 18472 37077
rect 25228 37068 25280 37120
rect 29736 37068 29788 37120
rect 31300 37068 31352 37120
rect 32404 37068 32456 37120
rect 34796 37068 34848 37120
rect 37096 37111 37148 37120
rect 37096 37077 37105 37111
rect 37105 37077 37139 37111
rect 37139 37077 37148 37111
rect 37096 37068 37148 37077
rect 37556 37068 37608 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 6920 36864 6972 36916
rect 8944 36907 8996 36916
rect 8944 36873 8953 36907
rect 8953 36873 8987 36907
rect 8987 36873 8996 36907
rect 8944 36864 8996 36873
rect 10232 36864 10284 36916
rect 11336 36864 11388 36916
rect 11980 36864 12032 36916
rect 12992 36864 13044 36916
rect 13912 36864 13964 36916
rect 16304 36864 16356 36916
rect 17868 36907 17920 36916
rect 17868 36873 17877 36907
rect 17877 36873 17911 36907
rect 17911 36873 17920 36907
rect 17868 36864 17920 36873
rect 21456 36864 21508 36916
rect 22560 36796 22612 36848
rect 26608 36839 26660 36848
rect 8208 36728 8260 36780
rect 9220 36728 9272 36780
rect 10876 36728 10928 36780
rect 14280 36728 14332 36780
rect 14648 36771 14700 36780
rect 14648 36737 14657 36771
rect 14657 36737 14691 36771
rect 14691 36737 14700 36771
rect 14648 36728 14700 36737
rect 18328 36771 18380 36780
rect 18328 36737 18337 36771
rect 18337 36737 18371 36771
rect 18371 36737 18380 36771
rect 18328 36728 18380 36737
rect 21916 36728 21968 36780
rect 22008 36728 22060 36780
rect 22652 36728 22704 36780
rect 26608 36805 26617 36839
rect 26617 36805 26651 36839
rect 26651 36805 26660 36839
rect 26608 36796 26660 36805
rect 23848 36728 23900 36780
rect 25688 36771 25740 36780
rect 25688 36737 25697 36771
rect 25697 36737 25731 36771
rect 25731 36737 25740 36771
rect 25688 36728 25740 36737
rect 9864 36635 9916 36644
rect 5540 36567 5592 36576
rect 5540 36533 5549 36567
rect 5549 36533 5583 36567
rect 5583 36533 5592 36567
rect 5540 36524 5592 36533
rect 6184 36567 6236 36576
rect 6184 36533 6193 36567
rect 6193 36533 6227 36567
rect 6227 36533 6236 36567
rect 6184 36524 6236 36533
rect 7104 36524 7156 36576
rect 9864 36601 9873 36635
rect 9873 36601 9907 36635
rect 9907 36601 9916 36635
rect 9864 36592 9916 36601
rect 10232 36592 10284 36644
rect 11428 36524 11480 36576
rect 14004 36592 14056 36644
rect 15568 36635 15620 36644
rect 15568 36601 15577 36635
rect 15577 36601 15611 36635
rect 15611 36601 15620 36635
rect 15568 36592 15620 36601
rect 15752 36592 15804 36644
rect 18420 36635 18472 36644
rect 18420 36601 18429 36635
rect 18429 36601 18463 36635
rect 18463 36601 18472 36635
rect 18420 36592 18472 36601
rect 19064 36592 19116 36644
rect 19892 36635 19944 36644
rect 19892 36601 19901 36635
rect 19901 36601 19935 36635
rect 19935 36601 19944 36635
rect 19892 36592 19944 36601
rect 21732 36592 21784 36644
rect 21916 36635 21968 36644
rect 21916 36601 21925 36635
rect 21925 36601 21959 36635
rect 21959 36601 21968 36635
rect 21916 36592 21968 36601
rect 21364 36524 21416 36576
rect 21824 36524 21876 36576
rect 24032 36592 24084 36644
rect 23572 36524 23624 36576
rect 25228 36660 25280 36712
rect 26792 36703 26844 36712
rect 26792 36669 26801 36703
rect 26801 36669 26835 36703
rect 26835 36669 26844 36703
rect 26792 36660 26844 36669
rect 27620 36660 27672 36712
rect 27988 36864 28040 36916
rect 29644 36864 29696 36916
rect 31116 36907 31168 36916
rect 31116 36873 31125 36907
rect 31125 36873 31159 36907
rect 31159 36873 31168 36907
rect 31116 36864 31168 36873
rect 32312 36864 32364 36916
rect 33784 36907 33836 36916
rect 33784 36873 33793 36907
rect 33793 36873 33827 36907
rect 33827 36873 33836 36907
rect 33784 36864 33836 36873
rect 35808 36864 35860 36916
rect 36176 36864 36228 36916
rect 40776 36864 40828 36916
rect 41512 36907 41564 36916
rect 41512 36873 41521 36907
rect 41521 36873 41555 36907
rect 41555 36873 41564 36907
rect 41512 36864 41564 36873
rect 41604 36864 41656 36916
rect 32404 36771 32456 36780
rect 29736 36703 29788 36712
rect 28540 36592 28592 36644
rect 28908 36592 28960 36644
rect 29736 36669 29745 36703
rect 29745 36669 29779 36703
rect 29779 36669 29788 36703
rect 29736 36660 29788 36669
rect 32404 36737 32413 36771
rect 32413 36737 32447 36771
rect 32447 36737 32456 36771
rect 32404 36728 32456 36737
rect 32128 36703 32180 36712
rect 32128 36669 32137 36703
rect 32137 36669 32171 36703
rect 32171 36669 32180 36703
rect 32128 36660 32180 36669
rect 32956 36660 33008 36712
rect 33784 36660 33836 36712
rect 38660 36796 38712 36848
rect 38752 36796 38804 36848
rect 37556 36771 37608 36780
rect 37556 36737 37565 36771
rect 37565 36737 37599 36771
rect 37599 36737 37608 36771
rect 37556 36728 37608 36737
rect 39120 36771 39172 36780
rect 39120 36737 39129 36771
rect 39129 36737 39163 36771
rect 39163 36737 39172 36771
rect 39120 36728 39172 36737
rect 40592 36771 40644 36780
rect 40592 36737 40601 36771
rect 40601 36737 40635 36771
rect 40635 36737 40644 36771
rect 40592 36728 40644 36737
rect 41788 36796 41840 36848
rect 35992 36703 36044 36712
rect 32404 36592 32456 36644
rect 32680 36592 32732 36644
rect 35992 36669 36001 36703
rect 36001 36669 36035 36703
rect 36035 36669 36044 36703
rect 35992 36660 36044 36669
rect 24676 36524 24728 36576
rect 27896 36524 27948 36576
rect 28356 36567 28408 36576
rect 28356 36533 28365 36567
rect 28365 36533 28399 36567
rect 28399 36533 28408 36567
rect 28356 36524 28408 36533
rect 29368 36567 29420 36576
rect 29368 36533 29377 36567
rect 29377 36533 29411 36567
rect 29411 36533 29420 36567
rect 29368 36524 29420 36533
rect 29460 36524 29512 36576
rect 35440 36524 35492 36576
rect 36636 36524 36688 36576
rect 36728 36524 36780 36576
rect 37096 36660 37148 36712
rect 37924 36660 37976 36712
rect 38292 36660 38344 36712
rect 40684 36635 40736 36644
rect 40684 36601 40693 36635
rect 40693 36601 40727 36635
rect 40727 36601 40736 36635
rect 40684 36592 40736 36601
rect 41972 36796 42024 36848
rect 42340 36728 42392 36780
rect 38936 36524 38988 36576
rect 39580 36567 39632 36576
rect 39580 36533 39589 36567
rect 39589 36533 39623 36567
rect 39623 36533 39632 36567
rect 39580 36524 39632 36533
rect 43352 36567 43404 36576
rect 43352 36533 43361 36567
rect 43361 36533 43395 36567
rect 43395 36533 43404 36567
rect 43352 36524 43404 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 6092 36295 6144 36304
rect 6092 36261 6101 36295
rect 6101 36261 6135 36295
rect 6135 36261 6144 36295
rect 6092 36252 6144 36261
rect 7196 36252 7248 36304
rect 7840 36252 7892 36304
rect 8208 36295 8260 36304
rect 8208 36261 8217 36295
rect 8217 36261 8251 36295
rect 8251 36261 8260 36295
rect 8208 36252 8260 36261
rect 9036 36252 9088 36304
rect 10140 36252 10192 36304
rect 11428 36320 11480 36372
rect 12900 36363 12952 36372
rect 12900 36329 12909 36363
rect 12909 36329 12943 36363
rect 12943 36329 12952 36363
rect 12900 36320 12952 36329
rect 14648 36320 14700 36372
rect 18420 36320 18472 36372
rect 18972 36363 19024 36372
rect 18972 36329 18981 36363
rect 18981 36329 19015 36363
rect 19015 36329 19024 36363
rect 18972 36320 19024 36329
rect 10876 36252 10928 36304
rect 11796 36295 11848 36304
rect 11796 36261 11805 36295
rect 11805 36261 11839 36295
rect 11839 36261 11848 36295
rect 11796 36252 11848 36261
rect 17684 36252 17736 36304
rect 5264 36184 5316 36236
rect 14004 36184 14056 36236
rect 16212 36227 16264 36236
rect 16212 36193 16221 36227
rect 16221 36193 16255 36227
rect 16255 36193 16264 36227
rect 16212 36184 16264 36193
rect 19248 36184 19300 36236
rect 20260 36320 20312 36372
rect 19892 36295 19944 36304
rect 19892 36261 19901 36295
rect 19901 36261 19935 36295
rect 19935 36261 19944 36295
rect 19892 36252 19944 36261
rect 21088 36252 21140 36304
rect 21916 36320 21968 36372
rect 23572 36320 23624 36372
rect 25044 36320 25096 36372
rect 25228 36363 25280 36372
rect 25228 36329 25237 36363
rect 25237 36329 25271 36363
rect 25271 36329 25280 36363
rect 25228 36320 25280 36329
rect 27620 36363 27672 36372
rect 27620 36329 27629 36363
rect 27629 36329 27663 36363
rect 27663 36329 27672 36363
rect 27620 36320 27672 36329
rect 29920 36320 29972 36372
rect 31576 36320 31628 36372
rect 32128 36320 32180 36372
rect 24308 36295 24360 36304
rect 24308 36261 24317 36295
rect 24317 36261 24351 36295
rect 24351 36261 24360 36295
rect 24308 36252 24360 36261
rect 26424 36252 26476 36304
rect 30564 36295 30616 36304
rect 30564 36261 30573 36295
rect 30573 36261 30607 36295
rect 30607 36261 30616 36295
rect 30564 36252 30616 36261
rect 32864 36295 32916 36304
rect 23020 36184 23072 36236
rect 28908 36227 28960 36236
rect 28908 36193 28917 36227
rect 28917 36193 28951 36227
rect 28951 36193 28960 36227
rect 28908 36184 28960 36193
rect 29092 36227 29144 36236
rect 29092 36193 29101 36227
rect 29101 36193 29135 36227
rect 29135 36193 29144 36227
rect 29092 36184 29144 36193
rect 32404 36227 32456 36236
rect 32404 36193 32413 36227
rect 32413 36193 32447 36227
rect 32447 36193 32456 36227
rect 32404 36184 32456 36193
rect 32864 36261 32873 36295
rect 32873 36261 32907 36295
rect 32907 36261 32916 36295
rect 35900 36320 35952 36372
rect 36268 36320 36320 36372
rect 37924 36363 37976 36372
rect 37924 36329 37933 36363
rect 37933 36329 37967 36363
rect 37967 36329 37976 36363
rect 37924 36320 37976 36329
rect 32864 36252 32916 36261
rect 38936 36252 38988 36304
rect 39212 36295 39264 36304
rect 39212 36261 39221 36295
rect 39221 36261 39255 36295
rect 39255 36261 39264 36295
rect 40776 36295 40828 36304
rect 39212 36252 39264 36261
rect 40776 36261 40785 36295
rect 40785 36261 40819 36295
rect 40819 36261 40828 36295
rect 40776 36252 40828 36261
rect 33048 36184 33100 36236
rect 33232 36184 33284 36236
rect 34612 36184 34664 36236
rect 36084 36227 36136 36236
rect 36084 36193 36093 36227
rect 36093 36193 36127 36227
rect 36127 36193 36136 36227
rect 36084 36184 36136 36193
rect 36544 36227 36596 36236
rect 36544 36193 36553 36227
rect 36553 36193 36587 36227
rect 36587 36193 36596 36227
rect 36544 36184 36596 36193
rect 36636 36184 36688 36236
rect 38476 36184 38528 36236
rect 41696 36184 41748 36236
rect 42708 36184 42760 36236
rect 43904 36184 43956 36236
rect 6000 36159 6052 36168
rect 6000 36125 6009 36159
rect 6009 36125 6043 36159
rect 6043 36125 6052 36159
rect 6000 36116 6052 36125
rect 8208 36116 8260 36168
rect 10416 36116 10468 36168
rect 11704 36159 11756 36168
rect 11704 36125 11713 36159
rect 11713 36125 11747 36159
rect 11747 36125 11756 36159
rect 11704 36116 11756 36125
rect 11980 36159 12032 36168
rect 11980 36125 11989 36159
rect 11989 36125 12023 36159
rect 12023 36125 12032 36159
rect 11980 36116 12032 36125
rect 15660 36116 15712 36168
rect 17408 36116 17460 36168
rect 20720 36116 20772 36168
rect 24492 36159 24544 36168
rect 19064 36048 19116 36100
rect 22008 36048 22060 36100
rect 24124 36048 24176 36100
rect 24492 36125 24501 36159
rect 24501 36125 24535 36159
rect 24535 36125 24544 36159
rect 24492 36116 24544 36125
rect 27528 36116 27580 36168
rect 29368 36159 29420 36168
rect 29368 36125 29377 36159
rect 29377 36125 29411 36159
rect 29411 36125 29420 36159
rect 29368 36116 29420 36125
rect 30472 36159 30524 36168
rect 30472 36125 30481 36159
rect 30481 36125 30515 36159
rect 30515 36125 30524 36159
rect 30472 36116 30524 36125
rect 36820 36159 36872 36168
rect 36820 36125 36829 36159
rect 36829 36125 36863 36159
rect 36863 36125 36872 36159
rect 36820 36116 36872 36125
rect 39396 36159 39448 36168
rect 39396 36125 39405 36159
rect 39405 36125 39439 36159
rect 39439 36125 39448 36159
rect 39396 36116 39448 36125
rect 40316 36116 40368 36168
rect 41328 36159 41380 36168
rect 41328 36125 41337 36159
rect 41337 36125 41371 36159
rect 41371 36125 41380 36159
rect 41328 36116 41380 36125
rect 43260 36116 43312 36168
rect 27252 36048 27304 36100
rect 29276 36048 29328 36100
rect 31024 36091 31076 36100
rect 31024 36057 31033 36091
rect 31033 36057 31067 36091
rect 31067 36057 31076 36091
rect 31024 36048 31076 36057
rect 32496 36048 32548 36100
rect 34060 36048 34112 36100
rect 41144 36048 41196 36100
rect 41696 36048 41748 36100
rect 41788 36048 41840 36100
rect 4620 36023 4672 36032
rect 4620 35989 4629 36023
rect 4629 35989 4663 36023
rect 4663 35989 4672 36023
rect 4620 35980 4672 35989
rect 7104 36023 7156 36032
rect 7104 35989 7113 36023
rect 7113 35989 7147 36023
rect 7147 35989 7156 36023
rect 7104 35980 7156 35989
rect 9864 36023 9916 36032
rect 9864 35989 9873 36023
rect 9873 35989 9907 36023
rect 9907 35989 9916 36023
rect 9864 35980 9916 35989
rect 13636 36023 13688 36032
rect 13636 35989 13645 36023
rect 13645 35989 13679 36023
rect 13679 35989 13688 36023
rect 13636 35980 13688 35989
rect 15568 36023 15620 36032
rect 15568 35989 15577 36023
rect 15577 35989 15611 36023
rect 15611 35989 15620 36023
rect 15568 35980 15620 35989
rect 16028 35980 16080 36032
rect 24032 36023 24084 36032
rect 24032 35989 24041 36023
rect 24041 35989 24075 36023
rect 24075 35989 24084 36023
rect 24032 35980 24084 35989
rect 34704 35980 34756 36032
rect 43076 35980 43128 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 5540 35819 5592 35828
rect 5540 35785 5549 35819
rect 5549 35785 5583 35819
rect 5583 35785 5592 35819
rect 5540 35776 5592 35785
rect 6092 35776 6144 35828
rect 10140 35819 10192 35828
rect 10140 35785 10149 35819
rect 10149 35785 10183 35819
rect 10183 35785 10192 35819
rect 10140 35776 10192 35785
rect 11704 35776 11756 35828
rect 16212 35819 16264 35828
rect 16212 35785 16221 35819
rect 16221 35785 16255 35819
rect 16255 35785 16264 35819
rect 16212 35776 16264 35785
rect 19248 35819 19300 35828
rect 19248 35785 19257 35819
rect 19257 35785 19291 35819
rect 19291 35785 19300 35819
rect 19248 35776 19300 35785
rect 21088 35776 21140 35828
rect 23020 35776 23072 35828
rect 30472 35776 30524 35828
rect 30564 35819 30616 35828
rect 30564 35785 30573 35819
rect 30573 35785 30607 35819
rect 30607 35785 30616 35819
rect 30564 35776 30616 35785
rect 31300 35776 31352 35828
rect 31576 35819 31628 35828
rect 31576 35785 31585 35819
rect 31585 35785 31619 35819
rect 31619 35785 31628 35819
rect 31576 35776 31628 35785
rect 32404 35776 32456 35828
rect 35808 35776 35860 35828
rect 37004 35776 37056 35828
rect 38476 35819 38528 35828
rect 38476 35785 38485 35819
rect 38485 35785 38519 35819
rect 38519 35785 38528 35819
rect 38476 35776 38528 35785
rect 38936 35819 38988 35828
rect 38936 35785 38945 35819
rect 38945 35785 38979 35819
rect 38979 35785 38988 35819
rect 38936 35776 38988 35785
rect 40316 35819 40368 35828
rect 40316 35785 40325 35819
rect 40325 35785 40359 35819
rect 40359 35785 40368 35819
rect 40316 35776 40368 35785
rect 40776 35819 40828 35828
rect 40776 35785 40785 35819
rect 40785 35785 40819 35819
rect 40819 35785 40828 35819
rect 40776 35776 40828 35785
rect 41696 35776 41748 35828
rect 6184 35708 6236 35760
rect 11796 35708 11848 35760
rect 15292 35708 15344 35760
rect 21640 35708 21692 35760
rect 23204 35708 23256 35760
rect 7196 35640 7248 35692
rect 8944 35640 8996 35692
rect 11980 35640 12032 35692
rect 13636 35683 13688 35692
rect 13636 35649 13645 35683
rect 13645 35649 13679 35683
rect 13679 35649 13688 35683
rect 13636 35640 13688 35649
rect 14280 35683 14332 35692
rect 14280 35649 14289 35683
rect 14289 35649 14323 35683
rect 14323 35649 14332 35683
rect 14280 35640 14332 35649
rect 22192 35683 22244 35692
rect 22192 35649 22201 35683
rect 22201 35649 22235 35683
rect 22235 35649 22244 35683
rect 22192 35640 22244 35649
rect 24308 35640 24360 35692
rect 26884 35640 26936 35692
rect 26976 35683 27028 35692
rect 26976 35649 26985 35683
rect 26985 35649 27019 35683
rect 27019 35649 27028 35683
rect 28908 35708 28960 35760
rect 33232 35708 33284 35760
rect 26976 35640 27028 35649
rect 4620 35615 4672 35624
rect 4620 35581 4629 35615
rect 4629 35581 4663 35615
rect 4663 35581 4672 35615
rect 4620 35572 4672 35581
rect 4160 35479 4212 35488
rect 4160 35445 4169 35479
rect 4169 35445 4203 35479
rect 4203 35445 4212 35479
rect 4160 35436 4212 35445
rect 4712 35436 4764 35488
rect 7104 35504 7156 35556
rect 9312 35504 9364 35556
rect 10416 35504 10468 35556
rect 10876 35547 10928 35556
rect 10876 35513 10885 35547
rect 10885 35513 10919 35547
rect 10919 35513 10928 35547
rect 10876 35504 10928 35513
rect 7840 35479 7892 35488
rect 7840 35445 7849 35479
rect 7849 35445 7883 35479
rect 7883 35445 7892 35479
rect 7840 35436 7892 35445
rect 8208 35479 8260 35488
rect 8208 35445 8217 35479
rect 8217 35445 8251 35479
rect 8251 35445 8260 35479
rect 8208 35436 8260 35445
rect 10692 35479 10744 35488
rect 10692 35445 10701 35479
rect 10701 35445 10735 35479
rect 10735 35445 10744 35479
rect 10692 35436 10744 35445
rect 12900 35436 12952 35488
rect 13452 35504 13504 35556
rect 13728 35547 13780 35556
rect 13728 35513 13737 35547
rect 13737 35513 13771 35547
rect 13771 35513 13780 35547
rect 13728 35504 13780 35513
rect 15292 35547 15344 35556
rect 15292 35513 15301 35547
rect 15301 35513 15335 35547
rect 15335 35513 15344 35547
rect 15292 35504 15344 35513
rect 29276 35615 29328 35624
rect 19892 35504 19944 35556
rect 21364 35547 21416 35556
rect 21364 35513 21373 35547
rect 21373 35513 21407 35547
rect 21407 35513 21416 35547
rect 21364 35504 21416 35513
rect 24032 35504 24084 35556
rect 24400 35547 24452 35556
rect 24400 35513 24409 35547
rect 24409 35513 24443 35547
rect 24443 35513 24452 35547
rect 24400 35504 24452 35513
rect 26332 35504 26384 35556
rect 14556 35479 14608 35488
rect 14556 35445 14565 35479
rect 14565 35445 14599 35479
rect 14599 35445 14608 35479
rect 14556 35436 14608 35445
rect 17224 35479 17276 35488
rect 17224 35445 17233 35479
rect 17233 35445 17267 35479
rect 17267 35445 17276 35479
rect 17224 35436 17276 35445
rect 17684 35479 17736 35488
rect 17684 35445 17693 35479
rect 17693 35445 17727 35479
rect 17727 35445 17736 35479
rect 17684 35436 17736 35445
rect 24124 35436 24176 35488
rect 26424 35436 26476 35488
rect 29276 35581 29285 35615
rect 29285 35581 29319 35615
rect 29319 35581 29328 35615
rect 29276 35572 29328 35581
rect 29552 35504 29604 35556
rect 31852 35547 31904 35556
rect 31852 35513 31861 35547
rect 31861 35513 31895 35547
rect 31895 35513 31904 35547
rect 31852 35504 31904 35513
rect 33324 35547 33376 35556
rect 33324 35513 33333 35547
rect 33333 35513 33367 35547
rect 33367 35513 33376 35547
rect 33324 35504 33376 35513
rect 33416 35547 33468 35556
rect 33416 35513 33425 35547
rect 33425 35513 33459 35547
rect 33459 35513 33468 35547
rect 36820 35640 36872 35692
rect 41236 35683 41288 35692
rect 41236 35649 41245 35683
rect 41245 35649 41279 35683
rect 41279 35649 41288 35683
rect 41236 35640 41288 35649
rect 43076 35683 43128 35692
rect 43076 35649 43085 35683
rect 43085 35649 43119 35683
rect 43119 35649 43128 35683
rect 43076 35640 43128 35649
rect 43260 35640 43312 35692
rect 35900 35615 35952 35624
rect 35900 35581 35909 35615
rect 35909 35581 35943 35615
rect 35943 35581 35952 35615
rect 35900 35572 35952 35581
rect 37280 35615 37332 35624
rect 33416 35504 33468 35513
rect 34244 35504 34296 35556
rect 37280 35581 37289 35615
rect 37289 35581 37323 35615
rect 37323 35581 37332 35615
rect 37280 35572 37332 35581
rect 38016 35572 38068 35624
rect 27528 35479 27580 35488
rect 27528 35445 27537 35479
rect 27537 35445 27571 35479
rect 27571 35445 27580 35479
rect 27528 35436 27580 35445
rect 28264 35436 28316 35488
rect 30196 35479 30248 35488
rect 30196 35445 30205 35479
rect 30205 35445 30239 35479
rect 30239 35445 30248 35479
rect 30196 35436 30248 35445
rect 33048 35479 33100 35488
rect 33048 35445 33057 35479
rect 33057 35445 33091 35479
rect 33091 35445 33100 35479
rect 37004 35504 37056 35556
rect 33048 35436 33100 35445
rect 34612 35436 34664 35488
rect 36544 35436 36596 35488
rect 39212 35504 39264 35556
rect 39120 35436 39172 35488
rect 41880 35436 41932 35488
rect 43904 35436 43956 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 4712 35275 4764 35284
rect 4712 35241 4721 35275
rect 4721 35241 4755 35275
rect 4755 35241 4764 35275
rect 4712 35232 4764 35241
rect 5264 35275 5316 35284
rect 5264 35241 5273 35275
rect 5273 35241 5307 35275
rect 5307 35241 5316 35275
rect 5264 35232 5316 35241
rect 6000 35275 6052 35284
rect 6000 35241 6009 35275
rect 6009 35241 6043 35275
rect 6043 35241 6052 35275
rect 6000 35232 6052 35241
rect 13084 35275 13136 35284
rect 13084 35241 13093 35275
rect 13093 35241 13127 35275
rect 13127 35241 13136 35275
rect 13084 35232 13136 35241
rect 14004 35275 14056 35284
rect 14004 35241 14013 35275
rect 14013 35241 14047 35275
rect 14047 35241 14056 35275
rect 14004 35232 14056 35241
rect 20720 35275 20772 35284
rect 6092 35164 6144 35216
rect 7932 35164 7984 35216
rect 8944 35164 8996 35216
rect 9312 35164 9364 35216
rect 10692 35164 10744 35216
rect 11704 35207 11756 35216
rect 11704 35173 11713 35207
rect 11713 35173 11747 35207
rect 11747 35173 11756 35207
rect 11704 35164 11756 35173
rect 13728 35164 13780 35216
rect 15660 35164 15712 35216
rect 17684 35164 17736 35216
rect 19156 35164 19208 35216
rect 20720 35241 20729 35275
rect 20729 35241 20763 35275
rect 20763 35241 20772 35275
rect 20720 35232 20772 35241
rect 21272 35275 21324 35284
rect 21272 35241 21281 35275
rect 21281 35241 21315 35275
rect 21315 35241 21324 35275
rect 21272 35232 21324 35241
rect 21364 35232 21416 35284
rect 22192 35232 22244 35284
rect 19892 35164 19944 35216
rect 24308 35207 24360 35216
rect 24308 35173 24317 35207
rect 24317 35173 24351 35207
rect 24351 35173 24360 35207
rect 24308 35164 24360 35173
rect 26976 35232 27028 35284
rect 29092 35232 29144 35284
rect 30472 35232 30524 35284
rect 26424 35164 26476 35216
rect 29552 35164 29604 35216
rect 29736 35164 29788 35216
rect 30196 35164 30248 35216
rect 33048 35232 33100 35284
rect 33416 35232 33468 35284
rect 37280 35275 37332 35284
rect 34704 35164 34756 35216
rect 35348 35207 35400 35216
rect 35348 35173 35357 35207
rect 35357 35173 35391 35207
rect 35391 35173 35400 35207
rect 35348 35164 35400 35173
rect 37280 35241 37289 35275
rect 37289 35241 37323 35275
rect 37323 35241 37332 35275
rect 37280 35232 37332 35241
rect 41236 35275 41288 35284
rect 41236 35241 41245 35275
rect 41245 35241 41279 35275
rect 41279 35241 41288 35275
rect 41236 35232 41288 35241
rect 35716 35164 35768 35216
rect 4160 35096 4212 35148
rect 11888 35096 11940 35148
rect 17224 35096 17276 35148
rect 22836 35096 22888 35148
rect 23204 35096 23256 35148
rect 29368 35139 29420 35148
rect 4068 35028 4120 35080
rect 6460 35028 6512 35080
rect 7932 35071 7984 35080
rect 7932 35037 7941 35071
rect 7941 35037 7975 35071
rect 7975 35037 7984 35071
rect 7932 35028 7984 35037
rect 8576 35028 8628 35080
rect 10416 35071 10468 35080
rect 10416 35037 10425 35071
rect 10425 35037 10459 35071
rect 10459 35037 10468 35071
rect 10416 35028 10468 35037
rect 12716 35071 12768 35080
rect 12716 35037 12725 35071
rect 12725 35037 12759 35071
rect 12759 35037 12768 35071
rect 12716 35028 12768 35037
rect 16580 35028 16632 35080
rect 18420 35071 18472 35080
rect 18420 35037 18429 35071
rect 18429 35037 18463 35071
rect 18463 35037 18472 35071
rect 18420 35028 18472 35037
rect 20536 35028 20588 35080
rect 21824 35028 21876 35080
rect 24216 35071 24268 35080
rect 24216 35037 24225 35071
rect 24225 35037 24259 35071
rect 24259 35037 24268 35071
rect 24216 35028 24268 35037
rect 26608 35071 26660 35080
rect 26608 35037 26617 35071
rect 26617 35037 26651 35071
rect 26651 35037 26660 35071
rect 26608 35028 26660 35037
rect 26884 35071 26936 35080
rect 26884 35037 26893 35071
rect 26893 35037 26927 35071
rect 26927 35037 26936 35071
rect 26884 35028 26936 35037
rect 29368 35105 29377 35139
rect 29377 35105 29411 35139
rect 29411 35105 29420 35139
rect 29368 35096 29420 35105
rect 30564 35096 30616 35148
rect 31852 35096 31904 35148
rect 38200 35164 38252 35216
rect 39212 35207 39264 35216
rect 39212 35173 39221 35207
rect 39221 35173 39255 35207
rect 39255 35173 39264 35207
rect 39212 35164 39264 35173
rect 41880 35207 41932 35216
rect 41880 35173 41889 35207
rect 41889 35173 41923 35207
rect 41923 35173 41932 35207
rect 41880 35164 41932 35173
rect 40592 35139 40644 35148
rect 40592 35105 40601 35139
rect 40601 35105 40635 35139
rect 40635 35105 40644 35139
rect 40592 35096 40644 35105
rect 43260 35139 43312 35148
rect 43260 35105 43269 35139
rect 43269 35105 43303 35139
rect 43303 35105 43312 35139
rect 43260 35096 43312 35105
rect 11152 34960 11204 35012
rect 16028 35003 16080 35012
rect 16028 34969 16037 35003
rect 16037 34969 16071 35003
rect 16071 34969 16080 35003
rect 16028 34960 16080 34969
rect 25780 34960 25832 35012
rect 29552 35028 29604 35080
rect 32220 35071 32272 35080
rect 32220 35037 32229 35071
rect 32229 35037 32263 35071
rect 32263 35037 32272 35071
rect 32220 35028 32272 35037
rect 33784 35071 33836 35080
rect 33784 35037 33793 35071
rect 33793 35037 33827 35071
rect 33827 35037 33836 35071
rect 33784 35028 33836 35037
rect 35624 35071 35676 35080
rect 32864 34960 32916 35012
rect 35624 35037 35633 35071
rect 35633 35037 35667 35071
rect 35667 35037 35676 35071
rect 35624 35028 35676 35037
rect 39120 35071 39172 35080
rect 39120 35037 39129 35071
rect 39129 35037 39163 35071
rect 39163 35037 39172 35071
rect 39120 35028 39172 35037
rect 40868 35028 40920 35080
rect 41788 35071 41840 35080
rect 41788 35037 41797 35071
rect 41797 35037 41831 35071
rect 41831 35037 41840 35071
rect 41788 35028 41840 35037
rect 42892 35028 42944 35080
rect 38844 35003 38896 35012
rect 38844 34969 38853 35003
rect 38853 34969 38887 35003
rect 38887 34969 38896 35003
rect 38844 34960 38896 34969
rect 41144 34960 41196 35012
rect 7196 34892 7248 34944
rect 8852 34935 8904 34944
rect 8852 34901 8861 34935
rect 8861 34901 8895 34935
rect 8895 34901 8904 34935
rect 8852 34892 8904 34901
rect 10876 34935 10928 34944
rect 10876 34901 10885 34935
rect 10885 34901 10919 34935
rect 10919 34901 10928 34935
rect 10876 34892 10928 34901
rect 16212 34892 16264 34944
rect 17408 34892 17460 34944
rect 18512 34892 18564 34944
rect 23756 34935 23808 34944
rect 23756 34901 23765 34935
rect 23765 34901 23799 34935
rect 23799 34901 23808 34935
rect 23756 34892 23808 34901
rect 26332 34935 26384 34944
rect 26332 34901 26341 34935
rect 26341 34901 26375 34935
rect 26375 34901 26384 34935
rect 26332 34892 26384 34901
rect 30012 34892 30064 34944
rect 33324 34935 33376 34944
rect 33324 34901 33333 34935
rect 33333 34901 33367 34935
rect 33367 34901 33376 34935
rect 33324 34892 33376 34901
rect 33968 34892 34020 34944
rect 36084 34892 36136 34944
rect 42524 34892 42576 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 8208 34688 8260 34740
rect 9312 34731 9364 34740
rect 9312 34697 9321 34731
rect 9321 34697 9355 34731
rect 9355 34697 9364 34731
rect 9312 34688 9364 34697
rect 10876 34688 10928 34740
rect 12900 34688 12952 34740
rect 10416 34663 10468 34672
rect 10416 34629 10425 34663
rect 10425 34629 10459 34663
rect 10459 34629 10468 34663
rect 10416 34620 10468 34629
rect 11152 34663 11204 34672
rect 11152 34629 11161 34663
rect 11161 34629 11195 34663
rect 11195 34629 11204 34663
rect 11152 34620 11204 34629
rect 7932 34552 7984 34604
rect 8760 34552 8812 34604
rect 9496 34552 9548 34604
rect 13636 34552 13688 34604
rect 15292 34688 15344 34740
rect 16580 34731 16632 34740
rect 16580 34697 16589 34731
rect 16589 34697 16623 34731
rect 16623 34697 16632 34731
rect 16580 34688 16632 34697
rect 17224 34688 17276 34740
rect 20260 34731 20312 34740
rect 20260 34697 20269 34731
rect 20269 34697 20303 34731
rect 20303 34697 20312 34731
rect 20260 34688 20312 34697
rect 21272 34731 21324 34740
rect 21272 34697 21281 34731
rect 21281 34697 21315 34731
rect 21315 34697 21324 34731
rect 22836 34731 22888 34740
rect 21272 34688 21324 34697
rect 15568 34620 15620 34672
rect 19156 34663 19208 34672
rect 19156 34629 19165 34663
rect 19165 34629 19199 34663
rect 19199 34629 19208 34663
rect 19156 34620 19208 34629
rect 22008 34620 22060 34672
rect 22836 34697 22845 34731
rect 22845 34697 22879 34731
rect 22879 34697 22888 34731
rect 22836 34688 22888 34697
rect 24308 34688 24360 34740
rect 23296 34620 23348 34672
rect 23848 34620 23900 34672
rect 24032 34620 24084 34672
rect 29368 34688 29420 34740
rect 31852 34688 31904 34740
rect 33784 34688 33836 34740
rect 33968 34688 34020 34740
rect 35348 34688 35400 34740
rect 37004 34688 37056 34740
rect 39212 34688 39264 34740
rect 41420 34731 41472 34740
rect 41420 34697 41429 34731
rect 41429 34697 41463 34731
rect 41463 34697 41472 34731
rect 41420 34688 41472 34697
rect 41880 34688 41932 34740
rect 26608 34620 26660 34672
rect 27252 34663 27304 34672
rect 27252 34629 27261 34663
rect 27261 34629 27295 34663
rect 27295 34629 27304 34663
rect 27252 34620 27304 34629
rect 29552 34620 29604 34672
rect 29736 34663 29788 34672
rect 29736 34629 29745 34663
rect 29745 34629 29779 34663
rect 29779 34629 29788 34663
rect 29736 34620 29788 34629
rect 16028 34595 16080 34604
rect 16028 34561 16037 34595
rect 16037 34561 16071 34595
rect 16071 34561 16080 34595
rect 16028 34552 16080 34561
rect 18420 34552 18472 34604
rect 24216 34552 24268 34604
rect 25872 34552 25924 34604
rect 30012 34552 30064 34604
rect 30840 34552 30892 34604
rect 31024 34595 31076 34604
rect 31024 34561 31033 34595
rect 31033 34561 31067 34595
rect 31067 34561 31076 34595
rect 31024 34552 31076 34561
rect 32680 34620 32732 34672
rect 32956 34620 33008 34672
rect 35624 34620 35676 34672
rect 35716 34663 35768 34672
rect 35716 34629 35725 34663
rect 35725 34629 35759 34663
rect 35759 34629 35768 34663
rect 35716 34620 35768 34629
rect 3332 34527 3384 34536
rect 3332 34493 3341 34527
rect 3341 34493 3375 34527
rect 3375 34493 3384 34527
rect 3332 34484 3384 34493
rect 4896 34484 4948 34536
rect 7288 34484 7340 34536
rect 12256 34484 12308 34536
rect 18236 34527 18288 34536
rect 18236 34493 18245 34527
rect 18245 34493 18279 34527
rect 18279 34493 18288 34527
rect 18236 34484 18288 34493
rect 18512 34527 18564 34536
rect 18512 34493 18521 34527
rect 18521 34493 18555 34527
rect 18555 34493 18564 34527
rect 18512 34484 18564 34493
rect 20260 34484 20312 34536
rect 4712 34348 4764 34400
rect 5356 34391 5408 34400
rect 5356 34357 5365 34391
rect 5365 34357 5399 34391
rect 5399 34357 5408 34391
rect 5356 34348 5408 34357
rect 6092 34391 6144 34400
rect 6092 34357 6101 34391
rect 6101 34357 6135 34391
rect 6135 34357 6144 34391
rect 6092 34348 6144 34357
rect 6460 34391 6512 34400
rect 6460 34357 6469 34391
rect 6469 34357 6503 34391
rect 6503 34357 6512 34391
rect 6460 34348 6512 34357
rect 7840 34348 7892 34400
rect 8300 34348 8352 34400
rect 9864 34416 9916 34468
rect 11796 34416 11848 34468
rect 13084 34416 13136 34468
rect 13728 34416 13780 34468
rect 15292 34416 15344 34468
rect 20076 34416 20128 34468
rect 20536 34459 20588 34468
rect 20536 34425 20545 34459
rect 20545 34425 20579 34459
rect 20579 34425 20588 34459
rect 20536 34416 20588 34425
rect 11888 34391 11940 34400
rect 11888 34357 11897 34391
rect 11897 34357 11931 34391
rect 11931 34357 11940 34391
rect 11888 34348 11940 34357
rect 12348 34348 12400 34400
rect 14188 34391 14240 34400
rect 14188 34357 14197 34391
rect 14197 34357 14231 34391
rect 14231 34357 14240 34391
rect 14188 34348 14240 34357
rect 21088 34348 21140 34400
rect 23756 34484 23808 34536
rect 26148 34527 26200 34536
rect 26148 34493 26157 34527
rect 26157 34493 26191 34527
rect 26191 34493 26200 34527
rect 26148 34484 26200 34493
rect 21824 34459 21876 34468
rect 21824 34425 21833 34459
rect 21833 34425 21867 34459
rect 21867 34425 21876 34459
rect 21824 34416 21876 34425
rect 21916 34459 21968 34468
rect 21916 34425 21925 34459
rect 21925 34425 21959 34459
rect 21959 34425 21968 34459
rect 21916 34416 21968 34425
rect 23848 34416 23900 34468
rect 26884 34416 26936 34468
rect 25596 34348 25648 34400
rect 26424 34391 26476 34400
rect 26424 34357 26433 34391
rect 26433 34357 26467 34391
rect 26467 34357 26476 34391
rect 26424 34348 26476 34357
rect 29552 34484 29604 34536
rect 30196 34416 30248 34468
rect 32220 34552 32272 34604
rect 28908 34348 28960 34400
rect 29184 34348 29236 34400
rect 31852 34348 31904 34400
rect 33600 34416 33652 34468
rect 35532 34484 35584 34536
rect 40592 34620 40644 34672
rect 38844 34595 38896 34604
rect 38844 34561 38853 34595
rect 38853 34561 38887 34595
rect 38887 34561 38896 34595
rect 38844 34552 38896 34561
rect 38936 34552 38988 34604
rect 36820 34484 36872 34536
rect 41420 34484 41472 34536
rect 37004 34348 37056 34400
rect 38844 34416 38896 34468
rect 39488 34459 39540 34468
rect 37924 34391 37976 34400
rect 37924 34357 37933 34391
rect 37933 34357 37967 34391
rect 37967 34357 37976 34391
rect 37924 34348 37976 34357
rect 38200 34391 38252 34400
rect 38200 34357 38209 34391
rect 38209 34357 38243 34391
rect 38243 34357 38252 34391
rect 38200 34348 38252 34357
rect 38660 34391 38712 34400
rect 38660 34357 38669 34391
rect 38669 34357 38703 34391
rect 38703 34357 38712 34391
rect 39488 34425 39497 34459
rect 39497 34425 39531 34459
rect 39531 34425 39540 34459
rect 39488 34416 39540 34425
rect 42616 34688 42668 34740
rect 43260 34688 43312 34740
rect 42524 34595 42576 34604
rect 42524 34561 42533 34595
rect 42533 34561 42567 34595
rect 42567 34561 42576 34595
rect 42524 34552 42576 34561
rect 42800 34595 42852 34604
rect 42800 34561 42809 34595
rect 42809 34561 42843 34595
rect 42843 34561 42852 34595
rect 42800 34552 42852 34561
rect 44364 34416 44416 34468
rect 38660 34348 38712 34357
rect 40776 34348 40828 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 7196 34144 7248 34196
rect 8576 34144 8628 34196
rect 8852 34144 8904 34196
rect 12256 34187 12308 34196
rect 12256 34153 12265 34187
rect 12265 34153 12299 34187
rect 12299 34153 12308 34187
rect 12256 34144 12308 34153
rect 14556 34144 14608 34196
rect 17408 34187 17460 34196
rect 17408 34153 17417 34187
rect 17417 34153 17451 34187
rect 17451 34153 17460 34187
rect 17408 34144 17460 34153
rect 18420 34187 18472 34196
rect 18420 34153 18429 34187
rect 18429 34153 18463 34187
rect 18463 34153 18472 34187
rect 18420 34144 18472 34153
rect 21824 34144 21876 34196
rect 24124 34144 24176 34196
rect 24216 34144 24268 34196
rect 25872 34144 25924 34196
rect 26608 34144 26660 34196
rect 26792 34144 26844 34196
rect 29368 34144 29420 34196
rect 30840 34187 30892 34196
rect 30840 34153 30849 34187
rect 30849 34153 30883 34187
rect 30883 34153 30892 34187
rect 30840 34144 30892 34153
rect 32220 34144 32272 34196
rect 32680 34187 32732 34196
rect 32680 34153 32689 34187
rect 32689 34153 32723 34187
rect 32723 34153 32732 34187
rect 32680 34144 32732 34153
rect 32956 34187 33008 34196
rect 32956 34153 32965 34187
rect 32965 34153 32999 34187
rect 32999 34153 33008 34187
rect 32956 34144 33008 34153
rect 34796 34144 34848 34196
rect 38660 34187 38712 34196
rect 38660 34153 38669 34187
rect 38669 34153 38703 34187
rect 38703 34153 38712 34187
rect 38660 34144 38712 34153
rect 39120 34187 39172 34196
rect 39120 34153 39129 34187
rect 39129 34153 39163 34187
rect 39163 34153 39172 34187
rect 39120 34144 39172 34153
rect 39396 34187 39448 34196
rect 39396 34153 39405 34187
rect 39405 34153 39439 34187
rect 39439 34153 39448 34187
rect 39396 34144 39448 34153
rect 41788 34187 41840 34196
rect 41788 34153 41797 34187
rect 41797 34153 41831 34187
rect 41831 34153 41840 34187
rect 41788 34144 41840 34153
rect 8300 34119 8352 34128
rect 8300 34085 8309 34119
rect 8309 34085 8343 34119
rect 8343 34085 8352 34119
rect 8300 34076 8352 34085
rect 9312 34076 9364 34128
rect 9588 34076 9640 34128
rect 11888 34076 11940 34128
rect 15292 34076 15344 34128
rect 19432 34119 19484 34128
rect 19432 34085 19441 34119
rect 19441 34085 19475 34119
rect 19475 34085 19484 34119
rect 19432 34076 19484 34085
rect 21272 34076 21324 34128
rect 21916 34119 21968 34128
rect 21916 34085 21925 34119
rect 21925 34085 21959 34119
rect 21959 34085 21968 34119
rect 21916 34076 21968 34085
rect 26884 34119 26936 34128
rect 26884 34085 26893 34119
rect 26893 34085 26927 34119
rect 26927 34085 26936 34119
rect 26884 34076 26936 34085
rect 29276 34119 29328 34128
rect 29276 34085 29285 34119
rect 29285 34085 29319 34119
rect 29319 34085 29328 34119
rect 29276 34076 29328 34085
rect 36820 34119 36872 34128
rect 36820 34085 36829 34119
rect 36829 34085 36863 34119
rect 36863 34085 36872 34119
rect 36820 34076 36872 34085
rect 37004 34076 37056 34128
rect 37832 34076 37884 34128
rect 40592 34119 40644 34128
rect 40592 34085 40601 34119
rect 40601 34085 40635 34119
rect 40635 34085 40644 34119
rect 40592 34076 40644 34085
rect 41144 34119 41196 34128
rect 41144 34085 41153 34119
rect 41153 34085 41187 34119
rect 41187 34085 41196 34119
rect 41144 34076 41196 34085
rect 42800 34076 42852 34128
rect 43536 34119 43588 34128
rect 43536 34085 43545 34119
rect 43545 34085 43579 34119
rect 43579 34085 43588 34119
rect 43536 34076 43588 34085
rect 4712 34051 4764 34060
rect 4712 34017 4721 34051
rect 4721 34017 4755 34051
rect 4755 34017 4764 34051
rect 4712 34008 4764 34017
rect 5172 34008 5224 34060
rect 5356 34008 5408 34060
rect 6184 34008 6236 34060
rect 8024 34008 8076 34060
rect 8484 34008 8536 34060
rect 14188 34008 14240 34060
rect 16212 34051 16264 34060
rect 16212 34017 16221 34051
rect 16221 34017 16255 34051
rect 16255 34017 16264 34051
rect 16212 34008 16264 34017
rect 17132 34051 17184 34060
rect 17132 34017 17141 34051
rect 17141 34017 17175 34051
rect 17175 34017 17184 34051
rect 17132 34008 17184 34017
rect 17684 34051 17736 34060
rect 17684 34017 17693 34051
rect 17693 34017 17727 34051
rect 17727 34017 17736 34051
rect 17684 34008 17736 34017
rect 21640 34051 21692 34060
rect 21640 34017 21649 34051
rect 21649 34017 21683 34051
rect 21683 34017 21692 34051
rect 21640 34008 21692 34017
rect 22376 34008 22428 34060
rect 23112 34008 23164 34060
rect 24676 34008 24728 34060
rect 25412 34051 25464 34060
rect 4988 33983 5040 33992
rect 4988 33949 4997 33983
rect 4997 33949 5031 33983
rect 5031 33949 5040 33983
rect 4988 33940 5040 33949
rect 9772 33983 9824 33992
rect 9772 33949 9781 33983
rect 9781 33949 9815 33983
rect 9815 33949 9824 33983
rect 9772 33940 9824 33949
rect 9864 33940 9916 33992
rect 11336 33983 11388 33992
rect 11336 33949 11345 33983
rect 11345 33949 11379 33983
rect 11379 33949 11388 33983
rect 11336 33940 11388 33949
rect 19340 33983 19392 33992
rect 19340 33949 19349 33983
rect 19349 33949 19383 33983
rect 19383 33949 19392 33983
rect 19340 33940 19392 33949
rect 20996 33983 21048 33992
rect 20996 33949 21005 33983
rect 21005 33949 21039 33983
rect 21039 33949 21048 33983
rect 20996 33940 21048 33949
rect 23020 33940 23072 33992
rect 25412 34017 25456 34051
rect 25456 34017 25464 34051
rect 28540 34051 28592 34060
rect 25412 34008 25464 34017
rect 28540 34017 28549 34051
rect 28549 34017 28583 34051
rect 28583 34017 28592 34051
rect 28540 34008 28592 34017
rect 28816 34008 28868 34060
rect 29092 34051 29144 34060
rect 29092 34017 29101 34051
rect 29101 34017 29135 34051
rect 29135 34017 29144 34051
rect 29092 34008 29144 34017
rect 32128 34008 32180 34060
rect 33508 34008 33560 34060
rect 34428 34051 34480 34060
rect 34428 34017 34437 34051
rect 34437 34017 34471 34051
rect 34471 34017 34480 34051
rect 34428 34008 34480 34017
rect 36360 34051 36412 34060
rect 36360 34017 36369 34051
rect 36369 34017 36403 34051
rect 36403 34017 36412 34051
rect 36360 34008 36412 34017
rect 36544 34051 36596 34060
rect 36544 34017 36553 34051
rect 36553 34017 36587 34051
rect 36587 34017 36596 34051
rect 36544 34008 36596 34017
rect 41236 34008 41288 34060
rect 42248 34051 42300 34060
rect 42248 34017 42292 34051
rect 42292 34017 42300 34051
rect 42248 34008 42300 34017
rect 26792 33983 26844 33992
rect 26792 33949 26801 33983
rect 26801 33949 26835 33983
rect 26835 33949 26844 33983
rect 26792 33940 26844 33949
rect 27068 33983 27120 33992
rect 27068 33949 27077 33983
rect 27077 33949 27111 33983
rect 27111 33949 27120 33983
rect 27068 33940 27120 33949
rect 30380 33983 30432 33992
rect 30380 33949 30389 33983
rect 30389 33949 30423 33983
rect 30423 33949 30432 33983
rect 30380 33940 30432 33949
rect 37740 33983 37792 33992
rect 37740 33949 37749 33983
rect 37749 33949 37783 33983
rect 37783 33949 37792 33983
rect 37740 33940 37792 33949
rect 40868 33940 40920 33992
rect 41512 33940 41564 33992
rect 43076 33940 43128 33992
rect 19892 33915 19944 33924
rect 19892 33881 19901 33915
rect 19901 33881 19935 33915
rect 19935 33881 19944 33915
rect 19892 33872 19944 33881
rect 42892 33872 42944 33924
rect 4068 33804 4120 33856
rect 7288 33847 7340 33856
rect 7288 33813 7297 33847
rect 7297 33813 7331 33847
rect 7331 33813 7340 33847
rect 7288 33804 7340 33813
rect 12716 33804 12768 33856
rect 13268 33804 13320 33856
rect 13636 33804 13688 33856
rect 23848 33804 23900 33856
rect 29552 33847 29604 33856
rect 29552 33813 29561 33847
rect 29561 33813 29595 33847
rect 29595 33813 29604 33847
rect 29552 33804 29604 33813
rect 31852 33804 31904 33856
rect 33140 33804 33192 33856
rect 35532 33804 35584 33856
rect 42708 33847 42760 33856
rect 42708 33813 42717 33847
rect 42717 33813 42751 33847
rect 42751 33813 42760 33847
rect 42708 33804 42760 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 3332 33600 3384 33652
rect 6184 33643 6236 33652
rect 6184 33609 6193 33643
rect 6193 33609 6227 33643
rect 6227 33609 6236 33643
rect 6184 33600 6236 33609
rect 7288 33600 7340 33652
rect 8024 33643 8076 33652
rect 8024 33609 8033 33643
rect 8033 33609 8067 33643
rect 8067 33609 8076 33643
rect 8024 33600 8076 33609
rect 8392 33600 8444 33652
rect 9772 33600 9824 33652
rect 11336 33600 11388 33652
rect 14188 33600 14240 33652
rect 16212 33600 16264 33652
rect 16580 33643 16632 33652
rect 16580 33609 16589 33643
rect 16589 33609 16623 33643
rect 16623 33609 16632 33643
rect 16580 33600 16632 33609
rect 17132 33643 17184 33652
rect 17132 33609 17141 33643
rect 17141 33609 17175 33643
rect 17175 33609 17184 33643
rect 17132 33600 17184 33609
rect 19432 33600 19484 33652
rect 20996 33600 21048 33652
rect 21272 33643 21324 33652
rect 21272 33609 21281 33643
rect 21281 33609 21315 33643
rect 21315 33609 21324 33643
rect 21272 33600 21324 33609
rect 22376 33600 22428 33652
rect 24308 33600 24360 33652
rect 24676 33643 24728 33652
rect 24676 33609 24685 33643
rect 24685 33609 24719 33643
rect 24719 33609 24728 33643
rect 24676 33600 24728 33609
rect 25412 33643 25464 33652
rect 25412 33609 25421 33643
rect 25421 33609 25455 33643
rect 25455 33609 25464 33643
rect 25412 33600 25464 33609
rect 27528 33600 27580 33652
rect 28540 33600 28592 33652
rect 30380 33600 30432 33652
rect 33508 33643 33560 33652
rect 9496 33575 9548 33584
rect 9496 33541 9505 33575
rect 9505 33541 9539 33575
rect 9539 33541 9548 33575
rect 9496 33532 9548 33541
rect 9588 33532 9640 33584
rect 19340 33532 19392 33584
rect 26976 33532 27028 33584
rect 4988 33507 5040 33516
rect 4988 33473 4997 33507
rect 4997 33473 5031 33507
rect 5031 33473 5040 33507
rect 4988 33464 5040 33473
rect 13636 33507 13688 33516
rect 13636 33473 13645 33507
rect 13645 33473 13679 33507
rect 13679 33473 13688 33507
rect 13636 33464 13688 33473
rect 21088 33464 21140 33516
rect 23940 33464 23992 33516
rect 3700 33439 3752 33448
rect 3700 33405 3709 33439
rect 3709 33405 3743 33439
rect 3743 33405 3752 33439
rect 3700 33396 3752 33405
rect 3976 33439 4028 33448
rect 3976 33405 3985 33439
rect 3985 33405 4019 33439
rect 4019 33405 4028 33439
rect 3976 33396 4028 33405
rect 6460 33396 6512 33448
rect 6828 33439 6880 33448
rect 6828 33405 6837 33439
rect 6837 33405 6871 33439
rect 6871 33405 6880 33439
rect 6828 33396 6880 33405
rect 9588 33396 9640 33448
rect 6092 33328 6144 33380
rect 7840 33328 7892 33380
rect 8852 33328 8904 33380
rect 11520 33396 11572 33448
rect 13360 33396 13412 33448
rect 13544 33396 13596 33448
rect 14648 33439 14700 33448
rect 14648 33405 14657 33439
rect 14657 33405 14691 33439
rect 14691 33405 14700 33439
rect 14648 33396 14700 33405
rect 18604 33439 18656 33448
rect 18604 33405 18613 33439
rect 18613 33405 18647 33439
rect 18647 33405 18656 33439
rect 18604 33396 18656 33405
rect 20904 33396 20956 33448
rect 23388 33439 23440 33448
rect 23388 33405 23397 33439
rect 23397 33405 23431 33439
rect 23431 33405 23440 33439
rect 23388 33396 23440 33405
rect 23848 33396 23900 33448
rect 24124 33439 24176 33448
rect 24124 33405 24133 33439
rect 24133 33405 24167 33439
rect 24167 33405 24176 33439
rect 24124 33396 24176 33405
rect 29644 33532 29696 33584
rect 26056 33439 26108 33448
rect 26056 33405 26065 33439
rect 26065 33405 26099 33439
rect 26099 33405 26108 33439
rect 26056 33396 26108 33405
rect 29460 33464 29512 33516
rect 33508 33609 33517 33643
rect 33517 33609 33551 33643
rect 33551 33609 33560 33643
rect 33508 33600 33560 33609
rect 34428 33643 34480 33652
rect 34428 33609 34437 33643
rect 34437 33609 34471 33643
rect 34471 33609 34480 33643
rect 34428 33600 34480 33609
rect 36360 33600 36412 33652
rect 37832 33643 37884 33652
rect 37832 33609 37841 33643
rect 37841 33609 37875 33643
rect 37875 33609 37884 33643
rect 37832 33600 37884 33609
rect 37924 33600 37976 33652
rect 38936 33600 38988 33652
rect 40592 33600 40644 33652
rect 41512 33643 41564 33652
rect 41512 33609 41521 33643
rect 41521 33609 41555 33643
rect 41555 33609 41564 33643
rect 41512 33600 41564 33609
rect 42248 33643 42300 33652
rect 42248 33609 42257 33643
rect 42257 33609 42291 33643
rect 42291 33609 42300 33643
rect 42248 33600 42300 33609
rect 31024 33507 31076 33516
rect 31024 33473 31033 33507
rect 31033 33473 31067 33507
rect 31067 33473 31076 33507
rect 31024 33464 31076 33473
rect 32956 33532 33008 33584
rect 33232 33532 33284 33584
rect 34612 33532 34664 33584
rect 32772 33507 32824 33516
rect 32772 33473 32781 33507
rect 32781 33473 32815 33507
rect 32815 33473 32824 33507
rect 32772 33464 32824 33473
rect 29184 33396 29236 33448
rect 11888 33371 11940 33380
rect 11888 33337 11897 33371
rect 11897 33337 11931 33371
rect 11931 33337 11940 33371
rect 11888 33328 11940 33337
rect 13728 33328 13780 33380
rect 15476 33328 15528 33380
rect 17684 33328 17736 33380
rect 18512 33328 18564 33380
rect 18696 33328 18748 33380
rect 19156 33328 19208 33380
rect 4712 33260 4764 33312
rect 8484 33260 8536 33312
rect 12440 33260 12492 33312
rect 20904 33303 20956 33312
rect 20904 33269 20913 33303
rect 20913 33269 20947 33303
rect 20947 33269 20956 33303
rect 20904 33260 20956 33269
rect 21272 33260 21324 33312
rect 25964 33328 26016 33380
rect 26884 33328 26936 33380
rect 27712 33328 27764 33380
rect 23756 33303 23808 33312
rect 23756 33269 23765 33303
rect 23765 33269 23799 33303
rect 23799 33269 23808 33303
rect 23756 33260 23808 33269
rect 29736 33260 29788 33312
rect 34060 33396 34112 33448
rect 37740 33464 37792 33516
rect 39396 33532 39448 33584
rect 42892 33532 42944 33584
rect 39212 33464 39264 33516
rect 39488 33507 39540 33516
rect 39488 33473 39497 33507
rect 39497 33473 39531 33507
rect 39531 33473 39540 33507
rect 39488 33464 39540 33473
rect 40776 33464 40828 33516
rect 42708 33507 42760 33516
rect 42708 33473 42717 33507
rect 42717 33473 42751 33507
rect 42751 33473 42760 33507
rect 42708 33464 42760 33473
rect 42800 33464 42852 33516
rect 44548 33507 44600 33516
rect 44548 33473 44557 33507
rect 44557 33473 44591 33507
rect 44591 33473 44600 33507
rect 44548 33464 44600 33473
rect 35256 33396 35308 33448
rect 30564 33328 30616 33380
rect 32128 33303 32180 33312
rect 32128 33269 32137 33303
rect 32137 33269 32171 33303
rect 32171 33269 32180 33303
rect 32128 33260 32180 33269
rect 35900 33328 35952 33380
rect 36544 33396 36596 33448
rect 36912 33328 36964 33380
rect 38936 33371 38988 33380
rect 38936 33337 38945 33371
rect 38945 33337 38979 33371
rect 38979 33337 38988 33371
rect 38936 33328 38988 33337
rect 40684 33371 40736 33380
rect 40684 33337 40693 33371
rect 40693 33337 40727 33371
rect 40727 33337 40736 33371
rect 42800 33371 42852 33380
rect 40684 33328 40736 33337
rect 42800 33337 42809 33371
rect 42809 33337 42843 33371
rect 42843 33337 42852 33371
rect 42800 33328 42852 33337
rect 43536 33328 43588 33380
rect 44088 33328 44140 33380
rect 33048 33260 33100 33312
rect 33416 33260 33468 33312
rect 35256 33260 35308 33312
rect 38108 33260 38160 33312
rect 39580 33260 39632 33312
rect 43996 33303 44048 33312
rect 43996 33269 44005 33303
rect 44005 33269 44039 33303
rect 44039 33269 44048 33303
rect 44364 33371 44416 33380
rect 44364 33337 44373 33371
rect 44373 33337 44407 33371
rect 44407 33337 44416 33371
rect 44364 33328 44416 33337
rect 43996 33260 44048 33269
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 4068 33056 4120 33108
rect 4988 33056 5040 33108
rect 7840 33099 7892 33108
rect 7840 33065 7849 33099
rect 7849 33065 7883 33099
rect 7883 33065 7892 33099
rect 7840 33056 7892 33065
rect 8484 33056 8536 33108
rect 9588 33056 9640 33108
rect 12348 33099 12400 33108
rect 12348 33065 12357 33099
rect 12357 33065 12391 33099
rect 12391 33065 12400 33099
rect 12348 33056 12400 33065
rect 13268 33099 13320 33108
rect 13268 33065 13277 33099
rect 13277 33065 13311 33099
rect 13311 33065 13320 33099
rect 13268 33056 13320 33065
rect 13452 33056 13504 33108
rect 14648 33099 14700 33108
rect 3976 32988 4028 33040
rect 3516 32920 3568 32972
rect 11428 32988 11480 33040
rect 11888 32988 11940 33040
rect 5172 32920 5224 32972
rect 6368 32963 6420 32972
rect 6368 32929 6377 32963
rect 6377 32929 6411 32963
rect 6411 32929 6420 32963
rect 6368 32920 6420 32929
rect 6828 32963 6880 32972
rect 6828 32929 6837 32963
rect 6837 32929 6871 32963
rect 6871 32929 6880 32963
rect 6828 32920 6880 32929
rect 13452 32963 13504 32972
rect 13452 32929 13461 32963
rect 13461 32929 13495 32963
rect 13495 32929 13504 32963
rect 13452 32920 13504 32929
rect 14648 33065 14657 33099
rect 14657 33065 14691 33099
rect 14691 33065 14700 33099
rect 14648 33056 14700 33065
rect 18604 33099 18656 33108
rect 18604 33065 18613 33099
rect 18613 33065 18647 33099
rect 18647 33065 18656 33099
rect 18604 33056 18656 33065
rect 19064 33099 19116 33108
rect 19064 33065 19073 33099
rect 19073 33065 19107 33099
rect 19107 33065 19116 33099
rect 20260 33099 20312 33108
rect 19064 33056 19116 33065
rect 15476 32988 15528 33040
rect 17408 32988 17460 33040
rect 18696 32988 18748 33040
rect 20260 33065 20269 33099
rect 20269 33065 20303 33099
rect 20303 33065 20312 33099
rect 20260 33056 20312 33065
rect 21640 33056 21692 33108
rect 22376 33056 22428 33108
rect 23480 33056 23532 33108
rect 19340 33031 19392 33040
rect 19340 32997 19349 33031
rect 19349 32997 19383 33031
rect 19383 32997 19392 33031
rect 19340 32988 19392 32997
rect 23296 32988 23348 33040
rect 26792 33056 26844 33108
rect 27712 33056 27764 33108
rect 29552 33056 29604 33108
rect 30656 33031 30708 33040
rect 30656 32997 30665 33031
rect 30665 32997 30699 33031
rect 30699 32997 30708 33031
rect 30656 32988 30708 32997
rect 32772 33056 32824 33108
rect 33048 33099 33100 33108
rect 33048 33065 33057 33099
rect 33057 33065 33091 33099
rect 33091 33065 33100 33099
rect 33048 33056 33100 33065
rect 33324 33056 33376 33108
rect 34152 33056 34204 33108
rect 38384 33056 38436 33108
rect 39856 33056 39908 33108
rect 42708 33056 42760 33108
rect 43076 33099 43128 33108
rect 32404 33031 32456 33040
rect 32404 32997 32413 33031
rect 32413 32997 32447 33031
rect 32447 32997 32456 33031
rect 32404 32988 32456 32997
rect 33508 32988 33560 33040
rect 36912 33031 36964 33040
rect 36912 32997 36921 33031
rect 36921 32997 36955 33031
rect 36955 32997 36964 33031
rect 36912 32988 36964 32997
rect 39028 33031 39080 33040
rect 39028 32997 39037 33031
rect 39037 32997 39071 33031
rect 39071 32997 39080 33031
rect 39028 32988 39080 32997
rect 40592 33031 40644 33040
rect 40592 32997 40601 33031
rect 40601 32997 40635 33031
rect 40635 32997 40644 33031
rect 40592 32988 40644 32997
rect 42800 33031 42852 33040
rect 42800 32997 42809 33031
rect 42809 32997 42843 33031
rect 42843 32997 42852 33031
rect 42800 32988 42852 32997
rect 43076 33065 43085 33099
rect 43085 33065 43119 33099
rect 43119 33065 43128 33099
rect 43076 33056 43128 33065
rect 44364 33056 44416 33108
rect 6276 32852 6328 32904
rect 7472 32895 7524 32904
rect 7472 32861 7481 32895
rect 7481 32861 7515 32895
rect 7515 32861 7524 32895
rect 7472 32852 7524 32861
rect 10416 32852 10468 32904
rect 11888 32852 11940 32904
rect 13544 32852 13596 32904
rect 15292 32895 15344 32904
rect 15292 32861 15301 32895
rect 15301 32861 15335 32895
rect 15335 32861 15344 32895
rect 15292 32852 15344 32861
rect 19892 32895 19944 32904
rect 3240 32716 3292 32768
rect 3976 32716 4028 32768
rect 5172 32759 5224 32768
rect 5172 32725 5181 32759
rect 5181 32725 5215 32759
rect 5215 32725 5224 32759
rect 5172 32716 5224 32725
rect 12992 32759 13044 32768
rect 12992 32725 13001 32759
rect 13001 32725 13035 32759
rect 13035 32725 13044 32759
rect 12992 32716 13044 32725
rect 17316 32759 17368 32768
rect 17316 32725 17325 32759
rect 17325 32725 17359 32759
rect 17359 32725 17368 32759
rect 19892 32861 19901 32895
rect 19901 32861 19935 32895
rect 19935 32861 19944 32895
rect 19892 32852 19944 32861
rect 20444 32852 20496 32904
rect 22100 32920 22152 32972
rect 24124 32920 24176 32972
rect 25596 32920 25648 32972
rect 22284 32852 22336 32904
rect 22836 32852 22888 32904
rect 23480 32852 23532 32904
rect 26240 32920 26292 32972
rect 28080 32920 28132 32972
rect 29184 32963 29236 32972
rect 29184 32929 29193 32963
rect 29193 32929 29227 32963
rect 29227 32929 29236 32963
rect 29184 32920 29236 32929
rect 29368 32963 29420 32972
rect 29368 32929 29377 32963
rect 29377 32929 29411 32963
rect 29411 32929 29420 32963
rect 29368 32920 29420 32929
rect 37740 32963 37792 32972
rect 37740 32929 37749 32963
rect 37749 32929 37783 32963
rect 37783 32929 37792 32963
rect 37740 32920 37792 32929
rect 38752 32920 38804 32972
rect 43352 32920 43404 32972
rect 43812 32920 43864 32972
rect 26332 32852 26384 32904
rect 19340 32784 19392 32836
rect 26700 32784 26752 32836
rect 29000 32784 29052 32836
rect 29552 32895 29604 32904
rect 29552 32861 29561 32895
rect 29561 32861 29595 32895
rect 29595 32861 29604 32895
rect 29552 32852 29604 32861
rect 30748 32852 30800 32904
rect 32312 32852 32364 32904
rect 33968 32895 34020 32904
rect 33968 32861 33977 32895
rect 33977 32861 34011 32895
rect 34011 32861 34020 32895
rect 33968 32852 34020 32861
rect 34244 32895 34296 32904
rect 34244 32861 34253 32895
rect 34253 32861 34287 32895
rect 34287 32861 34296 32895
rect 34244 32852 34296 32861
rect 35532 32895 35584 32904
rect 35532 32861 35541 32895
rect 35541 32861 35575 32895
rect 35575 32861 35584 32895
rect 35532 32852 35584 32861
rect 35808 32895 35860 32904
rect 35808 32861 35817 32895
rect 35817 32861 35851 32895
rect 35851 32861 35860 32895
rect 35808 32852 35860 32861
rect 38936 32895 38988 32904
rect 38936 32861 38945 32895
rect 38945 32861 38979 32895
rect 38979 32861 38988 32895
rect 38936 32852 38988 32861
rect 41236 32852 41288 32904
rect 43996 32852 44048 32904
rect 21364 32759 21416 32768
rect 17316 32716 17368 32725
rect 21364 32725 21373 32759
rect 21373 32725 21407 32759
rect 21407 32725 21416 32759
rect 21364 32716 21416 32725
rect 24124 32759 24176 32768
rect 24124 32725 24133 32759
rect 24133 32725 24167 32759
rect 24167 32725 24176 32759
rect 24124 32716 24176 32725
rect 25228 32759 25280 32768
rect 25228 32725 25237 32759
rect 25237 32725 25271 32759
rect 25271 32725 25280 32759
rect 25228 32716 25280 32725
rect 26516 32716 26568 32768
rect 26608 32716 26660 32768
rect 28816 32716 28868 32768
rect 29092 32716 29144 32768
rect 29920 32759 29972 32768
rect 29920 32725 29929 32759
rect 29929 32725 29963 32759
rect 29963 32725 29972 32759
rect 29920 32716 29972 32725
rect 33140 32784 33192 32836
rect 33784 32784 33836 32836
rect 36544 32827 36596 32836
rect 36544 32793 36553 32827
rect 36553 32793 36587 32827
rect 36587 32793 36596 32827
rect 36544 32784 36596 32793
rect 39212 32784 39264 32836
rect 35624 32716 35676 32768
rect 36728 32716 36780 32768
rect 38844 32716 38896 32768
rect 42064 32759 42116 32768
rect 42064 32725 42073 32759
rect 42073 32725 42107 32759
rect 42107 32725 42116 32759
rect 42064 32716 42116 32725
rect 44088 32716 44140 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 3240 32555 3292 32564
rect 3240 32521 3249 32555
rect 3249 32521 3283 32555
rect 3283 32521 3292 32555
rect 3240 32512 3292 32521
rect 5172 32555 5224 32564
rect 5172 32521 5181 32555
rect 5181 32521 5215 32555
rect 5215 32521 5224 32555
rect 5172 32512 5224 32521
rect 6368 32512 6420 32564
rect 8852 32555 8904 32564
rect 8852 32521 8861 32555
rect 8861 32521 8895 32555
rect 8895 32521 8904 32555
rect 8852 32512 8904 32521
rect 15476 32512 15528 32564
rect 17408 32555 17460 32564
rect 17408 32521 17417 32555
rect 17417 32521 17451 32555
rect 17451 32521 17460 32555
rect 17408 32512 17460 32521
rect 19340 32512 19392 32564
rect 8392 32444 8444 32496
rect 22284 32512 22336 32564
rect 22836 32555 22888 32564
rect 22836 32521 22845 32555
rect 22845 32521 22879 32555
rect 22879 32521 22888 32555
rect 22836 32512 22888 32521
rect 25964 32512 26016 32564
rect 26240 32512 26292 32564
rect 27712 32512 27764 32564
rect 29000 32555 29052 32564
rect 29000 32521 29009 32555
rect 29009 32521 29043 32555
rect 29043 32521 29052 32555
rect 29000 32512 29052 32521
rect 29644 32555 29696 32564
rect 29644 32521 29653 32555
rect 29653 32521 29687 32555
rect 29687 32521 29696 32555
rect 29644 32512 29696 32521
rect 30564 32512 30616 32564
rect 33508 32512 33560 32564
rect 35532 32512 35584 32564
rect 39028 32555 39080 32564
rect 39028 32521 39037 32555
rect 39037 32521 39071 32555
rect 39071 32521 39080 32555
rect 39028 32512 39080 32521
rect 39856 32555 39908 32564
rect 39856 32521 39865 32555
rect 39865 32521 39899 32555
rect 39899 32521 39908 32555
rect 39856 32512 39908 32521
rect 40408 32512 40460 32564
rect 4620 32419 4672 32428
rect 4620 32385 4629 32419
rect 4629 32385 4663 32419
rect 4663 32385 4672 32419
rect 4620 32376 4672 32385
rect 8300 32376 8352 32428
rect 14648 32419 14700 32428
rect 14648 32385 14657 32419
rect 14657 32385 14691 32419
rect 14691 32385 14700 32419
rect 14648 32376 14700 32385
rect 15292 32376 15344 32428
rect 22100 32444 22152 32496
rect 18604 32419 18656 32428
rect 3240 32308 3292 32360
rect 4528 32351 4580 32360
rect 4528 32317 4537 32351
rect 4537 32317 4571 32351
rect 4571 32317 4580 32351
rect 4528 32308 4580 32317
rect 5172 32308 5224 32360
rect 6184 32308 6236 32360
rect 7380 32308 7432 32360
rect 9680 32351 9732 32360
rect 9680 32317 9689 32351
rect 9689 32317 9723 32351
rect 9723 32317 9732 32351
rect 9680 32308 9732 32317
rect 11152 32308 11204 32360
rect 12992 32351 13044 32360
rect 12992 32317 13001 32351
rect 13001 32317 13035 32351
rect 13035 32317 13044 32351
rect 12992 32308 13044 32317
rect 14004 32351 14056 32360
rect 14004 32317 14013 32351
rect 14013 32317 14047 32351
rect 14047 32317 14056 32351
rect 14004 32308 14056 32317
rect 15660 32351 15712 32360
rect 7840 32283 7892 32292
rect 7840 32249 7849 32283
rect 7849 32249 7883 32283
rect 7883 32249 7892 32283
rect 7840 32240 7892 32249
rect 11428 32283 11480 32292
rect 11428 32249 11437 32283
rect 11437 32249 11471 32283
rect 11471 32249 11480 32283
rect 11428 32240 11480 32249
rect 11888 32283 11940 32292
rect 11888 32249 11897 32283
rect 11897 32249 11931 32283
rect 11931 32249 11940 32283
rect 11888 32240 11940 32249
rect 3516 32215 3568 32224
rect 3516 32181 3525 32215
rect 3525 32181 3559 32215
rect 3559 32181 3568 32215
rect 3516 32172 3568 32181
rect 6092 32172 6144 32224
rect 6276 32215 6328 32224
rect 6276 32181 6285 32215
rect 6285 32181 6319 32215
rect 6319 32181 6328 32215
rect 6276 32172 6328 32181
rect 10416 32172 10468 32224
rect 14188 32240 14240 32292
rect 15660 32317 15669 32351
rect 15669 32317 15703 32351
rect 15703 32317 15712 32351
rect 15660 32308 15712 32317
rect 18604 32385 18613 32419
rect 18613 32385 18647 32419
rect 18647 32385 18656 32419
rect 18604 32376 18656 32385
rect 20260 32376 20312 32428
rect 21732 32419 21784 32428
rect 21732 32385 21741 32419
rect 21741 32385 21775 32419
rect 21775 32385 21784 32419
rect 21732 32376 21784 32385
rect 26976 32444 27028 32496
rect 28080 32487 28132 32496
rect 28080 32453 28089 32487
rect 28089 32453 28123 32487
rect 28123 32453 28132 32487
rect 28080 32444 28132 32453
rect 32128 32444 32180 32496
rect 35624 32487 35676 32496
rect 35624 32453 35633 32487
rect 35633 32453 35667 32487
rect 35667 32453 35676 32487
rect 35624 32444 35676 32453
rect 42064 32444 42116 32496
rect 24216 32419 24268 32428
rect 24216 32385 24225 32419
rect 24225 32385 24259 32419
rect 24259 32385 24268 32419
rect 24216 32376 24268 32385
rect 26516 32376 26568 32428
rect 27528 32376 27580 32428
rect 29920 32376 29972 32428
rect 18512 32351 18564 32360
rect 18512 32317 18521 32351
rect 18521 32317 18555 32351
rect 18555 32317 18564 32351
rect 18512 32308 18564 32317
rect 25228 32351 25280 32360
rect 25228 32317 25237 32351
rect 25237 32317 25271 32351
rect 25271 32317 25280 32351
rect 25228 32308 25280 32317
rect 17868 32240 17920 32292
rect 19892 32283 19944 32292
rect 19892 32249 19901 32283
rect 19901 32249 19935 32283
rect 19935 32249 19944 32283
rect 20444 32283 20496 32292
rect 19892 32240 19944 32249
rect 20444 32249 20453 32283
rect 20453 32249 20487 32283
rect 20487 32249 20496 32283
rect 20444 32240 20496 32249
rect 21180 32240 21232 32292
rect 21456 32283 21508 32292
rect 21456 32249 21465 32283
rect 21465 32249 21499 32283
rect 21499 32249 21508 32283
rect 21456 32240 21508 32249
rect 24124 32240 24176 32292
rect 13452 32215 13504 32224
rect 13452 32181 13461 32215
rect 13461 32181 13495 32215
rect 13495 32181 13504 32215
rect 13452 32172 13504 32181
rect 22376 32215 22428 32224
rect 22376 32181 22385 32215
rect 22385 32181 22419 32215
rect 22419 32181 22428 32215
rect 22376 32172 22428 32181
rect 23020 32172 23072 32224
rect 23296 32172 23348 32224
rect 26700 32240 26752 32292
rect 29644 32240 29696 32292
rect 32404 32376 32456 32428
rect 33416 32376 33468 32428
rect 33784 32419 33836 32428
rect 33784 32385 33793 32419
rect 33793 32385 33827 32419
rect 33827 32385 33836 32419
rect 33784 32376 33836 32385
rect 31852 32351 31904 32360
rect 31852 32317 31861 32351
rect 31861 32317 31895 32351
rect 31895 32317 31904 32351
rect 31852 32308 31904 32317
rect 32036 32351 32088 32360
rect 32036 32317 32045 32351
rect 32045 32317 32079 32351
rect 32079 32317 32088 32351
rect 32036 32308 32088 32317
rect 40776 32376 40828 32428
rect 42432 32419 42484 32428
rect 42432 32385 42441 32419
rect 42441 32385 42475 32419
rect 42475 32385 42484 32419
rect 44548 32444 44600 32496
rect 42432 32376 42484 32385
rect 43536 32376 43588 32428
rect 30472 32240 30524 32292
rect 30656 32240 30708 32292
rect 28632 32215 28684 32224
rect 28632 32181 28641 32215
rect 28641 32181 28675 32215
rect 28675 32181 28684 32215
rect 28632 32172 28684 32181
rect 32312 32283 32364 32292
rect 32312 32249 32321 32283
rect 32321 32249 32355 32283
rect 32355 32249 32364 32283
rect 32312 32240 32364 32249
rect 33508 32240 33560 32292
rect 36452 32308 36504 32360
rect 37372 32351 37424 32360
rect 37372 32317 37381 32351
rect 37381 32317 37415 32351
rect 37415 32317 37424 32351
rect 37372 32308 37424 32317
rect 39856 32308 39908 32360
rect 33140 32172 33192 32224
rect 40408 32240 40460 32292
rect 41236 32283 41288 32292
rect 37832 32172 37884 32224
rect 38752 32172 38804 32224
rect 41236 32249 41245 32283
rect 41245 32249 41279 32283
rect 41279 32249 41288 32283
rect 41236 32240 41288 32249
rect 44088 32240 44140 32292
rect 43352 32215 43404 32224
rect 43352 32181 43361 32215
rect 43361 32181 43395 32215
rect 43395 32181 43404 32215
rect 43352 32172 43404 32181
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 9680 31968 9732 32020
rect 11244 31968 11296 32020
rect 14188 32011 14240 32020
rect 14188 31977 14197 32011
rect 14197 31977 14231 32011
rect 14231 31977 14240 32011
rect 14188 31968 14240 31977
rect 14832 31968 14884 32020
rect 15660 32011 15712 32020
rect 15660 31977 15669 32011
rect 15669 31977 15703 32011
rect 15703 31977 15712 32011
rect 15660 31968 15712 31977
rect 17316 32011 17368 32020
rect 17316 31977 17325 32011
rect 17325 31977 17359 32011
rect 17359 31977 17368 32011
rect 17316 31968 17368 31977
rect 22100 32011 22152 32020
rect 22100 31977 22109 32011
rect 22109 31977 22143 32011
rect 22143 31977 22152 32011
rect 22100 31968 22152 31977
rect 23020 32011 23072 32020
rect 23020 31977 23029 32011
rect 23029 31977 23063 32011
rect 23063 31977 23072 32011
rect 23020 31968 23072 31977
rect 24124 31968 24176 32020
rect 24492 31968 24544 32020
rect 27528 32011 27580 32020
rect 4896 31900 4948 31952
rect 12072 31900 12124 31952
rect 19432 31943 19484 31952
rect 19432 31909 19441 31943
rect 19441 31909 19475 31943
rect 19475 31909 19484 31943
rect 19432 31900 19484 31909
rect 21180 31900 21232 31952
rect 24584 31943 24636 31952
rect 3792 31832 3844 31884
rect 4528 31875 4580 31884
rect 4528 31841 4537 31875
rect 4537 31841 4571 31875
rect 4571 31841 4580 31875
rect 4528 31832 4580 31841
rect 5816 31832 5868 31884
rect 6368 31832 6420 31884
rect 7380 31875 7432 31884
rect 7380 31841 7389 31875
rect 7389 31841 7423 31875
rect 7423 31841 7432 31875
rect 7380 31832 7432 31841
rect 8392 31832 8444 31884
rect 9588 31832 9640 31884
rect 10140 31875 10192 31884
rect 10140 31841 10149 31875
rect 10149 31841 10183 31875
rect 10183 31841 10192 31875
rect 10140 31832 10192 31841
rect 11428 31875 11480 31884
rect 11428 31841 11437 31875
rect 11437 31841 11471 31875
rect 11471 31841 11480 31875
rect 11428 31832 11480 31841
rect 12256 31832 12308 31884
rect 13268 31832 13320 31884
rect 16488 31832 16540 31884
rect 17316 31875 17368 31884
rect 17316 31841 17325 31875
rect 17325 31841 17359 31875
rect 17359 31841 17368 31875
rect 17316 31832 17368 31841
rect 17868 31832 17920 31884
rect 21548 31832 21600 31884
rect 24584 31909 24593 31943
rect 24593 31909 24627 31943
rect 24627 31909 24636 31943
rect 24584 31900 24636 31909
rect 26700 31943 26752 31952
rect 26700 31909 26709 31943
rect 26709 31909 26743 31943
rect 26743 31909 26752 31943
rect 26700 31900 26752 31909
rect 27528 31977 27537 32011
rect 27537 31977 27571 32011
rect 27571 31977 27580 32011
rect 27528 31968 27580 31977
rect 29644 31968 29696 32020
rect 30472 32011 30524 32020
rect 30472 31977 30481 32011
rect 30481 31977 30515 32011
rect 30515 31977 30524 32011
rect 30472 31968 30524 31977
rect 30748 32011 30800 32020
rect 30748 31977 30757 32011
rect 30757 31977 30791 32011
rect 30791 31977 30800 32011
rect 30748 31968 30800 31977
rect 32312 32011 32364 32020
rect 32312 31977 32321 32011
rect 32321 31977 32355 32011
rect 32355 31977 32364 32011
rect 32312 31968 32364 31977
rect 33968 31968 34020 32020
rect 37372 32011 37424 32020
rect 37372 31977 37381 32011
rect 37381 31977 37415 32011
rect 37415 31977 37424 32011
rect 37372 31968 37424 31977
rect 40592 31968 40644 32020
rect 33416 31943 33468 31952
rect 33416 31909 33425 31943
rect 33425 31909 33459 31943
rect 33459 31909 33468 31943
rect 33416 31900 33468 31909
rect 33508 31900 33560 31952
rect 29552 31875 29604 31884
rect 29552 31841 29561 31875
rect 29561 31841 29595 31875
rect 29595 31841 29604 31875
rect 29552 31832 29604 31841
rect 32588 31832 32640 31884
rect 35348 31832 35400 31884
rect 35716 31832 35768 31884
rect 35992 31832 36044 31884
rect 37740 31900 37792 31952
rect 37832 31900 37884 31952
rect 38476 31900 38528 31952
rect 38936 31943 38988 31952
rect 38936 31909 38945 31943
rect 38945 31909 38979 31943
rect 38979 31909 38988 31943
rect 38936 31900 38988 31909
rect 39672 31900 39724 31952
rect 41512 31900 41564 31952
rect 44088 31900 44140 31952
rect 40408 31875 40460 31884
rect 7472 31807 7524 31816
rect 7472 31773 7481 31807
rect 7481 31773 7515 31807
rect 7515 31773 7524 31807
rect 7472 31764 7524 31773
rect 19340 31807 19392 31816
rect 19340 31773 19349 31807
rect 19349 31773 19383 31807
rect 19383 31773 19392 31807
rect 19340 31764 19392 31773
rect 7840 31696 7892 31748
rect 15292 31696 15344 31748
rect 16488 31696 16540 31748
rect 20444 31764 20496 31816
rect 22652 31807 22704 31816
rect 22652 31773 22661 31807
rect 22661 31773 22695 31807
rect 22695 31773 22704 31807
rect 22652 31764 22704 31773
rect 24492 31807 24544 31816
rect 24492 31773 24501 31807
rect 24501 31773 24535 31807
rect 24535 31773 24544 31807
rect 24492 31764 24544 31773
rect 26608 31807 26660 31816
rect 24216 31696 24268 31748
rect 26608 31773 26617 31807
rect 26617 31773 26651 31807
rect 26651 31773 26660 31807
rect 26608 31764 26660 31773
rect 26884 31764 26936 31816
rect 26240 31696 26292 31748
rect 31760 31764 31812 31816
rect 33600 31764 33652 31816
rect 33968 31807 34020 31816
rect 33968 31773 33977 31807
rect 33977 31773 34011 31807
rect 34011 31773 34020 31807
rect 33968 31764 34020 31773
rect 37740 31807 37792 31816
rect 33784 31696 33836 31748
rect 37740 31773 37749 31807
rect 37749 31773 37783 31807
rect 37783 31773 37792 31807
rect 37740 31764 37792 31773
rect 39488 31807 39540 31816
rect 39488 31773 39497 31807
rect 39497 31773 39531 31807
rect 39531 31773 39540 31807
rect 39488 31764 39540 31773
rect 40408 31841 40417 31875
rect 40417 31841 40451 31875
rect 40451 31841 40460 31875
rect 40408 31832 40460 31841
rect 41880 31764 41932 31816
rect 43444 31807 43496 31816
rect 43444 31773 43453 31807
rect 43453 31773 43487 31807
rect 43487 31773 43496 31807
rect 43444 31764 43496 31773
rect 34428 31696 34480 31748
rect 38568 31696 38620 31748
rect 41236 31696 41288 31748
rect 5172 31628 5224 31680
rect 6184 31671 6236 31680
rect 6184 31637 6193 31671
rect 6193 31637 6227 31671
rect 6227 31637 6236 31671
rect 6184 31628 6236 31637
rect 8300 31671 8352 31680
rect 8300 31637 8309 31671
rect 8309 31637 8343 31671
rect 8343 31637 8352 31671
rect 8300 31628 8352 31637
rect 12256 31628 12308 31680
rect 12992 31628 13044 31680
rect 14188 31628 14240 31680
rect 17868 31628 17920 31680
rect 18972 31671 19024 31680
rect 18972 31637 18981 31671
rect 18981 31637 19015 31671
rect 19015 31637 19024 31671
rect 18972 31628 19024 31637
rect 21364 31671 21416 31680
rect 21364 31637 21373 31671
rect 21373 31637 21407 31671
rect 21407 31637 21416 31671
rect 21364 31628 21416 31637
rect 25596 31628 25648 31680
rect 28632 31628 28684 31680
rect 29368 31671 29420 31680
rect 29368 31637 29377 31671
rect 29377 31637 29411 31671
rect 29411 31637 29420 31671
rect 29368 31628 29420 31637
rect 30472 31628 30524 31680
rect 32036 31628 32088 31680
rect 35348 31671 35400 31680
rect 35348 31637 35357 31671
rect 35357 31637 35391 31671
rect 35391 31637 35400 31671
rect 35348 31628 35400 31637
rect 36176 31628 36228 31680
rect 39396 31628 39448 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 4620 31424 4672 31476
rect 16488 31467 16540 31476
rect 16488 31433 16497 31467
rect 16497 31433 16531 31467
rect 16531 31433 16540 31467
rect 16488 31424 16540 31433
rect 19432 31424 19484 31476
rect 21548 31467 21600 31476
rect 21548 31433 21557 31467
rect 21557 31433 21591 31467
rect 21591 31433 21600 31467
rect 21548 31424 21600 31433
rect 24400 31424 24452 31476
rect 24584 31424 24636 31476
rect 25964 31467 26016 31476
rect 25964 31433 25973 31467
rect 25973 31433 26007 31467
rect 26007 31433 26016 31467
rect 25964 31424 26016 31433
rect 26608 31424 26660 31476
rect 29644 31424 29696 31476
rect 30288 31467 30340 31476
rect 30288 31433 30297 31467
rect 30297 31433 30331 31467
rect 30331 31433 30340 31467
rect 30288 31424 30340 31433
rect 32588 31424 32640 31476
rect 33968 31424 34020 31476
rect 34152 31467 34204 31476
rect 34152 31433 34161 31467
rect 34161 31433 34195 31467
rect 34195 31433 34204 31467
rect 34152 31424 34204 31433
rect 35992 31467 36044 31476
rect 35992 31433 36001 31467
rect 36001 31433 36035 31467
rect 36035 31433 36044 31467
rect 35992 31424 36044 31433
rect 36452 31424 36504 31476
rect 37740 31424 37792 31476
rect 39396 31467 39448 31476
rect 39396 31433 39405 31467
rect 39405 31433 39439 31467
rect 39439 31433 39448 31467
rect 39396 31424 39448 31433
rect 40776 31467 40828 31476
rect 40776 31433 40785 31467
rect 40785 31433 40819 31467
rect 40819 31433 40828 31467
rect 40776 31424 40828 31433
rect 41880 31467 41932 31476
rect 41880 31433 41889 31467
rect 41889 31433 41923 31467
rect 41923 31433 41932 31467
rect 41880 31424 41932 31433
rect 43444 31424 43496 31476
rect 43628 31424 43680 31476
rect 44088 31467 44140 31476
rect 44088 31433 44097 31467
rect 44097 31433 44131 31467
rect 44131 31433 44140 31467
rect 44088 31424 44140 31433
rect 7012 31288 7064 31340
rect 10140 31288 10192 31340
rect 13268 31288 13320 31340
rect 5172 31220 5224 31272
rect 10784 31263 10836 31272
rect 10784 31229 10793 31263
rect 10793 31229 10827 31263
rect 10827 31229 10836 31263
rect 10784 31220 10836 31229
rect 11152 31220 11204 31272
rect 14464 31263 14516 31272
rect 14464 31229 14473 31263
rect 14473 31229 14507 31263
rect 14507 31229 14516 31263
rect 14464 31220 14516 31229
rect 15292 31220 15344 31272
rect 18696 31356 18748 31408
rect 3792 31084 3844 31136
rect 4988 31084 5040 31136
rect 5356 31127 5408 31136
rect 5356 31093 5365 31127
rect 5365 31093 5399 31127
rect 5399 31093 5408 31127
rect 5356 31084 5408 31093
rect 6368 31084 6420 31136
rect 7012 31195 7064 31204
rect 7012 31161 7021 31195
rect 7021 31161 7055 31195
rect 7055 31161 7064 31195
rect 7012 31152 7064 31161
rect 8852 31195 8904 31204
rect 8852 31161 8861 31195
rect 8861 31161 8895 31195
rect 8895 31161 8904 31195
rect 8852 31152 8904 31161
rect 8944 31195 8996 31204
rect 8944 31161 8953 31195
rect 8953 31161 8987 31195
rect 8987 31161 8996 31195
rect 8944 31152 8996 31161
rect 9680 31152 9732 31204
rect 12532 31195 12584 31204
rect 12532 31161 12541 31195
rect 12541 31161 12575 31195
rect 12575 31161 12584 31195
rect 12532 31152 12584 31161
rect 13176 31195 13228 31204
rect 8392 31084 8444 31136
rect 9588 31084 9640 31136
rect 10140 31127 10192 31136
rect 10140 31093 10149 31127
rect 10149 31093 10183 31127
rect 10183 31093 10192 31127
rect 10140 31084 10192 31093
rect 10876 31127 10928 31136
rect 10876 31093 10885 31127
rect 10885 31093 10919 31127
rect 10919 31093 10928 31127
rect 10876 31084 10928 31093
rect 11428 31084 11480 31136
rect 13176 31161 13185 31195
rect 13185 31161 13219 31195
rect 13219 31161 13228 31195
rect 13176 31152 13228 31161
rect 12900 31084 12952 31136
rect 13912 31152 13964 31204
rect 17316 31152 17368 31204
rect 17776 31152 17828 31204
rect 19340 31356 19392 31408
rect 21732 31356 21784 31408
rect 32772 31356 32824 31408
rect 33140 31356 33192 31408
rect 22652 31331 22704 31340
rect 22652 31297 22661 31331
rect 22661 31297 22695 31331
rect 22695 31297 22704 31331
rect 22652 31288 22704 31297
rect 25228 31288 25280 31340
rect 26884 31331 26936 31340
rect 26884 31297 26893 31331
rect 26893 31297 26927 31331
rect 26927 31297 26936 31331
rect 26884 31288 26936 31297
rect 27160 31331 27212 31340
rect 27160 31297 27169 31331
rect 27169 31297 27203 31331
rect 27203 31297 27212 31331
rect 27160 31288 27212 31297
rect 29920 31331 29972 31340
rect 29920 31297 29929 31331
rect 29929 31297 29963 31331
rect 29963 31297 29972 31331
rect 29920 31288 29972 31297
rect 30380 31288 30432 31340
rect 31944 31331 31996 31340
rect 18972 31263 19024 31272
rect 18972 31229 18981 31263
rect 18981 31229 19015 31263
rect 19015 31229 19024 31263
rect 18972 31220 19024 31229
rect 21916 31263 21968 31272
rect 19248 31152 19300 31204
rect 17868 31084 17920 31136
rect 20904 31127 20956 31136
rect 20904 31093 20913 31127
rect 20913 31093 20947 31127
rect 20947 31093 20956 31127
rect 20904 31084 20956 31093
rect 21916 31229 21925 31263
rect 21925 31229 21959 31263
rect 21959 31229 21968 31263
rect 21916 31220 21968 31229
rect 22100 31220 22152 31272
rect 24584 31220 24636 31272
rect 29460 31263 29512 31272
rect 29460 31229 29469 31263
rect 29469 31229 29503 31263
rect 29503 31229 29512 31263
rect 29460 31220 29512 31229
rect 30472 31220 30524 31272
rect 31944 31297 31953 31331
rect 31953 31297 31987 31331
rect 31987 31297 31996 31331
rect 31944 31288 31996 31297
rect 34244 31288 34296 31340
rect 33416 31220 33468 31272
rect 34152 31220 34204 31272
rect 35440 31288 35492 31340
rect 25964 31152 26016 31204
rect 35992 31220 36044 31272
rect 36452 31263 36504 31272
rect 36452 31229 36461 31263
rect 36461 31229 36495 31263
rect 36495 31229 36504 31263
rect 36452 31220 36504 31229
rect 39672 31399 39724 31408
rect 39672 31365 39681 31399
rect 39681 31365 39715 31399
rect 39715 31365 39724 31399
rect 41512 31399 41564 31408
rect 39672 31356 39724 31365
rect 41512 31365 41521 31399
rect 41521 31365 41555 31399
rect 41555 31365 41564 31399
rect 41512 31356 41564 31365
rect 38476 31288 38528 31340
rect 38568 31288 38620 31340
rect 38292 31220 38344 31272
rect 39120 31220 39172 31272
rect 21640 31084 21692 31136
rect 22284 31084 22336 31136
rect 23020 31084 23072 31136
rect 23756 31084 23808 31136
rect 26700 31084 26752 31136
rect 31024 31127 31076 31136
rect 31024 31093 31033 31127
rect 31033 31093 31067 31127
rect 31067 31093 31076 31127
rect 31024 31084 31076 31093
rect 31576 31084 31628 31136
rect 39488 31152 39540 31204
rect 42156 31220 42208 31272
rect 43536 31288 43588 31340
rect 43628 31220 43680 31272
rect 33508 31127 33560 31136
rect 33508 31093 33517 31127
rect 33517 31093 33551 31127
rect 33551 31093 33560 31127
rect 33508 31084 33560 31093
rect 37832 31084 37884 31136
rect 41052 31127 41104 31136
rect 41052 31093 41061 31127
rect 41061 31093 41095 31127
rect 41095 31093 41104 31127
rect 41052 31084 41104 31093
rect 42708 31127 42760 31136
rect 42708 31093 42717 31127
rect 42717 31093 42751 31127
rect 42751 31093 42760 31127
rect 42708 31084 42760 31093
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 4620 30923 4672 30932
rect 4620 30889 4629 30923
rect 4629 30889 4663 30923
rect 4663 30889 4672 30923
rect 4620 30880 4672 30889
rect 5816 30880 5868 30932
rect 6184 30880 6236 30932
rect 7012 30880 7064 30932
rect 8852 30923 8904 30932
rect 5908 30812 5960 30864
rect 7840 30855 7892 30864
rect 7840 30821 7849 30855
rect 7849 30821 7883 30855
rect 7883 30821 7892 30855
rect 7840 30812 7892 30821
rect 8852 30889 8861 30923
rect 8861 30889 8895 30923
rect 8895 30889 8904 30923
rect 8852 30880 8904 30889
rect 12532 30923 12584 30932
rect 12532 30889 12541 30923
rect 12541 30889 12575 30923
rect 12575 30889 12584 30923
rect 12532 30880 12584 30889
rect 19248 30923 19300 30932
rect 19248 30889 19257 30923
rect 19257 30889 19291 30923
rect 19291 30889 19300 30923
rect 19248 30880 19300 30889
rect 24492 30880 24544 30932
rect 29552 30923 29604 30932
rect 29552 30889 29561 30923
rect 29561 30889 29595 30923
rect 29595 30889 29604 30923
rect 29552 30880 29604 30889
rect 31944 30923 31996 30932
rect 31944 30889 31953 30923
rect 31953 30889 31987 30923
rect 31987 30889 31996 30923
rect 31944 30880 31996 30889
rect 33968 30880 34020 30932
rect 35440 30880 35492 30932
rect 36452 30923 36504 30932
rect 36452 30889 36461 30923
rect 36461 30889 36495 30923
rect 36495 30889 36504 30923
rect 36452 30880 36504 30889
rect 38292 30923 38344 30932
rect 38292 30889 38301 30923
rect 38301 30889 38335 30923
rect 38335 30889 38344 30923
rect 38292 30880 38344 30889
rect 39212 30880 39264 30932
rect 8484 30812 8536 30864
rect 11244 30855 11296 30864
rect 11244 30821 11253 30855
rect 11253 30821 11287 30855
rect 11287 30821 11296 30855
rect 11244 30812 11296 30821
rect 12256 30855 12308 30864
rect 12256 30821 12265 30855
rect 12265 30821 12299 30855
rect 12299 30821 12308 30855
rect 12256 30812 12308 30821
rect 23848 30855 23900 30864
rect 23848 30821 23857 30855
rect 23857 30821 23891 30855
rect 23891 30821 23900 30855
rect 23848 30812 23900 30821
rect 26700 30855 26752 30864
rect 26700 30821 26709 30855
rect 26709 30821 26743 30855
rect 26743 30821 26752 30855
rect 26700 30812 26752 30821
rect 27252 30855 27304 30864
rect 27252 30821 27261 30855
rect 27261 30821 27295 30855
rect 27295 30821 27304 30855
rect 27252 30812 27304 30821
rect 32404 30855 32456 30864
rect 32404 30821 32413 30855
rect 32413 30821 32447 30855
rect 32447 30821 32456 30855
rect 32404 30812 32456 30821
rect 32772 30812 32824 30864
rect 33508 30812 33560 30864
rect 6092 30744 6144 30796
rect 7472 30744 7524 30796
rect 10048 30787 10100 30796
rect 10048 30753 10066 30787
rect 10066 30753 10100 30787
rect 10048 30744 10100 30753
rect 13268 30787 13320 30796
rect 13268 30753 13277 30787
rect 13277 30753 13311 30787
rect 13311 30753 13320 30787
rect 13268 30744 13320 30753
rect 13360 30744 13412 30796
rect 15476 30787 15528 30796
rect 15476 30753 15485 30787
rect 15485 30753 15519 30787
rect 15519 30753 15528 30787
rect 15476 30744 15528 30753
rect 17132 30787 17184 30796
rect 17132 30753 17141 30787
rect 17141 30753 17175 30787
rect 17175 30753 17184 30787
rect 17132 30744 17184 30753
rect 19892 30744 19944 30796
rect 21732 30744 21784 30796
rect 22744 30744 22796 30796
rect 24400 30744 24452 30796
rect 26240 30744 26292 30796
rect 29092 30744 29144 30796
rect 30196 30787 30248 30796
rect 30196 30753 30205 30787
rect 30205 30753 30239 30787
rect 30239 30753 30248 30787
rect 30196 30744 30248 30753
rect 30472 30787 30524 30796
rect 30472 30753 30481 30787
rect 30481 30753 30515 30787
rect 30515 30753 30524 30787
rect 30472 30744 30524 30753
rect 37740 30787 37792 30796
rect 37740 30753 37749 30787
rect 37749 30753 37783 30787
rect 37783 30753 37792 30787
rect 37740 30744 37792 30753
rect 38936 30744 38988 30796
rect 39764 30787 39816 30796
rect 39764 30753 39773 30787
rect 39773 30753 39807 30787
rect 39807 30753 39816 30787
rect 39764 30744 39816 30753
rect 41144 30787 41196 30796
rect 41144 30753 41153 30787
rect 41153 30753 41187 30787
rect 41187 30753 41196 30787
rect 41144 30744 41196 30753
rect 4896 30676 4948 30728
rect 6000 30719 6052 30728
rect 6000 30685 6009 30719
rect 6009 30685 6043 30719
rect 6043 30685 6052 30719
rect 6000 30676 6052 30685
rect 8116 30719 8168 30728
rect 8116 30685 8125 30719
rect 8125 30685 8159 30719
rect 8159 30685 8168 30719
rect 8116 30676 8168 30685
rect 10968 30719 11020 30728
rect 10968 30685 10977 30719
rect 10977 30685 11011 30719
rect 11011 30685 11020 30719
rect 10968 30676 11020 30685
rect 13820 30719 13872 30728
rect 13820 30685 13829 30719
rect 13829 30685 13863 30719
rect 13863 30685 13872 30719
rect 13820 30676 13872 30685
rect 14740 30676 14792 30728
rect 16948 30719 17000 30728
rect 16948 30685 16957 30719
rect 16957 30685 16991 30719
rect 16991 30685 17000 30719
rect 16948 30676 17000 30685
rect 18880 30719 18932 30728
rect 18880 30685 18889 30719
rect 18889 30685 18923 30719
rect 18923 30685 18932 30719
rect 18880 30676 18932 30685
rect 23940 30676 23992 30728
rect 24124 30719 24176 30728
rect 24124 30685 24133 30719
rect 24133 30685 24167 30719
rect 24167 30685 24176 30719
rect 24124 30676 24176 30685
rect 17776 30608 17828 30660
rect 21916 30651 21968 30660
rect 21916 30617 21925 30651
rect 21925 30617 21959 30651
rect 21959 30617 21968 30651
rect 30656 30719 30708 30728
rect 30656 30685 30665 30719
rect 30665 30685 30699 30719
rect 30699 30685 30708 30719
rect 30656 30676 30708 30685
rect 31944 30676 31996 30728
rect 33968 30719 34020 30728
rect 33968 30685 33977 30719
rect 33977 30685 34011 30719
rect 34011 30685 34020 30719
rect 33968 30676 34020 30685
rect 34244 30719 34296 30728
rect 34244 30685 34253 30719
rect 34253 30685 34287 30719
rect 34287 30685 34296 30719
rect 34244 30676 34296 30685
rect 34612 30676 34664 30728
rect 35808 30719 35860 30728
rect 35808 30685 35817 30719
rect 35817 30685 35851 30719
rect 35851 30685 35860 30719
rect 35808 30676 35860 30685
rect 21916 30608 21968 30617
rect 6736 30540 6788 30592
rect 7380 30540 7432 30592
rect 10140 30540 10192 30592
rect 10324 30540 10376 30592
rect 11152 30540 11204 30592
rect 18328 30583 18380 30592
rect 18328 30549 18337 30583
rect 18337 30549 18371 30583
rect 18371 30549 18380 30583
rect 18328 30540 18380 30549
rect 18788 30540 18840 30592
rect 23020 30540 23072 30592
rect 24584 30540 24636 30592
rect 30472 30608 30524 30660
rect 32956 30608 33008 30660
rect 36452 30608 36504 30660
rect 28172 30540 28224 30592
rect 35348 30540 35400 30592
rect 38844 30540 38896 30592
rect 39212 30583 39264 30592
rect 39212 30549 39221 30583
rect 39221 30549 39255 30583
rect 39255 30549 39264 30583
rect 39212 30540 39264 30549
rect 40960 30583 41012 30592
rect 40960 30549 40969 30583
rect 40969 30549 41003 30583
rect 41003 30549 41012 30583
rect 40960 30540 41012 30549
rect 41788 30540 41840 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 6000 30336 6052 30388
rect 10048 30379 10100 30388
rect 10048 30345 10057 30379
rect 10057 30345 10091 30379
rect 10091 30345 10100 30379
rect 10048 30336 10100 30345
rect 11520 30379 11572 30388
rect 11520 30345 11529 30379
rect 11529 30345 11563 30379
rect 11563 30345 11572 30379
rect 11520 30336 11572 30345
rect 15476 30379 15528 30388
rect 15476 30345 15485 30379
rect 15485 30345 15519 30379
rect 15519 30345 15528 30379
rect 15476 30336 15528 30345
rect 19248 30336 19300 30388
rect 21364 30379 21416 30388
rect 3056 30268 3108 30320
rect 3700 30268 3752 30320
rect 2964 29996 3016 30048
rect 5080 30175 5132 30184
rect 3148 30064 3200 30116
rect 3516 30064 3568 30116
rect 5080 30141 5089 30175
rect 5089 30141 5123 30175
rect 5123 30141 5132 30175
rect 5080 30132 5132 30141
rect 10784 30268 10836 30320
rect 12256 30268 12308 30320
rect 13268 30268 13320 30320
rect 7472 30243 7524 30252
rect 7472 30209 7481 30243
rect 7481 30209 7515 30243
rect 7515 30209 7524 30243
rect 7472 30200 7524 30209
rect 8116 30243 8168 30252
rect 8116 30209 8125 30243
rect 8125 30209 8159 30243
rect 8159 30209 8168 30243
rect 9036 30243 9088 30252
rect 8116 30200 8168 30209
rect 9036 30209 9045 30243
rect 9045 30209 9079 30243
rect 9079 30209 9088 30243
rect 9036 30200 9088 30209
rect 10876 30200 10928 30252
rect 13820 30200 13872 30252
rect 17868 30243 17920 30252
rect 17868 30209 17877 30243
rect 17877 30209 17911 30243
rect 17911 30209 17920 30243
rect 17868 30200 17920 30209
rect 18880 30200 18932 30252
rect 5264 30175 5316 30184
rect 5264 30141 5273 30175
rect 5273 30141 5307 30175
rect 5307 30141 5316 30175
rect 5264 30132 5316 30141
rect 14648 30132 14700 30184
rect 17684 30132 17736 30184
rect 18328 30175 18380 30184
rect 18328 30141 18337 30175
rect 18337 30141 18371 30175
rect 18371 30141 18380 30175
rect 18328 30132 18380 30141
rect 18788 30175 18840 30184
rect 18788 30141 18797 30175
rect 18797 30141 18831 30175
rect 18831 30141 18840 30175
rect 18788 30132 18840 30141
rect 3884 30064 3936 30116
rect 5908 30064 5960 30116
rect 7564 30107 7616 30116
rect 7564 30073 7573 30107
rect 7573 30073 7607 30107
rect 7607 30073 7616 30107
rect 7564 30064 7616 30073
rect 9496 30064 9548 30116
rect 9680 30107 9732 30116
rect 9680 30073 9689 30107
rect 9689 30073 9723 30107
rect 9723 30073 9732 30107
rect 9680 30064 9732 30073
rect 11244 30064 11296 30116
rect 13728 30064 13780 30116
rect 14096 30064 14148 30116
rect 15660 30107 15712 30116
rect 15660 30073 15669 30107
rect 15669 30073 15703 30107
rect 15703 30073 15712 30107
rect 15660 30064 15712 30073
rect 21364 30345 21373 30379
rect 21373 30345 21407 30379
rect 21407 30345 21416 30379
rect 21364 30336 21416 30345
rect 22744 30336 22796 30388
rect 23480 30379 23532 30388
rect 23480 30345 23489 30379
rect 23489 30345 23523 30379
rect 23523 30345 23532 30379
rect 23480 30336 23532 30345
rect 23848 30336 23900 30388
rect 23940 30336 23992 30388
rect 27252 30336 27304 30388
rect 28264 30336 28316 30388
rect 30288 30336 30340 30388
rect 31576 30379 31628 30388
rect 31576 30345 31585 30379
rect 31585 30345 31619 30379
rect 31619 30345 31628 30379
rect 31576 30336 31628 30345
rect 32404 30336 32456 30388
rect 33508 30336 33560 30388
rect 34152 30336 34204 30388
rect 36452 30379 36504 30388
rect 36452 30345 36461 30379
rect 36461 30345 36495 30379
rect 36495 30345 36504 30379
rect 36452 30336 36504 30345
rect 39672 30336 39724 30388
rect 26240 30311 26292 30320
rect 26240 30277 26249 30311
rect 26249 30277 26283 30311
rect 26283 30277 26292 30311
rect 26240 30268 26292 30277
rect 27160 30268 27212 30320
rect 30196 30311 30248 30320
rect 30196 30277 30205 30311
rect 30205 30277 30239 30311
rect 30239 30277 30248 30311
rect 30196 30268 30248 30277
rect 36912 30268 36964 30320
rect 24124 30243 24176 30252
rect 20444 30175 20496 30184
rect 20444 30141 20453 30175
rect 20453 30141 20487 30175
rect 20487 30141 20496 30175
rect 20444 30132 20496 30141
rect 24124 30209 24133 30243
rect 24133 30209 24167 30243
rect 24167 30209 24176 30243
rect 24124 30200 24176 30209
rect 26332 30200 26384 30252
rect 30656 30243 30708 30252
rect 30656 30209 30665 30243
rect 30665 30209 30699 30243
rect 30699 30209 30708 30243
rect 30656 30200 30708 30209
rect 33508 30200 33560 30252
rect 40960 30243 41012 30252
rect 40960 30209 40969 30243
rect 40969 30209 41003 30243
rect 41003 30209 41012 30243
rect 40960 30200 41012 30209
rect 25780 30132 25832 30184
rect 20996 30064 21048 30116
rect 23848 30107 23900 30116
rect 4620 29996 4672 30048
rect 4896 30039 4948 30048
rect 4896 30005 4905 30039
rect 4905 30005 4939 30039
rect 4939 30005 4948 30039
rect 4896 29996 4948 30005
rect 8484 30039 8536 30048
rect 8484 30005 8493 30039
rect 8493 30005 8527 30039
rect 8527 30005 8536 30039
rect 8484 29996 8536 30005
rect 10692 29996 10744 30048
rect 12992 29996 13044 30048
rect 17132 29996 17184 30048
rect 21732 30039 21784 30048
rect 21732 30005 21741 30039
rect 21741 30005 21775 30039
rect 21775 30005 21784 30039
rect 21732 29996 21784 30005
rect 23848 30073 23857 30107
rect 23857 30073 23891 30107
rect 23891 30073 23900 30107
rect 23848 30064 23900 30073
rect 24124 30064 24176 30116
rect 25780 29996 25832 30048
rect 28264 30132 28316 30184
rect 28540 30132 28592 30184
rect 26516 30064 26568 30116
rect 26056 29996 26108 30048
rect 28172 30064 28224 30116
rect 32864 30132 32916 30184
rect 30288 30064 30340 30116
rect 28080 29996 28132 30048
rect 29092 29996 29144 30048
rect 32496 30064 32548 30116
rect 35256 30175 35308 30184
rect 35256 30141 35265 30175
rect 35265 30141 35299 30175
rect 35299 30141 35308 30175
rect 35256 30132 35308 30141
rect 33508 30064 33560 30116
rect 36452 30132 36504 30184
rect 37280 30107 37332 30116
rect 37280 30073 37289 30107
rect 37289 30073 37323 30107
rect 37323 30073 37332 30107
rect 37280 30064 37332 30073
rect 38568 30175 38620 30184
rect 38568 30141 38577 30175
rect 38577 30141 38611 30175
rect 38611 30141 38620 30175
rect 38568 30132 38620 30141
rect 39212 30132 39264 30184
rect 37556 30064 37608 30116
rect 41328 30200 41380 30252
rect 43352 30200 43404 30252
rect 41972 30132 42024 30184
rect 35992 30039 36044 30048
rect 35992 30005 36001 30039
rect 36001 30005 36035 30039
rect 36035 30005 36044 30039
rect 35992 29996 36044 30005
rect 37740 30039 37792 30048
rect 37740 30005 37749 30039
rect 37749 30005 37783 30039
rect 37783 30005 37792 30039
rect 37740 29996 37792 30005
rect 38384 29996 38436 30048
rect 38936 30039 38988 30048
rect 38936 30005 38945 30039
rect 38945 30005 38979 30039
rect 38979 30005 38988 30039
rect 38936 29996 38988 30005
rect 39764 30039 39816 30048
rect 39764 30005 39773 30039
rect 39773 30005 39807 30039
rect 39807 30005 39816 30039
rect 39764 29996 39816 30005
rect 41880 30039 41932 30048
rect 41880 30005 41889 30039
rect 41889 30005 41923 30039
rect 41923 30005 41932 30039
rect 41880 29996 41932 30005
rect 42524 29996 42576 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 4896 29792 4948 29844
rect 5264 29835 5316 29844
rect 5264 29801 5273 29835
rect 5273 29801 5307 29835
rect 5307 29801 5316 29835
rect 5264 29792 5316 29801
rect 6000 29792 6052 29844
rect 7840 29792 7892 29844
rect 9036 29835 9088 29844
rect 9036 29801 9045 29835
rect 9045 29801 9079 29835
rect 9079 29801 9088 29835
rect 9036 29792 9088 29801
rect 10876 29792 10928 29844
rect 10968 29792 11020 29844
rect 13820 29835 13872 29844
rect 13820 29801 13829 29835
rect 13829 29801 13863 29835
rect 13863 29801 13872 29835
rect 13820 29792 13872 29801
rect 18880 29792 18932 29844
rect 20904 29792 20956 29844
rect 23480 29835 23532 29844
rect 23480 29801 23489 29835
rect 23489 29801 23523 29835
rect 23523 29801 23532 29835
rect 26332 29835 26384 29844
rect 23480 29792 23532 29801
rect 26332 29801 26341 29835
rect 26341 29801 26375 29835
rect 26375 29801 26384 29835
rect 26332 29792 26384 29801
rect 31944 29835 31996 29844
rect 31944 29801 31953 29835
rect 31953 29801 31987 29835
rect 31987 29801 31996 29835
rect 31944 29792 31996 29801
rect 34152 29835 34204 29844
rect 34152 29801 34161 29835
rect 34161 29801 34195 29835
rect 34195 29801 34204 29835
rect 34152 29792 34204 29801
rect 34612 29835 34664 29844
rect 34612 29801 34621 29835
rect 34621 29801 34655 29835
rect 34655 29801 34664 29835
rect 34612 29792 34664 29801
rect 35256 29792 35308 29844
rect 36084 29792 36136 29844
rect 37648 29792 37700 29844
rect 38200 29792 38252 29844
rect 41144 29792 41196 29844
rect 42524 29835 42576 29844
rect 42524 29801 42533 29835
rect 42533 29801 42567 29835
rect 42567 29801 42576 29835
rect 42524 29792 42576 29801
rect 4620 29724 4672 29776
rect 7564 29767 7616 29776
rect 7564 29733 7573 29767
rect 7573 29733 7607 29767
rect 7607 29733 7616 29767
rect 7564 29724 7616 29733
rect 7932 29724 7984 29776
rect 8852 29724 8904 29776
rect 12716 29724 12768 29776
rect 5080 29656 5132 29708
rect 5908 29656 5960 29708
rect 6276 29699 6328 29708
rect 6276 29665 6285 29699
rect 6285 29665 6319 29699
rect 6319 29665 6328 29699
rect 6276 29656 6328 29665
rect 10140 29656 10192 29708
rect 10784 29699 10836 29708
rect 10784 29665 10793 29699
rect 10793 29665 10827 29699
rect 10827 29665 10836 29699
rect 10784 29656 10836 29665
rect 11428 29656 11480 29708
rect 3884 29588 3936 29640
rect 6460 29588 6512 29640
rect 8208 29588 8260 29640
rect 12440 29631 12492 29640
rect 12440 29597 12449 29631
rect 12449 29597 12483 29631
rect 12483 29597 12492 29631
rect 12440 29588 12492 29597
rect 12532 29588 12584 29640
rect 13176 29724 13228 29776
rect 15476 29767 15528 29776
rect 15476 29733 15485 29767
rect 15485 29733 15519 29767
rect 15519 29733 15528 29767
rect 15476 29724 15528 29733
rect 16948 29724 17000 29776
rect 17408 29724 17460 29776
rect 22284 29724 22336 29776
rect 23112 29724 23164 29776
rect 24860 29724 24912 29776
rect 25780 29724 25832 29776
rect 26240 29724 26292 29776
rect 26700 29767 26752 29776
rect 26700 29733 26709 29767
rect 26709 29733 26743 29767
rect 26743 29733 26752 29767
rect 26700 29724 26752 29733
rect 28080 29724 28132 29776
rect 30196 29724 30248 29776
rect 30472 29724 30524 29776
rect 32864 29767 32916 29776
rect 13636 29656 13688 29708
rect 18696 29699 18748 29708
rect 18696 29665 18705 29699
rect 18705 29665 18739 29699
rect 18739 29665 18748 29699
rect 18696 29656 18748 29665
rect 18788 29656 18840 29708
rect 21088 29699 21140 29708
rect 21088 29665 21097 29699
rect 21097 29665 21131 29699
rect 21131 29665 21140 29699
rect 21088 29656 21140 29665
rect 21456 29656 21508 29708
rect 22100 29656 22152 29708
rect 24124 29656 24176 29708
rect 28172 29699 28224 29708
rect 28172 29665 28181 29699
rect 28181 29665 28215 29699
rect 28215 29665 28224 29699
rect 28172 29656 28224 29665
rect 28632 29699 28684 29708
rect 28632 29665 28641 29699
rect 28641 29665 28675 29699
rect 28675 29665 28684 29699
rect 28632 29656 28684 29665
rect 30564 29699 30616 29708
rect 30564 29665 30573 29699
rect 30573 29665 30607 29699
rect 30607 29665 30616 29699
rect 30564 29656 30616 29665
rect 31024 29656 31076 29708
rect 32496 29656 32548 29708
rect 32864 29733 32873 29767
rect 32873 29733 32907 29767
rect 32907 29733 32916 29767
rect 32864 29724 32916 29733
rect 33968 29724 34020 29776
rect 35992 29767 36044 29776
rect 35992 29733 36001 29767
rect 36001 29733 36035 29767
rect 36035 29733 36044 29767
rect 35992 29724 36044 29733
rect 32772 29656 32824 29708
rect 33508 29656 33560 29708
rect 36084 29699 36136 29708
rect 15384 29631 15436 29640
rect 15384 29597 15393 29631
rect 15393 29597 15427 29631
rect 15427 29597 15436 29631
rect 15384 29588 15436 29597
rect 16120 29588 16172 29640
rect 17592 29631 17644 29640
rect 17592 29597 17601 29631
rect 17601 29597 17635 29631
rect 17635 29597 17644 29631
rect 17592 29588 17644 29597
rect 18972 29631 19024 29640
rect 18972 29597 18981 29631
rect 18981 29597 19015 29631
rect 19015 29597 19024 29631
rect 18972 29588 19024 29597
rect 23388 29588 23440 29640
rect 23940 29588 23992 29640
rect 28908 29631 28960 29640
rect 28908 29597 28917 29631
rect 28917 29597 28951 29631
rect 28951 29597 28960 29631
rect 28908 29588 28960 29597
rect 31208 29631 31260 29640
rect 31208 29597 31217 29631
rect 31217 29597 31251 29631
rect 31251 29597 31260 29631
rect 31208 29588 31260 29597
rect 33876 29588 33928 29640
rect 36084 29665 36093 29699
rect 36093 29665 36127 29699
rect 36127 29665 36136 29699
rect 36084 29656 36136 29665
rect 38476 29724 38528 29776
rect 40592 29767 40644 29776
rect 40592 29733 40601 29767
rect 40601 29733 40635 29767
rect 40635 29733 40644 29767
rect 40592 29724 40644 29733
rect 43536 29767 43588 29776
rect 43536 29733 43545 29767
rect 43545 29733 43579 29767
rect 43579 29733 43588 29767
rect 43536 29724 43588 29733
rect 37556 29656 37608 29708
rect 41696 29656 41748 29708
rect 36820 29631 36872 29640
rect 36820 29597 36829 29631
rect 36829 29597 36863 29631
rect 36863 29597 36872 29631
rect 36820 29588 36872 29597
rect 37188 29588 37240 29640
rect 39672 29588 39724 29640
rect 18236 29520 18288 29572
rect 22468 29520 22520 29572
rect 23756 29520 23808 29572
rect 23848 29520 23900 29572
rect 27160 29563 27212 29572
rect 27160 29529 27169 29563
rect 27169 29529 27203 29563
rect 27203 29529 27212 29563
rect 27160 29520 27212 29529
rect 41144 29631 41196 29640
rect 41144 29597 41153 29631
rect 41153 29597 41187 29631
rect 41187 29597 41196 29631
rect 41144 29588 41196 29597
rect 43444 29631 43496 29640
rect 43444 29597 43453 29631
rect 43453 29597 43487 29631
rect 43487 29597 43496 29631
rect 43444 29588 43496 29597
rect 41236 29520 41288 29572
rect 42340 29520 42392 29572
rect 3148 29452 3200 29504
rect 4068 29452 4120 29504
rect 6920 29495 6972 29504
rect 6920 29461 6929 29495
rect 6929 29461 6963 29495
rect 6963 29461 6972 29495
rect 6920 29452 6972 29461
rect 11520 29452 11572 29504
rect 13176 29452 13228 29504
rect 13360 29495 13412 29504
rect 13360 29461 13369 29495
rect 13369 29461 13403 29495
rect 13403 29461 13412 29495
rect 13360 29452 13412 29461
rect 13728 29452 13780 29504
rect 20260 29452 20312 29504
rect 20444 29495 20496 29504
rect 20444 29461 20453 29495
rect 20453 29461 20487 29495
rect 20487 29461 20496 29495
rect 20444 29452 20496 29461
rect 25504 29495 25556 29504
rect 25504 29461 25513 29495
rect 25513 29461 25547 29495
rect 25547 29461 25556 29495
rect 25504 29452 25556 29461
rect 39580 29495 39632 29504
rect 39580 29461 39589 29495
rect 39589 29461 39623 29495
rect 39623 29461 39632 29495
rect 39580 29452 39632 29461
rect 40316 29495 40368 29504
rect 40316 29461 40325 29495
rect 40325 29461 40359 29495
rect 40359 29461 40368 29495
rect 40316 29452 40368 29461
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 5172 29291 5224 29300
rect 5172 29257 5181 29291
rect 5181 29257 5215 29291
rect 5215 29257 5224 29291
rect 5172 29248 5224 29257
rect 8208 29291 8260 29300
rect 8208 29257 8217 29291
rect 8217 29257 8251 29291
rect 8251 29257 8260 29291
rect 8208 29248 8260 29257
rect 10784 29291 10836 29300
rect 10784 29257 10793 29291
rect 10793 29257 10827 29291
rect 10827 29257 10836 29291
rect 10784 29248 10836 29257
rect 12992 29248 13044 29300
rect 11612 29180 11664 29232
rect 12716 29180 12768 29232
rect 7196 29155 7248 29164
rect 2964 29087 3016 29096
rect 2964 29053 2973 29087
rect 2973 29053 3007 29087
rect 3007 29053 3016 29087
rect 2964 29044 3016 29053
rect 3240 29087 3292 29096
rect 3240 29053 3249 29087
rect 3249 29053 3283 29087
rect 3283 29053 3292 29087
rect 3240 29044 3292 29053
rect 7196 29121 7205 29155
rect 7205 29121 7239 29155
rect 7239 29121 7248 29155
rect 7196 29112 7248 29121
rect 12808 29155 12860 29164
rect 12808 29121 12817 29155
rect 12817 29121 12851 29155
rect 12851 29121 12860 29155
rect 12808 29112 12860 29121
rect 10784 29044 10836 29096
rect 15476 29248 15528 29300
rect 17868 29291 17920 29300
rect 17868 29257 17877 29291
rect 17877 29257 17911 29291
rect 17911 29257 17920 29291
rect 17868 29248 17920 29257
rect 21456 29291 21508 29300
rect 21456 29257 21465 29291
rect 21465 29257 21499 29291
rect 21499 29257 21508 29291
rect 21456 29248 21508 29257
rect 23112 29291 23164 29300
rect 23112 29257 23121 29291
rect 23121 29257 23155 29291
rect 23155 29257 23164 29291
rect 23112 29248 23164 29257
rect 23388 29291 23440 29300
rect 23388 29257 23397 29291
rect 23397 29257 23431 29291
rect 23431 29257 23440 29291
rect 23388 29248 23440 29257
rect 23940 29291 23992 29300
rect 23940 29257 23949 29291
rect 23949 29257 23983 29291
rect 23983 29257 23992 29291
rect 23940 29248 23992 29257
rect 24584 29291 24636 29300
rect 24584 29257 24593 29291
rect 24593 29257 24627 29291
rect 24627 29257 24636 29291
rect 24584 29248 24636 29257
rect 24860 29291 24912 29300
rect 24860 29257 24869 29291
rect 24869 29257 24903 29291
rect 24903 29257 24912 29291
rect 24860 29248 24912 29257
rect 14648 29155 14700 29164
rect 14648 29121 14657 29155
rect 14657 29121 14691 29155
rect 14691 29121 14700 29155
rect 14648 29112 14700 29121
rect 15384 29112 15436 29164
rect 20444 29155 20496 29164
rect 20444 29121 20453 29155
rect 20453 29121 20487 29155
rect 20487 29121 20496 29155
rect 20444 29112 20496 29121
rect 18880 29087 18932 29096
rect 4528 28976 4580 29028
rect 6920 29019 6972 29028
rect 3976 28908 4028 28960
rect 6920 28985 6929 29019
rect 6929 28985 6963 29019
rect 6963 28985 6972 29019
rect 6920 28976 6972 28985
rect 5816 28951 5868 28960
rect 5816 28917 5825 28951
rect 5825 28917 5859 28951
rect 5859 28917 5868 28951
rect 5816 28908 5868 28917
rect 5908 28908 5960 28960
rect 8484 28976 8536 29028
rect 9128 29019 9180 29028
rect 9128 28985 9137 29019
rect 9137 28985 9171 29019
rect 9171 28985 9180 29019
rect 9128 28976 9180 28985
rect 7932 28951 7984 28960
rect 7932 28917 7941 28951
rect 7941 28917 7975 28951
rect 7975 28917 7984 28951
rect 7932 28908 7984 28917
rect 8944 28951 8996 28960
rect 8944 28917 8953 28951
rect 8953 28917 8987 28951
rect 8987 28917 8996 28951
rect 9864 28976 9916 29028
rect 12532 29019 12584 29028
rect 12532 28985 12541 29019
rect 12541 28985 12575 29019
rect 12575 28985 12584 29019
rect 12532 28976 12584 28985
rect 10140 28951 10192 28960
rect 8944 28908 8996 28917
rect 10140 28917 10149 28951
rect 10149 28917 10183 28951
rect 10183 28917 10192 28951
rect 10140 28908 10192 28917
rect 10876 28908 10928 28960
rect 11428 28951 11480 28960
rect 11428 28917 11437 28951
rect 11437 28917 11471 28951
rect 11471 28917 11480 28951
rect 11428 28908 11480 28917
rect 13820 28976 13872 29028
rect 18880 29053 18889 29087
rect 18889 29053 18923 29087
rect 18923 29053 18932 29087
rect 18880 29044 18932 29053
rect 20168 29087 20220 29096
rect 20168 29053 20177 29087
rect 20177 29053 20211 29087
rect 20211 29053 20220 29087
rect 20168 29044 20220 29053
rect 20260 29044 20312 29096
rect 21732 29044 21784 29096
rect 22008 29087 22060 29096
rect 14740 28976 14792 29028
rect 16488 29019 16540 29028
rect 16488 28985 16497 29019
rect 16497 28985 16531 29019
rect 16531 28985 16540 29019
rect 16488 28976 16540 28985
rect 15476 28908 15528 28960
rect 17224 28976 17276 29028
rect 17500 29019 17552 29028
rect 17500 28985 17509 29019
rect 17509 28985 17543 29019
rect 17543 28985 17552 29019
rect 17500 28976 17552 28985
rect 17040 28908 17092 28960
rect 18696 28908 18748 28960
rect 19432 28908 19484 28960
rect 21088 28951 21140 28960
rect 21088 28917 21097 28951
rect 21097 28917 21131 28951
rect 21131 28917 21140 28951
rect 21088 28908 21140 28917
rect 21180 28908 21232 28960
rect 22008 29053 22017 29087
rect 22017 29053 22051 29087
rect 22051 29053 22060 29087
rect 22008 29044 22060 29053
rect 22100 29044 22152 29096
rect 26424 29248 26476 29300
rect 26700 29291 26752 29300
rect 26700 29257 26709 29291
rect 26709 29257 26743 29291
rect 26743 29257 26752 29291
rect 26700 29248 26752 29257
rect 28080 29291 28132 29300
rect 28080 29257 28089 29291
rect 28089 29257 28123 29291
rect 28123 29257 28132 29291
rect 28080 29248 28132 29257
rect 30196 29291 30248 29300
rect 30196 29257 30205 29291
rect 30205 29257 30239 29291
rect 30239 29257 30248 29291
rect 30196 29248 30248 29257
rect 32404 29248 32456 29300
rect 32496 29291 32548 29300
rect 32496 29257 32505 29291
rect 32505 29257 32539 29291
rect 32539 29257 32548 29291
rect 32772 29291 32824 29300
rect 32496 29248 32548 29257
rect 32772 29257 32781 29291
rect 32781 29257 32815 29291
rect 32815 29257 32824 29291
rect 32772 29248 32824 29257
rect 34612 29248 34664 29300
rect 37556 29291 37608 29300
rect 37556 29257 37565 29291
rect 37565 29257 37599 29291
rect 37599 29257 37608 29291
rect 37556 29248 37608 29257
rect 39580 29248 39632 29300
rect 40592 29248 40644 29300
rect 41880 29248 41932 29300
rect 43536 29248 43588 29300
rect 39672 29223 39724 29232
rect 39672 29189 39681 29223
rect 39681 29189 39715 29223
rect 39715 29189 39724 29223
rect 39672 29180 39724 29189
rect 25504 29112 25556 29164
rect 25872 29112 25924 29164
rect 31208 29155 31260 29164
rect 27160 29087 27212 29096
rect 27160 29053 27169 29087
rect 27169 29053 27203 29087
rect 27203 29053 27212 29087
rect 27160 29044 27212 29053
rect 31208 29121 31217 29155
rect 31217 29121 31251 29155
rect 31251 29121 31260 29155
rect 31208 29112 31260 29121
rect 32956 29112 33008 29164
rect 33416 29112 33468 29164
rect 37188 29155 37240 29164
rect 37188 29121 37197 29155
rect 37197 29121 37231 29155
rect 37231 29121 37240 29155
rect 37188 29112 37240 29121
rect 37280 29112 37332 29164
rect 38108 29155 38160 29164
rect 38108 29121 38117 29155
rect 38117 29121 38151 29155
rect 38151 29121 38160 29155
rect 38108 29112 38160 29121
rect 40040 29112 40092 29164
rect 41236 29112 41288 29164
rect 42524 29180 42576 29232
rect 42432 29155 42484 29164
rect 42432 29121 42441 29155
rect 42441 29121 42475 29155
rect 42475 29121 42484 29155
rect 42432 29112 42484 29121
rect 43444 29112 43496 29164
rect 34152 29044 34204 29096
rect 35256 29087 35308 29096
rect 35256 29053 35265 29087
rect 35265 29053 35299 29087
rect 35299 29053 35308 29087
rect 35256 29044 35308 29053
rect 35992 29044 36044 29096
rect 36912 29044 36964 29096
rect 37556 29044 37608 29096
rect 28264 28976 28316 29028
rect 28632 28976 28684 29028
rect 30564 29019 30616 29028
rect 30564 28985 30573 29019
rect 30573 28985 30607 29019
rect 30607 28985 30616 29019
rect 30564 28976 30616 28985
rect 25412 28908 25464 28960
rect 28080 28908 28132 28960
rect 29460 28951 29512 28960
rect 29460 28917 29469 28951
rect 29469 28917 29503 28951
rect 29503 28917 29512 28951
rect 29460 28908 29512 28917
rect 30380 28908 30432 28960
rect 33508 28976 33560 29028
rect 35716 29019 35768 29028
rect 31116 28951 31168 28960
rect 31116 28917 31125 28951
rect 31125 28917 31159 28951
rect 31159 28917 31168 28951
rect 31116 28908 31168 28917
rect 34152 28951 34204 28960
rect 34152 28917 34161 28951
rect 34161 28917 34195 28951
rect 34195 28917 34204 28951
rect 34152 28908 34204 28917
rect 35716 28985 35725 29019
rect 35725 28985 35759 29019
rect 35759 28985 35768 29019
rect 35716 28976 35768 28985
rect 36084 29019 36136 29028
rect 36084 28985 36093 29019
rect 36093 28985 36127 29019
rect 36127 28985 36136 29019
rect 36084 28976 36136 28985
rect 37648 28908 37700 28960
rect 38200 28908 38252 28960
rect 38568 28908 38620 28960
rect 41236 29019 41288 29028
rect 41236 28985 41245 29019
rect 41245 28985 41279 29019
rect 41279 28985 41288 29019
rect 41236 28976 41288 28985
rect 41972 28976 42024 29028
rect 41144 28908 41196 28960
rect 41696 28908 41748 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 6920 28704 6972 28756
rect 4068 28636 4120 28688
rect 5172 28636 5224 28688
rect 4620 28568 4672 28620
rect 6460 28636 6512 28688
rect 6552 28679 6604 28688
rect 6552 28645 6561 28679
rect 6561 28645 6595 28679
rect 6595 28645 6604 28679
rect 7932 28704 7984 28756
rect 9496 28704 9548 28756
rect 12164 28704 12216 28756
rect 12808 28704 12860 28756
rect 6552 28636 6604 28645
rect 7196 28636 7248 28688
rect 9128 28636 9180 28688
rect 9864 28679 9916 28688
rect 9864 28645 9873 28679
rect 9873 28645 9907 28679
rect 9907 28645 9916 28679
rect 9864 28636 9916 28645
rect 11520 28679 11572 28688
rect 11520 28645 11529 28679
rect 11529 28645 11563 28679
rect 11563 28645 11572 28679
rect 11520 28636 11572 28645
rect 11612 28679 11664 28688
rect 11612 28645 11621 28679
rect 11621 28645 11655 28679
rect 11655 28645 11664 28679
rect 11612 28636 11664 28645
rect 12532 28636 12584 28688
rect 13912 28636 13964 28688
rect 14648 28636 14700 28688
rect 16120 28704 16172 28756
rect 22100 28747 22152 28756
rect 22100 28713 22109 28747
rect 22109 28713 22143 28747
rect 22143 28713 22152 28747
rect 22100 28704 22152 28713
rect 26240 28747 26292 28756
rect 26240 28713 26249 28747
rect 26249 28713 26283 28747
rect 26283 28713 26292 28747
rect 26240 28704 26292 28713
rect 31208 28704 31260 28756
rect 35440 28704 35492 28756
rect 36912 28747 36964 28756
rect 36912 28713 36921 28747
rect 36921 28713 36955 28747
rect 36955 28713 36964 28747
rect 36912 28704 36964 28713
rect 38108 28747 38160 28756
rect 38108 28713 38117 28747
rect 38117 28713 38151 28747
rect 38151 28713 38160 28747
rect 38108 28704 38160 28713
rect 40132 28704 40184 28756
rect 41144 28747 41196 28756
rect 16488 28636 16540 28688
rect 16764 28636 16816 28688
rect 17500 28636 17552 28688
rect 20076 28636 20128 28688
rect 27160 28679 27212 28688
rect 27160 28645 27169 28679
rect 27169 28645 27203 28679
rect 27203 28645 27212 28679
rect 27160 28636 27212 28645
rect 30380 28636 30432 28688
rect 33416 28679 33468 28688
rect 33416 28645 33425 28679
rect 33425 28645 33459 28679
rect 33459 28645 33468 28679
rect 33416 28636 33468 28645
rect 35256 28679 35308 28688
rect 35256 28645 35265 28679
rect 35265 28645 35299 28679
rect 35299 28645 35308 28679
rect 35256 28636 35308 28645
rect 38200 28636 38252 28688
rect 38476 28636 38528 28688
rect 40040 28679 40092 28688
rect 40040 28645 40049 28679
rect 40049 28645 40083 28679
rect 40083 28645 40092 28679
rect 40040 28636 40092 28645
rect 41144 28713 41153 28747
rect 41153 28713 41187 28747
rect 41187 28713 41196 28747
rect 41144 28704 41196 28713
rect 41788 28679 41840 28688
rect 41788 28645 41797 28679
rect 41797 28645 41831 28679
rect 41831 28645 41840 28679
rect 41788 28636 41840 28645
rect 41880 28679 41932 28688
rect 41880 28645 41889 28679
rect 41889 28645 41923 28679
rect 41923 28645 41932 28679
rect 41880 28636 41932 28645
rect 42800 28636 42852 28688
rect 7656 28568 7708 28620
rect 12440 28568 12492 28620
rect 14924 28568 14976 28620
rect 18144 28568 18196 28620
rect 18972 28568 19024 28620
rect 19340 28568 19392 28620
rect 20260 28568 20312 28620
rect 21456 28611 21508 28620
rect 3884 28500 3936 28552
rect 6460 28543 6512 28552
rect 6460 28509 6469 28543
rect 6469 28509 6503 28543
rect 6503 28509 6512 28543
rect 6460 28500 6512 28509
rect 9312 28500 9364 28552
rect 11980 28500 12032 28552
rect 12532 28500 12584 28552
rect 13728 28543 13780 28552
rect 13728 28509 13737 28543
rect 13737 28509 13771 28543
rect 13771 28509 13780 28543
rect 13728 28500 13780 28509
rect 14372 28500 14424 28552
rect 16580 28500 16632 28552
rect 17224 28543 17276 28552
rect 17224 28509 17233 28543
rect 17233 28509 17267 28543
rect 17267 28509 17276 28543
rect 17224 28500 17276 28509
rect 17684 28500 17736 28552
rect 21456 28577 21465 28611
rect 21465 28577 21499 28611
rect 21499 28577 21508 28611
rect 21456 28568 21508 28577
rect 22468 28611 22520 28620
rect 22468 28577 22477 28611
rect 22477 28577 22511 28611
rect 22511 28577 22520 28611
rect 22468 28568 22520 28577
rect 23112 28568 23164 28620
rect 25412 28611 25464 28620
rect 25412 28577 25421 28611
rect 25421 28577 25455 28611
rect 25455 28577 25464 28611
rect 25412 28568 25464 28577
rect 21180 28500 21232 28552
rect 21548 28543 21600 28552
rect 21548 28509 21557 28543
rect 21557 28509 21591 28543
rect 21591 28509 21600 28543
rect 21548 28500 21600 28509
rect 23204 28543 23256 28552
rect 23204 28509 23213 28543
rect 23213 28509 23247 28543
rect 23247 28509 23256 28543
rect 23204 28500 23256 28509
rect 20168 28432 20220 28484
rect 25228 28500 25280 28552
rect 27528 28568 27580 28620
rect 27988 28611 28040 28620
rect 27988 28577 27997 28611
rect 27997 28577 28031 28611
rect 28031 28577 28040 28611
rect 27988 28568 28040 28577
rect 28264 28611 28316 28620
rect 28264 28577 28273 28611
rect 28273 28577 28307 28611
rect 28307 28577 28316 28611
rect 28264 28568 28316 28577
rect 31024 28611 31076 28620
rect 31024 28577 31033 28611
rect 31033 28577 31067 28611
rect 31067 28577 31076 28611
rect 31024 28568 31076 28577
rect 32956 28568 33008 28620
rect 34612 28568 34664 28620
rect 35624 28568 35676 28620
rect 35992 28568 36044 28620
rect 36820 28568 36872 28620
rect 38844 28568 38896 28620
rect 27160 28500 27212 28552
rect 29184 28500 29236 28552
rect 33324 28543 33376 28552
rect 33324 28509 33333 28543
rect 33333 28509 33367 28543
rect 33367 28509 33376 28543
rect 33324 28500 33376 28509
rect 33692 28543 33744 28552
rect 33692 28509 33701 28543
rect 33701 28509 33735 28543
rect 33735 28509 33744 28543
rect 33692 28500 33744 28509
rect 36452 28543 36504 28552
rect 36452 28509 36461 28543
rect 36461 28509 36495 28543
rect 36495 28509 36504 28543
rect 36452 28500 36504 28509
rect 40684 28500 40736 28552
rect 42524 28500 42576 28552
rect 39948 28432 40000 28484
rect 41236 28432 41288 28484
rect 3240 28364 3292 28416
rect 5356 28364 5408 28416
rect 8208 28364 8260 28416
rect 15292 28364 15344 28416
rect 16028 28364 16080 28416
rect 18236 28364 18288 28416
rect 24216 28364 24268 28416
rect 28264 28364 28316 28416
rect 30196 28407 30248 28416
rect 30196 28373 30205 28407
rect 30205 28373 30239 28407
rect 30239 28373 30248 28407
rect 30196 28364 30248 28373
rect 30472 28407 30524 28416
rect 30472 28373 30481 28407
rect 30481 28373 30515 28407
rect 30515 28373 30524 28407
rect 30472 28364 30524 28373
rect 31208 28407 31260 28416
rect 31208 28373 31217 28407
rect 31217 28373 31251 28407
rect 31251 28373 31260 28407
rect 31208 28364 31260 28373
rect 32496 28364 32548 28416
rect 33140 28364 33192 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 5172 28203 5224 28212
rect 5172 28169 5181 28203
rect 5181 28169 5215 28203
rect 5215 28169 5224 28203
rect 5172 28160 5224 28169
rect 6552 28160 6604 28212
rect 7656 28203 7708 28212
rect 7656 28169 7665 28203
rect 7665 28169 7699 28203
rect 7699 28169 7708 28203
rect 7656 28160 7708 28169
rect 9312 28203 9364 28212
rect 9312 28169 9321 28203
rect 9321 28169 9355 28203
rect 9355 28169 9364 28203
rect 9312 28160 9364 28169
rect 9864 28160 9916 28212
rect 11520 28160 11572 28212
rect 13636 28160 13688 28212
rect 13912 28160 13964 28212
rect 14372 28203 14424 28212
rect 14372 28169 14381 28203
rect 14381 28169 14415 28203
rect 14415 28169 14424 28203
rect 14372 28160 14424 28169
rect 6460 28092 6512 28144
rect 8760 28135 8812 28144
rect 8760 28101 8769 28135
rect 8769 28101 8803 28135
rect 8803 28101 8812 28135
rect 8760 28092 8812 28101
rect 4068 28067 4120 28076
rect 4068 28033 4077 28067
rect 4077 28033 4111 28067
rect 4111 28033 4120 28067
rect 4068 28024 4120 28033
rect 8208 28067 8260 28076
rect 8208 28033 8217 28067
rect 8217 28033 8251 28067
rect 8251 28033 8260 28067
rect 8208 28024 8260 28033
rect 2964 27956 3016 28008
rect 3792 27999 3844 28008
rect 3792 27965 3801 27999
rect 3801 27965 3835 27999
rect 3835 27965 3844 27999
rect 3792 27956 3844 27965
rect 3884 27956 3936 28008
rect 5172 27956 5224 28008
rect 7564 27956 7616 28008
rect 7932 27888 7984 27940
rect 11612 28092 11664 28144
rect 10876 28067 10928 28076
rect 10876 28033 10885 28067
rect 10885 28033 10919 28067
rect 10919 28033 10928 28067
rect 10876 28024 10928 28033
rect 12164 28024 12216 28076
rect 13820 28024 13872 28076
rect 15660 28160 15712 28212
rect 16764 28203 16816 28212
rect 16764 28169 16773 28203
rect 16773 28169 16807 28203
rect 16807 28169 16816 28203
rect 16764 28160 16816 28169
rect 17132 28203 17184 28212
rect 17132 28169 17141 28203
rect 17141 28169 17175 28203
rect 17175 28169 17184 28203
rect 17132 28160 17184 28169
rect 18144 28160 18196 28212
rect 21640 28160 21692 28212
rect 27160 28203 27212 28212
rect 27160 28169 27169 28203
rect 27169 28169 27203 28203
rect 27203 28169 27212 28203
rect 27160 28160 27212 28169
rect 27252 28160 27304 28212
rect 27528 28203 27580 28212
rect 27528 28169 27537 28203
rect 27537 28169 27571 28203
rect 27571 28169 27580 28203
rect 27528 28160 27580 28169
rect 32956 28160 33008 28212
rect 33324 28160 33376 28212
rect 35624 28160 35676 28212
rect 38844 28203 38896 28212
rect 38844 28169 38853 28203
rect 38853 28169 38887 28203
rect 38887 28169 38896 28203
rect 38844 28160 38896 28169
rect 40132 28203 40184 28212
rect 40132 28169 40141 28203
rect 40141 28169 40175 28203
rect 40175 28169 40184 28203
rect 40132 28160 40184 28169
rect 42800 28203 42852 28212
rect 42800 28169 42809 28203
rect 42809 28169 42843 28203
rect 42843 28169 42852 28203
rect 42800 28160 42852 28169
rect 16948 28092 17000 28144
rect 20996 28092 21048 28144
rect 21180 28135 21232 28144
rect 21180 28101 21189 28135
rect 21189 28101 21223 28135
rect 21223 28101 21232 28135
rect 21180 28092 21232 28101
rect 21456 28092 21508 28144
rect 23112 28135 23164 28144
rect 23112 28101 23121 28135
rect 23121 28101 23155 28135
rect 23155 28101 23164 28135
rect 23112 28092 23164 28101
rect 25136 28092 25188 28144
rect 16120 28067 16172 28076
rect 16120 28033 16129 28067
rect 16129 28033 16163 28067
rect 16163 28033 16172 28067
rect 16120 28024 16172 28033
rect 12808 27999 12860 28008
rect 12808 27965 12817 27999
rect 12817 27965 12851 27999
rect 12851 27965 12860 27999
rect 12808 27956 12860 27965
rect 17040 28024 17092 28076
rect 19064 28024 19116 28076
rect 22284 28024 22336 28076
rect 22468 28024 22520 28076
rect 25228 28024 25280 28076
rect 18236 27999 18288 28008
rect 18236 27965 18245 27999
rect 18245 27965 18279 27999
rect 18279 27965 18288 27999
rect 18236 27956 18288 27965
rect 10692 27931 10744 27940
rect 10692 27897 10701 27931
rect 10701 27897 10735 27931
rect 10735 27897 10744 27931
rect 10692 27888 10744 27897
rect 4620 27863 4672 27872
rect 4620 27829 4629 27863
rect 4629 27829 4663 27863
rect 4663 27829 4672 27863
rect 4620 27820 4672 27829
rect 7840 27820 7892 27872
rect 9680 27863 9732 27872
rect 9680 27829 9689 27863
rect 9689 27829 9723 27863
rect 9723 27829 9732 27863
rect 9680 27820 9732 27829
rect 9956 27863 10008 27872
rect 9956 27829 9965 27863
rect 9965 27829 9999 27863
rect 9999 27829 10008 27863
rect 9956 27820 10008 27829
rect 12532 27888 12584 27940
rect 14096 27888 14148 27940
rect 12900 27820 12952 27872
rect 14924 27863 14976 27872
rect 14924 27829 14933 27863
rect 14933 27829 14967 27863
rect 14967 27829 14976 27863
rect 14924 27820 14976 27829
rect 15660 27888 15712 27940
rect 17868 27888 17920 27940
rect 20352 27888 20404 27940
rect 21088 27956 21140 28008
rect 25044 27999 25096 28008
rect 21456 27888 21508 27940
rect 21824 27931 21876 27940
rect 21824 27897 21833 27931
rect 21833 27897 21867 27931
rect 21867 27897 21876 27931
rect 21824 27888 21876 27897
rect 21916 27931 21968 27940
rect 21916 27897 21925 27931
rect 21925 27897 21959 27931
rect 21959 27897 21968 27931
rect 21916 27888 21968 27897
rect 16028 27820 16080 27872
rect 18972 27820 19024 27872
rect 24124 27820 24176 27872
rect 25044 27965 25053 27999
rect 25053 27965 25087 27999
rect 25087 27965 25096 27999
rect 25044 27956 25096 27965
rect 25412 28092 25464 28144
rect 29460 28092 29512 28144
rect 34612 28135 34664 28144
rect 34612 28101 34621 28135
rect 34621 28101 34655 28135
rect 34655 28101 34664 28135
rect 34612 28092 34664 28101
rect 25504 28067 25556 28076
rect 25504 28033 25513 28067
rect 25513 28033 25547 28067
rect 25547 28033 25556 28067
rect 25504 28024 25556 28033
rect 28908 28024 28960 28076
rect 30472 28024 30524 28076
rect 27528 27956 27580 28008
rect 27804 27999 27856 28008
rect 27804 27965 27813 27999
rect 27813 27965 27847 27999
rect 27847 27965 27856 27999
rect 27804 27956 27856 27965
rect 28264 27956 28316 28008
rect 32496 27956 32548 28008
rect 34152 27956 34204 28008
rect 35808 28092 35860 28144
rect 38016 28092 38068 28144
rect 35716 28024 35768 28076
rect 36636 28024 36688 28076
rect 38292 27956 38344 28008
rect 29736 27888 29788 27940
rect 31116 27888 31168 27940
rect 38476 27931 38528 27940
rect 38476 27897 38485 27931
rect 38485 27897 38519 27931
rect 38519 27897 38528 27931
rect 38476 27888 38528 27897
rect 40408 27956 40460 28008
rect 41052 27956 41104 28008
rect 39764 27888 39816 27940
rect 25596 27820 25648 27872
rect 28356 27820 28408 27872
rect 30932 27820 30984 27872
rect 31024 27863 31076 27872
rect 31024 27829 31033 27863
rect 31033 27829 31067 27863
rect 31067 27829 31076 27863
rect 31024 27820 31076 27829
rect 33416 27820 33468 27872
rect 33784 27820 33836 27872
rect 36176 27863 36228 27872
rect 36176 27829 36185 27863
rect 36185 27829 36219 27863
rect 36219 27829 36228 27863
rect 36176 27820 36228 27829
rect 38016 27863 38068 27872
rect 38016 27829 38025 27863
rect 38025 27829 38059 27863
rect 38059 27829 38068 27863
rect 38016 27820 38068 27829
rect 39580 27820 39632 27872
rect 39672 27863 39724 27872
rect 39672 27829 39681 27863
rect 39681 27829 39715 27863
rect 39715 27829 39724 27863
rect 39672 27820 39724 27829
rect 41512 27820 41564 27872
rect 42524 27931 42576 27940
rect 42524 27897 42533 27931
rect 42533 27897 42567 27931
rect 42567 27897 42576 27931
rect 42524 27888 42576 27897
rect 44824 27820 44876 27872
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 4620 27616 4672 27668
rect 6460 27616 6512 27668
rect 9772 27659 9824 27668
rect 9772 27625 9781 27659
rect 9781 27625 9815 27659
rect 9815 27625 9824 27659
rect 9772 27616 9824 27625
rect 10876 27659 10928 27668
rect 10876 27625 10885 27659
rect 10885 27625 10919 27659
rect 10919 27625 10928 27659
rect 10876 27616 10928 27625
rect 15292 27616 15344 27668
rect 3976 27548 4028 27600
rect 4804 27548 4856 27600
rect 7840 27548 7892 27600
rect 8484 27548 8536 27600
rect 8760 27591 8812 27600
rect 8760 27557 8769 27591
rect 8769 27557 8803 27591
rect 8803 27557 8812 27591
rect 8760 27548 8812 27557
rect 12808 27548 12860 27600
rect 16580 27616 16632 27668
rect 18236 27659 18288 27668
rect 18236 27625 18245 27659
rect 18245 27625 18279 27659
rect 18279 27625 18288 27659
rect 18236 27616 18288 27625
rect 19340 27659 19392 27668
rect 19340 27625 19349 27659
rect 19349 27625 19383 27659
rect 19383 27625 19392 27659
rect 19340 27616 19392 27625
rect 20352 27659 20404 27668
rect 20352 27625 20361 27659
rect 20361 27625 20395 27659
rect 20395 27625 20404 27659
rect 20352 27616 20404 27625
rect 21180 27616 21232 27668
rect 21916 27616 21968 27668
rect 23204 27616 23256 27668
rect 23664 27659 23716 27668
rect 23664 27625 23673 27659
rect 23673 27625 23707 27659
rect 23707 27625 23716 27659
rect 23664 27616 23716 27625
rect 25044 27659 25096 27668
rect 25044 27625 25053 27659
rect 25053 27625 25087 27659
rect 25087 27625 25096 27659
rect 25044 27616 25096 27625
rect 25412 27659 25464 27668
rect 25412 27625 25421 27659
rect 25421 27625 25455 27659
rect 25455 27625 25464 27659
rect 25412 27616 25464 27625
rect 27620 27616 27672 27668
rect 27804 27616 27856 27668
rect 29184 27659 29236 27668
rect 29184 27625 29193 27659
rect 29193 27625 29227 27659
rect 29227 27625 29236 27659
rect 29184 27616 29236 27625
rect 29736 27659 29788 27668
rect 29736 27625 29745 27659
rect 29745 27625 29779 27659
rect 29779 27625 29788 27659
rect 29736 27616 29788 27625
rect 35992 27616 36044 27668
rect 36636 27659 36688 27668
rect 36636 27625 36645 27659
rect 36645 27625 36679 27659
rect 36679 27625 36688 27659
rect 36636 27616 36688 27625
rect 15476 27591 15528 27600
rect 15476 27557 15485 27591
rect 15485 27557 15519 27591
rect 15519 27557 15528 27591
rect 17040 27591 17092 27600
rect 15476 27548 15528 27557
rect 17040 27557 17049 27591
rect 17049 27557 17083 27591
rect 17083 27557 17092 27591
rect 17040 27548 17092 27557
rect 17592 27591 17644 27600
rect 17592 27557 17601 27591
rect 17601 27557 17635 27591
rect 17635 27557 17644 27591
rect 17592 27548 17644 27557
rect 24492 27548 24544 27600
rect 32312 27591 32364 27600
rect 32312 27557 32321 27591
rect 32321 27557 32355 27591
rect 32355 27557 32364 27591
rect 32312 27548 32364 27557
rect 33784 27548 33836 27600
rect 4068 27523 4120 27532
rect 4068 27489 4077 27523
rect 4077 27489 4111 27523
rect 4111 27489 4120 27523
rect 4068 27480 4120 27489
rect 5632 27480 5684 27532
rect 6368 27480 6420 27532
rect 7012 27480 7064 27532
rect 9864 27523 9916 27532
rect 9864 27489 9873 27523
rect 9873 27489 9907 27523
rect 9907 27489 9916 27523
rect 9864 27480 9916 27489
rect 12256 27523 12308 27532
rect 6828 27412 6880 27464
rect 9588 27412 9640 27464
rect 12256 27489 12265 27523
rect 12265 27489 12299 27523
rect 12299 27489 12308 27523
rect 12256 27480 12308 27489
rect 12716 27523 12768 27532
rect 12716 27489 12725 27523
rect 12725 27489 12759 27523
rect 12759 27489 12768 27523
rect 12716 27480 12768 27489
rect 13728 27523 13780 27532
rect 13728 27489 13737 27523
rect 13737 27489 13771 27523
rect 13771 27489 13780 27523
rect 13728 27480 13780 27489
rect 19064 27480 19116 27532
rect 19892 27480 19944 27532
rect 26148 27480 26200 27532
rect 27344 27480 27396 27532
rect 27988 27523 28040 27532
rect 27988 27489 27997 27523
rect 27997 27489 28031 27523
rect 28031 27489 28040 27523
rect 27988 27480 28040 27489
rect 28264 27523 28316 27532
rect 28264 27489 28273 27523
rect 28273 27489 28307 27523
rect 28307 27489 28316 27523
rect 28264 27480 28316 27489
rect 35348 27523 35400 27532
rect 35348 27489 35357 27523
rect 35357 27489 35391 27523
rect 35391 27489 35400 27523
rect 35348 27480 35400 27489
rect 35716 27480 35768 27532
rect 39212 27616 39264 27668
rect 41788 27616 41840 27668
rect 38016 27548 38068 27600
rect 38292 27591 38344 27600
rect 38292 27557 38301 27591
rect 38301 27557 38335 27591
rect 38335 27557 38344 27591
rect 39764 27591 39816 27600
rect 38292 27548 38344 27557
rect 39764 27557 39773 27591
rect 39773 27557 39807 27591
rect 39807 27557 39816 27591
rect 39764 27548 39816 27557
rect 39856 27591 39908 27600
rect 39856 27557 39865 27591
rect 39865 27557 39899 27591
rect 39899 27557 39908 27591
rect 39856 27548 39908 27557
rect 41512 27548 41564 27600
rect 42432 27591 42484 27600
rect 42432 27557 42441 27591
rect 42441 27557 42475 27591
rect 42475 27557 42484 27591
rect 42432 27548 42484 27557
rect 43904 27480 43956 27532
rect 16028 27455 16080 27464
rect 16028 27421 16037 27455
rect 16037 27421 16071 27455
rect 16071 27421 16080 27455
rect 16028 27412 16080 27421
rect 12808 27344 12860 27396
rect 16856 27344 16908 27396
rect 21088 27412 21140 27464
rect 24032 27455 24084 27464
rect 24032 27421 24041 27455
rect 24041 27421 24075 27455
rect 24075 27421 24084 27455
rect 24032 27412 24084 27421
rect 24308 27455 24360 27464
rect 24308 27421 24317 27455
rect 24317 27421 24351 27455
rect 24351 27421 24360 27455
rect 24308 27412 24360 27421
rect 29000 27412 29052 27464
rect 32220 27455 32272 27464
rect 32220 27421 32229 27455
rect 32229 27421 32263 27455
rect 32263 27421 32272 27455
rect 32220 27412 32272 27421
rect 24400 27344 24452 27396
rect 25964 27344 26016 27396
rect 31024 27344 31076 27396
rect 31116 27344 31168 27396
rect 33416 27412 33468 27464
rect 34428 27455 34480 27464
rect 34428 27421 34437 27455
rect 34437 27421 34471 27455
rect 34471 27421 34480 27455
rect 34428 27412 34480 27421
rect 35900 27455 35952 27464
rect 35900 27421 35909 27455
rect 35909 27421 35943 27455
rect 35943 27421 35952 27455
rect 35900 27412 35952 27421
rect 38568 27455 38620 27464
rect 38568 27421 38577 27455
rect 38577 27421 38611 27455
rect 38611 27421 38620 27455
rect 38568 27412 38620 27421
rect 40040 27455 40092 27464
rect 40040 27421 40049 27455
rect 40049 27421 40083 27455
rect 40083 27421 40092 27455
rect 40040 27412 40092 27421
rect 32772 27344 32824 27396
rect 40776 27387 40828 27396
rect 40776 27353 40785 27387
rect 40785 27353 40819 27387
rect 40819 27353 40828 27387
rect 40776 27344 40828 27353
rect 42432 27344 42484 27396
rect 3976 27276 4028 27328
rect 7564 27276 7616 27328
rect 12716 27276 12768 27328
rect 13452 27276 13504 27328
rect 14188 27319 14240 27328
rect 14188 27285 14197 27319
rect 14197 27285 14231 27319
rect 14231 27285 14240 27319
rect 14188 27276 14240 27285
rect 17960 27276 18012 27328
rect 21916 27276 21968 27328
rect 25596 27276 25648 27328
rect 30564 27276 30616 27328
rect 30840 27319 30892 27328
rect 30840 27285 30849 27319
rect 30849 27285 30883 27319
rect 30883 27285 30892 27319
rect 30840 27276 30892 27285
rect 32680 27276 32732 27328
rect 34428 27276 34480 27328
rect 35992 27276 36044 27328
rect 37832 27276 37884 27328
rect 38660 27276 38712 27328
rect 43168 27276 43220 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 5172 27115 5224 27124
rect 5172 27081 5181 27115
rect 5181 27081 5215 27115
rect 5215 27081 5224 27115
rect 5172 27072 5224 27081
rect 7012 27072 7064 27124
rect 7656 27072 7708 27124
rect 7840 27072 7892 27124
rect 10784 27115 10836 27124
rect 10784 27081 10793 27115
rect 10793 27081 10827 27115
rect 10827 27081 10836 27115
rect 10784 27072 10836 27081
rect 12164 27115 12216 27124
rect 12164 27081 12173 27115
rect 12173 27081 12207 27115
rect 12207 27081 12216 27115
rect 12164 27072 12216 27081
rect 12624 27072 12676 27124
rect 14096 27115 14148 27124
rect 14096 27081 14105 27115
rect 14105 27081 14139 27115
rect 14139 27081 14148 27115
rect 14096 27072 14148 27081
rect 15292 27072 15344 27124
rect 17040 27072 17092 27124
rect 19064 27115 19116 27124
rect 19064 27081 19073 27115
rect 19073 27081 19107 27115
rect 19107 27081 19116 27115
rect 19064 27072 19116 27081
rect 24492 27072 24544 27124
rect 26976 27072 27028 27124
rect 27988 27072 28040 27124
rect 29000 27115 29052 27124
rect 29000 27081 29009 27115
rect 29009 27081 29043 27115
rect 29043 27081 29052 27115
rect 29000 27072 29052 27081
rect 29736 27115 29788 27124
rect 29736 27081 29745 27115
rect 29745 27081 29779 27115
rect 29779 27081 29788 27115
rect 29736 27072 29788 27081
rect 30564 27115 30616 27124
rect 30564 27081 30573 27115
rect 30573 27081 30607 27115
rect 30607 27081 30616 27115
rect 30564 27072 30616 27081
rect 30932 27072 30984 27124
rect 32496 27072 32548 27124
rect 33416 27115 33468 27124
rect 33416 27081 33425 27115
rect 33425 27081 33459 27115
rect 33459 27081 33468 27115
rect 33416 27072 33468 27081
rect 36452 27072 36504 27124
rect 8484 27004 8536 27056
rect 9680 27004 9732 27056
rect 6828 26979 6880 26988
rect 4252 26911 4304 26920
rect 4252 26877 4261 26911
rect 4261 26877 4295 26911
rect 4295 26877 4304 26911
rect 4252 26868 4304 26877
rect 6828 26945 6837 26979
rect 6837 26945 6871 26979
rect 6871 26945 6880 26979
rect 6828 26936 6880 26945
rect 9772 26936 9824 26988
rect 11980 26936 12032 26988
rect 12808 26979 12860 26988
rect 12808 26945 12817 26979
rect 12817 26945 12851 26979
rect 12851 26945 12860 26979
rect 12808 26936 12860 26945
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 15476 26979 15528 26988
rect 15476 26945 15485 26979
rect 15485 26945 15519 26979
rect 15519 26945 15528 26979
rect 15476 26936 15528 26945
rect 7748 26868 7800 26920
rect 9588 26868 9640 26920
rect 12256 26868 12308 26920
rect 17592 26936 17644 26988
rect 18144 26979 18196 26988
rect 18144 26945 18153 26979
rect 18153 26945 18187 26979
rect 18187 26945 18196 26979
rect 18144 26936 18196 26945
rect 18420 26979 18472 26988
rect 18420 26945 18429 26979
rect 18429 26945 18463 26979
rect 18463 26945 18472 26979
rect 18420 26936 18472 26945
rect 17960 26868 18012 26920
rect 23940 27004 23992 27056
rect 24860 27004 24912 27056
rect 30196 27004 30248 27056
rect 32312 27004 32364 27056
rect 21548 26979 21600 26988
rect 21548 26945 21557 26979
rect 21557 26945 21591 26979
rect 21591 26945 21600 26979
rect 21548 26936 21600 26945
rect 23664 26979 23716 26988
rect 23664 26945 23673 26979
rect 23673 26945 23707 26979
rect 23707 26945 23716 26979
rect 23664 26936 23716 26945
rect 26884 26979 26936 26988
rect 26884 26945 26893 26979
rect 26893 26945 26927 26979
rect 26927 26945 26936 26979
rect 26884 26936 26936 26945
rect 27344 26979 27396 26988
rect 27344 26945 27353 26979
rect 27353 26945 27387 26979
rect 27387 26945 27396 26979
rect 27344 26936 27396 26945
rect 30840 26979 30892 26988
rect 30840 26945 30849 26979
rect 30849 26945 30883 26979
rect 30883 26945 30892 26979
rect 30840 26936 30892 26945
rect 31116 26979 31168 26988
rect 31116 26945 31125 26979
rect 31125 26945 31159 26979
rect 31159 26945 31168 26979
rect 31116 26936 31168 26945
rect 32680 26936 32732 26988
rect 32772 26979 32824 26988
rect 32772 26945 32781 26979
rect 32781 26945 32815 26979
rect 32815 26945 32824 26979
rect 38016 27072 38068 27124
rect 39764 27072 39816 27124
rect 43168 27115 43220 27124
rect 43168 27081 43177 27115
rect 43177 27081 43211 27115
rect 43211 27081 43220 27115
rect 43168 27072 43220 27081
rect 43904 27072 43956 27124
rect 38292 27004 38344 27056
rect 41512 27047 41564 27056
rect 41512 27013 41521 27047
rect 41521 27013 41555 27047
rect 41555 27013 41564 27047
rect 41512 27004 41564 27013
rect 42340 27047 42392 27056
rect 42340 27013 42349 27047
rect 42349 27013 42383 27047
rect 42383 27013 42392 27047
rect 42340 27004 42392 27013
rect 32772 26936 32824 26945
rect 38568 26979 38620 26988
rect 38568 26945 38577 26979
rect 38577 26945 38611 26979
rect 38611 26945 38620 26979
rect 38568 26936 38620 26945
rect 41604 26936 41656 26988
rect 4804 26800 4856 26852
rect 5448 26800 5500 26852
rect 6920 26800 6972 26852
rect 10600 26800 10652 26852
rect 12532 26843 12584 26852
rect 12532 26809 12541 26843
rect 12541 26809 12575 26843
rect 12575 26809 12584 26843
rect 12532 26800 12584 26809
rect 12624 26843 12676 26852
rect 12624 26809 12633 26843
rect 12633 26809 12667 26843
rect 12667 26809 12676 26843
rect 12624 26800 12676 26809
rect 14096 26800 14148 26852
rect 18236 26843 18288 26852
rect 18236 26809 18245 26843
rect 18245 26809 18279 26843
rect 18279 26809 18288 26843
rect 19892 26843 19944 26852
rect 18236 26800 18288 26809
rect 19892 26809 19901 26843
rect 19901 26809 19935 26843
rect 19935 26809 19944 26843
rect 26056 26868 26108 26920
rect 26240 26911 26292 26920
rect 26240 26877 26249 26911
rect 26249 26877 26283 26911
rect 26283 26877 26292 26911
rect 26608 26911 26660 26920
rect 26240 26868 26292 26877
rect 26608 26877 26617 26911
rect 26617 26877 26651 26911
rect 26651 26877 26660 26911
rect 26608 26868 26660 26877
rect 26792 26911 26844 26920
rect 26792 26877 26801 26911
rect 26801 26877 26835 26911
rect 26835 26877 26844 26911
rect 26792 26868 26844 26877
rect 27712 26868 27764 26920
rect 28816 26868 28868 26920
rect 19892 26800 19944 26809
rect 5632 26732 5684 26784
rect 8760 26775 8812 26784
rect 8760 26741 8769 26775
rect 8769 26741 8803 26775
rect 8803 26741 8812 26775
rect 8760 26732 8812 26741
rect 12348 26732 12400 26784
rect 13728 26732 13780 26784
rect 15936 26732 15988 26784
rect 17316 26732 17368 26784
rect 20904 26732 20956 26784
rect 21180 26732 21232 26784
rect 23664 26800 23716 26852
rect 25780 26800 25832 26852
rect 27344 26800 27396 26852
rect 29736 26800 29788 26852
rect 22468 26775 22520 26784
rect 22468 26741 22477 26775
rect 22477 26741 22511 26775
rect 22511 26741 22520 26775
rect 22468 26732 22520 26741
rect 27804 26732 27856 26784
rect 35440 26911 35492 26920
rect 35440 26877 35449 26911
rect 35449 26877 35483 26911
rect 35483 26877 35492 26911
rect 35440 26868 35492 26877
rect 35716 26911 35768 26920
rect 35716 26877 35725 26911
rect 35725 26877 35759 26911
rect 35759 26877 35768 26911
rect 35716 26868 35768 26877
rect 40868 26868 40920 26920
rect 41328 26868 41380 26920
rect 42984 26868 43036 26920
rect 30288 26732 30340 26784
rect 30564 26732 30616 26784
rect 32496 26843 32548 26852
rect 32496 26809 32505 26843
rect 32505 26809 32539 26843
rect 32539 26809 32548 26843
rect 32496 26800 32548 26809
rect 36084 26800 36136 26852
rect 33784 26775 33836 26784
rect 33784 26741 33793 26775
rect 33793 26741 33827 26775
rect 33827 26741 33836 26775
rect 33784 26732 33836 26741
rect 36176 26732 36228 26784
rect 38660 26843 38712 26852
rect 38660 26809 38669 26843
rect 38669 26809 38703 26843
rect 38703 26809 38712 26843
rect 38660 26800 38712 26809
rect 39948 26800 40000 26852
rect 41512 26800 41564 26852
rect 39764 26775 39816 26784
rect 39764 26741 39773 26775
rect 39773 26741 39807 26775
rect 39807 26741 39816 26775
rect 39764 26732 39816 26741
rect 41052 26732 41104 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 4068 26528 4120 26580
rect 4252 26528 4304 26580
rect 5816 26571 5868 26580
rect 5816 26537 5825 26571
rect 5825 26537 5859 26571
rect 5859 26537 5868 26571
rect 5816 26528 5868 26537
rect 6920 26528 6972 26580
rect 7564 26571 7616 26580
rect 7564 26537 7573 26571
rect 7573 26537 7607 26571
rect 7607 26537 7616 26571
rect 7564 26528 7616 26537
rect 3792 26392 3844 26444
rect 4712 26460 4764 26512
rect 10140 26528 10192 26580
rect 12256 26528 12308 26580
rect 10324 26460 10376 26512
rect 10600 26503 10652 26512
rect 10600 26469 10603 26503
rect 10603 26469 10637 26503
rect 10637 26469 10652 26503
rect 10600 26460 10652 26469
rect 12532 26528 12584 26580
rect 13912 26528 13964 26580
rect 16856 26571 16908 26580
rect 16856 26537 16865 26571
rect 16865 26537 16899 26571
rect 16899 26537 16908 26571
rect 16856 26528 16908 26537
rect 18144 26528 18196 26580
rect 21088 26571 21140 26580
rect 21088 26537 21097 26571
rect 21097 26537 21131 26571
rect 21131 26537 21140 26571
rect 21088 26528 21140 26537
rect 21548 26528 21600 26580
rect 24032 26571 24084 26580
rect 24032 26537 24041 26571
rect 24041 26537 24075 26571
rect 24075 26537 24084 26571
rect 24032 26528 24084 26537
rect 24492 26528 24544 26580
rect 28632 26528 28684 26580
rect 14188 26460 14240 26512
rect 15476 26503 15528 26512
rect 15476 26469 15485 26503
rect 15485 26469 15519 26503
rect 15519 26469 15528 26503
rect 15476 26460 15528 26469
rect 16028 26503 16080 26512
rect 16028 26469 16037 26503
rect 16037 26469 16071 26503
rect 16071 26469 16080 26503
rect 16028 26460 16080 26469
rect 17500 26460 17552 26512
rect 22468 26460 22520 26512
rect 25780 26460 25832 26512
rect 27344 26460 27396 26512
rect 33324 26528 33376 26580
rect 35348 26571 35400 26580
rect 35348 26537 35357 26571
rect 35357 26537 35391 26571
rect 35391 26537 35400 26571
rect 35348 26528 35400 26537
rect 35716 26571 35768 26580
rect 35716 26537 35725 26571
rect 35725 26537 35759 26571
rect 35759 26537 35768 26571
rect 35716 26528 35768 26537
rect 36176 26528 36228 26580
rect 32036 26460 32088 26512
rect 4620 26435 4672 26444
rect 4620 26401 4629 26435
rect 4629 26401 4663 26435
rect 4663 26401 4672 26435
rect 4620 26392 4672 26401
rect 5632 26435 5684 26444
rect 5632 26401 5641 26435
rect 5641 26401 5675 26435
rect 5675 26401 5684 26435
rect 5632 26392 5684 26401
rect 8576 26435 8628 26444
rect 8576 26401 8585 26435
rect 8585 26401 8619 26435
rect 8619 26401 8628 26435
rect 8576 26392 8628 26401
rect 12256 26392 12308 26444
rect 13544 26435 13596 26444
rect 13544 26401 13553 26435
rect 13553 26401 13587 26435
rect 13587 26401 13596 26435
rect 13544 26392 13596 26401
rect 14004 26435 14056 26444
rect 14004 26401 14013 26435
rect 14013 26401 14047 26435
rect 14047 26401 14056 26435
rect 14004 26392 14056 26401
rect 19064 26435 19116 26444
rect 6920 26324 6972 26376
rect 10232 26367 10284 26376
rect 10232 26333 10241 26367
rect 10241 26333 10275 26367
rect 10275 26333 10284 26367
rect 10232 26324 10284 26333
rect 13728 26324 13780 26376
rect 15844 26324 15896 26376
rect 17224 26324 17276 26376
rect 18420 26324 18472 26376
rect 9956 26256 10008 26308
rect 19064 26401 19073 26435
rect 19073 26401 19107 26435
rect 19107 26401 19116 26435
rect 19064 26392 19116 26401
rect 21272 26392 21324 26444
rect 30748 26392 30800 26444
rect 32128 26392 32180 26444
rect 33784 26460 33836 26512
rect 38292 26460 38344 26512
rect 39580 26503 39632 26512
rect 39580 26469 39589 26503
rect 39589 26469 39623 26503
rect 39623 26469 39632 26503
rect 39580 26460 39632 26469
rect 41052 26528 41104 26580
rect 43076 26528 43128 26580
rect 39764 26460 39816 26512
rect 40776 26460 40828 26512
rect 41604 26503 41656 26512
rect 41604 26469 41613 26503
rect 41613 26469 41647 26503
rect 41647 26469 41656 26503
rect 41604 26460 41656 26469
rect 41880 26503 41932 26512
rect 41880 26469 41889 26503
rect 41889 26469 41923 26503
rect 41923 26469 41932 26503
rect 41880 26460 41932 26469
rect 42432 26503 42484 26512
rect 42432 26469 42441 26503
rect 42441 26469 42475 26503
rect 42475 26469 42484 26503
rect 42432 26460 42484 26469
rect 43536 26503 43588 26512
rect 43536 26469 43545 26503
rect 43545 26469 43579 26503
rect 43579 26469 43588 26503
rect 43536 26460 43588 26469
rect 34796 26435 34848 26444
rect 34796 26401 34805 26435
rect 34805 26401 34839 26435
rect 34839 26401 34848 26435
rect 34796 26392 34848 26401
rect 35900 26435 35952 26444
rect 35900 26401 35909 26435
rect 35909 26401 35943 26435
rect 35943 26401 35952 26435
rect 35900 26392 35952 26401
rect 22928 26324 22980 26376
rect 25596 26324 25648 26376
rect 26884 26367 26936 26376
rect 26884 26333 26893 26367
rect 26893 26333 26927 26367
rect 26927 26333 26936 26367
rect 26884 26324 26936 26333
rect 29092 26324 29144 26376
rect 33140 26324 33192 26376
rect 38476 26324 38528 26376
rect 41788 26367 41840 26376
rect 41788 26333 41797 26367
rect 41797 26333 41831 26367
rect 41831 26333 41840 26367
rect 41788 26324 41840 26333
rect 22836 26256 22888 26308
rect 25136 26299 25188 26308
rect 9864 26231 9916 26240
rect 9864 26197 9873 26231
rect 9873 26197 9907 26231
rect 9907 26197 9916 26231
rect 9864 26188 9916 26197
rect 12532 26188 12584 26240
rect 12716 26231 12768 26240
rect 12716 26197 12725 26231
rect 12725 26197 12759 26231
rect 12759 26197 12768 26231
rect 12716 26188 12768 26197
rect 14556 26231 14608 26240
rect 14556 26197 14565 26231
rect 14565 26197 14599 26231
rect 14599 26197 14608 26231
rect 14556 26188 14608 26197
rect 19984 26231 20036 26240
rect 19984 26197 19993 26231
rect 19993 26197 20027 26231
rect 20027 26197 20036 26231
rect 19984 26188 20036 26197
rect 21824 26231 21876 26240
rect 21824 26197 21833 26231
rect 21833 26197 21867 26231
rect 21867 26197 21876 26231
rect 21824 26188 21876 26197
rect 22284 26188 22336 26240
rect 25136 26265 25145 26299
rect 25145 26265 25179 26299
rect 25179 26265 25188 26299
rect 25136 26256 25188 26265
rect 27528 26256 27580 26308
rect 31116 26256 31168 26308
rect 32220 26256 32272 26308
rect 33876 26299 33928 26308
rect 33876 26265 33885 26299
rect 33885 26265 33919 26299
rect 33919 26265 33928 26299
rect 33876 26256 33928 26265
rect 38568 26299 38620 26308
rect 38568 26265 38577 26299
rect 38577 26265 38611 26299
rect 38611 26265 38620 26299
rect 38568 26256 38620 26265
rect 40316 26256 40368 26308
rect 42524 26256 42576 26308
rect 28264 26188 28316 26240
rect 31300 26231 31352 26240
rect 31300 26197 31309 26231
rect 31309 26197 31343 26231
rect 31343 26197 31352 26231
rect 31300 26188 31352 26197
rect 32680 26231 32732 26240
rect 32680 26197 32689 26231
rect 32689 26197 32723 26231
rect 32723 26197 32732 26231
rect 32680 26188 32732 26197
rect 33416 26188 33468 26240
rect 37740 26188 37792 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 4712 26027 4764 26036
rect 4712 25993 4721 26027
rect 4721 25993 4755 26027
rect 4755 25993 4764 26027
rect 4712 25984 4764 25993
rect 4804 25984 4856 26036
rect 5356 26027 5408 26036
rect 5356 25993 5365 26027
rect 5365 25993 5399 26027
rect 5399 25993 5408 26027
rect 5356 25984 5408 25993
rect 6828 25984 6880 26036
rect 3976 25916 4028 25968
rect 5632 25848 5684 25900
rect 4344 25780 4396 25832
rect 6828 25712 6880 25764
rect 7656 25780 7708 25832
rect 12164 25984 12216 26036
rect 13544 26027 13596 26036
rect 13544 25993 13553 26027
rect 13553 25993 13587 26027
rect 13587 25993 13596 26027
rect 13544 25984 13596 25993
rect 14096 26027 14148 26036
rect 14096 25993 14105 26027
rect 14105 25993 14139 26027
rect 14139 25993 14148 26027
rect 14096 25984 14148 25993
rect 14924 25984 14976 26036
rect 15476 26027 15528 26036
rect 15476 25993 15485 26027
rect 15485 25993 15519 26027
rect 15519 25993 15528 26027
rect 15476 25984 15528 25993
rect 15936 26027 15988 26036
rect 15936 25993 15945 26027
rect 15945 25993 15979 26027
rect 15979 25993 15988 26027
rect 15936 25984 15988 25993
rect 17224 25984 17276 26036
rect 17500 26027 17552 26036
rect 17500 25993 17509 26027
rect 17509 25993 17543 26027
rect 17543 25993 17552 26027
rect 17500 25984 17552 25993
rect 18236 25984 18288 26036
rect 19064 26027 19116 26036
rect 19064 25993 19073 26027
rect 19073 25993 19107 26027
rect 19107 25993 19116 26027
rect 19064 25984 19116 25993
rect 21272 25984 21324 26036
rect 22468 25984 22520 26036
rect 22928 25984 22980 26036
rect 24492 25984 24544 26036
rect 25596 26027 25648 26036
rect 25596 25993 25605 26027
rect 25605 25993 25639 26027
rect 25639 25993 25648 26027
rect 25596 25984 25648 25993
rect 26884 25984 26936 26036
rect 28632 26027 28684 26036
rect 28632 25993 28641 26027
rect 28641 25993 28675 26027
rect 28675 25993 28684 26027
rect 28632 25984 28684 25993
rect 33784 26027 33836 26036
rect 33784 25993 33793 26027
rect 33793 25993 33827 26027
rect 33827 25993 33836 26027
rect 33784 25984 33836 25993
rect 34796 25984 34848 26036
rect 35348 26027 35400 26036
rect 35348 25993 35357 26027
rect 35357 25993 35391 26027
rect 35391 25993 35400 26027
rect 35348 25984 35400 25993
rect 37740 26027 37792 26036
rect 37740 25993 37749 26027
rect 37749 25993 37783 26027
rect 37783 25993 37792 26027
rect 37740 25984 37792 25993
rect 39580 25984 39632 26036
rect 41788 25984 41840 26036
rect 42340 25984 42392 26036
rect 43076 26027 43128 26036
rect 43076 25993 43085 26027
rect 43085 25993 43119 26027
rect 43119 25993 43128 26027
rect 43076 25984 43128 25993
rect 10600 25959 10652 25968
rect 10600 25925 10609 25959
rect 10609 25925 10643 25959
rect 10643 25925 10652 25959
rect 10600 25916 10652 25925
rect 3056 25644 3108 25696
rect 3700 25687 3752 25696
rect 3700 25653 3709 25687
rect 3709 25653 3743 25687
rect 3743 25653 3752 25687
rect 3700 25644 3752 25653
rect 4620 25644 4672 25696
rect 6000 25687 6052 25696
rect 6000 25653 6009 25687
rect 6009 25653 6043 25687
rect 6043 25653 6052 25687
rect 6000 25644 6052 25653
rect 6920 25687 6972 25696
rect 6920 25653 6929 25687
rect 6929 25653 6963 25687
rect 6963 25653 6972 25687
rect 6920 25644 6972 25653
rect 8576 25848 8628 25900
rect 11152 25848 11204 25900
rect 8208 25687 8260 25696
rect 8208 25653 8217 25687
rect 8217 25653 8251 25687
rect 8251 25653 8260 25687
rect 8208 25644 8260 25653
rect 9956 25780 10008 25832
rect 10232 25755 10284 25764
rect 10232 25721 10241 25755
rect 10241 25721 10275 25755
rect 10275 25721 10284 25755
rect 10232 25712 10284 25721
rect 9864 25644 9916 25696
rect 12532 25780 12584 25832
rect 21824 25916 21876 25968
rect 22284 25959 22336 25968
rect 22284 25925 22293 25959
rect 22293 25925 22327 25959
rect 22327 25925 22336 25959
rect 22284 25916 22336 25925
rect 24676 25916 24728 25968
rect 25228 25916 25280 25968
rect 26608 25916 26660 25968
rect 30840 25916 30892 25968
rect 32036 25916 32088 25968
rect 32312 25916 32364 25968
rect 33140 25916 33192 25968
rect 38568 25959 38620 25968
rect 38568 25925 38577 25959
rect 38577 25925 38611 25959
rect 38611 25925 38620 25959
rect 38568 25916 38620 25925
rect 42248 25959 42300 25968
rect 42248 25925 42257 25959
rect 42257 25925 42291 25959
rect 42291 25925 42300 25959
rect 42248 25916 42300 25925
rect 14556 25848 14608 25900
rect 19984 25848 20036 25900
rect 21732 25848 21784 25900
rect 27344 25848 27396 25900
rect 31300 25891 31352 25900
rect 31300 25857 31309 25891
rect 31309 25857 31343 25891
rect 31343 25857 31352 25891
rect 31300 25848 31352 25857
rect 31576 25891 31628 25900
rect 31576 25857 31585 25891
rect 31585 25857 31619 25891
rect 31619 25857 31628 25891
rect 31576 25848 31628 25857
rect 33692 25848 33744 25900
rect 14740 25712 14792 25764
rect 17316 25780 17368 25832
rect 18052 25780 18104 25832
rect 26608 25823 26660 25832
rect 26608 25789 26617 25823
rect 26617 25789 26651 25823
rect 26651 25789 26660 25823
rect 26608 25780 26660 25789
rect 26792 25780 26844 25832
rect 28264 25780 28316 25832
rect 28356 25780 28408 25832
rect 31024 25780 31076 25832
rect 34060 25780 34112 25832
rect 37832 25848 37884 25900
rect 38384 25848 38436 25900
rect 38476 25848 38528 25900
rect 36084 25823 36136 25832
rect 36084 25789 36093 25823
rect 36093 25789 36127 25823
rect 36127 25789 36136 25823
rect 36084 25780 36136 25789
rect 40960 25823 41012 25832
rect 40960 25789 40969 25823
rect 40969 25789 41003 25823
rect 41003 25789 41012 25823
rect 40960 25780 41012 25789
rect 42708 25780 42760 25832
rect 44640 25823 44692 25832
rect 44640 25789 44649 25823
rect 44649 25789 44683 25823
rect 44683 25789 44692 25823
rect 44640 25780 44692 25789
rect 11888 25687 11940 25696
rect 11888 25653 11897 25687
rect 11897 25653 11931 25687
rect 11931 25653 11940 25687
rect 11888 25644 11940 25653
rect 12256 25687 12308 25696
rect 12256 25653 12265 25687
rect 12265 25653 12299 25687
rect 12299 25653 12308 25687
rect 12256 25644 12308 25653
rect 13176 25644 13228 25696
rect 17132 25687 17184 25696
rect 17132 25653 17141 25687
rect 17141 25653 17175 25687
rect 17175 25653 17184 25687
rect 17132 25644 17184 25653
rect 21180 25712 21232 25764
rect 21732 25755 21784 25764
rect 21732 25721 21741 25755
rect 21741 25721 21775 25755
rect 21775 25721 21784 25755
rect 21732 25712 21784 25721
rect 21824 25755 21876 25764
rect 21824 25721 21833 25755
rect 21833 25721 21867 25755
rect 21867 25721 21876 25755
rect 24216 25755 24268 25764
rect 21824 25712 21876 25721
rect 24216 25721 24225 25755
rect 24225 25721 24259 25755
rect 24259 25721 24268 25755
rect 24216 25712 24268 25721
rect 24492 25712 24544 25764
rect 27160 25755 27212 25764
rect 27160 25721 27169 25755
rect 27169 25721 27203 25755
rect 27203 25721 27212 25755
rect 27160 25712 27212 25721
rect 32864 25755 32916 25764
rect 18880 25644 18932 25696
rect 22928 25644 22980 25696
rect 24032 25644 24084 25696
rect 27988 25687 28040 25696
rect 27988 25653 27997 25687
rect 27997 25653 28031 25687
rect 28031 25653 28040 25687
rect 27988 25644 28040 25653
rect 29092 25687 29144 25696
rect 29092 25653 29101 25687
rect 29101 25653 29135 25687
rect 29135 25653 29144 25687
rect 29092 25644 29144 25653
rect 29644 25644 29696 25696
rect 30656 25644 30708 25696
rect 30748 25644 30800 25696
rect 31208 25644 31260 25696
rect 32864 25721 32873 25755
rect 32873 25721 32907 25755
rect 32907 25721 32916 25755
rect 32864 25712 32916 25721
rect 33140 25712 33192 25764
rect 33876 25712 33928 25764
rect 35164 25712 35216 25764
rect 36176 25712 36228 25764
rect 37740 25712 37792 25764
rect 41696 25755 41748 25764
rect 34704 25644 34756 25696
rect 37004 25687 37056 25696
rect 37004 25653 37013 25687
rect 37013 25653 37047 25687
rect 37047 25653 37056 25687
rect 37004 25644 37056 25653
rect 37372 25687 37424 25696
rect 37372 25653 37381 25687
rect 37381 25653 37415 25687
rect 37415 25653 37424 25687
rect 37372 25644 37424 25653
rect 39764 25644 39816 25696
rect 40776 25644 40828 25696
rect 41696 25721 41705 25755
rect 41705 25721 41739 25755
rect 41739 25721 41748 25755
rect 41696 25712 41748 25721
rect 41604 25644 41656 25696
rect 41880 25712 41932 25764
rect 43536 25712 43588 25764
rect 43076 25644 43128 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 4344 25483 4396 25492
rect 4344 25449 4353 25483
rect 4353 25449 4387 25483
rect 4387 25449 4396 25483
rect 4344 25440 4396 25449
rect 6920 25440 6972 25492
rect 7472 25440 7524 25492
rect 8760 25440 8812 25492
rect 10232 25440 10284 25492
rect 11888 25440 11940 25492
rect 17684 25483 17736 25492
rect 17684 25449 17693 25483
rect 17693 25449 17727 25483
rect 17727 25449 17736 25483
rect 17684 25440 17736 25449
rect 18052 25483 18104 25492
rect 18052 25449 18061 25483
rect 18061 25449 18095 25483
rect 18095 25449 18104 25483
rect 18052 25440 18104 25449
rect 21180 25440 21232 25492
rect 24216 25483 24268 25492
rect 24216 25449 24225 25483
rect 24225 25449 24259 25483
rect 24259 25449 24268 25483
rect 24216 25440 24268 25449
rect 27160 25483 27212 25492
rect 27160 25449 27169 25483
rect 27169 25449 27203 25483
rect 27203 25449 27212 25483
rect 27160 25440 27212 25449
rect 3884 25372 3936 25424
rect 2228 25304 2280 25356
rect 2964 25347 3016 25356
rect 2964 25313 2973 25347
rect 2973 25313 3007 25347
rect 3007 25313 3016 25347
rect 2964 25304 3016 25313
rect 6000 25415 6052 25424
rect 5540 25304 5592 25356
rect 6000 25381 6009 25415
rect 6009 25381 6043 25415
rect 6043 25381 6052 25415
rect 6000 25372 6052 25381
rect 6828 25415 6880 25424
rect 6828 25381 6837 25415
rect 6837 25381 6871 25415
rect 6871 25381 6880 25415
rect 6828 25372 6880 25381
rect 8300 25372 8352 25424
rect 10416 25415 10468 25424
rect 10416 25381 10425 25415
rect 10425 25381 10459 25415
rect 10459 25381 10468 25415
rect 10416 25372 10468 25381
rect 12348 25415 12400 25424
rect 12348 25381 12357 25415
rect 12357 25381 12391 25415
rect 12391 25381 12400 25415
rect 12348 25372 12400 25381
rect 12716 25372 12768 25424
rect 6368 25304 6420 25356
rect 7656 25347 7708 25356
rect 7656 25313 7665 25347
rect 7665 25313 7699 25347
rect 7699 25313 7708 25347
rect 7656 25304 7708 25313
rect 9956 25347 10008 25356
rect 2136 25143 2188 25152
rect 2136 25109 2145 25143
rect 2145 25109 2179 25143
rect 2179 25109 2188 25143
rect 2136 25100 2188 25109
rect 3240 25100 3292 25152
rect 6736 25236 6788 25288
rect 9956 25313 9965 25347
rect 9965 25313 9999 25347
rect 9999 25313 10008 25347
rect 9956 25304 10008 25313
rect 11796 25347 11848 25356
rect 11796 25313 11805 25347
rect 11805 25313 11839 25347
rect 11839 25313 11848 25347
rect 11796 25304 11848 25313
rect 11980 25347 12032 25356
rect 11980 25313 11989 25347
rect 11989 25313 12023 25347
rect 12023 25313 12032 25347
rect 11980 25304 12032 25313
rect 13544 25347 13596 25356
rect 13544 25313 13553 25347
rect 13553 25313 13587 25347
rect 13587 25313 13596 25347
rect 13544 25304 13596 25313
rect 14556 25372 14608 25424
rect 19984 25415 20036 25424
rect 19984 25381 19993 25415
rect 19993 25381 20027 25415
rect 20027 25381 20036 25415
rect 19984 25372 20036 25381
rect 24032 25372 24084 25424
rect 24308 25372 24360 25424
rect 24492 25372 24544 25424
rect 14464 25347 14516 25356
rect 14464 25313 14473 25347
rect 14473 25313 14507 25347
rect 14507 25313 14516 25347
rect 14464 25304 14516 25313
rect 14832 25304 14884 25356
rect 15292 25347 15344 25356
rect 15292 25313 15301 25347
rect 15301 25313 15335 25347
rect 15335 25313 15344 25347
rect 15292 25304 15344 25313
rect 16488 25347 16540 25356
rect 16488 25313 16497 25347
rect 16497 25313 16531 25347
rect 16531 25313 16540 25347
rect 16488 25304 16540 25313
rect 17500 25347 17552 25356
rect 17500 25313 17509 25347
rect 17509 25313 17543 25347
rect 17543 25313 17552 25347
rect 17500 25304 17552 25313
rect 19432 25347 19484 25356
rect 19432 25313 19441 25347
rect 19441 25313 19475 25347
rect 19475 25313 19484 25347
rect 19432 25304 19484 25313
rect 20352 25304 20404 25356
rect 23572 25304 23624 25356
rect 30656 25440 30708 25492
rect 32496 25440 32548 25492
rect 36084 25440 36136 25492
rect 38384 25483 38436 25492
rect 38384 25449 38393 25483
rect 38393 25449 38427 25483
rect 38427 25449 38436 25483
rect 38384 25440 38436 25449
rect 41604 25483 41656 25492
rect 41604 25449 41613 25483
rect 41613 25449 41647 25483
rect 41647 25449 41656 25483
rect 41604 25440 41656 25449
rect 41696 25440 41748 25492
rect 43076 25440 43128 25492
rect 44548 25483 44600 25492
rect 44548 25449 44557 25483
rect 44557 25449 44591 25483
rect 44591 25449 44600 25483
rect 44548 25440 44600 25449
rect 27344 25372 27396 25424
rect 27988 25372 28040 25424
rect 29092 25415 29144 25424
rect 29092 25381 29101 25415
rect 29101 25381 29135 25415
rect 29135 25381 29144 25415
rect 29092 25372 29144 25381
rect 29184 25415 29236 25424
rect 29184 25381 29193 25415
rect 29193 25381 29227 25415
rect 29227 25381 29236 25415
rect 33416 25415 33468 25424
rect 29184 25372 29236 25381
rect 33416 25381 33425 25415
rect 33425 25381 33459 25415
rect 33459 25381 33468 25415
rect 33416 25372 33468 25381
rect 35256 25372 35308 25424
rect 36176 25415 36228 25424
rect 36176 25381 36185 25415
rect 36185 25381 36219 25415
rect 36219 25381 36228 25415
rect 36176 25372 36228 25381
rect 37004 25372 37056 25424
rect 39764 25415 39816 25424
rect 39764 25381 39773 25415
rect 39773 25381 39807 25415
rect 39807 25381 39816 25415
rect 39764 25372 39816 25381
rect 40316 25415 40368 25424
rect 40316 25381 40325 25415
rect 40325 25381 40359 25415
rect 40359 25381 40368 25415
rect 40316 25372 40368 25381
rect 30656 25347 30708 25356
rect 30656 25313 30665 25347
rect 30665 25313 30699 25347
rect 30699 25313 30708 25347
rect 30656 25304 30708 25313
rect 31760 25304 31812 25356
rect 32128 25347 32180 25356
rect 32128 25313 32172 25347
rect 32172 25313 32180 25347
rect 32128 25304 32180 25313
rect 38844 25304 38896 25356
rect 17132 25236 17184 25288
rect 20260 25236 20312 25288
rect 22100 25236 22152 25288
rect 25044 25236 25096 25288
rect 32864 25236 32916 25288
rect 33692 25279 33744 25288
rect 33692 25245 33701 25279
rect 33701 25245 33735 25279
rect 33735 25245 33744 25279
rect 33692 25236 33744 25245
rect 34704 25236 34756 25288
rect 35164 25236 35216 25288
rect 39304 25236 39356 25288
rect 13728 25168 13780 25220
rect 21732 25168 21784 25220
rect 23204 25168 23256 25220
rect 24860 25168 24912 25220
rect 24952 25168 25004 25220
rect 29644 25211 29696 25220
rect 29644 25177 29653 25211
rect 29653 25177 29687 25211
rect 29687 25177 29696 25211
rect 29644 25168 29696 25177
rect 31024 25168 31076 25220
rect 4988 25143 5040 25152
rect 4988 25109 4997 25143
rect 4997 25109 5031 25143
rect 5031 25109 5040 25143
rect 4988 25100 5040 25109
rect 8944 25100 8996 25152
rect 14556 25100 14608 25152
rect 21272 25100 21324 25152
rect 28448 25143 28500 25152
rect 28448 25109 28457 25143
rect 28457 25109 28491 25143
rect 28491 25109 28500 25143
rect 28448 25100 28500 25109
rect 31208 25143 31260 25152
rect 31208 25109 31217 25143
rect 31217 25109 31251 25143
rect 31251 25109 31260 25143
rect 31208 25100 31260 25109
rect 31668 25143 31720 25152
rect 31668 25109 31677 25143
rect 31677 25109 31711 25143
rect 31711 25109 31720 25143
rect 31668 25100 31720 25109
rect 32772 25100 32824 25152
rect 35808 25168 35860 25220
rect 36360 25211 36412 25220
rect 36360 25177 36369 25211
rect 36369 25177 36403 25211
rect 36403 25177 36412 25211
rect 41972 25304 42024 25356
rect 42064 25304 42116 25356
rect 43260 25347 43312 25356
rect 43260 25313 43269 25347
rect 43269 25313 43303 25347
rect 43303 25313 43312 25347
rect 43260 25304 43312 25313
rect 44640 25304 44692 25356
rect 42340 25236 42392 25288
rect 36360 25168 36412 25177
rect 34520 25100 34572 25152
rect 36176 25100 36228 25152
rect 39212 25100 39264 25152
rect 41052 25143 41104 25152
rect 41052 25109 41061 25143
rect 41061 25109 41095 25143
rect 41095 25109 41104 25143
rect 41052 25100 41104 25109
rect 41144 25100 41196 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 3884 24939 3936 24948
rect 3884 24905 3893 24939
rect 3893 24905 3927 24939
rect 3927 24905 3936 24939
rect 3884 24896 3936 24905
rect 9956 24896 10008 24948
rect 12256 24896 12308 24948
rect 13544 24896 13596 24948
rect 17868 24896 17920 24948
rect 19432 24896 19484 24948
rect 21180 24896 21232 24948
rect 22100 24939 22152 24948
rect 22100 24905 22109 24939
rect 22109 24905 22143 24939
rect 22143 24905 22152 24939
rect 22100 24896 22152 24905
rect 23020 24939 23072 24948
rect 23020 24905 23029 24939
rect 23029 24905 23063 24939
rect 23063 24905 23072 24939
rect 23020 24896 23072 24905
rect 23572 24896 23624 24948
rect 24492 24896 24544 24948
rect 25044 24939 25096 24948
rect 25044 24905 25053 24939
rect 25053 24905 25087 24939
rect 25087 24905 25096 24939
rect 25044 24896 25096 24905
rect 112 24828 164 24880
rect 6368 24828 6420 24880
rect 11796 24828 11848 24880
rect 17500 24871 17552 24880
rect 17500 24837 17509 24871
rect 17509 24837 17543 24871
rect 17543 24837 17552 24871
rect 17500 24828 17552 24837
rect 2228 24760 2280 24812
rect 4988 24760 5040 24812
rect 3608 24692 3660 24744
rect 3792 24692 3844 24744
rect 2412 24667 2464 24676
rect 2412 24633 2421 24667
rect 2421 24633 2455 24667
rect 2455 24633 2464 24667
rect 2412 24624 2464 24633
rect 4160 24692 4212 24744
rect 5264 24692 5316 24744
rect 4528 24624 4580 24676
rect 8208 24760 8260 24812
rect 7472 24735 7524 24744
rect 7472 24701 7481 24735
rect 7481 24701 7515 24735
rect 7515 24701 7524 24735
rect 7472 24692 7524 24701
rect 7932 24692 7984 24744
rect 13636 24760 13688 24812
rect 20260 24803 20312 24812
rect 8944 24735 8996 24744
rect 8576 24624 8628 24676
rect 5540 24599 5592 24608
rect 5540 24565 5549 24599
rect 5549 24565 5583 24599
rect 5583 24565 5592 24599
rect 5540 24556 5592 24565
rect 5908 24599 5960 24608
rect 5908 24565 5917 24599
rect 5917 24565 5951 24599
rect 5951 24565 5960 24599
rect 5908 24556 5960 24565
rect 6644 24599 6696 24608
rect 6644 24565 6653 24599
rect 6653 24565 6687 24599
rect 6687 24565 6696 24599
rect 6644 24556 6696 24565
rect 8116 24556 8168 24608
rect 8944 24701 8953 24735
rect 8953 24701 8987 24735
rect 8987 24701 8996 24735
rect 8944 24692 8996 24701
rect 8760 24624 8812 24676
rect 11980 24692 12032 24744
rect 12440 24692 12492 24744
rect 14464 24735 14516 24744
rect 14464 24701 14473 24735
rect 14473 24701 14507 24735
rect 14507 24701 14516 24735
rect 14464 24692 14516 24701
rect 14648 24735 14700 24744
rect 14648 24701 14657 24735
rect 14657 24701 14691 24735
rect 14691 24701 14700 24735
rect 14648 24692 14700 24701
rect 14924 24735 14976 24744
rect 14924 24701 14933 24735
rect 14933 24701 14967 24735
rect 14967 24701 14976 24735
rect 14924 24692 14976 24701
rect 12072 24624 12124 24676
rect 17132 24692 17184 24744
rect 17776 24692 17828 24744
rect 19800 24735 19852 24744
rect 19800 24701 19809 24735
rect 19809 24701 19843 24735
rect 19843 24701 19852 24735
rect 19800 24692 19852 24701
rect 20260 24769 20269 24803
rect 20269 24769 20303 24803
rect 20303 24769 20312 24803
rect 20260 24760 20312 24769
rect 21272 24760 21324 24812
rect 22284 24760 22336 24812
rect 24308 24871 24360 24880
rect 24308 24837 24317 24871
rect 24317 24837 24351 24871
rect 24351 24837 24360 24871
rect 24308 24828 24360 24837
rect 24860 24828 24912 24880
rect 20352 24692 20404 24744
rect 28540 24896 28592 24948
rect 29092 24939 29144 24948
rect 29092 24905 29101 24939
rect 29101 24905 29135 24939
rect 29135 24905 29144 24939
rect 29092 24896 29144 24905
rect 27344 24871 27396 24880
rect 27344 24837 27353 24871
rect 27353 24837 27387 24871
rect 27387 24837 27396 24871
rect 27344 24828 27396 24837
rect 29184 24828 29236 24880
rect 33416 24896 33468 24948
rect 35900 24939 35952 24948
rect 35900 24905 35909 24939
rect 35909 24905 35943 24939
rect 35943 24905 35952 24939
rect 35900 24896 35952 24905
rect 39304 24939 39356 24948
rect 39304 24905 39313 24939
rect 39313 24905 39347 24939
rect 39347 24905 39356 24939
rect 39304 24896 39356 24905
rect 39764 24896 39816 24948
rect 41972 24939 42024 24948
rect 41972 24905 41981 24939
rect 41981 24905 42015 24939
rect 42015 24905 42024 24939
rect 41972 24896 42024 24905
rect 43260 24896 43312 24948
rect 34336 24828 34388 24880
rect 36360 24828 36412 24880
rect 38752 24828 38804 24880
rect 43996 24828 44048 24880
rect 28448 24760 28500 24812
rect 29644 24803 29696 24812
rect 26056 24692 26108 24744
rect 29644 24769 29653 24803
rect 29653 24769 29687 24803
rect 29687 24769 29696 24803
rect 29644 24760 29696 24769
rect 31668 24760 31720 24812
rect 32128 24803 32180 24812
rect 32128 24769 32137 24803
rect 32137 24769 32171 24803
rect 32171 24769 32180 24803
rect 32128 24760 32180 24769
rect 32496 24803 32548 24812
rect 32496 24769 32505 24803
rect 32505 24769 32539 24803
rect 32539 24769 32548 24803
rect 32496 24760 32548 24769
rect 33140 24803 33192 24812
rect 33140 24769 33149 24803
rect 33149 24769 33183 24803
rect 33183 24769 33192 24803
rect 33140 24760 33192 24769
rect 34428 24760 34480 24812
rect 36820 24803 36872 24812
rect 36820 24769 36829 24803
rect 36829 24769 36863 24803
rect 36863 24769 36872 24803
rect 36820 24760 36872 24769
rect 39948 24760 40000 24812
rect 16488 24624 16540 24676
rect 17684 24624 17736 24676
rect 21180 24667 21232 24676
rect 21180 24633 21189 24667
rect 21189 24633 21223 24667
rect 21223 24633 21232 24667
rect 21180 24624 21232 24633
rect 21272 24667 21324 24676
rect 21272 24633 21281 24667
rect 21281 24633 21315 24667
rect 21315 24633 21324 24667
rect 23848 24667 23900 24676
rect 21272 24624 21324 24633
rect 23848 24633 23857 24667
rect 23857 24633 23891 24667
rect 23891 24633 23900 24667
rect 23848 24624 23900 24633
rect 31576 24735 31628 24744
rect 31576 24701 31585 24735
rect 31585 24701 31619 24735
rect 31619 24701 31628 24735
rect 38016 24735 38068 24744
rect 31576 24692 31628 24701
rect 38016 24701 38025 24735
rect 38025 24701 38059 24735
rect 38059 24701 38068 24735
rect 38016 24692 38068 24701
rect 10692 24599 10744 24608
rect 10692 24565 10701 24599
rect 10701 24565 10735 24599
rect 10735 24565 10744 24599
rect 10692 24556 10744 24565
rect 11244 24599 11296 24608
rect 11244 24565 11253 24599
rect 11253 24565 11287 24599
rect 11287 24565 11296 24599
rect 11244 24556 11296 24565
rect 14188 24556 14240 24608
rect 15292 24556 15344 24608
rect 17408 24556 17460 24608
rect 22928 24556 22980 24608
rect 26608 24556 26660 24608
rect 27712 24624 27764 24676
rect 29368 24667 29420 24676
rect 29368 24633 29377 24667
rect 29377 24633 29411 24667
rect 29411 24633 29420 24667
rect 29368 24624 29420 24633
rect 29092 24556 29144 24608
rect 31300 24624 31352 24676
rect 32588 24667 32640 24676
rect 32588 24633 32597 24667
rect 32597 24633 32631 24667
rect 32631 24633 32640 24667
rect 32588 24624 32640 24633
rect 30564 24556 30616 24608
rect 30656 24556 30708 24608
rect 31392 24556 31444 24608
rect 32128 24556 32180 24608
rect 34152 24624 34204 24676
rect 34520 24624 34572 24676
rect 35256 24624 35308 24676
rect 36912 24624 36964 24676
rect 37648 24624 37700 24676
rect 40408 24692 40460 24744
rect 42708 24692 42760 24744
rect 41052 24667 41104 24676
rect 41052 24633 41061 24667
rect 41061 24633 41095 24667
rect 41095 24633 41104 24667
rect 41052 24624 41104 24633
rect 37556 24599 37608 24608
rect 37556 24565 37565 24599
rect 37565 24565 37599 24599
rect 37599 24565 37608 24599
rect 37556 24556 37608 24565
rect 38844 24599 38896 24608
rect 38844 24565 38853 24599
rect 38853 24565 38887 24599
rect 38887 24565 38896 24599
rect 38844 24556 38896 24565
rect 39764 24556 39816 24608
rect 41788 24624 41840 24676
rect 41328 24556 41380 24608
rect 41420 24556 41472 24608
rect 44272 24667 44324 24676
rect 44272 24633 44281 24667
rect 44281 24633 44315 24667
rect 44315 24633 44324 24667
rect 44272 24624 44324 24633
rect 43168 24556 43220 24608
rect 43536 24556 43588 24608
rect 44640 24599 44692 24608
rect 44640 24565 44649 24599
rect 44649 24565 44683 24599
rect 44683 24565 44692 24599
rect 44640 24556 44692 24565
rect 44732 24556 44784 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 2228 24395 2280 24404
rect 2228 24361 2237 24395
rect 2237 24361 2271 24395
rect 2271 24361 2280 24395
rect 2228 24352 2280 24361
rect 2964 24352 3016 24404
rect 3424 24352 3476 24404
rect 3700 24352 3752 24404
rect 6644 24352 6696 24404
rect 9956 24352 10008 24404
rect 1492 24216 1544 24268
rect 3976 24284 4028 24336
rect 6368 24327 6420 24336
rect 6368 24293 6377 24327
rect 6377 24293 6411 24327
rect 6411 24293 6420 24327
rect 6368 24284 6420 24293
rect 6736 24327 6788 24336
rect 6736 24293 6745 24327
rect 6745 24293 6779 24327
rect 6779 24293 6788 24327
rect 6736 24284 6788 24293
rect 2136 24216 2188 24268
rect 2964 24259 3016 24268
rect 2964 24225 2973 24259
rect 2973 24225 3007 24259
rect 3007 24225 3016 24259
rect 2964 24216 3016 24225
rect 2504 24080 2556 24132
rect 4160 24148 4212 24200
rect 4620 24148 4672 24200
rect 4068 24012 4120 24064
rect 4528 24080 4580 24132
rect 5816 24216 5868 24268
rect 6000 24216 6052 24268
rect 7196 24259 7248 24268
rect 7196 24225 7205 24259
rect 7205 24225 7239 24259
rect 7239 24225 7248 24259
rect 7196 24216 7248 24225
rect 7380 24259 7432 24268
rect 7380 24225 7389 24259
rect 7389 24225 7423 24259
rect 7423 24225 7432 24259
rect 7380 24216 7432 24225
rect 8576 24259 8628 24268
rect 8576 24225 8585 24259
rect 8585 24225 8619 24259
rect 8619 24225 8628 24259
rect 8576 24216 8628 24225
rect 10692 24352 10744 24404
rect 11152 24395 11204 24404
rect 11152 24361 11161 24395
rect 11161 24361 11195 24395
rect 11195 24361 11204 24395
rect 11152 24352 11204 24361
rect 12532 24395 12584 24404
rect 12532 24361 12541 24395
rect 12541 24361 12575 24395
rect 12575 24361 12584 24395
rect 12532 24352 12584 24361
rect 14556 24395 14608 24404
rect 11244 24284 11296 24336
rect 13636 24327 13688 24336
rect 13636 24293 13645 24327
rect 13645 24293 13679 24327
rect 13679 24293 13688 24327
rect 14188 24327 14240 24336
rect 13636 24284 13688 24293
rect 14188 24293 14197 24327
rect 14197 24293 14231 24327
rect 14231 24293 14240 24327
rect 14188 24284 14240 24293
rect 14556 24361 14565 24395
rect 14565 24361 14599 24395
rect 14599 24361 14608 24395
rect 14556 24352 14608 24361
rect 15660 24327 15712 24336
rect 15660 24293 15663 24327
rect 15663 24293 15697 24327
rect 15697 24293 15712 24327
rect 15660 24284 15712 24293
rect 17132 24284 17184 24336
rect 18788 24284 18840 24336
rect 11060 24259 11112 24268
rect 11060 24225 11069 24259
rect 11069 24225 11103 24259
rect 11103 24225 11112 24259
rect 11060 24216 11112 24225
rect 12440 24259 12492 24268
rect 10140 24148 10192 24200
rect 12440 24225 12449 24259
rect 12449 24225 12483 24259
rect 12483 24225 12492 24259
rect 12440 24216 12492 24225
rect 13820 24259 13872 24268
rect 13820 24225 13829 24259
rect 13829 24225 13863 24259
rect 13863 24225 13872 24259
rect 13820 24216 13872 24225
rect 12348 24148 12400 24200
rect 17776 24216 17828 24268
rect 17960 24259 18012 24268
rect 17960 24225 17969 24259
rect 17969 24225 18003 24259
rect 18003 24225 18012 24259
rect 17960 24216 18012 24225
rect 20076 24352 20128 24404
rect 20352 24352 20404 24404
rect 24124 24352 24176 24404
rect 27712 24395 27764 24404
rect 19892 24284 19944 24336
rect 21088 24284 21140 24336
rect 22836 24327 22888 24336
rect 22836 24293 22845 24327
rect 22845 24293 22879 24327
rect 22879 24293 22888 24327
rect 22836 24284 22888 24293
rect 23848 24284 23900 24336
rect 19064 24216 19116 24268
rect 15292 24191 15344 24200
rect 15292 24157 15301 24191
rect 15301 24157 15335 24191
rect 15335 24157 15344 24191
rect 15292 24148 15344 24157
rect 17316 24191 17368 24200
rect 17316 24157 17325 24191
rect 17325 24157 17359 24191
rect 17359 24157 17368 24191
rect 17316 24148 17368 24157
rect 20904 24148 20956 24200
rect 21916 24148 21968 24200
rect 22928 24148 22980 24200
rect 27712 24361 27721 24395
rect 27721 24361 27755 24395
rect 27755 24361 27764 24395
rect 28908 24395 28960 24404
rect 27712 24352 27764 24361
rect 28908 24361 28917 24395
rect 28917 24361 28951 24395
rect 28951 24361 28960 24395
rect 28908 24352 28960 24361
rect 29368 24352 29420 24404
rect 34520 24352 34572 24404
rect 34704 24395 34756 24404
rect 34704 24361 34713 24395
rect 34713 24361 34747 24395
rect 34747 24361 34756 24395
rect 34704 24352 34756 24361
rect 42064 24352 42116 24404
rect 43996 24352 44048 24404
rect 24768 24327 24820 24336
rect 24768 24293 24777 24327
rect 24777 24293 24811 24327
rect 24811 24293 24820 24327
rect 24768 24284 24820 24293
rect 27344 24284 27396 24336
rect 30564 24284 30616 24336
rect 32404 24284 32456 24336
rect 33416 24284 33468 24336
rect 34612 24284 34664 24336
rect 36912 24284 36964 24336
rect 37372 24284 37424 24336
rect 39304 24284 39356 24336
rect 26516 24259 26568 24268
rect 26516 24225 26525 24259
rect 26525 24225 26559 24259
rect 26559 24225 26568 24259
rect 26516 24216 26568 24225
rect 5724 24123 5776 24132
rect 5724 24089 5733 24123
rect 5733 24089 5767 24123
rect 5767 24089 5776 24123
rect 5724 24080 5776 24089
rect 7564 24080 7616 24132
rect 10692 24080 10744 24132
rect 13728 24080 13780 24132
rect 14648 24080 14700 24132
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 27988 24191 28040 24200
rect 27988 24157 27997 24191
rect 27997 24157 28031 24191
rect 28031 24157 28040 24191
rect 27988 24148 28040 24157
rect 30564 24191 30616 24200
rect 30564 24157 30573 24191
rect 30573 24157 30607 24191
rect 30607 24157 30616 24191
rect 30564 24148 30616 24157
rect 30748 24148 30800 24200
rect 31300 24148 31352 24200
rect 32588 24148 32640 24200
rect 34244 24216 34296 24268
rect 35808 24216 35860 24268
rect 36360 24259 36412 24268
rect 36360 24225 36404 24259
rect 36404 24225 36412 24259
rect 36360 24216 36412 24225
rect 37648 24216 37700 24268
rect 41328 24284 41380 24336
rect 43628 24284 43680 24336
rect 44916 24259 44968 24268
rect 44916 24225 44925 24259
rect 44925 24225 44959 24259
rect 44959 24225 44968 24259
rect 44916 24216 44968 24225
rect 31576 24080 31628 24132
rect 32680 24080 32732 24132
rect 39120 24148 39172 24200
rect 39764 24148 39816 24200
rect 41512 24148 41564 24200
rect 43260 24148 43312 24200
rect 43444 24191 43496 24200
rect 43444 24157 43453 24191
rect 43453 24157 43487 24191
rect 43487 24157 43496 24191
rect 43444 24148 43496 24157
rect 35256 24080 35308 24132
rect 35440 24123 35492 24132
rect 35440 24089 35449 24123
rect 35449 24089 35483 24123
rect 35483 24089 35492 24123
rect 35440 24080 35492 24089
rect 37648 24080 37700 24132
rect 38108 24080 38160 24132
rect 41880 24080 41932 24132
rect 43812 24148 43864 24200
rect 5080 24055 5132 24064
rect 5080 24021 5089 24055
rect 5089 24021 5123 24055
rect 5123 24021 5132 24055
rect 5080 24012 5132 24021
rect 7656 24012 7708 24064
rect 8760 24055 8812 24064
rect 8760 24021 8769 24055
rect 8769 24021 8803 24055
rect 8803 24021 8812 24055
rect 8760 24012 8812 24021
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 14464 24012 14516 24064
rect 16212 24055 16264 24064
rect 16212 24021 16221 24055
rect 16221 24021 16255 24055
rect 16255 24021 16264 24055
rect 16212 24012 16264 24021
rect 23848 24055 23900 24064
rect 23848 24021 23857 24055
rect 23857 24021 23891 24055
rect 23891 24021 23900 24055
rect 23848 24012 23900 24021
rect 26700 24055 26752 24064
rect 26700 24021 26709 24055
rect 26709 24021 26743 24055
rect 26743 24021 26752 24055
rect 26700 24012 26752 24021
rect 27068 24055 27120 24064
rect 27068 24021 27077 24055
rect 27077 24021 27111 24055
rect 27111 24021 27120 24055
rect 27068 24012 27120 24021
rect 29092 24012 29144 24064
rect 31484 24055 31536 24064
rect 31484 24021 31493 24055
rect 31493 24021 31527 24055
rect 31527 24021 31536 24055
rect 31484 24012 31536 24021
rect 36636 24012 36688 24064
rect 36912 24055 36964 24064
rect 36912 24021 36921 24055
rect 36921 24021 36955 24055
rect 36955 24021 36964 24055
rect 38200 24055 38252 24064
rect 36912 24012 36964 24021
rect 38200 24021 38209 24055
rect 38209 24021 38243 24055
rect 38243 24021 38252 24055
rect 38200 24012 38252 24021
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 2412 23851 2464 23860
rect 2412 23817 2421 23851
rect 2421 23817 2455 23851
rect 2455 23817 2464 23851
rect 2412 23808 2464 23817
rect 3424 23851 3476 23860
rect 3424 23817 3433 23851
rect 3433 23817 3467 23851
rect 3467 23817 3476 23851
rect 3424 23808 3476 23817
rect 3976 23808 4028 23860
rect 8116 23808 8168 23860
rect 8576 23851 8628 23860
rect 8576 23817 8585 23851
rect 8585 23817 8619 23851
rect 8619 23817 8628 23851
rect 8576 23808 8628 23817
rect 11060 23808 11112 23860
rect 12440 23808 12492 23860
rect 13820 23808 13872 23860
rect 14740 23851 14792 23860
rect 14740 23817 14749 23851
rect 14749 23817 14783 23851
rect 14783 23817 14792 23851
rect 14740 23808 14792 23817
rect 15292 23808 15344 23860
rect 17408 23808 17460 23860
rect 3148 23740 3200 23792
rect 4068 23740 4120 23792
rect 5172 23740 5224 23792
rect 5724 23740 5776 23792
rect 4620 23672 4672 23724
rect 5632 23672 5684 23724
rect 7748 23715 7800 23724
rect 7748 23681 7754 23715
rect 7754 23681 7800 23715
rect 7748 23672 7800 23681
rect 7840 23672 7892 23724
rect 8944 23715 8996 23724
rect 8944 23681 8953 23715
rect 8953 23681 8987 23715
rect 8987 23681 8996 23715
rect 8944 23672 8996 23681
rect 2964 23647 3016 23656
rect 2964 23613 2973 23647
rect 2973 23613 3007 23647
rect 3007 23613 3016 23647
rect 2964 23604 3016 23613
rect 5080 23604 5132 23656
rect 5264 23647 5316 23656
rect 5264 23613 5273 23647
rect 5273 23613 5307 23647
rect 5307 23613 5316 23647
rect 5264 23604 5316 23613
rect 5540 23604 5592 23656
rect 6644 23604 6696 23656
rect 6736 23604 6788 23656
rect 7564 23647 7616 23656
rect 7564 23613 7573 23647
rect 7573 23613 7607 23647
rect 7607 23613 7616 23647
rect 7564 23604 7616 23613
rect 8392 23604 8444 23656
rect 9128 23647 9180 23656
rect 9128 23613 9137 23647
rect 9137 23613 9171 23647
rect 9171 23613 9180 23647
rect 9128 23604 9180 23613
rect 9220 23647 9272 23656
rect 9220 23613 9229 23647
rect 9229 23613 9263 23647
rect 9263 23613 9272 23647
rect 10140 23672 10192 23724
rect 14924 23672 14976 23724
rect 9220 23604 9272 23613
rect 9496 23604 9548 23656
rect 10784 23604 10836 23656
rect 11244 23647 11296 23656
rect 11244 23613 11253 23647
rect 11253 23613 11287 23647
rect 11287 23613 11296 23647
rect 11244 23604 11296 23613
rect 3332 23536 3384 23588
rect 4252 23536 4304 23588
rect 7104 23536 7156 23588
rect 8300 23579 8352 23588
rect 8300 23545 8309 23579
rect 8309 23545 8343 23579
rect 8343 23545 8352 23579
rect 8300 23536 8352 23545
rect 13728 23604 13780 23656
rect 17960 23808 18012 23860
rect 22836 23808 22888 23860
rect 19064 23783 19116 23792
rect 19064 23749 19073 23783
rect 19073 23749 19107 23783
rect 19107 23749 19116 23783
rect 19064 23740 19116 23749
rect 25136 23783 25188 23792
rect 25136 23749 25145 23783
rect 25145 23749 25179 23783
rect 25179 23749 25188 23783
rect 25136 23740 25188 23749
rect 21180 23715 21232 23724
rect 21180 23681 21189 23715
rect 21189 23681 21223 23715
rect 21223 23681 21232 23715
rect 21180 23672 21232 23681
rect 27804 23808 27856 23860
rect 27988 23808 28040 23860
rect 28356 23851 28408 23860
rect 28356 23817 28365 23851
rect 28365 23817 28399 23851
rect 28399 23817 28408 23851
rect 28356 23808 28408 23817
rect 28908 23808 28960 23860
rect 31208 23808 31260 23860
rect 31392 23808 31444 23860
rect 34244 23851 34296 23860
rect 26516 23783 26568 23792
rect 26516 23749 26525 23783
rect 26525 23749 26559 23783
rect 26559 23749 26568 23783
rect 26516 23740 26568 23749
rect 27344 23740 27396 23792
rect 18788 23604 18840 23656
rect 20168 23604 20220 23656
rect 23112 23604 23164 23656
rect 30564 23740 30616 23792
rect 32404 23740 32456 23792
rect 34244 23817 34253 23851
rect 34253 23817 34287 23851
rect 34287 23817 34296 23851
rect 34244 23808 34296 23817
rect 34612 23851 34664 23860
rect 34612 23817 34621 23851
rect 34621 23817 34655 23851
rect 34655 23817 34664 23851
rect 34612 23808 34664 23817
rect 36360 23851 36412 23860
rect 36360 23817 36369 23851
rect 36369 23817 36403 23851
rect 36403 23817 36412 23851
rect 36360 23808 36412 23817
rect 37648 23808 37700 23860
rect 41420 23808 41472 23860
rect 41512 23808 41564 23860
rect 42064 23808 42116 23860
rect 42524 23808 42576 23860
rect 27988 23715 28040 23724
rect 27988 23681 27997 23715
rect 27997 23681 28031 23715
rect 28031 23681 28040 23715
rect 27988 23672 28040 23681
rect 31484 23672 31536 23724
rect 31576 23715 31628 23724
rect 31576 23681 31585 23715
rect 31585 23681 31619 23715
rect 31619 23681 31628 23715
rect 37464 23740 37516 23792
rect 31576 23672 31628 23681
rect 34612 23672 34664 23724
rect 35440 23715 35492 23724
rect 35440 23681 35449 23715
rect 35449 23681 35483 23715
rect 35483 23681 35492 23715
rect 35440 23672 35492 23681
rect 36636 23672 36688 23724
rect 38108 23715 38160 23724
rect 38108 23681 38117 23715
rect 38117 23681 38151 23715
rect 38151 23681 38160 23715
rect 38108 23672 38160 23681
rect 43444 23740 43496 23792
rect 38568 23672 38620 23724
rect 39120 23672 39172 23724
rect 41144 23672 41196 23724
rect 43168 23715 43220 23724
rect 43168 23681 43177 23715
rect 43177 23681 43211 23715
rect 43211 23681 43220 23715
rect 43168 23672 43220 23681
rect 43260 23672 43312 23724
rect 27068 23604 27120 23656
rect 27344 23604 27396 23656
rect 28816 23604 28868 23656
rect 30840 23604 30892 23656
rect 44916 23808 44968 23860
rect 45468 23851 45520 23860
rect 45468 23817 45477 23851
rect 45477 23817 45511 23851
rect 45511 23817 45520 23851
rect 45468 23808 45520 23817
rect 1492 23468 1544 23520
rect 2320 23468 2372 23520
rect 4896 23468 4948 23520
rect 5080 23468 5132 23520
rect 5908 23468 5960 23520
rect 6000 23511 6052 23520
rect 6000 23477 6009 23511
rect 6009 23477 6043 23511
rect 6043 23477 6052 23511
rect 6644 23511 6696 23520
rect 6000 23468 6052 23477
rect 6644 23477 6653 23511
rect 6653 23477 6687 23511
rect 6687 23477 6696 23511
rect 6644 23468 6696 23477
rect 10232 23468 10284 23520
rect 13820 23536 13872 23588
rect 14556 23536 14608 23588
rect 14740 23536 14792 23588
rect 15660 23536 15712 23588
rect 18236 23536 18288 23588
rect 20720 23579 20772 23588
rect 20720 23545 20729 23579
rect 20729 23545 20763 23579
rect 20763 23545 20772 23579
rect 20720 23536 20772 23545
rect 17408 23468 17460 23520
rect 17960 23468 18012 23520
rect 18604 23468 18656 23520
rect 21088 23468 21140 23520
rect 22836 23468 22888 23520
rect 23848 23468 23900 23520
rect 24768 23536 24820 23588
rect 27436 23579 27488 23588
rect 27436 23545 27445 23579
rect 27445 23545 27479 23579
rect 27479 23545 27488 23579
rect 27436 23536 27488 23545
rect 33324 23579 33376 23588
rect 33324 23545 33333 23579
rect 33333 23545 33367 23579
rect 33367 23545 33376 23579
rect 33324 23536 33376 23545
rect 33416 23579 33468 23588
rect 33416 23545 33425 23579
rect 33425 23545 33459 23579
rect 33459 23545 33468 23579
rect 33416 23536 33468 23545
rect 34152 23536 34204 23588
rect 34796 23536 34848 23588
rect 29736 23511 29788 23520
rect 29736 23477 29745 23511
rect 29745 23477 29779 23511
rect 29779 23477 29788 23511
rect 29736 23468 29788 23477
rect 30840 23468 30892 23520
rect 34336 23468 34388 23520
rect 34704 23468 34756 23520
rect 36268 23468 36320 23520
rect 37464 23536 37516 23588
rect 38200 23579 38252 23588
rect 38200 23545 38209 23579
rect 38209 23545 38243 23579
rect 38243 23545 38252 23579
rect 38200 23536 38252 23545
rect 39672 23536 39724 23588
rect 40408 23536 40460 23588
rect 41328 23536 41380 23588
rect 41696 23579 41748 23588
rect 41696 23545 41705 23579
rect 41705 23545 41739 23579
rect 41739 23545 41748 23579
rect 41696 23536 41748 23545
rect 39304 23511 39356 23520
rect 39304 23477 39313 23511
rect 39313 23477 39347 23511
rect 39347 23477 39356 23511
rect 39304 23468 39356 23477
rect 42892 23511 42944 23520
rect 42892 23477 42901 23511
rect 42901 23477 42935 23511
rect 42935 23477 42944 23511
rect 43628 23536 43680 23588
rect 42892 23468 42944 23477
rect 44180 23468 44232 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 2504 23307 2556 23316
rect 2504 23273 2513 23307
rect 2513 23273 2547 23307
rect 2547 23273 2556 23307
rect 2504 23264 2556 23273
rect 2872 23264 2924 23316
rect 5172 23264 5224 23316
rect 5816 23264 5868 23316
rect 7840 23264 7892 23316
rect 8208 23264 8260 23316
rect 9220 23307 9272 23316
rect 9220 23273 9229 23307
rect 9229 23273 9263 23307
rect 9263 23273 9272 23307
rect 9220 23264 9272 23273
rect 10692 23307 10744 23316
rect 3976 23196 4028 23248
rect 4252 23239 4304 23248
rect 4252 23205 4261 23239
rect 4261 23205 4295 23239
rect 4295 23205 4304 23239
rect 4252 23196 4304 23205
rect 5264 23196 5316 23248
rect 2320 23171 2372 23180
rect 2320 23137 2329 23171
rect 2329 23137 2363 23171
rect 2363 23137 2372 23171
rect 2320 23128 2372 23137
rect 2412 23128 2464 23180
rect 4712 23128 4764 23180
rect 5540 23128 5592 23180
rect 6644 23196 6696 23248
rect 7380 23196 7432 23248
rect 9496 23196 9548 23248
rect 10692 23273 10701 23307
rect 10701 23273 10735 23307
rect 10735 23273 10744 23307
rect 10692 23264 10744 23273
rect 12348 23307 12400 23316
rect 12348 23273 12357 23307
rect 12357 23273 12391 23307
rect 12391 23273 12400 23307
rect 12348 23264 12400 23273
rect 13636 23264 13688 23316
rect 14924 23264 14976 23316
rect 20720 23307 20772 23316
rect 20720 23273 20729 23307
rect 20729 23273 20763 23307
rect 20763 23273 20772 23307
rect 20720 23264 20772 23273
rect 27988 23264 28040 23316
rect 29092 23264 29144 23316
rect 31300 23307 31352 23316
rect 31300 23273 31309 23307
rect 31309 23273 31343 23307
rect 31343 23273 31352 23307
rect 31300 23264 31352 23273
rect 32496 23307 32548 23316
rect 32496 23273 32505 23307
rect 32505 23273 32539 23307
rect 32539 23273 32548 23307
rect 32496 23264 32548 23273
rect 33416 23264 33468 23316
rect 35256 23307 35308 23316
rect 35256 23273 35265 23307
rect 35265 23273 35299 23307
rect 35299 23273 35308 23307
rect 35256 23264 35308 23273
rect 36636 23264 36688 23316
rect 43168 23307 43220 23316
rect 43168 23273 43177 23307
rect 43177 23273 43211 23307
rect 43211 23273 43220 23307
rect 43168 23264 43220 23273
rect 43352 23264 43404 23316
rect 6736 23171 6788 23180
rect 6736 23137 6745 23171
rect 6745 23137 6779 23171
rect 6779 23137 6788 23171
rect 6736 23128 6788 23137
rect 7104 23128 7156 23180
rect 7288 23128 7340 23180
rect 8208 23171 8260 23180
rect 8208 23137 8217 23171
rect 8217 23137 8251 23171
rect 8251 23137 8260 23171
rect 8208 23128 8260 23137
rect 8392 23171 8444 23180
rect 8392 23137 8401 23171
rect 8401 23137 8435 23171
rect 8435 23137 8444 23171
rect 8392 23128 8444 23137
rect 9220 23128 9272 23180
rect 9680 23171 9732 23180
rect 9680 23137 9689 23171
rect 9689 23137 9723 23171
rect 9723 23137 9732 23171
rect 9680 23128 9732 23137
rect 11152 23196 11204 23248
rect 11060 23171 11112 23180
rect 11060 23137 11069 23171
rect 11069 23137 11103 23171
rect 11103 23137 11112 23171
rect 11060 23128 11112 23137
rect 15108 23196 15160 23248
rect 17316 23196 17368 23248
rect 18604 23239 18656 23248
rect 18604 23205 18613 23239
rect 18613 23205 18647 23239
rect 18647 23205 18656 23239
rect 18604 23196 18656 23205
rect 20812 23196 20864 23248
rect 23296 23196 23348 23248
rect 23848 23196 23900 23248
rect 24768 23196 24820 23248
rect 28448 23196 28500 23248
rect 31484 23196 31536 23248
rect 33508 23196 33560 23248
rect 34704 23196 34756 23248
rect 36268 23239 36320 23248
rect 36268 23205 36277 23239
rect 36277 23205 36311 23239
rect 36311 23205 36320 23239
rect 36268 23196 36320 23205
rect 38568 23239 38620 23248
rect 38568 23205 38577 23239
rect 38577 23205 38611 23239
rect 38611 23205 38620 23239
rect 38568 23196 38620 23205
rect 39304 23196 39356 23248
rect 41328 23239 41380 23248
rect 41328 23205 41337 23239
rect 41337 23205 41371 23239
rect 41371 23205 41380 23239
rect 41328 23196 41380 23205
rect 41880 23239 41932 23248
rect 41880 23205 41889 23239
rect 41889 23205 41923 23239
rect 41923 23205 41932 23239
rect 41880 23196 41932 23205
rect 43628 23196 43680 23248
rect 13176 23128 13228 23180
rect 13452 23171 13504 23180
rect 13452 23137 13461 23171
rect 13461 23137 13495 23171
rect 13495 23137 13504 23171
rect 13452 23128 13504 23137
rect 13636 23171 13688 23180
rect 13636 23137 13645 23171
rect 13645 23137 13679 23171
rect 13679 23137 13688 23171
rect 13636 23128 13688 23137
rect 16212 23128 16264 23180
rect 21272 23128 21324 23180
rect 22100 23128 22152 23180
rect 26608 23128 26660 23180
rect 27068 23128 27120 23180
rect 27436 23128 27488 23180
rect 28172 23128 28224 23180
rect 29736 23171 29788 23180
rect 29736 23137 29745 23171
rect 29745 23137 29779 23171
rect 29779 23137 29788 23171
rect 29736 23128 29788 23137
rect 30288 23128 30340 23180
rect 38292 23171 38344 23180
rect 4988 23060 5040 23112
rect 6000 23103 6052 23112
rect 6000 23069 6009 23103
rect 6009 23069 6043 23103
rect 6043 23069 6052 23103
rect 6000 23060 6052 23069
rect 5172 23035 5224 23044
rect 5172 23001 5181 23035
rect 5181 23001 5215 23035
rect 5215 23001 5224 23035
rect 5172 22992 5224 23001
rect 2872 22924 2924 22976
rect 3148 22924 3200 22976
rect 3332 22967 3384 22976
rect 3332 22933 3341 22967
rect 3341 22933 3375 22967
rect 3375 22933 3384 22967
rect 3332 22924 3384 22933
rect 3792 22967 3844 22976
rect 3792 22933 3801 22967
rect 3801 22933 3835 22967
rect 3835 22933 3844 22967
rect 3792 22924 3844 22933
rect 4068 22924 4120 22976
rect 5632 22924 5684 22976
rect 5908 22967 5960 22976
rect 5908 22933 5917 22967
rect 5917 22933 5951 22967
rect 5951 22933 5960 22967
rect 5908 22924 5960 22933
rect 6828 22924 6880 22976
rect 12072 23060 12124 23112
rect 13912 23103 13964 23112
rect 13912 23069 13921 23103
rect 13921 23069 13955 23103
rect 13955 23069 13964 23103
rect 13912 23060 13964 23069
rect 7196 22992 7248 23044
rect 9864 22992 9916 23044
rect 16764 22992 16816 23044
rect 18236 23060 18288 23112
rect 18788 23060 18840 23112
rect 23020 23103 23072 23112
rect 23020 23069 23029 23103
rect 23029 23069 23063 23103
rect 23063 23069 23072 23103
rect 23020 23060 23072 23069
rect 24584 23103 24636 23112
rect 17868 22992 17920 23044
rect 21916 22992 21968 23044
rect 24584 23069 24593 23103
rect 24593 23069 24627 23103
rect 24627 23069 24636 23103
rect 24584 23060 24636 23069
rect 24860 23103 24912 23112
rect 24860 23069 24869 23103
rect 24869 23069 24903 23103
rect 24903 23069 24912 23103
rect 24860 23060 24912 23069
rect 27344 23060 27396 23112
rect 32128 23103 32180 23112
rect 32128 23069 32137 23103
rect 32137 23069 32171 23103
rect 32171 23069 32180 23103
rect 32128 23060 32180 23069
rect 33324 23103 33376 23112
rect 33324 23069 33333 23103
rect 33333 23069 33367 23103
rect 33367 23069 33376 23103
rect 33324 23060 33376 23069
rect 33968 23103 34020 23112
rect 33968 23069 33977 23103
rect 33977 23069 34011 23103
rect 34011 23069 34020 23103
rect 33968 23060 34020 23069
rect 34152 23060 34204 23112
rect 25228 22992 25280 23044
rect 8392 22924 8444 22976
rect 18696 22924 18748 22976
rect 20076 22924 20128 22976
rect 27160 22967 27212 22976
rect 27160 22933 27169 22967
rect 27169 22933 27203 22967
rect 27203 22933 27212 22967
rect 27160 22924 27212 22933
rect 27344 22924 27396 22976
rect 28264 22992 28316 23044
rect 34796 22992 34848 23044
rect 35808 23060 35860 23112
rect 36176 23103 36228 23112
rect 36176 23069 36185 23103
rect 36185 23069 36219 23103
rect 36219 23069 36228 23103
rect 36176 23060 36228 23069
rect 38292 23137 38301 23171
rect 38301 23137 38335 23171
rect 38335 23137 38344 23171
rect 38844 23171 38896 23180
rect 38292 23128 38344 23137
rect 38844 23137 38853 23171
rect 38853 23137 38887 23171
rect 38887 23137 38896 23171
rect 38844 23128 38896 23137
rect 44916 23171 44968 23180
rect 44916 23137 44925 23171
rect 44925 23137 44959 23171
rect 44959 23137 44968 23171
rect 44916 23128 44968 23137
rect 38108 23060 38160 23112
rect 39396 23103 39448 23112
rect 39396 23069 39405 23103
rect 39405 23069 39439 23103
rect 39439 23069 39448 23103
rect 39396 23060 39448 23069
rect 40500 23060 40552 23112
rect 40776 23060 40828 23112
rect 41696 23060 41748 23112
rect 42064 23060 42116 23112
rect 43444 23103 43496 23112
rect 36820 22992 36872 23044
rect 43444 23069 43453 23103
rect 43453 23069 43487 23103
rect 43487 23069 43496 23103
rect 43444 23060 43496 23069
rect 28908 22924 28960 22976
rect 29276 22967 29328 22976
rect 29276 22933 29285 22967
rect 29285 22933 29319 22967
rect 29319 22933 29328 22967
rect 29276 22924 29328 22933
rect 30472 22967 30524 22976
rect 30472 22933 30481 22967
rect 30481 22933 30515 22967
rect 30515 22933 30524 22967
rect 30472 22924 30524 22933
rect 37188 22924 37240 22976
rect 42892 22924 42944 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 3976 22763 4028 22772
rect 3976 22729 3985 22763
rect 3985 22729 4019 22763
rect 4019 22729 4028 22763
rect 3976 22720 4028 22729
rect 4712 22720 4764 22772
rect 6000 22720 6052 22772
rect 7012 22763 7064 22772
rect 7012 22729 7021 22763
rect 7021 22729 7055 22763
rect 7055 22729 7064 22763
rect 7012 22720 7064 22729
rect 7288 22763 7340 22772
rect 7288 22729 7297 22763
rect 7297 22729 7331 22763
rect 7331 22729 7340 22763
rect 7288 22720 7340 22729
rect 7840 22763 7892 22772
rect 7840 22729 7849 22763
rect 7849 22729 7883 22763
rect 7883 22729 7892 22763
rect 7840 22720 7892 22729
rect 8208 22763 8260 22772
rect 8208 22729 8217 22763
rect 8217 22729 8251 22763
rect 8251 22729 8260 22763
rect 8208 22720 8260 22729
rect 9496 22720 9548 22772
rect 11152 22720 11204 22772
rect 16212 22720 16264 22772
rect 16764 22763 16816 22772
rect 16764 22729 16773 22763
rect 16773 22729 16807 22763
rect 16807 22729 16816 22763
rect 16764 22720 16816 22729
rect 17316 22720 17368 22772
rect 21088 22720 21140 22772
rect 21272 22763 21324 22772
rect 21272 22729 21281 22763
rect 21281 22729 21315 22763
rect 21315 22729 21324 22763
rect 21272 22720 21324 22729
rect 23020 22720 23072 22772
rect 24584 22720 24636 22772
rect 26240 22763 26292 22772
rect 26240 22729 26249 22763
rect 26249 22729 26283 22763
rect 26283 22729 26292 22763
rect 26240 22720 26292 22729
rect 26608 22763 26660 22772
rect 26608 22729 26617 22763
rect 26617 22729 26651 22763
rect 26651 22729 26660 22763
rect 26608 22720 26660 22729
rect 28172 22720 28224 22772
rect 29000 22720 29052 22772
rect 33508 22720 33560 22772
rect 33968 22720 34020 22772
rect 34704 22763 34756 22772
rect 34704 22729 34713 22763
rect 34713 22729 34747 22763
rect 34747 22729 34756 22763
rect 34704 22720 34756 22729
rect 34796 22720 34848 22772
rect 35808 22763 35860 22772
rect 35808 22729 35817 22763
rect 35817 22729 35851 22763
rect 35851 22729 35860 22763
rect 35808 22720 35860 22729
rect 37556 22720 37608 22772
rect 38108 22763 38160 22772
rect 38108 22729 38117 22763
rect 38117 22729 38151 22763
rect 38151 22729 38160 22763
rect 38108 22720 38160 22729
rect 40500 22720 40552 22772
rect 41052 22720 41104 22772
rect 41328 22763 41380 22772
rect 41328 22729 41337 22763
rect 41337 22729 41371 22763
rect 41371 22729 41380 22763
rect 41328 22720 41380 22729
rect 43444 22720 43496 22772
rect 3608 22652 3660 22704
rect 5632 22695 5684 22704
rect 5632 22661 5641 22695
rect 5641 22661 5675 22695
rect 5675 22661 5684 22695
rect 5632 22652 5684 22661
rect 5908 22652 5960 22704
rect 11520 22652 11572 22704
rect 12900 22652 12952 22704
rect 18328 22652 18380 22704
rect 18972 22652 19024 22704
rect 21916 22652 21968 22704
rect 23296 22652 23348 22704
rect 2872 22627 2924 22636
rect 2872 22593 2881 22627
rect 2881 22593 2915 22627
rect 2915 22593 2924 22627
rect 2872 22584 2924 22593
rect 2320 22516 2372 22568
rect 4620 22584 4672 22636
rect 3976 22448 4028 22500
rect 6828 22559 6880 22568
rect 6828 22525 6837 22559
rect 6837 22525 6871 22559
rect 6871 22525 6880 22559
rect 6828 22516 6880 22525
rect 8116 22516 8168 22568
rect 13728 22584 13780 22636
rect 14740 22584 14792 22636
rect 5172 22491 5224 22500
rect 5172 22457 5181 22491
rect 5181 22457 5215 22491
rect 5215 22457 5224 22491
rect 5172 22448 5224 22457
rect 7840 22448 7892 22500
rect 10692 22516 10744 22568
rect 13360 22559 13412 22568
rect 13360 22525 13369 22559
rect 13369 22525 13403 22559
rect 13403 22525 13412 22559
rect 13360 22516 13412 22525
rect 15108 22559 15160 22568
rect 15108 22525 15117 22559
rect 15117 22525 15151 22559
rect 15151 22525 15160 22559
rect 19248 22584 19300 22636
rect 26424 22652 26476 22704
rect 26700 22652 26752 22704
rect 15108 22516 15160 22525
rect 18696 22559 18748 22568
rect 18696 22525 18705 22559
rect 18705 22525 18739 22559
rect 18739 22525 18748 22559
rect 18696 22516 18748 22525
rect 20260 22516 20312 22568
rect 24768 22584 24820 22636
rect 28356 22584 28408 22636
rect 38292 22652 38344 22704
rect 39028 22652 39080 22704
rect 31484 22584 31536 22636
rect 38016 22584 38068 22636
rect 9128 22491 9180 22500
rect 9128 22457 9137 22491
rect 9137 22457 9171 22491
rect 9171 22457 9180 22491
rect 9128 22448 9180 22457
rect 10600 22491 10652 22500
rect 10600 22457 10609 22491
rect 10609 22457 10643 22491
rect 10643 22457 10652 22491
rect 10600 22448 10652 22457
rect 11060 22448 11112 22500
rect 13452 22448 13504 22500
rect 18052 22491 18104 22500
rect 18052 22457 18061 22491
rect 18061 22457 18095 22491
rect 18095 22457 18104 22491
rect 18052 22448 18104 22457
rect 21640 22448 21692 22500
rect 22100 22516 22152 22568
rect 24676 22559 24728 22568
rect 22928 22448 22980 22500
rect 24676 22525 24685 22559
rect 24685 22525 24719 22559
rect 24719 22525 24728 22559
rect 24676 22516 24728 22525
rect 26240 22516 26292 22568
rect 26792 22559 26844 22568
rect 26792 22525 26801 22559
rect 26801 22525 26835 22559
rect 26835 22525 26844 22559
rect 26792 22516 26844 22525
rect 27160 22559 27212 22568
rect 27160 22525 27169 22559
rect 27169 22525 27203 22559
rect 27203 22525 27212 22559
rect 27160 22516 27212 22525
rect 28448 22516 28500 22568
rect 29276 22559 29328 22568
rect 29276 22525 29285 22559
rect 29285 22525 29319 22559
rect 29319 22525 29328 22559
rect 29276 22516 29328 22525
rect 29828 22516 29880 22568
rect 30472 22559 30524 22568
rect 30472 22525 30481 22559
rect 30481 22525 30515 22559
rect 30515 22525 30524 22559
rect 30472 22516 30524 22525
rect 31024 22559 31076 22568
rect 31024 22525 31033 22559
rect 31033 22525 31067 22559
rect 31067 22525 31076 22559
rect 31024 22516 31076 22525
rect 33600 22516 33652 22568
rect 1952 22423 2004 22432
rect 1952 22389 1961 22423
rect 1961 22389 1995 22423
rect 1995 22389 2004 22423
rect 1952 22380 2004 22389
rect 9680 22380 9732 22432
rect 10140 22423 10192 22432
rect 10140 22389 10149 22423
rect 10149 22389 10183 22423
rect 10183 22389 10192 22423
rect 10140 22380 10192 22389
rect 11796 22423 11848 22432
rect 11796 22389 11805 22423
rect 11805 22389 11839 22423
rect 11839 22389 11848 22423
rect 11796 22380 11848 22389
rect 13728 22423 13780 22432
rect 13728 22389 13737 22423
rect 13737 22389 13771 22423
rect 13771 22389 13780 22423
rect 13728 22380 13780 22389
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 14280 22380 14332 22389
rect 15568 22380 15620 22432
rect 18604 22380 18656 22432
rect 21824 22423 21876 22432
rect 21824 22389 21833 22423
rect 21833 22389 21867 22423
rect 21867 22389 21876 22423
rect 21824 22380 21876 22389
rect 23848 22423 23900 22432
rect 23848 22389 23857 22423
rect 23857 22389 23891 22423
rect 23891 22389 23900 22423
rect 23848 22380 23900 22389
rect 25780 22380 25832 22432
rect 29920 22448 29972 22500
rect 28448 22380 28500 22432
rect 30288 22423 30340 22432
rect 30288 22389 30297 22423
rect 30297 22389 30331 22423
rect 30331 22389 30340 22423
rect 30288 22380 30340 22389
rect 32496 22380 32548 22432
rect 32956 22380 33008 22432
rect 34244 22380 34296 22432
rect 36728 22559 36780 22568
rect 34612 22448 34664 22500
rect 36728 22525 36737 22559
rect 36737 22525 36771 22559
rect 36771 22525 36780 22559
rect 36728 22516 36780 22525
rect 37188 22516 37240 22568
rect 38384 22559 38436 22568
rect 38384 22525 38393 22559
rect 38393 22525 38427 22559
rect 38427 22525 38436 22559
rect 38384 22516 38436 22525
rect 39396 22584 39448 22636
rect 40408 22516 40460 22568
rect 43168 22627 43220 22636
rect 43168 22593 43177 22627
rect 43177 22593 43211 22627
rect 43211 22593 43220 22627
rect 43168 22584 43220 22593
rect 44180 22584 44232 22636
rect 40868 22448 40920 22500
rect 36176 22380 36228 22432
rect 39304 22380 39356 22432
rect 40316 22380 40368 22432
rect 43812 22491 43864 22500
rect 41144 22380 41196 22432
rect 41880 22380 41932 22432
rect 42892 22380 42944 22432
rect 43812 22457 43821 22491
rect 43821 22457 43855 22491
rect 43855 22457 43864 22491
rect 43812 22448 43864 22457
rect 43628 22380 43680 22432
rect 44916 22423 44968 22432
rect 44916 22389 44925 22423
rect 44925 22389 44959 22423
rect 44959 22389 44968 22423
rect 44916 22380 44968 22389
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 4620 22219 4672 22228
rect 4620 22185 4629 22219
rect 4629 22185 4663 22219
rect 4663 22185 4672 22219
rect 4620 22176 4672 22185
rect 5448 22176 5500 22228
rect 6736 22176 6788 22228
rect 8392 22176 8444 22228
rect 9588 22176 9640 22228
rect 10692 22219 10744 22228
rect 10692 22185 10701 22219
rect 10701 22185 10735 22219
rect 10735 22185 10744 22219
rect 10692 22176 10744 22185
rect 13912 22176 13964 22228
rect 18696 22176 18748 22228
rect 23480 22176 23532 22228
rect 24768 22176 24820 22228
rect 26792 22219 26844 22228
rect 3792 22108 3844 22160
rect 7196 22108 7248 22160
rect 13360 22151 13412 22160
rect 13360 22117 13369 22151
rect 13369 22117 13403 22151
rect 13403 22117 13412 22151
rect 13360 22108 13412 22117
rect 15200 22108 15252 22160
rect 17316 22108 17368 22160
rect 17868 22151 17920 22160
rect 17868 22117 17877 22151
rect 17877 22117 17911 22151
rect 17911 22117 17920 22151
rect 17868 22108 17920 22117
rect 18052 22108 18104 22160
rect 18788 22151 18840 22160
rect 18788 22117 18797 22151
rect 18797 22117 18831 22151
rect 18831 22117 18840 22151
rect 18788 22108 18840 22117
rect 21088 22151 21140 22160
rect 21088 22117 21097 22151
rect 21097 22117 21131 22151
rect 21131 22117 21140 22151
rect 21088 22108 21140 22117
rect 21732 22108 21784 22160
rect 26792 22185 26801 22219
rect 26801 22185 26835 22219
rect 26835 22185 26844 22219
rect 26792 22176 26844 22185
rect 28540 22176 28592 22228
rect 31116 22176 31168 22228
rect 33324 22176 33376 22228
rect 38384 22219 38436 22228
rect 25780 22108 25832 22160
rect 28724 22108 28776 22160
rect 29276 22108 29328 22160
rect 30380 22108 30432 22160
rect 2136 22083 2188 22092
rect 2136 22049 2145 22083
rect 2145 22049 2179 22083
rect 2179 22049 2188 22083
rect 2136 22040 2188 22049
rect 4068 22040 4120 22092
rect 8300 22040 8352 22092
rect 9680 22083 9732 22092
rect 9680 22049 9689 22083
rect 9689 22049 9723 22083
rect 9723 22049 9732 22083
rect 9680 22040 9732 22049
rect 11796 22040 11848 22092
rect 12624 22083 12676 22092
rect 12624 22049 12633 22083
rect 12633 22049 12667 22083
rect 12667 22049 12676 22083
rect 12624 22040 12676 22049
rect 5172 22015 5224 22024
rect 5172 21981 5181 22015
rect 5181 21981 5215 22015
rect 5215 21981 5224 22015
rect 5172 21972 5224 21981
rect 7012 22015 7064 22024
rect 7012 21981 7021 22015
rect 7021 21981 7055 22015
rect 7055 21981 7064 22015
rect 7012 21972 7064 21981
rect 14280 22040 14332 22092
rect 19248 22040 19300 22092
rect 3516 21904 3568 21956
rect 7564 21947 7616 21956
rect 7564 21913 7573 21947
rect 7573 21913 7607 21947
rect 7607 21913 7616 21947
rect 7564 21904 7616 21913
rect 10140 21904 10192 21956
rect 11612 21904 11664 21956
rect 13084 21904 13136 21956
rect 13636 21947 13688 21956
rect 13636 21913 13645 21947
rect 13645 21913 13679 21947
rect 13679 21913 13688 21947
rect 13636 21904 13688 21913
rect 16120 21972 16172 22024
rect 18604 21972 18656 22024
rect 20996 22015 21048 22024
rect 20996 21981 21005 22015
rect 21005 21981 21039 22015
rect 21039 21981 21048 22015
rect 20996 21972 21048 21981
rect 22928 22015 22980 22024
rect 22928 21981 22937 22015
rect 22937 21981 22971 22015
rect 22971 21981 22980 22015
rect 22928 21972 22980 21981
rect 24768 22015 24820 22024
rect 24768 21981 24777 22015
rect 24777 21981 24811 22015
rect 24811 21981 24820 22015
rect 24768 21972 24820 21981
rect 25044 22015 25096 22024
rect 25044 21981 25053 22015
rect 25053 21981 25087 22015
rect 25087 21981 25096 22015
rect 25044 21972 25096 21981
rect 16028 21904 16080 21956
rect 19432 21904 19484 21956
rect 26976 22040 27028 22092
rect 27528 22040 27580 22092
rect 29092 22040 29144 22092
rect 31024 22083 31076 22092
rect 31024 22049 31033 22083
rect 31033 22049 31067 22083
rect 31067 22049 31076 22083
rect 31024 22040 31076 22049
rect 32128 22108 32180 22160
rect 38384 22185 38393 22219
rect 38393 22185 38427 22219
rect 38427 22185 38436 22219
rect 38384 22176 38436 22185
rect 41880 22176 41932 22228
rect 42340 22176 42392 22228
rect 43168 22219 43220 22228
rect 43168 22185 43177 22219
rect 43177 22185 43211 22219
rect 43211 22185 43220 22219
rect 43168 22176 43220 22185
rect 34520 22108 34572 22160
rect 36176 22151 36228 22160
rect 36176 22117 36185 22151
rect 36185 22117 36219 22151
rect 36219 22117 36228 22151
rect 36176 22108 36228 22117
rect 36268 22151 36320 22160
rect 36268 22117 36277 22151
rect 36277 22117 36311 22151
rect 36311 22117 36320 22151
rect 36268 22108 36320 22117
rect 41696 22108 41748 22160
rect 33140 22040 33192 22092
rect 37832 22083 37884 22092
rect 37832 22049 37850 22083
rect 37850 22049 37884 22083
rect 37832 22040 37884 22049
rect 38292 22040 38344 22092
rect 39212 22083 39264 22092
rect 2688 21836 2740 21888
rect 4988 21879 5040 21888
rect 4988 21845 4997 21879
rect 4997 21845 5031 21879
rect 5031 21845 5040 21879
rect 4988 21836 5040 21845
rect 10232 21836 10284 21888
rect 10600 21836 10652 21888
rect 13360 21836 13412 21888
rect 20260 21836 20312 21888
rect 22100 21879 22152 21888
rect 22100 21845 22109 21879
rect 22109 21845 22143 21879
rect 22143 21845 22152 21879
rect 22100 21836 22152 21845
rect 25504 21836 25556 21888
rect 28172 21972 28224 22024
rect 28448 22015 28500 22024
rect 28448 21981 28457 22015
rect 28457 21981 28491 22015
rect 28491 21981 28500 22015
rect 28448 21972 28500 21981
rect 33876 22015 33928 22024
rect 29552 21904 29604 21956
rect 33876 21981 33885 22015
rect 33885 21981 33919 22015
rect 33919 21981 33928 22015
rect 33876 21972 33928 21981
rect 34152 22015 34204 22024
rect 34152 21981 34161 22015
rect 34161 21981 34195 22015
rect 34195 21981 34204 22015
rect 34152 21972 34204 21981
rect 36820 22015 36872 22024
rect 36820 21981 36829 22015
rect 36829 21981 36863 22015
rect 36863 21981 36872 22015
rect 36820 21972 36872 21981
rect 38200 21972 38252 22024
rect 39212 22049 39221 22083
rect 39221 22049 39255 22083
rect 39255 22049 39264 22083
rect 39212 22040 39264 22049
rect 42984 22040 43036 22092
rect 43352 22083 43404 22092
rect 43352 22049 43396 22083
rect 43396 22049 43404 22083
rect 43352 22040 43404 22049
rect 44824 22040 44876 22092
rect 39488 22015 39540 22024
rect 39488 21981 39497 22015
rect 39497 21981 39531 22015
rect 39531 21981 39540 22015
rect 39488 21972 39540 21981
rect 41328 22015 41380 22024
rect 41328 21981 41337 22015
rect 41337 21981 41371 22015
rect 41371 21981 41380 22015
rect 41328 21972 41380 21981
rect 40592 21904 40644 21956
rect 40960 21904 41012 21956
rect 41788 21972 41840 22024
rect 43812 21972 43864 22024
rect 43996 21972 44048 22024
rect 27344 21836 27396 21888
rect 27528 21836 27580 21888
rect 27988 21836 28040 21888
rect 28356 21879 28408 21888
rect 28356 21845 28365 21879
rect 28365 21845 28399 21879
rect 28399 21845 28408 21879
rect 28356 21836 28408 21845
rect 29276 21836 29328 21888
rect 35348 21879 35400 21888
rect 35348 21845 35357 21879
rect 35357 21845 35391 21879
rect 35391 21845 35400 21879
rect 35348 21836 35400 21845
rect 36912 21836 36964 21888
rect 40500 21879 40552 21888
rect 40500 21845 40509 21879
rect 40509 21845 40543 21879
rect 40543 21845 40552 21879
rect 40500 21836 40552 21845
rect 43904 21836 43956 21888
rect 44548 21879 44600 21888
rect 44548 21845 44557 21879
rect 44557 21845 44591 21879
rect 44591 21845 44600 21879
rect 44548 21836 44600 21845
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 3332 21632 3384 21684
rect 3516 21675 3568 21684
rect 3516 21641 3525 21675
rect 3525 21641 3559 21675
rect 3559 21641 3568 21675
rect 3516 21632 3568 21641
rect 4068 21675 4120 21684
rect 4068 21641 4077 21675
rect 4077 21641 4111 21675
rect 4111 21641 4120 21675
rect 4068 21632 4120 21641
rect 5448 21632 5500 21684
rect 8300 21632 8352 21684
rect 8392 21675 8444 21684
rect 8392 21641 8401 21675
rect 8401 21641 8435 21675
rect 8435 21641 8444 21675
rect 11796 21675 11848 21684
rect 8392 21632 8444 21641
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 12624 21632 12676 21684
rect 15200 21675 15252 21684
rect 15200 21641 15209 21675
rect 15209 21641 15243 21675
rect 15243 21641 15252 21675
rect 15200 21632 15252 21641
rect 17868 21632 17920 21684
rect 19248 21675 19300 21684
rect 19248 21641 19257 21675
rect 19257 21641 19291 21675
rect 19291 21641 19300 21675
rect 19248 21632 19300 21641
rect 19432 21632 19484 21684
rect 4988 21496 5040 21548
rect 1400 21292 1452 21344
rect 2136 21428 2188 21480
rect 3516 21428 3568 21480
rect 4712 21360 4764 21412
rect 5448 21360 5500 21412
rect 8116 21428 8168 21480
rect 9404 21564 9456 21616
rect 10968 21564 11020 21616
rect 14004 21564 14056 21616
rect 18052 21564 18104 21616
rect 9680 21539 9732 21548
rect 9680 21505 9689 21539
rect 9689 21505 9723 21539
rect 9723 21505 9732 21539
rect 9680 21496 9732 21505
rect 13912 21539 13964 21548
rect 13912 21505 13921 21539
rect 13921 21505 13955 21539
rect 13955 21505 13964 21539
rect 13912 21496 13964 21505
rect 16028 21539 16080 21548
rect 16028 21505 16037 21539
rect 16037 21505 16071 21539
rect 16071 21505 16080 21539
rect 16028 21496 16080 21505
rect 18512 21496 18564 21548
rect 18604 21539 18656 21548
rect 18604 21505 18613 21539
rect 18613 21505 18647 21539
rect 18647 21505 18656 21539
rect 18604 21496 18656 21505
rect 7564 21403 7616 21412
rect 5540 21335 5592 21344
rect 5540 21301 5549 21335
rect 5549 21301 5583 21335
rect 5583 21301 5592 21335
rect 5540 21292 5592 21301
rect 6736 21292 6788 21344
rect 7564 21369 7573 21403
rect 7573 21369 7607 21403
rect 7607 21369 7616 21403
rect 7564 21360 7616 21369
rect 8392 21360 8444 21412
rect 10876 21403 10928 21412
rect 10876 21369 10885 21403
rect 10885 21369 10919 21403
rect 10919 21369 10928 21403
rect 10876 21360 10928 21369
rect 10968 21403 11020 21412
rect 10968 21369 10977 21403
rect 10977 21369 11011 21403
rect 11011 21369 11020 21403
rect 10968 21360 11020 21369
rect 12072 21360 12124 21412
rect 13636 21428 13688 21480
rect 21088 21632 21140 21684
rect 21640 21675 21692 21684
rect 21640 21641 21649 21675
rect 21649 21641 21683 21675
rect 21683 21641 21692 21675
rect 21640 21632 21692 21641
rect 23296 21632 23348 21684
rect 25504 21675 25556 21684
rect 25504 21641 25513 21675
rect 25513 21641 25547 21675
rect 25547 21641 25556 21675
rect 25504 21632 25556 21641
rect 25964 21632 26016 21684
rect 26976 21675 27028 21684
rect 26976 21641 26985 21675
rect 26985 21641 27019 21675
rect 27019 21641 27028 21675
rect 26976 21632 27028 21641
rect 27896 21632 27948 21684
rect 28724 21632 28776 21684
rect 21732 21564 21784 21616
rect 27804 21607 27856 21616
rect 20260 21539 20312 21548
rect 20260 21505 20269 21539
rect 20269 21505 20303 21539
rect 20303 21505 20312 21539
rect 20260 21496 20312 21505
rect 22836 21496 22888 21548
rect 27804 21573 27813 21607
rect 27813 21573 27847 21607
rect 27847 21573 27856 21607
rect 27804 21564 27856 21573
rect 29276 21564 29328 21616
rect 29552 21607 29604 21616
rect 29552 21573 29561 21607
rect 29561 21573 29595 21607
rect 29595 21573 29604 21607
rect 29552 21564 29604 21573
rect 12164 21335 12216 21344
rect 12164 21301 12173 21335
rect 12173 21301 12207 21335
rect 12207 21301 12216 21335
rect 12164 21292 12216 21301
rect 12256 21292 12308 21344
rect 13084 21292 13136 21344
rect 20076 21428 20128 21480
rect 21732 21428 21784 21480
rect 15752 21403 15804 21412
rect 15752 21369 15761 21403
rect 15761 21369 15795 21403
rect 15795 21369 15804 21403
rect 15752 21360 15804 21369
rect 18236 21403 18288 21412
rect 14832 21335 14884 21344
rect 14832 21301 14841 21335
rect 14841 21301 14875 21335
rect 14875 21301 14884 21335
rect 14832 21292 14884 21301
rect 15568 21335 15620 21344
rect 15568 21301 15577 21335
rect 15577 21301 15611 21335
rect 15611 21301 15620 21335
rect 18236 21369 18245 21403
rect 18245 21369 18279 21403
rect 18279 21369 18288 21403
rect 18236 21360 18288 21369
rect 21640 21360 21692 21412
rect 23480 21428 23532 21480
rect 23296 21360 23348 21412
rect 25044 21496 25096 21548
rect 25596 21539 25648 21548
rect 25596 21505 25605 21539
rect 25605 21505 25639 21539
rect 25639 21505 25648 21539
rect 25596 21496 25648 21505
rect 27528 21496 27580 21548
rect 28448 21496 28500 21548
rect 29644 21539 29696 21548
rect 29644 21505 29653 21539
rect 29653 21505 29687 21539
rect 29687 21505 29696 21539
rect 29644 21496 29696 21505
rect 33600 21496 33652 21548
rect 33876 21632 33928 21684
rect 43352 21675 43404 21684
rect 43352 21641 43361 21675
rect 43361 21641 43395 21675
rect 43395 21641 43404 21675
rect 43352 21632 43404 21641
rect 37464 21607 37516 21616
rect 37464 21573 37473 21607
rect 37473 21573 37507 21607
rect 37507 21573 37516 21607
rect 37464 21564 37516 21573
rect 35348 21539 35400 21548
rect 35348 21505 35357 21539
rect 35357 21505 35391 21539
rect 35391 21505 35400 21539
rect 35348 21496 35400 21505
rect 35624 21539 35676 21548
rect 35624 21505 35633 21539
rect 35633 21505 35667 21539
rect 35667 21505 35676 21539
rect 35624 21496 35676 21505
rect 36360 21496 36412 21548
rect 36912 21539 36964 21548
rect 36912 21505 36921 21539
rect 36921 21505 36955 21539
rect 36955 21505 36964 21539
rect 36912 21496 36964 21505
rect 40500 21539 40552 21548
rect 40500 21505 40509 21539
rect 40509 21505 40543 21539
rect 40543 21505 40552 21539
rect 40500 21496 40552 21505
rect 42340 21539 42392 21548
rect 42340 21505 42349 21539
rect 42349 21505 42383 21539
rect 42383 21505 42392 21539
rect 42340 21496 42392 21505
rect 43260 21496 43312 21548
rect 43904 21539 43956 21548
rect 43904 21505 43913 21539
rect 43913 21505 43947 21539
rect 43947 21505 43956 21539
rect 43904 21496 43956 21505
rect 25136 21428 25188 21480
rect 27988 21428 28040 21480
rect 28172 21428 28224 21480
rect 32128 21471 32180 21480
rect 32128 21437 32137 21471
rect 32137 21437 32171 21471
rect 32171 21437 32180 21471
rect 32128 21428 32180 21437
rect 32588 21471 32640 21480
rect 32588 21437 32597 21471
rect 32597 21437 32631 21471
rect 32631 21437 32640 21471
rect 32588 21428 32640 21437
rect 38292 21428 38344 21480
rect 23756 21403 23808 21412
rect 23756 21369 23765 21403
rect 23765 21369 23799 21403
rect 23799 21369 23808 21403
rect 23756 21360 23808 21369
rect 24216 21360 24268 21412
rect 26516 21360 26568 21412
rect 27528 21403 27580 21412
rect 27528 21369 27537 21403
rect 27537 21369 27571 21403
rect 27571 21369 27580 21403
rect 27528 21360 27580 21369
rect 29184 21360 29236 21412
rect 30380 21360 30432 21412
rect 32864 21403 32916 21412
rect 32864 21369 32873 21403
rect 32873 21369 32907 21403
rect 32907 21369 32916 21403
rect 32864 21360 32916 21369
rect 33140 21360 33192 21412
rect 35164 21360 35216 21412
rect 25136 21335 25188 21344
rect 15568 21292 15620 21301
rect 25136 21301 25145 21335
rect 25145 21301 25179 21335
rect 25179 21301 25188 21335
rect 25136 21292 25188 21301
rect 27436 21335 27488 21344
rect 27436 21301 27445 21335
rect 27445 21301 27479 21335
rect 27479 21301 27488 21335
rect 27436 21292 27488 21301
rect 27804 21292 27856 21344
rect 28356 21292 28408 21344
rect 31116 21292 31168 21344
rect 31668 21292 31720 21344
rect 34520 21335 34572 21344
rect 34520 21301 34529 21335
rect 34529 21301 34563 21335
rect 34563 21301 34572 21335
rect 34520 21292 34572 21301
rect 36268 21335 36320 21344
rect 36268 21301 36277 21335
rect 36277 21301 36311 21335
rect 36311 21301 36320 21335
rect 36268 21292 36320 21301
rect 37648 21360 37700 21412
rect 39212 21428 39264 21480
rect 43996 21403 44048 21412
rect 38200 21292 38252 21344
rect 40316 21335 40368 21344
rect 40316 21301 40325 21335
rect 40325 21301 40359 21335
rect 40359 21301 40368 21335
rect 40316 21292 40368 21301
rect 41420 21335 41472 21344
rect 41420 21301 41429 21335
rect 41429 21301 41463 21335
rect 41463 21301 41472 21335
rect 41420 21292 41472 21301
rect 41696 21335 41748 21344
rect 41696 21301 41705 21335
rect 41705 21301 41739 21335
rect 41739 21301 41748 21335
rect 41696 21292 41748 21301
rect 43996 21369 44005 21403
rect 44005 21369 44039 21403
rect 44039 21369 44048 21403
rect 43996 21360 44048 21369
rect 44824 21335 44876 21344
rect 44824 21301 44833 21335
rect 44833 21301 44867 21335
rect 44867 21301 44876 21335
rect 44824 21292 44876 21301
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 5172 21131 5224 21140
rect 5172 21097 5181 21131
rect 5181 21097 5215 21131
rect 5215 21097 5224 21131
rect 5172 21088 5224 21097
rect 7012 21088 7064 21140
rect 12164 21088 12216 21140
rect 14280 21131 14332 21140
rect 14280 21097 14289 21131
rect 14289 21097 14323 21131
rect 14323 21097 14332 21131
rect 14280 21088 14332 21097
rect 15752 21131 15804 21140
rect 15752 21097 15761 21131
rect 15761 21097 15795 21131
rect 15795 21097 15804 21131
rect 15752 21088 15804 21097
rect 16120 21131 16172 21140
rect 16120 21097 16129 21131
rect 16129 21097 16163 21131
rect 16163 21097 16172 21131
rect 16120 21088 16172 21097
rect 18512 21131 18564 21140
rect 18512 21097 18521 21131
rect 18521 21097 18555 21131
rect 18555 21097 18564 21131
rect 18512 21088 18564 21097
rect 20076 21088 20128 21140
rect 21732 21131 21784 21140
rect 21732 21097 21741 21131
rect 21741 21097 21775 21131
rect 21775 21097 21784 21131
rect 21732 21088 21784 21097
rect 22928 21131 22980 21140
rect 22928 21097 22937 21131
rect 22937 21097 22971 21131
rect 22971 21097 22980 21131
rect 22928 21088 22980 21097
rect 23756 21131 23808 21140
rect 23756 21097 23765 21131
rect 23765 21097 23799 21131
rect 23799 21097 23808 21131
rect 23756 21088 23808 21097
rect 24768 21088 24820 21140
rect 28816 21088 28868 21140
rect 32588 21088 32640 21140
rect 4988 21020 5040 21072
rect 10784 21020 10836 21072
rect 11612 21063 11664 21072
rect 11612 21029 11621 21063
rect 11621 21029 11655 21063
rect 11655 21029 11664 21063
rect 11612 21020 11664 21029
rect 17316 21063 17368 21072
rect 17316 21029 17325 21063
rect 17325 21029 17359 21063
rect 17359 21029 17368 21063
rect 17316 21020 17368 21029
rect 25872 21020 25924 21072
rect 32496 21020 32548 21072
rect 34520 21088 34572 21140
rect 35348 21088 35400 21140
rect 36912 21088 36964 21140
rect 41328 21088 41380 21140
rect 43996 21088 44048 21140
rect 36176 21063 36228 21072
rect 36176 21029 36185 21063
rect 36185 21029 36219 21063
rect 36219 21029 36228 21063
rect 36176 21020 36228 21029
rect 39212 21020 39264 21072
rect 40316 21020 40368 21072
rect 41052 21020 41104 21072
rect 41696 21020 41748 21072
rect 42064 21063 42116 21072
rect 42064 21029 42073 21063
rect 42073 21029 42107 21063
rect 42107 21029 42116 21063
rect 42064 21020 42116 21029
rect 43536 21063 43588 21072
rect 43536 21029 43545 21063
rect 43545 21029 43579 21063
rect 43579 21029 43588 21063
rect 43536 21020 43588 21029
rect 43812 21020 43864 21072
rect 3884 20952 3936 21004
rect 4620 20995 4672 21004
rect 4620 20961 4629 20995
rect 4629 20961 4663 20995
rect 4663 20961 4672 20995
rect 4620 20952 4672 20961
rect 5540 20952 5592 21004
rect 7104 20952 7156 21004
rect 7748 20995 7800 21004
rect 7748 20961 7757 20995
rect 7757 20961 7791 20995
rect 7791 20961 7800 20995
rect 7748 20952 7800 20961
rect 8208 20995 8260 21004
rect 8208 20961 8217 20995
rect 8217 20961 8251 20995
rect 8251 20961 8260 20995
rect 8208 20952 8260 20961
rect 12900 20952 12952 21004
rect 13084 20952 13136 21004
rect 14832 20952 14884 21004
rect 15292 20995 15344 21004
rect 15292 20961 15336 20995
rect 15336 20961 15344 20995
rect 15292 20952 15344 20961
rect 18328 20952 18380 21004
rect 19064 20952 19116 21004
rect 21916 20995 21968 21004
rect 21916 20961 21925 20995
rect 21925 20961 21959 20995
rect 21959 20961 21968 20995
rect 21916 20952 21968 20961
rect 22100 20995 22152 21004
rect 22100 20961 22109 20995
rect 22109 20961 22143 20995
rect 22143 20961 22152 20995
rect 22100 20952 22152 20961
rect 23204 20995 23256 21004
rect 23204 20961 23213 20995
rect 23213 20961 23247 20995
rect 23247 20961 23256 20995
rect 23204 20952 23256 20961
rect 25412 20952 25464 21004
rect 26516 20995 26568 21004
rect 26516 20961 26525 20995
rect 26525 20961 26559 20995
rect 26559 20961 26568 20995
rect 26516 20952 26568 20961
rect 27896 20952 27948 21004
rect 29092 20995 29144 21004
rect 29092 20961 29101 20995
rect 29101 20961 29135 20995
rect 29135 20961 29144 20995
rect 29092 20952 29144 20961
rect 30656 20995 30708 21004
rect 30656 20961 30665 20995
rect 30665 20961 30699 20995
rect 30699 20961 30708 20995
rect 30656 20952 30708 20961
rect 32312 20952 32364 21004
rect 32772 20952 32824 21004
rect 32864 20952 32916 21004
rect 33416 20952 33468 21004
rect 35256 20952 35308 21004
rect 39488 20952 39540 21004
rect 45468 20952 45520 21004
rect 10508 20884 10560 20936
rect 12256 20884 12308 20936
rect 13544 20927 13596 20936
rect 13544 20893 13553 20927
rect 13553 20893 13587 20927
rect 13587 20893 13596 20927
rect 13544 20884 13596 20893
rect 16948 20884 17000 20936
rect 18972 20884 19024 20936
rect 25136 20884 25188 20936
rect 12072 20859 12124 20868
rect 12072 20825 12081 20859
rect 12081 20825 12115 20859
rect 12115 20825 12124 20859
rect 12072 20816 12124 20825
rect 7012 20791 7064 20800
rect 7012 20757 7021 20791
rect 7021 20757 7055 20791
rect 7055 20757 7064 20791
rect 7012 20748 7064 20757
rect 13360 20748 13412 20800
rect 17960 20816 18012 20868
rect 20996 20816 21048 20868
rect 22100 20816 22152 20868
rect 24308 20816 24360 20868
rect 25596 20884 25648 20936
rect 28816 20884 28868 20936
rect 27068 20816 27120 20868
rect 29000 20816 29052 20868
rect 29276 20859 29328 20868
rect 29276 20825 29282 20859
rect 29282 20825 29328 20859
rect 29276 20816 29328 20825
rect 29552 20884 29604 20936
rect 30564 20884 30616 20936
rect 36084 20927 36136 20936
rect 31024 20816 31076 20868
rect 36084 20893 36093 20927
rect 36093 20893 36127 20927
rect 36127 20893 36136 20927
rect 36084 20884 36136 20893
rect 36360 20927 36412 20936
rect 36360 20893 36369 20927
rect 36369 20893 36403 20927
rect 36403 20893 36412 20927
rect 36360 20884 36412 20893
rect 32772 20816 32824 20868
rect 38200 20884 38252 20936
rect 40776 20884 40828 20936
rect 42616 20884 42668 20936
rect 38476 20859 38528 20868
rect 38476 20825 38485 20859
rect 38485 20825 38519 20859
rect 38519 20825 38528 20859
rect 38476 20816 38528 20825
rect 18236 20791 18288 20800
rect 18236 20757 18245 20791
rect 18245 20757 18279 20791
rect 18279 20757 18288 20791
rect 18236 20748 18288 20757
rect 21272 20791 21324 20800
rect 21272 20757 21281 20791
rect 21281 20757 21315 20791
rect 21315 20757 21324 20791
rect 21272 20748 21324 20757
rect 25504 20748 25556 20800
rect 25872 20791 25924 20800
rect 25872 20757 25881 20791
rect 25881 20757 25915 20791
rect 25915 20757 25924 20791
rect 25872 20748 25924 20757
rect 26608 20748 26660 20800
rect 26792 20791 26844 20800
rect 26792 20757 26801 20791
rect 26801 20757 26835 20791
rect 26835 20757 26844 20791
rect 26792 20748 26844 20757
rect 27620 20791 27672 20800
rect 27620 20757 27629 20791
rect 27629 20757 27663 20791
rect 27663 20757 27672 20791
rect 27620 20748 27672 20757
rect 27988 20791 28040 20800
rect 27988 20757 27997 20791
rect 27997 20757 28031 20791
rect 28031 20757 28040 20791
rect 27988 20748 28040 20757
rect 29092 20748 29144 20800
rect 29368 20791 29420 20800
rect 29368 20757 29377 20791
rect 29377 20757 29411 20791
rect 29411 20757 29420 20791
rect 29368 20748 29420 20757
rect 31944 20748 31996 20800
rect 32128 20748 32180 20800
rect 39304 20748 39356 20800
rect 41052 20748 41104 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 3884 20544 3936 20596
rect 4712 20544 4764 20596
rect 5540 20544 5592 20596
rect 7656 20587 7708 20596
rect 7656 20553 7665 20587
rect 7665 20553 7699 20587
rect 7699 20553 7708 20587
rect 7656 20544 7708 20553
rect 10876 20544 10928 20596
rect 12256 20544 12308 20596
rect 12900 20544 12952 20596
rect 13636 20587 13688 20596
rect 13636 20553 13645 20587
rect 13645 20553 13679 20587
rect 13679 20553 13688 20587
rect 13636 20544 13688 20553
rect 15292 20587 15344 20596
rect 15292 20553 15301 20587
rect 15301 20553 15335 20587
rect 15335 20553 15344 20587
rect 15292 20544 15344 20553
rect 19064 20587 19116 20596
rect 19064 20553 19073 20587
rect 19073 20553 19107 20587
rect 19107 20553 19116 20587
rect 19064 20544 19116 20553
rect 22100 20544 22152 20596
rect 23204 20544 23256 20596
rect 26516 20544 26568 20596
rect 27160 20544 27212 20596
rect 29184 20544 29236 20596
rect 30656 20587 30708 20596
rect 30656 20553 30665 20587
rect 30665 20553 30699 20587
rect 30699 20553 30708 20587
rect 30656 20544 30708 20553
rect 30748 20544 30800 20596
rect 31484 20587 31536 20596
rect 31484 20553 31493 20587
rect 31493 20553 31527 20587
rect 31527 20553 31536 20587
rect 31484 20544 31536 20553
rect 31944 20587 31996 20596
rect 31944 20553 31953 20587
rect 31953 20553 31987 20587
rect 31987 20553 31996 20587
rect 31944 20544 31996 20553
rect 36084 20544 36136 20596
rect 36176 20544 36228 20596
rect 37924 20544 37976 20596
rect 38108 20587 38160 20596
rect 38108 20553 38117 20587
rect 38117 20553 38151 20587
rect 38151 20553 38160 20587
rect 38108 20544 38160 20553
rect 39488 20544 39540 20596
rect 40776 20587 40828 20596
rect 40776 20553 40785 20587
rect 40785 20553 40819 20587
rect 40819 20553 40828 20587
rect 40776 20544 40828 20553
rect 41052 20587 41104 20596
rect 41052 20553 41061 20587
rect 41061 20553 41095 20587
rect 41095 20553 41104 20587
rect 41052 20544 41104 20553
rect 42616 20587 42668 20596
rect 42616 20553 42625 20587
rect 42625 20553 42659 20587
rect 42659 20553 42668 20587
rect 42616 20544 42668 20553
rect 43536 20544 43588 20596
rect 3240 20476 3292 20528
rect 21916 20476 21968 20528
rect 26792 20476 26844 20528
rect 2780 20340 2832 20392
rect 3976 20408 4028 20460
rect 4620 20408 4672 20460
rect 3792 20340 3844 20392
rect 4712 20272 4764 20324
rect 6736 20408 6788 20460
rect 11612 20408 11664 20460
rect 12072 20408 12124 20460
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 18604 20408 18656 20460
rect 20076 20408 20128 20460
rect 24216 20451 24268 20460
rect 24216 20417 24225 20451
rect 24225 20417 24259 20451
rect 24259 20417 24268 20451
rect 24216 20408 24268 20417
rect 25872 20451 25924 20460
rect 25872 20417 25881 20451
rect 25881 20417 25915 20451
rect 25915 20417 25924 20451
rect 25872 20408 25924 20417
rect 7656 20340 7708 20392
rect 8208 20383 8260 20392
rect 8208 20349 8217 20383
rect 8217 20349 8251 20383
rect 8251 20349 8260 20383
rect 8208 20340 8260 20349
rect 5724 20272 5776 20324
rect 8300 20272 8352 20324
rect 5172 20247 5224 20256
rect 5172 20213 5181 20247
rect 5181 20213 5215 20247
rect 5215 20213 5224 20247
rect 5172 20204 5224 20213
rect 9312 20383 9364 20392
rect 9312 20349 9321 20383
rect 9321 20349 9355 20383
rect 9355 20349 9364 20383
rect 9312 20340 9364 20349
rect 8852 20247 8904 20256
rect 8852 20213 8861 20247
rect 8861 20213 8895 20247
rect 8895 20213 8904 20247
rect 8852 20204 8904 20213
rect 13360 20340 13412 20392
rect 13636 20272 13688 20324
rect 10784 20204 10836 20256
rect 12716 20247 12768 20256
rect 12716 20213 12725 20247
rect 12725 20213 12759 20247
rect 12759 20213 12768 20247
rect 12716 20204 12768 20213
rect 12992 20247 13044 20256
rect 12992 20213 13001 20247
rect 13001 20213 13035 20247
rect 13035 20213 13044 20247
rect 12992 20204 13044 20213
rect 21272 20383 21324 20392
rect 21272 20349 21281 20383
rect 21281 20349 21315 20383
rect 21315 20349 21324 20383
rect 21272 20340 21324 20349
rect 23020 20340 23072 20392
rect 18236 20315 18288 20324
rect 15476 20204 15528 20256
rect 16396 20247 16448 20256
rect 16396 20213 16405 20247
rect 16405 20213 16439 20247
rect 16439 20213 16448 20247
rect 16396 20204 16448 20213
rect 16580 20204 16632 20256
rect 17316 20204 17368 20256
rect 18236 20281 18245 20315
rect 18245 20281 18279 20315
rect 18279 20281 18288 20315
rect 18236 20272 18288 20281
rect 18788 20315 18840 20324
rect 18788 20281 18797 20315
rect 18797 20281 18831 20315
rect 18831 20281 18840 20315
rect 18788 20272 18840 20281
rect 20352 20315 20404 20324
rect 19432 20204 19484 20256
rect 20352 20281 20361 20315
rect 20361 20281 20395 20315
rect 20395 20281 20404 20315
rect 20352 20272 20404 20281
rect 22652 20204 22704 20256
rect 25136 20204 25188 20256
rect 26608 20340 26660 20392
rect 27068 20383 27120 20392
rect 27068 20349 27077 20383
rect 27077 20349 27111 20383
rect 27111 20349 27120 20383
rect 27068 20340 27120 20349
rect 28724 20340 28776 20392
rect 29276 20476 29328 20528
rect 29552 20519 29604 20528
rect 29552 20485 29561 20519
rect 29561 20485 29595 20519
rect 29595 20485 29604 20519
rect 31116 20519 31168 20528
rect 29552 20476 29604 20485
rect 31116 20485 31125 20519
rect 31125 20485 31159 20519
rect 31159 20485 31168 20519
rect 31116 20476 31168 20485
rect 31300 20476 31352 20528
rect 33784 20476 33836 20528
rect 39028 20476 39080 20528
rect 29644 20451 29696 20460
rect 29644 20417 29653 20451
rect 29653 20417 29687 20451
rect 29687 20417 29696 20451
rect 29644 20408 29696 20417
rect 25412 20272 25464 20324
rect 26332 20204 26384 20256
rect 27896 20204 27948 20256
rect 28264 20204 28316 20256
rect 29092 20272 29144 20324
rect 29644 20272 29696 20324
rect 30012 20315 30064 20324
rect 30012 20281 30021 20315
rect 30021 20281 30055 20315
rect 30055 20281 30064 20315
rect 30012 20272 30064 20281
rect 28724 20247 28776 20256
rect 28724 20213 28733 20247
rect 28733 20213 28767 20247
rect 28767 20213 28776 20247
rect 28724 20204 28776 20213
rect 34152 20408 34204 20460
rect 31024 20340 31076 20392
rect 35900 20340 35952 20392
rect 36084 20340 36136 20392
rect 38476 20408 38528 20460
rect 42064 20476 42116 20528
rect 42800 20476 42852 20528
rect 44456 20451 44508 20460
rect 44456 20417 44465 20451
rect 44465 20417 44499 20451
rect 44499 20417 44508 20451
rect 44456 20408 44508 20417
rect 45468 20451 45520 20460
rect 45468 20417 45477 20451
rect 45477 20417 45511 20451
rect 45511 20417 45520 20451
rect 45468 20408 45520 20417
rect 37004 20383 37056 20392
rect 37004 20349 37022 20383
rect 37022 20349 37056 20383
rect 37004 20340 37056 20349
rect 33784 20315 33836 20324
rect 32496 20204 32548 20256
rect 32956 20204 33008 20256
rect 33784 20281 33793 20315
rect 33793 20281 33827 20315
rect 33827 20281 33836 20315
rect 33784 20272 33836 20281
rect 35164 20247 35216 20256
rect 35164 20213 35173 20247
rect 35173 20213 35207 20247
rect 35207 20213 35216 20247
rect 35164 20204 35216 20213
rect 37280 20204 37332 20256
rect 37740 20247 37792 20256
rect 37740 20213 37749 20247
rect 37749 20213 37783 20247
rect 37783 20213 37792 20247
rect 38476 20272 38528 20324
rect 40960 20272 41012 20324
rect 41420 20315 41472 20324
rect 41420 20281 41429 20315
rect 41429 20281 41463 20315
rect 41463 20281 41472 20315
rect 41972 20315 42024 20324
rect 41420 20272 41472 20281
rect 41972 20281 41981 20315
rect 41981 20281 42015 20315
rect 42015 20281 42024 20315
rect 41972 20272 42024 20281
rect 43536 20272 43588 20324
rect 37740 20204 37792 20213
rect 40316 20204 40368 20256
rect 45008 20247 45060 20256
rect 45008 20213 45017 20247
rect 45017 20213 45051 20247
rect 45051 20213 45060 20247
rect 45008 20204 45060 20213
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 2780 20043 2832 20052
rect 2780 20009 2789 20043
rect 2789 20009 2823 20043
rect 2823 20009 2832 20043
rect 2780 20000 2832 20009
rect 3792 20043 3844 20052
rect 3792 20009 3801 20043
rect 3801 20009 3835 20043
rect 3835 20009 3844 20043
rect 3792 20000 3844 20009
rect 4712 20043 4764 20052
rect 4712 20009 4721 20043
rect 4721 20009 4755 20043
rect 4755 20009 4764 20043
rect 4712 20000 4764 20009
rect 7748 20043 7800 20052
rect 7748 20009 7757 20043
rect 7757 20009 7791 20043
rect 7791 20009 7800 20043
rect 7748 20000 7800 20009
rect 8300 20043 8352 20052
rect 8300 20009 8309 20043
rect 8309 20009 8343 20043
rect 8343 20009 8352 20043
rect 8300 20000 8352 20009
rect 9312 20043 9364 20052
rect 9312 20009 9321 20043
rect 9321 20009 9355 20043
rect 9355 20009 9364 20043
rect 9312 20000 9364 20009
rect 10508 20043 10560 20052
rect 10508 20009 10517 20043
rect 10517 20009 10551 20043
rect 10551 20009 10560 20043
rect 10508 20000 10560 20009
rect 13268 20000 13320 20052
rect 13636 20000 13688 20052
rect 16396 20000 16448 20052
rect 16948 20043 17000 20052
rect 16948 20009 16957 20043
rect 16957 20009 16991 20043
rect 16991 20009 17000 20043
rect 16948 20000 17000 20009
rect 18144 20043 18196 20052
rect 18144 20009 18153 20043
rect 18153 20009 18187 20043
rect 18187 20009 18196 20043
rect 18144 20000 18196 20009
rect 20076 20043 20128 20052
rect 20076 20009 20085 20043
rect 20085 20009 20119 20043
rect 20119 20009 20128 20043
rect 20076 20000 20128 20009
rect 26792 20000 26844 20052
rect 27528 20000 27580 20052
rect 28080 20000 28132 20052
rect 28816 20043 28868 20052
rect 28816 20009 28825 20043
rect 28825 20009 28859 20043
rect 28859 20009 28868 20043
rect 28816 20000 28868 20009
rect 29000 20000 29052 20052
rect 30748 20043 30800 20052
rect 6736 19975 6788 19984
rect 6736 19941 6745 19975
rect 6745 19941 6779 19975
rect 6779 19941 6788 19975
rect 6736 19932 6788 19941
rect 10324 19932 10376 19984
rect 13360 19932 13412 19984
rect 15476 19975 15528 19984
rect 15476 19941 15485 19975
rect 15485 19941 15519 19975
rect 15519 19941 15528 19975
rect 15476 19932 15528 19941
rect 15568 19975 15620 19984
rect 15568 19941 15577 19975
rect 15577 19941 15611 19975
rect 15611 19941 15620 19975
rect 15568 19932 15620 19941
rect 18052 19932 18104 19984
rect 25504 19932 25556 19984
rect 3792 19864 3844 19916
rect 7932 19864 7984 19916
rect 8852 19864 8904 19916
rect 9128 19864 9180 19916
rect 9680 19907 9732 19916
rect 9680 19873 9689 19907
rect 9689 19873 9723 19907
rect 9723 19873 9732 19907
rect 9680 19864 9732 19873
rect 11060 19864 11112 19916
rect 11888 19907 11940 19916
rect 11888 19873 11897 19907
rect 11897 19873 11931 19907
rect 11931 19873 11940 19907
rect 11888 19864 11940 19873
rect 12348 19907 12400 19916
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12992 19907 13044 19916
rect 12348 19864 12400 19873
rect 12992 19873 13001 19907
rect 13001 19873 13035 19907
rect 13035 19873 13044 19907
rect 12992 19864 13044 19873
rect 13544 19864 13596 19916
rect 20996 19907 21048 19916
rect 20996 19873 21005 19907
rect 21005 19873 21039 19907
rect 21039 19873 21048 19907
rect 20996 19864 21048 19873
rect 23204 19864 23256 19916
rect 25320 19907 25372 19916
rect 25320 19873 25329 19907
rect 25329 19873 25363 19907
rect 25363 19873 25372 19907
rect 27436 19932 27488 19984
rect 28264 19932 28316 19984
rect 29184 19932 29236 19984
rect 30748 20009 30757 20043
rect 30757 20009 30791 20043
rect 30791 20009 30800 20043
rect 30748 20000 30800 20009
rect 31576 20000 31628 20052
rect 31944 20000 31996 20052
rect 32496 20000 32548 20052
rect 33416 20043 33468 20052
rect 33416 20009 33425 20043
rect 33425 20009 33459 20043
rect 33459 20009 33468 20043
rect 33416 20000 33468 20009
rect 34060 20000 34112 20052
rect 40960 20043 41012 20052
rect 40960 20009 40969 20043
rect 40969 20009 41003 20043
rect 41003 20009 41012 20043
rect 40960 20000 41012 20009
rect 41420 20000 41472 20052
rect 31116 19932 31168 19984
rect 25320 19864 25372 19873
rect 27252 19864 27304 19916
rect 4620 19796 4672 19848
rect 5540 19796 5592 19848
rect 6552 19728 6604 19780
rect 7564 19796 7616 19848
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 16948 19796 17000 19848
rect 10232 19728 10284 19780
rect 18604 19796 18656 19848
rect 18972 19796 19024 19848
rect 22652 19796 22704 19848
rect 28080 19907 28132 19916
rect 28080 19873 28089 19907
rect 28089 19873 28123 19907
rect 28123 19873 28132 19907
rect 28080 19864 28132 19873
rect 28540 19864 28592 19916
rect 29460 19907 29512 19916
rect 29460 19873 29466 19907
rect 29466 19873 29512 19907
rect 29460 19864 29512 19873
rect 31024 19864 31076 19916
rect 31300 19864 31352 19916
rect 33600 19932 33652 19984
rect 36268 19975 36320 19984
rect 36268 19941 36277 19975
rect 36277 19941 36311 19975
rect 36311 19941 36320 19975
rect 36268 19932 36320 19941
rect 37280 19932 37332 19984
rect 37832 19975 37884 19984
rect 37832 19941 37841 19975
rect 37841 19941 37875 19975
rect 37875 19941 37884 19975
rect 37832 19932 37884 19941
rect 37924 19975 37976 19984
rect 37924 19941 37933 19975
rect 37933 19941 37967 19975
rect 37967 19941 37976 19975
rect 37924 19932 37976 19941
rect 39212 19932 39264 19984
rect 41788 19975 41840 19984
rect 39304 19907 39356 19916
rect 39304 19873 39313 19907
rect 39313 19873 39347 19907
rect 39347 19873 39356 19907
rect 39304 19864 39356 19873
rect 41788 19941 41797 19975
rect 41797 19941 41831 19975
rect 41831 19941 41840 19975
rect 41788 19932 41840 19941
rect 43720 20000 43772 20052
rect 45008 20000 45060 20052
rect 43628 19975 43680 19984
rect 43628 19941 43637 19975
rect 43637 19941 43671 19975
rect 43671 19941 43680 19975
rect 43628 19932 43680 19941
rect 44456 19932 44508 19984
rect 45008 19907 45060 19916
rect 45008 19873 45017 19907
rect 45017 19873 45051 19907
rect 45051 19873 45060 19907
rect 45008 19864 45060 19873
rect 17868 19728 17920 19780
rect 28448 19796 28500 19848
rect 28816 19796 28868 19848
rect 29736 19796 29788 19848
rect 32220 19839 32272 19848
rect 32220 19805 32229 19839
rect 32229 19805 32263 19839
rect 32263 19805 32272 19839
rect 32220 19796 32272 19805
rect 34796 19796 34848 19848
rect 35624 19796 35676 19848
rect 36176 19839 36228 19848
rect 36176 19805 36185 19839
rect 36185 19805 36219 19839
rect 36219 19805 36228 19839
rect 36176 19796 36228 19805
rect 36820 19839 36872 19848
rect 36820 19805 36829 19839
rect 36829 19805 36863 19839
rect 36863 19805 36872 19839
rect 36820 19796 36872 19805
rect 37464 19796 37516 19848
rect 41512 19796 41564 19848
rect 41972 19839 42024 19848
rect 33232 19728 33284 19780
rect 33784 19728 33836 19780
rect 4068 19660 4120 19712
rect 4804 19660 4856 19712
rect 5264 19703 5316 19712
rect 5264 19669 5273 19703
rect 5273 19669 5307 19703
rect 5307 19669 5316 19703
rect 5264 19660 5316 19669
rect 6368 19703 6420 19712
rect 6368 19669 6377 19703
rect 6377 19669 6411 19703
rect 6411 19669 6420 19703
rect 6368 19660 6420 19669
rect 8852 19660 8904 19712
rect 10508 19660 10560 19712
rect 12440 19660 12492 19712
rect 19708 19703 19760 19712
rect 19708 19669 19717 19703
rect 19717 19669 19751 19703
rect 19751 19669 19760 19703
rect 19708 19660 19760 19669
rect 21180 19703 21232 19712
rect 21180 19669 21189 19703
rect 21189 19669 21223 19703
rect 21223 19669 21232 19703
rect 21180 19660 21232 19669
rect 24308 19703 24360 19712
rect 24308 19669 24317 19703
rect 24317 19669 24351 19703
rect 24351 19669 24360 19703
rect 24308 19660 24360 19669
rect 25412 19660 25464 19712
rect 26884 19703 26936 19712
rect 26884 19669 26893 19703
rect 26893 19669 26927 19703
rect 26927 19669 26936 19703
rect 26884 19660 26936 19669
rect 29092 19703 29144 19712
rect 29092 19669 29101 19703
rect 29101 19669 29135 19703
rect 29135 19669 29144 19703
rect 29092 19660 29144 19669
rect 29368 19660 29420 19712
rect 30748 19660 30800 19712
rect 34428 19660 34480 19712
rect 36176 19660 36228 19712
rect 41972 19805 41981 19839
rect 41981 19805 42015 19839
rect 42015 19805 42024 19839
rect 41972 19796 42024 19805
rect 42892 19796 42944 19848
rect 43812 19839 43864 19848
rect 43812 19805 43821 19839
rect 43821 19805 43855 19839
rect 43855 19805 43864 19839
rect 43812 19796 43864 19805
rect 42064 19728 42116 19780
rect 40500 19703 40552 19712
rect 40500 19669 40509 19703
rect 40509 19669 40543 19703
rect 40543 19669 40552 19703
rect 40500 19660 40552 19669
rect 40592 19660 40644 19712
rect 41880 19660 41932 19712
rect 44548 19660 44600 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 3792 19499 3844 19508
rect 3792 19465 3801 19499
rect 3801 19465 3835 19499
rect 3835 19465 3844 19499
rect 3792 19456 3844 19465
rect 5172 19456 5224 19508
rect 5540 19499 5592 19508
rect 5540 19465 5549 19499
rect 5549 19465 5583 19499
rect 5583 19465 5592 19499
rect 5540 19456 5592 19465
rect 7012 19456 7064 19508
rect 7932 19499 7984 19508
rect 7932 19465 7941 19499
rect 7941 19465 7975 19499
rect 7975 19465 7984 19499
rect 7932 19456 7984 19465
rect 9680 19499 9732 19508
rect 9680 19465 9689 19499
rect 9689 19465 9723 19499
rect 9723 19465 9732 19499
rect 9680 19456 9732 19465
rect 12348 19456 12400 19508
rect 13360 19456 13412 19508
rect 14004 19456 14056 19508
rect 15476 19456 15528 19508
rect 16580 19499 16632 19508
rect 16580 19465 16589 19499
rect 16589 19465 16623 19499
rect 16623 19465 16632 19499
rect 16580 19456 16632 19465
rect 18052 19456 18104 19508
rect 18236 19456 18288 19508
rect 20996 19456 21048 19508
rect 21180 19456 21232 19508
rect 22652 19456 22704 19508
rect 27252 19456 27304 19508
rect 28264 19456 28316 19508
rect 29368 19456 29420 19508
rect 29460 19456 29512 19508
rect 29644 19499 29696 19508
rect 29644 19465 29653 19499
rect 29653 19465 29687 19499
rect 29687 19465 29696 19499
rect 29644 19456 29696 19465
rect 30932 19456 30984 19508
rect 32956 19456 33008 19508
rect 33600 19499 33652 19508
rect 33600 19465 33609 19499
rect 33609 19465 33643 19499
rect 33643 19465 33652 19499
rect 33600 19456 33652 19465
rect 36268 19499 36320 19508
rect 36268 19465 36277 19499
rect 36277 19465 36311 19499
rect 36311 19465 36320 19499
rect 36268 19456 36320 19465
rect 4712 19388 4764 19440
rect 6736 19388 6788 19440
rect 11888 19431 11940 19440
rect 11888 19397 11897 19431
rect 11897 19397 11931 19431
rect 11931 19397 11940 19431
rect 11888 19388 11940 19397
rect 15568 19388 15620 19440
rect 16120 19388 16172 19440
rect 2964 19320 3016 19372
rect 8852 19363 8904 19372
rect 8852 19329 8861 19363
rect 8861 19329 8895 19363
rect 8895 19329 8904 19363
rect 8852 19320 8904 19329
rect 12716 19320 12768 19372
rect 2872 19252 2924 19304
rect 4344 19295 4396 19304
rect 4344 19261 4353 19295
rect 4353 19261 4387 19295
rect 4387 19261 4396 19295
rect 4344 19252 4396 19261
rect 9588 19252 9640 19304
rect 9956 19295 10008 19304
rect 9956 19261 9965 19295
rect 9965 19261 9999 19295
rect 9999 19261 10008 19295
rect 9956 19252 10008 19261
rect 10508 19295 10560 19304
rect 10508 19261 10517 19295
rect 10517 19261 10551 19295
rect 10551 19261 10560 19295
rect 10508 19252 10560 19261
rect 11612 19252 11664 19304
rect 6368 19184 6420 19236
rect 7012 19227 7064 19236
rect 7012 19193 7021 19227
rect 7021 19193 7055 19227
rect 7055 19193 7064 19227
rect 7564 19227 7616 19236
rect 7012 19184 7064 19193
rect 7564 19193 7573 19227
rect 7573 19193 7607 19227
rect 7607 19193 7616 19227
rect 7564 19184 7616 19193
rect 8300 19184 8352 19236
rect 4712 19159 4764 19168
rect 4712 19125 4721 19159
rect 4721 19125 4755 19159
rect 4755 19125 4764 19159
rect 4712 19116 4764 19125
rect 5448 19116 5500 19168
rect 9404 19184 9456 19236
rect 10692 19227 10744 19236
rect 10692 19193 10701 19227
rect 10701 19193 10735 19227
rect 10735 19193 10744 19227
rect 10692 19184 10744 19193
rect 11060 19159 11112 19168
rect 11060 19125 11069 19159
rect 11069 19125 11103 19159
rect 11103 19125 11112 19159
rect 11060 19116 11112 19125
rect 12256 19184 12308 19236
rect 14096 19227 14148 19236
rect 14096 19193 14105 19227
rect 14105 19193 14139 19227
rect 14139 19193 14148 19227
rect 14096 19184 14148 19193
rect 14004 19116 14056 19168
rect 18972 19388 19024 19440
rect 18788 19363 18840 19372
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 19708 19363 19760 19372
rect 18788 19320 18840 19329
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 20352 19363 20404 19372
rect 20352 19329 20361 19363
rect 20361 19329 20395 19363
rect 20395 19329 20404 19363
rect 20352 19320 20404 19329
rect 21364 19320 21416 19372
rect 21548 19363 21600 19372
rect 21548 19329 21557 19363
rect 21557 19329 21591 19363
rect 21591 19329 21600 19363
rect 21548 19320 21600 19329
rect 24216 19320 24268 19372
rect 26792 19388 26844 19440
rect 30656 19388 30708 19440
rect 32128 19388 32180 19440
rect 37648 19456 37700 19508
rect 37832 19456 37884 19508
rect 39304 19456 39356 19508
rect 41788 19499 41840 19508
rect 41788 19465 41797 19499
rect 41797 19465 41831 19499
rect 41831 19465 41840 19499
rect 41788 19456 41840 19465
rect 43536 19456 43588 19508
rect 43720 19499 43772 19508
rect 43720 19465 43729 19499
rect 43729 19465 43763 19499
rect 43763 19465 43772 19499
rect 43720 19456 43772 19465
rect 36820 19388 36872 19440
rect 37924 19431 37976 19440
rect 37924 19397 37933 19431
rect 37933 19397 37967 19431
rect 37967 19397 37976 19431
rect 37924 19388 37976 19397
rect 29736 19363 29788 19372
rect 29736 19329 29745 19363
rect 29745 19329 29779 19363
rect 29779 19329 29788 19363
rect 29736 19320 29788 19329
rect 32312 19320 32364 19372
rect 40500 19363 40552 19372
rect 40500 19329 40509 19363
rect 40509 19329 40543 19363
rect 40543 19329 40552 19363
rect 40500 19320 40552 19329
rect 41512 19320 41564 19372
rect 42432 19363 42484 19372
rect 42432 19329 42441 19363
rect 42441 19329 42475 19363
rect 42475 19329 42484 19363
rect 42432 19320 42484 19329
rect 15752 19227 15804 19236
rect 15752 19193 15761 19227
rect 15761 19193 15795 19227
rect 15795 19193 15804 19227
rect 15752 19184 15804 19193
rect 18144 19227 18196 19236
rect 18144 19193 18153 19227
rect 18153 19193 18187 19227
rect 18187 19193 18196 19227
rect 18144 19184 18196 19193
rect 18236 19227 18288 19236
rect 18236 19193 18245 19227
rect 18245 19193 18279 19227
rect 18279 19193 18288 19227
rect 18236 19184 18288 19193
rect 21180 19116 21232 19168
rect 27528 19295 27580 19304
rect 27528 19261 27537 19295
rect 27537 19261 27571 19295
rect 27571 19261 27580 19295
rect 27528 19252 27580 19261
rect 27712 19252 27764 19304
rect 29092 19252 29144 19304
rect 30932 19295 30984 19304
rect 30932 19261 30976 19295
rect 30976 19261 30984 19295
rect 31944 19295 31996 19304
rect 30932 19252 30984 19261
rect 31944 19261 31953 19295
rect 31953 19261 31987 19295
rect 31987 19261 31996 19295
rect 31944 19252 31996 19261
rect 32956 19252 33008 19304
rect 34428 19252 34480 19304
rect 37556 19252 37608 19304
rect 39212 19252 39264 19304
rect 26148 19227 26200 19236
rect 26148 19193 26157 19227
rect 26157 19193 26191 19227
rect 26191 19193 26200 19227
rect 26148 19184 26200 19193
rect 30104 19227 30156 19236
rect 30104 19193 30113 19227
rect 30113 19193 30147 19227
rect 30147 19193 30156 19227
rect 30104 19184 30156 19193
rect 32036 19184 32088 19236
rect 32496 19184 32548 19236
rect 35348 19184 35400 19236
rect 36912 19227 36964 19236
rect 36912 19193 36921 19227
rect 36921 19193 36955 19227
rect 36955 19193 36964 19227
rect 36912 19184 36964 19193
rect 23112 19159 23164 19168
rect 23112 19125 23121 19159
rect 23121 19125 23155 19159
rect 23155 19125 23164 19159
rect 23112 19116 23164 19125
rect 24400 19159 24452 19168
rect 24400 19125 24409 19159
rect 24409 19125 24443 19159
rect 24443 19125 24452 19159
rect 24400 19116 24452 19125
rect 25320 19116 25372 19168
rect 26424 19159 26476 19168
rect 26424 19125 26433 19159
rect 26433 19125 26467 19159
rect 26467 19125 26476 19159
rect 26424 19116 26476 19125
rect 27528 19116 27580 19168
rect 27988 19159 28040 19168
rect 27988 19125 27997 19159
rect 27997 19125 28031 19159
rect 28031 19125 28040 19159
rect 27988 19116 28040 19125
rect 28448 19159 28500 19168
rect 28448 19125 28457 19159
rect 28457 19125 28491 19159
rect 28491 19125 28500 19159
rect 28448 19116 28500 19125
rect 31300 19116 31352 19168
rect 31392 19159 31444 19168
rect 31392 19125 31401 19159
rect 31401 19125 31435 19159
rect 31435 19125 31444 19159
rect 31392 19116 31444 19125
rect 32404 19116 32456 19168
rect 33324 19116 33376 19168
rect 36636 19159 36688 19168
rect 36636 19125 36645 19159
rect 36645 19125 36679 19159
rect 36679 19125 36688 19159
rect 40316 19159 40368 19168
rect 36636 19116 36688 19125
rect 40316 19125 40325 19159
rect 40325 19125 40359 19159
rect 40359 19125 40368 19159
rect 40316 19116 40368 19125
rect 43444 19116 43496 19168
rect 43996 19116 44048 19168
rect 45008 19159 45060 19168
rect 45008 19125 45017 19159
rect 45017 19125 45051 19159
rect 45051 19125 45060 19159
rect 45008 19116 45060 19125
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 2872 18955 2924 18964
rect 2872 18921 2881 18955
rect 2881 18921 2915 18955
rect 2915 18921 2924 18955
rect 2872 18912 2924 18921
rect 4344 18912 4396 18964
rect 6552 18955 6604 18964
rect 6552 18921 6561 18955
rect 6561 18921 6595 18955
rect 6595 18921 6604 18955
rect 6552 18912 6604 18921
rect 7104 18912 7156 18964
rect 9956 18955 10008 18964
rect 9956 18921 9965 18955
rect 9965 18921 9999 18955
rect 9999 18921 10008 18955
rect 9956 18912 10008 18921
rect 10876 18955 10928 18964
rect 10876 18921 10885 18955
rect 10885 18921 10919 18955
rect 10919 18921 10928 18955
rect 10876 18912 10928 18921
rect 12256 18912 12308 18964
rect 13544 18955 13596 18964
rect 13544 18921 13553 18955
rect 13553 18921 13587 18955
rect 13587 18921 13596 18955
rect 13544 18912 13596 18921
rect 14096 18955 14148 18964
rect 14096 18921 14105 18955
rect 14105 18921 14139 18955
rect 14139 18921 14148 18955
rect 14096 18912 14148 18921
rect 14372 18955 14424 18964
rect 14372 18921 14381 18955
rect 14381 18921 14415 18955
rect 14415 18921 14424 18955
rect 14372 18912 14424 18921
rect 17960 18912 18012 18964
rect 18144 18955 18196 18964
rect 18144 18921 18153 18955
rect 18153 18921 18187 18955
rect 18187 18921 18196 18955
rect 18144 18912 18196 18921
rect 18604 18912 18656 18964
rect 20996 18912 21048 18964
rect 21364 18955 21416 18964
rect 21364 18921 21373 18955
rect 21373 18921 21407 18955
rect 21407 18921 21416 18955
rect 21364 18912 21416 18921
rect 27620 18912 27672 18964
rect 29276 18955 29328 18964
rect 13268 18844 13320 18896
rect 14004 18844 14056 18896
rect 15752 18844 15804 18896
rect 17224 18887 17276 18896
rect 17224 18853 17233 18887
rect 17233 18853 17267 18887
rect 17267 18853 17276 18887
rect 17224 18844 17276 18853
rect 17316 18887 17368 18896
rect 17316 18853 17325 18887
rect 17325 18853 17359 18887
rect 17359 18853 17368 18887
rect 17868 18887 17920 18896
rect 17316 18844 17368 18853
rect 17868 18853 17877 18887
rect 17877 18853 17911 18887
rect 17911 18853 17920 18887
rect 19340 18887 19392 18896
rect 17868 18844 17920 18853
rect 19340 18853 19349 18887
rect 19349 18853 19383 18887
rect 19383 18853 19392 18887
rect 19340 18844 19392 18853
rect 19432 18887 19484 18896
rect 19432 18853 19441 18887
rect 19441 18853 19475 18887
rect 19475 18853 19484 18887
rect 19432 18844 19484 18853
rect 20536 18844 20588 18896
rect 21548 18844 21600 18896
rect 23020 18887 23072 18896
rect 23020 18853 23029 18887
rect 23029 18853 23063 18887
rect 23063 18853 23072 18887
rect 23020 18844 23072 18853
rect 29276 18921 29285 18955
rect 29285 18921 29319 18955
rect 29319 18921 29328 18955
rect 29276 18912 29328 18921
rect 29644 18912 29696 18964
rect 31576 18955 31628 18964
rect 31576 18921 31585 18955
rect 31585 18921 31619 18955
rect 31619 18921 31628 18955
rect 31576 18912 31628 18921
rect 32220 18955 32272 18964
rect 32220 18921 32229 18955
rect 32229 18921 32263 18955
rect 32263 18921 32272 18955
rect 32220 18912 32272 18921
rect 33600 18912 33652 18964
rect 34796 18955 34848 18964
rect 28908 18844 28960 18896
rect 4712 18776 4764 18828
rect 5080 18776 5132 18828
rect 5724 18819 5776 18828
rect 5724 18785 5733 18819
rect 5733 18785 5767 18819
rect 5767 18785 5776 18819
rect 5724 18776 5776 18785
rect 8576 18819 8628 18828
rect 8576 18785 8620 18819
rect 8620 18785 8628 18819
rect 8576 18776 8628 18785
rect 11060 18776 11112 18828
rect 14372 18776 14424 18828
rect 16764 18776 16816 18828
rect 21732 18776 21784 18828
rect 7380 18708 7432 18760
rect 10416 18708 10468 18760
rect 10692 18708 10744 18760
rect 13452 18708 13504 18760
rect 23664 18776 23716 18828
rect 25412 18819 25464 18828
rect 25412 18785 25421 18819
rect 25421 18785 25455 18819
rect 25455 18785 25464 18819
rect 25412 18776 25464 18785
rect 26608 18819 26660 18828
rect 26608 18785 26617 18819
rect 26617 18785 26651 18819
rect 26651 18785 26660 18819
rect 26608 18776 26660 18785
rect 23020 18708 23072 18760
rect 24216 18751 24268 18760
rect 24216 18717 24225 18751
rect 24225 18717 24259 18751
rect 24259 18717 24268 18751
rect 24216 18708 24268 18717
rect 26976 18751 27028 18760
rect 26976 18717 26985 18751
rect 26985 18717 27019 18751
rect 27019 18717 27028 18751
rect 26976 18708 27028 18717
rect 28632 18776 28684 18828
rect 30288 18776 30340 18828
rect 31116 18776 31168 18828
rect 32128 18776 32180 18828
rect 32220 18776 32272 18828
rect 32404 18819 32456 18828
rect 32404 18785 32413 18819
rect 32413 18785 32447 18819
rect 32447 18785 32456 18819
rect 32404 18776 32456 18785
rect 32588 18819 32640 18828
rect 32588 18785 32597 18819
rect 32597 18785 32631 18819
rect 32631 18785 32640 18819
rect 34796 18921 34805 18955
rect 34805 18921 34839 18955
rect 34839 18921 34848 18955
rect 34796 18912 34848 18921
rect 36636 18912 36688 18964
rect 39212 18912 39264 18964
rect 42800 18912 42852 18964
rect 34428 18887 34480 18896
rect 34428 18853 34437 18887
rect 34437 18853 34471 18887
rect 34471 18853 34480 18887
rect 34428 18844 34480 18853
rect 35348 18844 35400 18896
rect 37924 18887 37976 18896
rect 37924 18853 37933 18887
rect 37933 18853 37967 18887
rect 37967 18853 37976 18887
rect 37924 18844 37976 18853
rect 40316 18844 40368 18896
rect 42432 18887 42484 18896
rect 42432 18853 42441 18887
rect 42441 18853 42475 18887
rect 42475 18853 42484 18887
rect 42432 18844 42484 18853
rect 43536 18887 43588 18896
rect 43536 18853 43545 18887
rect 43545 18853 43579 18887
rect 43579 18853 43588 18887
rect 43536 18844 43588 18853
rect 32588 18776 32640 18785
rect 28540 18751 28592 18760
rect 28540 18717 28549 18751
rect 28549 18717 28583 18751
rect 28583 18717 28592 18751
rect 28540 18708 28592 18717
rect 32312 18708 32364 18760
rect 34704 18776 34756 18828
rect 36176 18776 36228 18828
rect 41880 18776 41932 18828
rect 12440 18640 12492 18692
rect 14096 18640 14148 18692
rect 26424 18640 26476 18692
rect 32220 18640 32272 18692
rect 37924 18708 37976 18760
rect 36912 18683 36964 18692
rect 36912 18649 36921 18683
rect 36921 18649 36955 18683
rect 36955 18649 36964 18683
rect 36912 18640 36964 18649
rect 7196 18572 7248 18624
rect 8300 18572 8352 18624
rect 8484 18572 8536 18624
rect 11244 18572 11296 18624
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16028 18572 16080 18581
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 23756 18615 23808 18624
rect 23756 18581 23765 18615
rect 23765 18581 23799 18615
rect 23799 18581 23808 18615
rect 23756 18572 23808 18581
rect 24308 18615 24360 18624
rect 24308 18581 24317 18615
rect 24317 18581 24351 18615
rect 24351 18581 24360 18615
rect 24308 18572 24360 18581
rect 25136 18572 25188 18624
rect 26884 18615 26936 18624
rect 26884 18581 26893 18615
rect 26893 18581 26927 18615
rect 26927 18581 26936 18615
rect 26884 18572 26936 18581
rect 27068 18615 27120 18624
rect 27068 18581 27077 18615
rect 27077 18581 27111 18615
rect 27111 18581 27120 18615
rect 27068 18572 27120 18581
rect 28448 18615 28500 18624
rect 28448 18581 28457 18615
rect 28457 18581 28491 18615
rect 28491 18581 28500 18615
rect 28448 18572 28500 18581
rect 29368 18572 29420 18624
rect 30196 18615 30248 18624
rect 30196 18581 30205 18615
rect 30205 18581 30239 18615
rect 30239 18581 30248 18615
rect 30196 18572 30248 18581
rect 31944 18615 31996 18624
rect 31944 18581 31953 18615
rect 31953 18581 31987 18615
rect 31987 18581 31996 18615
rect 31944 18572 31996 18581
rect 35256 18572 35308 18624
rect 39580 18572 39632 18624
rect 43260 18708 43312 18760
rect 43720 18751 43772 18760
rect 43720 18717 43729 18751
rect 43729 18717 43763 18751
rect 43763 18717 43772 18751
rect 43720 18708 43772 18717
rect 42340 18640 42392 18692
rect 40132 18572 40184 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 5080 18368 5132 18420
rect 7196 18368 7248 18420
rect 7380 18411 7432 18420
rect 7380 18377 7389 18411
rect 7389 18377 7423 18411
rect 7423 18377 7432 18411
rect 7380 18368 7432 18377
rect 9772 18368 9824 18420
rect 11244 18411 11296 18420
rect 11244 18377 11253 18411
rect 11253 18377 11287 18411
rect 11287 18377 11296 18411
rect 11244 18368 11296 18377
rect 13452 18411 13504 18420
rect 13452 18377 13461 18411
rect 13461 18377 13495 18411
rect 13495 18377 13504 18411
rect 13452 18368 13504 18377
rect 13820 18411 13872 18420
rect 13820 18377 13829 18411
rect 13829 18377 13863 18411
rect 13863 18377 13872 18411
rect 13820 18368 13872 18377
rect 14464 18368 14516 18420
rect 15936 18368 15988 18420
rect 17316 18411 17368 18420
rect 17316 18377 17325 18411
rect 17325 18377 17359 18411
rect 17359 18377 17368 18411
rect 17316 18368 17368 18377
rect 19432 18411 19484 18420
rect 19432 18377 19441 18411
rect 19441 18377 19475 18411
rect 19475 18377 19484 18411
rect 19432 18368 19484 18377
rect 21272 18368 21324 18420
rect 4620 18232 4672 18284
rect 4068 18207 4120 18216
rect 4068 18173 4077 18207
rect 4077 18173 4111 18207
rect 4111 18173 4120 18207
rect 4068 18164 4120 18173
rect 5724 18300 5776 18352
rect 6736 18300 6788 18352
rect 5448 18164 5500 18216
rect 23756 18300 23808 18352
rect 24768 18300 24820 18352
rect 8484 18232 8536 18284
rect 8852 18275 8904 18284
rect 8852 18241 8861 18275
rect 8861 18241 8895 18275
rect 8895 18241 8904 18275
rect 8852 18232 8904 18241
rect 9772 18207 9824 18216
rect 9772 18173 9781 18207
rect 9781 18173 9815 18207
rect 9815 18173 9824 18207
rect 9772 18164 9824 18173
rect 12256 18232 12308 18284
rect 10508 18164 10560 18216
rect 11244 18164 11296 18216
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 13820 18164 13872 18216
rect 14648 18164 14700 18216
rect 19432 18232 19484 18284
rect 15936 18207 15988 18216
rect 15936 18173 15945 18207
rect 15945 18173 15979 18207
rect 15979 18173 15988 18207
rect 15936 18164 15988 18173
rect 16028 18164 16080 18216
rect 21732 18275 21784 18284
rect 21732 18241 21741 18275
rect 21741 18241 21775 18275
rect 21775 18241 21784 18275
rect 21732 18232 21784 18241
rect 23480 18275 23532 18284
rect 23480 18241 23489 18275
rect 23489 18241 23523 18275
rect 23523 18241 23532 18275
rect 23480 18232 23532 18241
rect 24400 18232 24452 18284
rect 25044 18232 25096 18284
rect 26516 18368 26568 18420
rect 26884 18368 26936 18420
rect 28448 18368 28500 18420
rect 30196 18368 30248 18420
rect 30288 18368 30340 18420
rect 33508 18368 33560 18420
rect 33600 18368 33652 18420
rect 35348 18411 35400 18420
rect 25320 18300 25372 18352
rect 29552 18343 29604 18352
rect 10416 18139 10468 18148
rect 10416 18105 10425 18139
rect 10425 18105 10459 18139
rect 10459 18105 10468 18139
rect 10416 18096 10468 18105
rect 13176 18139 13228 18148
rect 13176 18105 13185 18139
rect 13185 18105 13219 18139
rect 13219 18105 13228 18139
rect 13176 18096 13228 18105
rect 15292 18096 15344 18148
rect 18236 18096 18288 18148
rect 20628 18139 20680 18148
rect 20628 18105 20637 18139
rect 20637 18105 20671 18139
rect 20671 18105 20680 18139
rect 20628 18096 20680 18105
rect 7104 18071 7156 18080
rect 7104 18037 7113 18071
rect 7113 18037 7147 18071
rect 7147 18037 7156 18071
rect 7104 18028 7156 18037
rect 10324 18028 10376 18080
rect 10876 18028 10928 18080
rect 14372 18028 14424 18080
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 16212 18028 16264 18037
rect 16764 18028 16816 18080
rect 17868 18028 17920 18080
rect 18512 18028 18564 18080
rect 20444 18071 20496 18080
rect 20444 18037 20453 18071
rect 20453 18037 20487 18071
rect 20487 18037 20496 18071
rect 25228 18207 25280 18216
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 23664 18139 23716 18148
rect 23664 18105 23673 18139
rect 23673 18105 23707 18139
rect 23707 18105 23716 18139
rect 23664 18096 23716 18105
rect 25136 18096 25188 18148
rect 22008 18071 22060 18080
rect 20444 18028 20496 18037
rect 22008 18037 22017 18071
rect 22017 18037 22051 18071
rect 22051 18037 22060 18071
rect 22008 18028 22060 18037
rect 22100 18028 22152 18080
rect 23020 18028 23072 18080
rect 23204 18028 23256 18080
rect 24768 18071 24820 18080
rect 24768 18037 24777 18071
rect 24777 18037 24811 18071
rect 24811 18037 24820 18071
rect 24768 18028 24820 18037
rect 25044 18071 25096 18080
rect 25044 18037 25053 18071
rect 25053 18037 25087 18071
rect 25087 18037 25096 18071
rect 26976 18232 27028 18284
rect 27988 18275 28040 18284
rect 27988 18241 27997 18275
rect 27997 18241 28031 18275
rect 28031 18241 28040 18275
rect 27988 18232 28040 18241
rect 28540 18232 28592 18284
rect 29552 18309 29561 18343
rect 29561 18309 29595 18343
rect 29595 18309 29604 18343
rect 29552 18300 29604 18309
rect 31116 18343 31168 18352
rect 31116 18309 31125 18343
rect 31125 18309 31159 18343
rect 31159 18309 31168 18343
rect 31116 18300 31168 18309
rect 34060 18300 34112 18352
rect 35348 18377 35357 18411
rect 35357 18377 35391 18411
rect 35391 18377 35400 18411
rect 35348 18368 35400 18377
rect 37832 18368 37884 18420
rect 38108 18368 38160 18420
rect 39304 18368 39356 18420
rect 41880 18368 41932 18420
rect 40040 18300 40092 18352
rect 43536 18368 43588 18420
rect 43260 18300 43312 18352
rect 29920 18232 29972 18284
rect 31944 18275 31996 18284
rect 27160 18164 27212 18216
rect 28632 18164 28684 18216
rect 29276 18207 29328 18216
rect 29276 18173 29285 18207
rect 29285 18173 29319 18207
rect 29319 18173 29328 18207
rect 31944 18241 31953 18275
rect 31953 18241 31987 18275
rect 31987 18241 31996 18275
rect 31944 18232 31996 18241
rect 33048 18232 33100 18284
rect 34152 18232 34204 18284
rect 39580 18275 39632 18284
rect 39580 18241 39589 18275
rect 39589 18241 39623 18275
rect 39623 18241 39632 18275
rect 39580 18232 39632 18241
rect 42340 18232 42392 18284
rect 42800 18232 42852 18284
rect 29276 18164 29328 18173
rect 31484 18164 31536 18216
rect 31852 18207 31904 18216
rect 31852 18173 31861 18207
rect 31861 18173 31895 18207
rect 31895 18173 31904 18207
rect 31852 18164 31904 18173
rect 26700 18096 26752 18148
rect 27620 18139 27672 18148
rect 27620 18105 27629 18139
rect 27629 18105 27663 18139
rect 27663 18105 27672 18139
rect 27620 18096 27672 18105
rect 29184 18096 29236 18148
rect 25872 18071 25924 18080
rect 25044 18028 25096 18037
rect 25872 18037 25881 18071
rect 25881 18037 25915 18071
rect 25915 18037 25924 18071
rect 25872 18028 25924 18037
rect 26240 18028 26292 18080
rect 26976 18028 27028 18080
rect 27896 18028 27948 18080
rect 31116 18096 31168 18148
rect 32680 18096 32732 18148
rect 33048 18139 33100 18148
rect 33048 18105 33057 18139
rect 33057 18105 33091 18139
rect 33091 18105 33100 18139
rect 33048 18096 33100 18105
rect 35348 18096 35400 18148
rect 35808 18096 35860 18148
rect 29920 18071 29972 18080
rect 29920 18037 29929 18071
rect 29929 18037 29963 18071
rect 29963 18037 29972 18071
rect 29920 18028 29972 18037
rect 30288 18071 30340 18080
rect 30288 18037 30297 18071
rect 30297 18037 30331 18071
rect 30331 18037 30340 18071
rect 30288 18028 30340 18037
rect 32404 18028 32456 18080
rect 32772 18028 32824 18080
rect 34704 18071 34756 18080
rect 34704 18037 34713 18071
rect 34713 18037 34747 18071
rect 34747 18037 34756 18071
rect 34704 18028 34756 18037
rect 38660 18164 38712 18216
rect 39028 18164 39080 18216
rect 39212 18164 39264 18216
rect 40500 18207 40552 18216
rect 40500 18173 40509 18207
rect 40509 18173 40543 18207
rect 40543 18173 40552 18207
rect 40500 18164 40552 18173
rect 37924 18096 37976 18148
rect 42340 18139 42392 18148
rect 37648 18028 37700 18080
rect 38476 18028 38528 18080
rect 38660 18071 38712 18080
rect 38660 18037 38669 18071
rect 38669 18037 38703 18071
rect 38703 18037 38712 18071
rect 38660 18028 38712 18037
rect 39672 18028 39724 18080
rect 40316 18028 40368 18080
rect 42340 18105 42349 18139
rect 42349 18105 42383 18139
rect 42383 18105 42392 18139
rect 42340 18096 42392 18105
rect 42432 18139 42484 18148
rect 42432 18105 42441 18139
rect 42441 18105 42475 18139
rect 42475 18105 42484 18139
rect 42432 18096 42484 18105
rect 42064 18028 42116 18080
rect 43720 18232 43772 18284
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 2872 17824 2924 17876
rect 4068 17824 4120 17876
rect 6368 17824 6420 17876
rect 8484 17824 8536 17876
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 9772 17867 9824 17876
rect 8576 17824 8628 17833
rect 9772 17833 9781 17867
rect 9781 17833 9815 17867
rect 9815 17833 9824 17867
rect 9772 17824 9824 17833
rect 10416 17824 10468 17876
rect 11796 17867 11848 17876
rect 11796 17833 11805 17867
rect 11805 17833 11839 17867
rect 11839 17833 11848 17867
rect 11796 17824 11848 17833
rect 14648 17867 14700 17876
rect 14648 17833 14657 17867
rect 14657 17833 14691 17867
rect 14691 17833 14700 17867
rect 14648 17824 14700 17833
rect 15660 17867 15712 17876
rect 15660 17833 15669 17867
rect 15669 17833 15703 17867
rect 15703 17833 15712 17867
rect 15660 17824 15712 17833
rect 17224 17824 17276 17876
rect 17684 17824 17736 17876
rect 19340 17867 19392 17876
rect 19340 17833 19349 17867
rect 19349 17833 19383 17867
rect 19383 17833 19392 17867
rect 19340 17824 19392 17833
rect 3792 17688 3844 17740
rect 4620 17731 4672 17740
rect 4620 17697 4629 17731
rect 4629 17697 4663 17731
rect 4663 17697 4672 17731
rect 4620 17688 4672 17697
rect 5264 17688 5316 17740
rect 7748 17756 7800 17808
rect 12808 17756 12860 17808
rect 7564 17731 7616 17740
rect 7564 17697 7573 17731
rect 7573 17697 7607 17731
rect 7607 17697 7616 17731
rect 7564 17688 7616 17697
rect 9956 17731 10008 17740
rect 9956 17697 9965 17731
rect 9965 17697 9999 17731
rect 9999 17697 10008 17731
rect 9956 17688 10008 17697
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 11980 17731 12032 17740
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 12164 17731 12216 17740
rect 12164 17697 12173 17731
rect 12173 17697 12207 17731
rect 12207 17697 12216 17731
rect 12164 17688 12216 17697
rect 12900 17688 12952 17740
rect 13544 17731 13596 17740
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 14188 17688 14240 17740
rect 18880 17756 18932 17808
rect 25136 17824 25188 17876
rect 25320 17867 25372 17876
rect 25320 17833 25329 17867
rect 25329 17833 25363 17867
rect 25363 17833 25372 17867
rect 25320 17824 25372 17833
rect 25412 17824 25464 17876
rect 28448 17824 28500 17876
rect 21088 17799 21140 17808
rect 21088 17765 21097 17799
rect 21097 17765 21131 17799
rect 21131 17765 21140 17799
rect 21088 17756 21140 17765
rect 16856 17688 16908 17740
rect 17868 17688 17920 17740
rect 17960 17688 18012 17740
rect 18512 17688 18564 17740
rect 19432 17731 19484 17740
rect 19432 17697 19441 17731
rect 19441 17697 19475 17731
rect 19475 17697 19484 17731
rect 19432 17688 19484 17697
rect 19616 17731 19668 17740
rect 19616 17697 19625 17731
rect 19625 17697 19659 17731
rect 19659 17697 19668 17731
rect 19616 17688 19668 17697
rect 23204 17756 23256 17808
rect 24768 17756 24820 17808
rect 27160 17756 27212 17808
rect 29552 17824 29604 17876
rect 31024 17867 31076 17876
rect 31024 17833 31033 17867
rect 31033 17833 31067 17867
rect 31067 17833 31076 17867
rect 31024 17824 31076 17833
rect 31484 17867 31536 17876
rect 31484 17833 31493 17867
rect 31493 17833 31527 17867
rect 31527 17833 31536 17867
rect 31484 17824 31536 17833
rect 31852 17867 31904 17876
rect 31852 17833 31861 17867
rect 31861 17833 31895 17867
rect 31895 17833 31904 17867
rect 31852 17824 31904 17833
rect 32588 17824 32640 17876
rect 35256 17824 35308 17876
rect 35808 17824 35860 17876
rect 37924 17867 37976 17876
rect 37924 17833 37933 17867
rect 37933 17833 37967 17867
rect 37967 17833 37976 17867
rect 37924 17824 37976 17833
rect 28908 17756 28960 17808
rect 25228 17688 25280 17740
rect 26148 17688 26200 17740
rect 26516 17731 26568 17740
rect 26516 17697 26525 17731
rect 26525 17697 26559 17731
rect 26559 17697 26568 17731
rect 26516 17688 26568 17697
rect 26792 17688 26844 17740
rect 27896 17688 27948 17740
rect 29644 17731 29696 17740
rect 29644 17697 29653 17731
rect 29653 17697 29687 17731
rect 29687 17697 29696 17731
rect 29644 17688 29696 17697
rect 30012 17731 30064 17740
rect 30012 17697 30021 17731
rect 30021 17697 30055 17731
rect 30055 17697 30064 17731
rect 30012 17688 30064 17697
rect 32312 17731 32364 17740
rect 32312 17697 32321 17731
rect 32321 17697 32355 17731
rect 32355 17697 32364 17731
rect 32312 17688 32364 17697
rect 34704 17756 34756 17808
rect 40132 17824 40184 17876
rect 40500 17824 40552 17876
rect 42340 17824 42392 17876
rect 33416 17688 33468 17740
rect 33784 17731 33836 17740
rect 7748 17663 7800 17672
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 7748 17620 7800 17629
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 20352 17620 20404 17672
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 21180 17620 21232 17672
rect 24032 17663 24084 17672
rect 24032 17629 24041 17663
rect 24041 17629 24075 17663
rect 24075 17629 24084 17663
rect 24032 17620 24084 17629
rect 30104 17620 30156 17672
rect 33784 17697 33793 17731
rect 33793 17697 33827 17731
rect 33827 17697 33836 17731
rect 33784 17688 33836 17697
rect 39212 17756 39264 17808
rect 36268 17688 36320 17740
rect 38384 17688 38436 17740
rect 38844 17688 38896 17740
rect 39488 17688 39540 17740
rect 40040 17688 40092 17740
rect 41972 17688 42024 17740
rect 42432 17688 42484 17740
rect 12716 17552 12768 17604
rect 18236 17552 18288 17604
rect 19340 17552 19392 17604
rect 26608 17552 26660 17604
rect 30932 17552 30984 17604
rect 35256 17620 35308 17672
rect 35348 17620 35400 17672
rect 37556 17620 37608 17672
rect 42064 17620 42116 17672
rect 14648 17484 14700 17536
rect 18144 17484 18196 17536
rect 22008 17484 22060 17536
rect 23204 17484 23256 17536
rect 23940 17527 23992 17536
rect 23940 17493 23949 17527
rect 23949 17493 23983 17527
rect 23983 17493 23992 17527
rect 23940 17484 23992 17493
rect 32496 17527 32548 17536
rect 32496 17493 32505 17527
rect 32505 17493 32539 17527
rect 32539 17493 32548 17527
rect 32496 17484 32548 17493
rect 38384 17552 38436 17604
rect 34336 17484 34388 17536
rect 36728 17484 36780 17536
rect 36912 17527 36964 17536
rect 36912 17493 36921 17527
rect 36921 17493 36955 17527
rect 36955 17493 36964 17527
rect 36912 17484 36964 17493
rect 37372 17484 37424 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 2964 17280 3016 17332
rect 3792 17280 3844 17332
rect 3976 17323 4028 17332
rect 3976 17289 3985 17323
rect 3985 17289 4019 17323
rect 4019 17289 4028 17323
rect 3976 17280 4028 17289
rect 5264 17280 5316 17332
rect 7840 17280 7892 17332
rect 9956 17280 10008 17332
rect 12164 17280 12216 17332
rect 13544 17323 13596 17332
rect 13544 17289 13553 17323
rect 13553 17289 13587 17323
rect 13587 17289 13596 17323
rect 13544 17280 13596 17289
rect 14188 17323 14240 17332
rect 14188 17289 14197 17323
rect 14197 17289 14231 17323
rect 14231 17289 14240 17323
rect 14188 17280 14240 17289
rect 16212 17280 16264 17332
rect 16856 17323 16908 17332
rect 16856 17289 16865 17323
rect 16865 17289 16899 17323
rect 16899 17289 16908 17323
rect 16856 17280 16908 17289
rect 11980 17212 12032 17264
rect 3976 17076 4028 17128
rect 4620 17119 4672 17128
rect 4620 17085 4629 17119
rect 4629 17085 4663 17119
rect 4663 17085 4672 17119
rect 7656 17144 7708 17196
rect 4620 17076 4672 17085
rect 4804 17008 4856 17060
rect 3240 16983 3292 16992
rect 3240 16949 3249 16983
rect 3249 16949 3283 16983
rect 3283 16949 3292 16983
rect 3240 16940 3292 16949
rect 7564 17076 7616 17128
rect 7656 17051 7708 17060
rect 7656 17017 7665 17051
rect 7665 17017 7699 17051
rect 7699 17017 7708 17051
rect 7656 17008 7708 17017
rect 9680 17076 9732 17128
rect 10784 17119 10836 17128
rect 9404 17008 9456 17060
rect 10784 17085 10793 17119
rect 10793 17085 10827 17119
rect 10827 17085 10836 17119
rect 10784 17076 10836 17085
rect 11888 17076 11940 17128
rect 19432 17280 19484 17332
rect 21088 17280 21140 17332
rect 22744 17280 22796 17332
rect 23204 17280 23256 17332
rect 25228 17280 25280 17332
rect 26792 17280 26844 17332
rect 28632 17323 28684 17332
rect 28632 17289 28641 17323
rect 28641 17289 28675 17323
rect 28675 17289 28684 17323
rect 28632 17280 28684 17289
rect 29276 17280 29328 17332
rect 32496 17280 32548 17332
rect 33140 17280 33192 17332
rect 33784 17280 33836 17332
rect 34704 17323 34756 17332
rect 34704 17289 34713 17323
rect 34713 17289 34747 17323
rect 34747 17289 34756 17323
rect 34704 17280 34756 17289
rect 34796 17280 34848 17332
rect 35348 17280 35400 17332
rect 19156 17212 19208 17264
rect 20996 17212 21048 17264
rect 23940 17255 23992 17264
rect 23940 17221 23949 17255
rect 23949 17221 23983 17255
rect 23983 17221 23992 17255
rect 23940 17212 23992 17221
rect 24768 17212 24820 17264
rect 32312 17212 32364 17264
rect 32956 17212 33008 17264
rect 36268 17255 36320 17264
rect 36268 17221 36277 17255
rect 36277 17221 36311 17255
rect 36311 17221 36320 17255
rect 36268 17212 36320 17221
rect 36636 17212 36688 17264
rect 38200 17212 38252 17264
rect 38844 17212 38896 17264
rect 39212 17212 39264 17264
rect 40040 17212 40092 17264
rect 20536 17187 20588 17196
rect 12992 17076 13044 17128
rect 14004 17119 14056 17128
rect 10140 17008 10192 17060
rect 14004 17085 14013 17119
rect 14013 17085 14047 17119
rect 14047 17085 14056 17119
rect 14004 17076 14056 17085
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 21180 17187 21232 17196
rect 21180 17153 21189 17187
rect 21189 17153 21223 17187
rect 21223 17153 21232 17187
rect 21180 17144 21232 17153
rect 6092 16940 6144 16992
rect 9588 16983 9640 16992
rect 9588 16949 9597 16983
rect 9597 16949 9631 16983
rect 9631 16949 9640 16983
rect 9588 16940 9640 16949
rect 10876 16940 10928 16992
rect 12532 16983 12584 16992
rect 12532 16949 12541 16983
rect 12541 16949 12575 16983
rect 12575 16949 12584 16983
rect 12532 16940 12584 16949
rect 14556 16940 14608 16992
rect 15660 17008 15712 17060
rect 18236 17119 18288 17128
rect 18236 17085 18245 17119
rect 18245 17085 18279 17119
rect 18279 17085 18288 17119
rect 18236 17076 18288 17085
rect 19892 17076 19944 17128
rect 22836 17119 22888 17128
rect 22836 17085 22845 17119
rect 22845 17085 22879 17119
rect 22879 17085 22888 17119
rect 22836 17076 22888 17085
rect 24492 17119 24544 17128
rect 24492 17085 24501 17119
rect 24501 17085 24535 17119
rect 24535 17085 24544 17119
rect 24492 17076 24544 17085
rect 26240 17076 26292 17128
rect 26700 17144 26752 17196
rect 29644 17144 29696 17196
rect 30104 17187 30156 17196
rect 30104 17153 30113 17187
rect 30113 17153 30147 17187
rect 30147 17153 30156 17187
rect 30104 17144 30156 17153
rect 31944 17187 31996 17196
rect 31944 17153 31953 17187
rect 31953 17153 31987 17187
rect 31987 17153 31996 17187
rect 31944 17144 31996 17153
rect 33324 17144 33376 17196
rect 36912 17144 36964 17196
rect 38476 17187 38528 17196
rect 38476 17153 38485 17187
rect 38485 17153 38519 17187
rect 38519 17153 38528 17187
rect 38476 17144 38528 17153
rect 27160 17076 27212 17128
rect 28264 17076 28316 17128
rect 29920 17076 29972 17128
rect 32680 17076 32732 17128
rect 33232 17076 33284 17128
rect 19616 17008 19668 17060
rect 20628 17051 20680 17060
rect 20628 17017 20637 17051
rect 20637 17017 20671 17051
rect 20671 17017 20680 17051
rect 20628 17008 20680 17017
rect 24124 17008 24176 17060
rect 24308 17051 24360 17060
rect 24308 17017 24317 17051
rect 24317 17017 24351 17051
rect 24351 17017 24360 17051
rect 24308 17008 24360 17017
rect 26516 17008 26568 17060
rect 28540 17008 28592 17060
rect 16120 16983 16172 16992
rect 16120 16949 16129 16983
rect 16129 16949 16163 16983
rect 16163 16949 16172 16983
rect 16120 16940 16172 16949
rect 16212 16940 16264 16992
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 17868 16983 17920 16992
rect 17868 16949 17877 16983
rect 17877 16949 17911 16983
rect 17911 16949 17920 16983
rect 17868 16940 17920 16949
rect 18328 16983 18380 16992
rect 18328 16949 18337 16983
rect 18337 16949 18371 16983
rect 18371 16949 18380 16983
rect 18328 16940 18380 16949
rect 18512 16940 18564 16992
rect 31392 17008 31444 17060
rect 31760 17008 31812 17060
rect 32588 17051 32640 17060
rect 26424 16983 26476 16992
rect 26424 16949 26433 16983
rect 26433 16949 26467 16983
rect 26467 16949 26476 16983
rect 26424 16940 26476 16949
rect 27896 16940 27948 16992
rect 28356 16983 28408 16992
rect 28356 16949 28365 16983
rect 28365 16949 28399 16983
rect 28399 16949 28408 16983
rect 28356 16940 28408 16949
rect 29644 16983 29696 16992
rect 29644 16949 29653 16983
rect 29653 16949 29687 16983
rect 29687 16949 29696 16983
rect 29644 16940 29696 16949
rect 30288 16940 30340 16992
rect 32588 17017 32597 17051
rect 32597 17017 32631 17051
rect 32631 17017 32640 17051
rect 32588 17008 32640 17017
rect 32312 16940 32364 16992
rect 32956 16940 33008 16992
rect 41972 17280 42024 17332
rect 43536 17119 43588 17128
rect 34336 17008 34388 17060
rect 35992 17051 36044 17060
rect 35992 17017 36001 17051
rect 36001 17017 36035 17051
rect 36035 17017 36044 17051
rect 35992 17008 36044 17017
rect 36636 17051 36688 17060
rect 36636 17017 36645 17051
rect 36645 17017 36679 17051
rect 36679 17017 36688 17051
rect 36636 17008 36688 17017
rect 37188 17051 37240 17060
rect 37188 17017 37197 17051
rect 37197 17017 37231 17051
rect 37231 17017 37240 17051
rect 37188 17008 37240 17017
rect 34612 16940 34664 16992
rect 36452 16940 36504 16992
rect 38200 17051 38252 17060
rect 38200 17017 38209 17051
rect 38209 17017 38243 17051
rect 38243 17017 38252 17051
rect 38200 17008 38252 17017
rect 38568 17008 38620 17060
rect 43536 17085 43545 17119
rect 43545 17085 43579 17119
rect 43579 17085 43588 17119
rect 43536 17076 43588 17085
rect 39488 16983 39540 16992
rect 39488 16949 39497 16983
rect 39497 16949 39531 16983
rect 39531 16949 39540 16983
rect 39488 16940 39540 16949
rect 40316 16940 40368 16992
rect 40868 17008 40920 17060
rect 41144 16940 41196 16992
rect 44088 16940 44140 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 7656 16736 7708 16788
rect 9404 16779 9456 16788
rect 9404 16745 9413 16779
rect 9413 16745 9447 16779
rect 9447 16745 9456 16779
rect 9404 16736 9456 16745
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 12164 16779 12216 16788
rect 12164 16745 12173 16779
rect 12173 16745 12207 16779
rect 12207 16745 12216 16779
rect 12164 16736 12216 16745
rect 12992 16779 13044 16788
rect 12992 16745 13001 16779
rect 13001 16745 13035 16779
rect 13035 16745 13044 16779
rect 12992 16736 13044 16745
rect 7104 16668 7156 16720
rect 9496 16668 9548 16720
rect 10324 16668 10376 16720
rect 14188 16736 14240 16788
rect 15292 16736 15344 16788
rect 18236 16736 18288 16788
rect 19432 16779 19484 16788
rect 17500 16711 17552 16720
rect 17500 16677 17509 16711
rect 17509 16677 17543 16711
rect 17543 16677 17552 16711
rect 17500 16668 17552 16677
rect 19432 16745 19441 16779
rect 19441 16745 19475 16779
rect 19475 16745 19484 16779
rect 19432 16736 19484 16745
rect 20536 16779 20588 16788
rect 20536 16745 20545 16779
rect 20545 16745 20579 16779
rect 20579 16745 20588 16779
rect 20536 16736 20588 16745
rect 21088 16736 21140 16788
rect 22744 16779 22796 16788
rect 22744 16745 22753 16779
rect 22753 16745 22787 16779
rect 22787 16745 22796 16779
rect 22744 16736 22796 16745
rect 26608 16779 26660 16788
rect 26608 16745 26617 16779
rect 26617 16745 26651 16779
rect 26651 16745 26660 16779
rect 26608 16736 26660 16745
rect 27620 16779 27672 16788
rect 27620 16745 27629 16779
rect 27629 16745 27663 16779
rect 27663 16745 27672 16779
rect 27620 16736 27672 16745
rect 28264 16779 28316 16788
rect 28264 16745 28273 16779
rect 28273 16745 28307 16779
rect 28307 16745 28316 16779
rect 28264 16736 28316 16745
rect 29736 16779 29788 16788
rect 23204 16711 23256 16720
rect 23204 16677 23213 16711
rect 23213 16677 23247 16711
rect 23247 16677 23256 16711
rect 23204 16668 23256 16677
rect 26700 16668 26752 16720
rect 2688 16643 2740 16652
rect 2688 16609 2697 16643
rect 2697 16609 2731 16643
rect 2731 16609 2740 16643
rect 2688 16600 2740 16609
rect 3240 16600 3292 16652
rect 3332 16600 3384 16652
rect 3976 16600 4028 16652
rect 4620 16643 4672 16652
rect 4620 16609 4629 16643
rect 4629 16609 4663 16643
rect 4663 16609 4672 16643
rect 4620 16600 4672 16609
rect 5080 16600 5132 16652
rect 5908 16600 5960 16652
rect 6092 16643 6144 16652
rect 6092 16609 6101 16643
rect 6101 16609 6135 16643
rect 6135 16609 6144 16643
rect 6092 16600 6144 16609
rect 7564 16600 7616 16652
rect 7748 16600 7800 16652
rect 9772 16600 9824 16652
rect 11796 16643 11848 16652
rect 11796 16609 11805 16643
rect 11805 16609 11839 16643
rect 11839 16609 11848 16643
rect 11796 16600 11848 16609
rect 13820 16600 13872 16652
rect 14648 16600 14700 16652
rect 15568 16643 15620 16652
rect 15568 16609 15586 16643
rect 15586 16609 15620 16643
rect 15568 16600 15620 16609
rect 16120 16600 16172 16652
rect 18512 16643 18564 16652
rect 3148 16575 3200 16584
rect 3148 16541 3157 16575
rect 3157 16541 3191 16575
rect 3191 16541 3200 16575
rect 3148 16532 3200 16541
rect 4896 16532 4948 16584
rect 6368 16575 6420 16584
rect 6368 16541 6377 16575
rect 6377 16541 6411 16575
rect 6411 16541 6420 16575
rect 6368 16532 6420 16541
rect 14004 16532 14056 16584
rect 16212 16532 16264 16584
rect 18512 16609 18521 16643
rect 18521 16609 18555 16643
rect 18555 16609 18564 16643
rect 18512 16600 18564 16609
rect 21088 16600 21140 16652
rect 22100 16600 22152 16652
rect 24492 16643 24544 16652
rect 24492 16609 24501 16643
rect 24501 16609 24535 16643
rect 24535 16609 24544 16643
rect 24492 16600 24544 16609
rect 26332 16600 26384 16652
rect 27252 16668 27304 16720
rect 28908 16668 28960 16720
rect 18052 16532 18104 16584
rect 19892 16575 19944 16584
rect 19892 16541 19901 16575
rect 19901 16541 19935 16575
rect 19935 16541 19944 16575
rect 19892 16532 19944 16541
rect 21180 16532 21232 16584
rect 22560 16532 22612 16584
rect 27160 16600 27212 16652
rect 28356 16600 28408 16652
rect 29736 16745 29745 16779
rect 29745 16745 29779 16779
rect 29779 16745 29788 16779
rect 29736 16736 29788 16745
rect 30012 16736 30064 16788
rect 31300 16736 31352 16788
rect 31944 16779 31996 16788
rect 31944 16745 31953 16779
rect 31953 16745 31987 16779
rect 31987 16745 31996 16779
rect 31944 16736 31996 16745
rect 33416 16779 33468 16788
rect 33416 16745 33425 16779
rect 33425 16745 33459 16779
rect 33459 16745 33468 16779
rect 33416 16736 33468 16745
rect 34336 16779 34388 16788
rect 34336 16745 34345 16779
rect 34345 16745 34379 16779
rect 34379 16745 34388 16779
rect 34336 16736 34388 16745
rect 40316 16779 40368 16788
rect 40316 16745 40325 16779
rect 40325 16745 40359 16779
rect 40359 16745 40368 16779
rect 40316 16736 40368 16745
rect 30288 16668 30340 16720
rect 32220 16711 32272 16720
rect 32220 16677 32229 16711
rect 32229 16677 32263 16711
rect 32263 16677 32272 16711
rect 32220 16668 32272 16677
rect 32312 16711 32364 16720
rect 32312 16677 32321 16711
rect 32321 16677 32355 16711
rect 32355 16677 32364 16711
rect 32312 16668 32364 16677
rect 36176 16668 36228 16720
rect 36728 16668 36780 16720
rect 37464 16668 37516 16720
rect 38016 16668 38068 16720
rect 38476 16711 38528 16720
rect 38476 16677 38485 16711
rect 38485 16677 38519 16711
rect 38519 16677 38528 16711
rect 38476 16668 38528 16677
rect 40868 16711 40920 16720
rect 40868 16677 40877 16711
rect 40877 16677 40911 16711
rect 40911 16677 40920 16711
rect 40868 16668 40920 16677
rect 41052 16668 41104 16720
rect 43168 16668 43220 16720
rect 43628 16668 43680 16720
rect 35256 16600 35308 16652
rect 39304 16643 39356 16652
rect 39304 16609 39313 16643
rect 39313 16609 39347 16643
rect 39347 16609 39356 16643
rect 39304 16600 39356 16609
rect 45008 16600 45060 16652
rect 30196 16575 30248 16584
rect 30196 16541 30205 16575
rect 30205 16541 30239 16575
rect 30239 16541 30248 16575
rect 30196 16532 30248 16541
rect 32496 16575 32548 16584
rect 32496 16541 32505 16575
rect 32505 16541 32539 16575
rect 32539 16541 32548 16575
rect 32496 16532 32548 16541
rect 33968 16575 34020 16584
rect 33968 16541 33977 16575
rect 33977 16541 34011 16575
rect 34011 16541 34020 16575
rect 33968 16532 34020 16541
rect 23572 16464 23624 16516
rect 24308 16464 24360 16516
rect 27896 16464 27948 16516
rect 42248 16464 42300 16516
rect 8576 16439 8628 16448
rect 8576 16405 8585 16439
rect 8585 16405 8619 16439
rect 8619 16405 8628 16439
rect 8576 16396 8628 16405
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 12716 16396 12768 16405
rect 15476 16396 15528 16448
rect 15844 16396 15896 16448
rect 22100 16439 22152 16448
rect 22100 16405 22109 16439
rect 22109 16405 22143 16439
rect 22143 16405 22152 16439
rect 22100 16396 22152 16405
rect 29000 16439 29052 16448
rect 29000 16405 29009 16439
rect 29009 16405 29043 16439
rect 29043 16405 29052 16439
rect 29000 16396 29052 16405
rect 31116 16439 31168 16448
rect 31116 16405 31125 16439
rect 31125 16405 31159 16439
rect 31159 16405 31168 16439
rect 31116 16396 31168 16405
rect 36360 16396 36412 16448
rect 36636 16439 36688 16448
rect 36636 16405 36645 16439
rect 36645 16405 36679 16439
rect 36679 16405 36688 16439
rect 36636 16396 36688 16405
rect 39488 16439 39540 16448
rect 39488 16405 39497 16439
rect 39497 16405 39531 16439
rect 39531 16405 39540 16439
rect 39488 16396 39540 16405
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 2688 16192 2740 16244
rect 3240 16192 3292 16244
rect 3700 16235 3752 16244
rect 3700 16201 3709 16235
rect 3709 16201 3743 16235
rect 3743 16201 3752 16235
rect 3700 16192 3752 16201
rect 3976 16192 4028 16244
rect 5908 16235 5960 16244
rect 5908 16201 5917 16235
rect 5917 16201 5951 16235
rect 5951 16201 5960 16235
rect 5908 16192 5960 16201
rect 6092 16192 6144 16244
rect 7748 16192 7800 16244
rect 13820 16235 13872 16244
rect 13820 16201 13829 16235
rect 13829 16201 13863 16235
rect 13863 16201 13872 16235
rect 15568 16235 15620 16244
rect 13820 16192 13872 16201
rect 15568 16201 15577 16235
rect 15577 16201 15611 16235
rect 15611 16201 15620 16235
rect 15568 16192 15620 16201
rect 20444 16192 20496 16244
rect 21088 16235 21140 16244
rect 21088 16201 21097 16235
rect 21097 16201 21131 16235
rect 21131 16201 21140 16235
rect 21088 16192 21140 16201
rect 23204 16192 23256 16244
rect 25872 16192 25924 16244
rect 27252 16235 27304 16244
rect 27252 16201 27261 16235
rect 27261 16201 27295 16235
rect 27295 16201 27304 16235
rect 27252 16192 27304 16201
rect 28908 16192 28960 16244
rect 18052 16124 18104 16176
rect 23572 16124 23624 16176
rect 24492 16124 24544 16176
rect 3148 16056 3200 16108
rect 7656 16056 7708 16108
rect 9588 16099 9640 16108
rect 9588 16065 9597 16099
rect 9597 16065 9631 16099
rect 9631 16065 9640 16099
rect 9588 16056 9640 16065
rect 12532 16056 12584 16108
rect 14280 16099 14332 16108
rect 14280 16065 14289 16099
rect 14289 16065 14323 16099
rect 14323 16065 14332 16099
rect 14280 16056 14332 16065
rect 18512 16056 18564 16108
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 4712 15988 4764 15997
rect 18144 15988 18196 16040
rect 18236 15988 18288 16040
rect 4988 15852 5040 15904
rect 6460 15920 6512 15972
rect 7656 15920 7708 15972
rect 9496 15963 9548 15972
rect 9496 15929 9505 15963
rect 9505 15929 9539 15963
rect 9539 15929 9548 15963
rect 9496 15920 9548 15929
rect 10324 15920 10376 15972
rect 12164 15963 12216 15972
rect 12164 15929 12173 15963
rect 12173 15929 12207 15963
rect 12207 15929 12216 15963
rect 12164 15920 12216 15929
rect 13544 15920 13596 15972
rect 14556 15920 14608 15972
rect 17868 15920 17920 15972
rect 26056 16056 26108 16108
rect 26424 16056 26476 16108
rect 26516 16056 26568 16108
rect 28632 16099 28684 16108
rect 19892 15988 19944 16040
rect 20904 15920 20956 15972
rect 22100 15963 22152 15972
rect 22100 15929 22109 15963
rect 22109 15929 22143 15963
rect 22143 15929 22152 15963
rect 22100 15920 22152 15929
rect 27160 15988 27212 16040
rect 28632 16065 28641 16099
rect 28641 16065 28675 16099
rect 28675 16065 28684 16099
rect 28632 16056 28684 16065
rect 31116 16192 31168 16244
rect 31576 16192 31628 16244
rect 32312 16192 32364 16244
rect 33140 16235 33192 16244
rect 33140 16201 33149 16235
rect 33149 16201 33183 16235
rect 33183 16201 33192 16235
rect 35256 16235 35308 16244
rect 33140 16192 33192 16201
rect 35256 16201 35265 16235
rect 35265 16201 35299 16235
rect 35299 16201 35308 16235
rect 35256 16192 35308 16201
rect 36176 16192 36228 16244
rect 39304 16192 39356 16244
rect 29644 16124 29696 16176
rect 30196 16056 30248 16108
rect 31300 16056 31352 16108
rect 32312 16056 32364 16108
rect 32496 16056 32548 16108
rect 29736 16031 29788 16040
rect 29736 15997 29745 16031
rect 29745 15997 29779 16031
rect 29779 15997 29788 16031
rect 29736 15988 29788 15997
rect 33968 16099 34020 16108
rect 33508 16031 33560 16040
rect 33508 15997 33517 16031
rect 33517 15997 33551 16031
rect 33551 15997 33560 16031
rect 33508 15988 33560 15997
rect 33968 16065 33977 16099
rect 33977 16065 34011 16099
rect 34011 16065 34020 16099
rect 33968 16056 34020 16065
rect 38568 16124 38620 16176
rect 42156 16124 42208 16176
rect 37188 16099 37240 16108
rect 34060 15988 34112 16040
rect 37188 16065 37197 16099
rect 37197 16065 37231 16099
rect 37231 16065 37240 16099
rect 37188 16056 37240 16065
rect 40316 16056 40368 16108
rect 42064 16056 42116 16108
rect 44088 16099 44140 16108
rect 44088 16065 44097 16099
rect 44097 16065 44131 16099
rect 44131 16065 44140 16099
rect 44088 16056 44140 16065
rect 38568 15988 38620 16040
rect 23756 15963 23808 15972
rect 5816 15852 5868 15904
rect 8484 15895 8536 15904
rect 8484 15861 8493 15895
rect 8493 15861 8527 15895
rect 8527 15861 8536 15895
rect 8484 15852 8536 15861
rect 10508 15852 10560 15904
rect 12256 15852 12308 15904
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 20168 15852 20220 15904
rect 23756 15929 23765 15963
rect 23765 15929 23799 15963
rect 23799 15929 23808 15963
rect 23756 15920 23808 15929
rect 23848 15963 23900 15972
rect 23848 15929 23857 15963
rect 23857 15929 23891 15963
rect 23891 15929 23900 15963
rect 23848 15920 23900 15929
rect 24584 15920 24636 15972
rect 26332 15920 26384 15972
rect 31484 15920 31536 15972
rect 31576 15963 31628 15972
rect 31576 15929 31585 15963
rect 31585 15929 31619 15963
rect 31619 15929 31628 15963
rect 31576 15920 31628 15929
rect 31760 15920 31812 15972
rect 34336 15920 34388 15972
rect 36544 15963 36596 15972
rect 36544 15929 36553 15963
rect 36553 15929 36587 15963
rect 36587 15929 36596 15963
rect 36544 15920 36596 15929
rect 25320 15852 25372 15904
rect 30288 15895 30340 15904
rect 30288 15861 30297 15895
rect 30297 15861 30331 15895
rect 30331 15861 30340 15895
rect 30288 15852 30340 15861
rect 34520 15852 34572 15904
rect 36176 15852 36228 15904
rect 36360 15852 36412 15904
rect 39672 15920 39724 15972
rect 40316 15920 40368 15972
rect 41052 15920 41104 15972
rect 37832 15852 37884 15904
rect 38016 15852 38068 15904
rect 42616 15895 42668 15904
rect 42616 15861 42625 15895
rect 42625 15861 42659 15895
rect 42659 15861 42668 15895
rect 42616 15852 42668 15861
rect 43628 15852 43680 15904
rect 45008 15895 45060 15904
rect 45008 15861 45017 15895
rect 45017 15861 45051 15895
rect 45051 15861 45060 15895
rect 45008 15852 45060 15861
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 4712 15648 4764 15700
rect 7656 15691 7708 15700
rect 7656 15657 7665 15691
rect 7665 15657 7699 15691
rect 7699 15657 7708 15691
rect 7656 15648 7708 15657
rect 9772 15648 9824 15700
rect 10876 15648 10928 15700
rect 11796 15691 11848 15700
rect 11796 15657 11805 15691
rect 11805 15657 11839 15691
rect 11839 15657 11848 15691
rect 11796 15648 11848 15657
rect 12532 15648 12584 15700
rect 14280 15691 14332 15700
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 22560 15691 22612 15700
rect 22560 15657 22569 15691
rect 22569 15657 22603 15691
rect 22603 15657 22612 15691
rect 22560 15648 22612 15657
rect 23756 15691 23808 15700
rect 23756 15657 23765 15691
rect 23765 15657 23799 15691
rect 23799 15657 23808 15691
rect 23756 15648 23808 15657
rect 26056 15691 26108 15700
rect 26056 15657 26065 15691
rect 26065 15657 26099 15691
rect 26099 15657 26108 15691
rect 26056 15648 26108 15657
rect 29736 15648 29788 15700
rect 32220 15648 32272 15700
rect 36452 15648 36504 15700
rect 36544 15648 36596 15700
rect 37464 15691 37516 15700
rect 37464 15657 37473 15691
rect 37473 15657 37507 15691
rect 37507 15657 37516 15691
rect 37464 15648 37516 15657
rect 37832 15648 37884 15700
rect 38568 15691 38620 15700
rect 38568 15657 38577 15691
rect 38577 15657 38611 15691
rect 38611 15657 38620 15691
rect 38568 15648 38620 15657
rect 42064 15648 42116 15700
rect 43168 15691 43220 15700
rect 43168 15657 43177 15691
rect 43177 15657 43211 15691
rect 43211 15657 43220 15691
rect 43168 15648 43220 15657
rect 44088 15648 44140 15700
rect 3700 15580 3752 15632
rect 3884 15512 3936 15564
rect 4620 15580 4672 15632
rect 6460 15580 6512 15632
rect 9864 15623 9916 15632
rect 9864 15589 9873 15623
rect 9873 15589 9907 15623
rect 9907 15589 9916 15623
rect 9864 15580 9916 15589
rect 13544 15580 13596 15632
rect 15844 15623 15896 15632
rect 15844 15589 15853 15623
rect 15853 15589 15887 15623
rect 15887 15589 15896 15623
rect 15844 15580 15896 15589
rect 15936 15623 15988 15632
rect 15936 15589 15945 15623
rect 15945 15589 15979 15623
rect 15979 15589 15988 15623
rect 15936 15580 15988 15589
rect 18052 15580 18104 15632
rect 19892 15623 19944 15632
rect 6368 15555 6420 15564
rect 6368 15521 6377 15555
rect 6377 15521 6411 15555
rect 6411 15521 6420 15555
rect 6368 15512 6420 15521
rect 8484 15512 8536 15564
rect 12256 15512 12308 15564
rect 13176 15512 13228 15564
rect 18236 15512 18288 15564
rect 18604 15512 18656 15564
rect 19340 15555 19392 15564
rect 19340 15521 19349 15555
rect 19349 15521 19383 15555
rect 19383 15521 19392 15555
rect 19340 15512 19392 15521
rect 19892 15589 19901 15623
rect 19901 15589 19935 15623
rect 19935 15589 19944 15623
rect 19892 15580 19944 15589
rect 23204 15580 23256 15632
rect 24124 15580 24176 15632
rect 25320 15580 25372 15632
rect 26332 15580 26384 15632
rect 29276 15623 29328 15632
rect 29276 15589 29285 15623
rect 29285 15589 29319 15623
rect 29319 15589 29328 15623
rect 29276 15580 29328 15589
rect 31576 15580 31628 15632
rect 32036 15580 32088 15632
rect 32588 15580 32640 15632
rect 41052 15623 41104 15632
rect 41052 15589 41061 15623
rect 41061 15589 41095 15623
rect 41095 15589 41104 15623
rect 41052 15580 41104 15589
rect 43628 15580 43680 15632
rect 21732 15512 21784 15564
rect 26608 15512 26660 15564
rect 30840 15512 30892 15564
rect 34152 15555 34204 15564
rect 34152 15521 34161 15555
rect 34161 15521 34195 15555
rect 34195 15521 34204 15555
rect 34152 15512 34204 15521
rect 34612 15512 34664 15564
rect 35072 15555 35124 15564
rect 35072 15521 35081 15555
rect 35081 15521 35115 15555
rect 35115 15521 35124 15555
rect 35072 15512 35124 15521
rect 36268 15512 36320 15564
rect 38200 15512 38252 15564
rect 38752 15555 38804 15564
rect 38752 15521 38761 15555
rect 38761 15521 38795 15555
rect 38795 15521 38804 15555
rect 38752 15512 38804 15521
rect 39488 15512 39540 15564
rect 44824 15512 44876 15564
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 15384 15444 15436 15496
rect 16672 15444 16724 15496
rect 22744 15487 22796 15496
rect 22744 15453 22753 15487
rect 22753 15453 22787 15487
rect 22787 15453 22796 15487
rect 22744 15444 22796 15453
rect 23388 15487 23440 15496
rect 23388 15453 23397 15487
rect 23397 15453 23431 15487
rect 23431 15453 23440 15487
rect 23388 15444 23440 15453
rect 24584 15487 24636 15496
rect 24584 15453 24593 15487
rect 24593 15453 24627 15487
rect 24627 15453 24636 15487
rect 24584 15444 24636 15453
rect 29368 15444 29420 15496
rect 31944 15444 31996 15496
rect 32956 15444 33008 15496
rect 33508 15444 33560 15496
rect 40960 15487 41012 15496
rect 40960 15453 40969 15487
rect 40969 15453 41003 15487
rect 41003 15453 41012 15487
rect 40960 15444 41012 15453
rect 44456 15444 44508 15496
rect 10140 15376 10192 15428
rect 11520 15376 11572 15428
rect 7564 15308 7616 15360
rect 8852 15351 8904 15360
rect 8852 15317 8861 15351
rect 8861 15317 8895 15351
rect 8895 15317 8904 15351
rect 8852 15308 8904 15317
rect 12072 15308 12124 15360
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 14004 15351 14056 15360
rect 14004 15317 14013 15351
rect 14013 15317 14047 15351
rect 14047 15317 14056 15351
rect 14004 15308 14056 15317
rect 32588 15376 32640 15428
rect 43720 15376 43772 15428
rect 22376 15308 22428 15360
rect 25228 15351 25280 15360
rect 25228 15317 25237 15351
rect 25237 15317 25271 15351
rect 25271 15317 25280 15351
rect 25228 15308 25280 15317
rect 26884 15308 26936 15360
rect 31760 15308 31812 15360
rect 34796 15308 34848 15360
rect 35348 15308 35400 15360
rect 36544 15308 36596 15360
rect 36636 15351 36688 15360
rect 36636 15317 36645 15351
rect 36645 15317 36679 15351
rect 36679 15317 36688 15351
rect 40040 15351 40092 15360
rect 36636 15308 36688 15317
rect 40040 15317 40049 15351
rect 40049 15317 40083 15351
rect 40083 15317 40092 15351
rect 40040 15308 40092 15317
rect 40592 15351 40644 15360
rect 40592 15317 40601 15351
rect 40601 15317 40635 15351
rect 40635 15317 40644 15351
rect 40592 15308 40644 15317
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 3700 15104 3752 15156
rect 3884 15147 3936 15156
rect 3884 15113 3893 15147
rect 3893 15113 3927 15147
rect 3927 15113 3936 15147
rect 3884 15104 3936 15113
rect 6276 15104 6328 15156
rect 8484 15104 8536 15156
rect 10140 15147 10192 15156
rect 10140 15113 10149 15147
rect 10149 15113 10183 15147
rect 10183 15113 10192 15147
rect 10140 15104 10192 15113
rect 12256 15104 12308 15156
rect 13176 15104 13228 15156
rect 18052 15104 18104 15156
rect 18604 15147 18656 15156
rect 18604 15113 18613 15147
rect 18613 15113 18647 15147
rect 18647 15113 18656 15147
rect 18604 15104 18656 15113
rect 22744 15104 22796 15156
rect 26608 15104 26660 15156
rect 29368 15104 29420 15156
rect 30840 15104 30892 15156
rect 7104 15036 7156 15088
rect 9864 15036 9916 15088
rect 12440 15036 12492 15088
rect 4620 14968 4672 15020
rect 6460 15011 6512 15020
rect 6460 14977 6469 15011
rect 6469 14977 6503 15011
rect 6503 14977 6512 15011
rect 6460 14968 6512 14977
rect 10048 14968 10100 15020
rect 10876 14968 10928 15020
rect 11152 15011 11204 15020
rect 11152 14977 11161 15011
rect 11161 14977 11195 15011
rect 11195 14977 11204 15011
rect 11152 14968 11204 14977
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 16948 15036 17000 15088
rect 23756 15036 23808 15088
rect 23848 15036 23900 15088
rect 26884 15036 26936 15088
rect 29276 15036 29328 15088
rect 15108 15011 15160 15020
rect 15108 14977 15117 15011
rect 15117 14977 15151 15011
rect 15151 14977 15160 15011
rect 15108 14968 15160 14977
rect 15476 14968 15528 15020
rect 16396 15011 16448 15020
rect 16396 14977 16405 15011
rect 16405 14977 16439 15011
rect 16439 14977 16448 15011
rect 16396 14968 16448 14977
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 19340 14968 19392 15020
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 24032 14968 24084 15020
rect 25228 15011 25280 15020
rect 25228 14977 25237 15011
rect 25237 14977 25271 15011
rect 25271 14977 25280 15011
rect 25228 14968 25280 14977
rect 25872 15011 25924 15020
rect 25872 14977 25881 15011
rect 25881 14977 25915 15011
rect 25915 14977 25924 15011
rect 25872 14968 25924 14977
rect 31668 15104 31720 15156
rect 32036 15104 32088 15156
rect 33140 15104 33192 15156
rect 5816 14900 5868 14952
rect 13360 14900 13412 14952
rect 4988 14832 5040 14884
rect 8852 14875 8904 14884
rect 8852 14841 8861 14875
rect 8861 14841 8895 14875
rect 8895 14841 8904 14875
rect 8852 14832 8904 14841
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 6920 14764 6972 14816
rect 8484 14764 8536 14816
rect 10600 14832 10652 14884
rect 13820 14832 13872 14884
rect 13544 14807 13596 14816
rect 13544 14773 13553 14807
rect 13553 14773 13587 14807
rect 13587 14773 13596 14807
rect 13544 14764 13596 14773
rect 18328 14900 18380 14952
rect 19892 14943 19944 14952
rect 19892 14909 19901 14943
rect 19901 14909 19935 14943
rect 19935 14909 19944 14943
rect 19892 14900 19944 14909
rect 22928 14943 22980 14952
rect 22928 14909 22937 14943
rect 22937 14909 22971 14943
rect 22971 14909 22980 14943
rect 22928 14900 22980 14909
rect 23204 14900 23256 14952
rect 28264 14900 28316 14952
rect 30564 14900 30616 14952
rect 31668 14900 31720 14952
rect 32956 14900 33008 14952
rect 33876 15104 33928 15156
rect 34612 15079 34664 15088
rect 34612 15045 34621 15079
rect 34621 15045 34655 15079
rect 34655 15045 34664 15079
rect 34612 15036 34664 15045
rect 36268 15079 36320 15088
rect 36268 15045 36277 15079
rect 36277 15045 36311 15079
rect 36311 15045 36320 15079
rect 36268 15036 36320 15045
rect 35256 15011 35308 15020
rect 35256 14977 35265 15011
rect 35265 14977 35299 15011
rect 35299 14977 35308 15011
rect 35256 14968 35308 14977
rect 36544 15011 36596 15020
rect 36544 14977 36553 15011
rect 36553 14977 36587 15011
rect 36587 14977 36596 15011
rect 36544 14968 36596 14977
rect 36820 15011 36872 15020
rect 36820 14977 36829 15011
rect 36829 14977 36863 15011
rect 36863 14977 36872 15011
rect 36820 14968 36872 14977
rect 38752 15104 38804 15156
rect 40316 15147 40368 15156
rect 40316 15113 40325 15147
rect 40325 15113 40359 15147
rect 40359 15113 40368 15147
rect 40316 15104 40368 15113
rect 43628 15104 43680 15156
rect 44456 15147 44508 15156
rect 44456 15113 44465 15147
rect 44465 15113 44499 15147
rect 44499 15113 44508 15147
rect 44456 15104 44508 15113
rect 38200 15079 38252 15088
rect 38200 15045 38209 15079
rect 38209 15045 38243 15079
rect 38243 15045 38252 15079
rect 38200 15036 38252 15045
rect 40592 15011 40644 15020
rect 40592 14977 40601 15011
rect 40601 14977 40635 15011
rect 40635 14977 40644 15011
rect 40592 14968 40644 14977
rect 44732 14968 44784 15020
rect 39120 14900 39172 14952
rect 40040 14900 40092 14952
rect 42524 14943 42576 14952
rect 42524 14909 42533 14943
rect 42533 14909 42567 14943
rect 42567 14909 42576 14943
rect 42524 14900 42576 14909
rect 14832 14875 14884 14884
rect 14832 14841 14841 14875
rect 14841 14841 14875 14875
rect 14875 14841 14884 14875
rect 14832 14832 14884 14841
rect 16856 14832 16908 14884
rect 20076 14832 20128 14884
rect 23296 14832 23348 14884
rect 25320 14875 25372 14884
rect 25320 14841 25329 14875
rect 25329 14841 25363 14875
rect 25363 14841 25372 14875
rect 25320 14832 25372 14841
rect 26792 14875 26844 14884
rect 26792 14841 26801 14875
rect 26801 14841 26835 14875
rect 26835 14841 26844 14875
rect 26792 14832 26844 14841
rect 26884 14875 26936 14884
rect 26884 14841 26893 14875
rect 26893 14841 26927 14875
rect 26927 14841 26936 14875
rect 26884 14832 26936 14841
rect 15936 14764 15988 14816
rect 20812 14807 20864 14816
rect 20812 14773 20821 14807
rect 20821 14773 20855 14807
rect 20855 14773 20864 14807
rect 20812 14764 20864 14773
rect 21732 14807 21784 14816
rect 21732 14773 21741 14807
rect 21741 14773 21775 14807
rect 21775 14773 21784 14807
rect 21732 14764 21784 14773
rect 26332 14764 26384 14816
rect 30288 14832 30340 14884
rect 34980 14875 35032 14884
rect 34980 14841 34989 14875
rect 34989 14841 35023 14875
rect 35023 14841 35032 14875
rect 34980 14832 35032 14841
rect 35348 14832 35400 14884
rect 36636 14875 36688 14884
rect 36636 14841 36645 14875
rect 36645 14841 36679 14875
rect 36679 14841 36688 14875
rect 36636 14832 36688 14841
rect 39580 14832 39632 14884
rect 40316 14832 40368 14884
rect 30196 14807 30248 14816
rect 30196 14773 30205 14807
rect 30205 14773 30239 14807
rect 30239 14773 30248 14807
rect 30196 14764 30248 14773
rect 32680 14764 32732 14816
rect 33968 14764 34020 14816
rect 34152 14807 34204 14816
rect 34152 14773 34161 14807
rect 34161 14773 34195 14807
rect 34195 14773 34204 14807
rect 34152 14764 34204 14773
rect 41696 14832 41748 14884
rect 43536 14875 43588 14884
rect 43536 14841 43545 14875
rect 43545 14841 43579 14875
rect 43579 14841 43588 14875
rect 43536 14832 43588 14841
rect 43628 14875 43680 14884
rect 43628 14841 43637 14875
rect 43637 14841 43671 14875
rect 43671 14841 43680 14875
rect 44180 14875 44232 14884
rect 43628 14832 43680 14841
rect 44180 14841 44189 14875
rect 44189 14841 44223 14875
rect 44223 14841 44232 14875
rect 44180 14832 44232 14841
rect 44824 14875 44876 14884
rect 44824 14841 44833 14875
rect 44833 14841 44867 14875
rect 44867 14841 44876 14875
rect 44824 14832 44876 14841
rect 46940 14832 46992 14884
rect 44916 14764 44968 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 6828 14560 6880 14612
rect 4988 14492 5040 14544
rect 12072 14560 12124 14612
rect 14832 14603 14884 14612
rect 10508 14535 10560 14544
rect 10508 14501 10517 14535
rect 10517 14501 10551 14535
rect 10551 14501 10560 14535
rect 10508 14492 10560 14501
rect 10600 14535 10652 14544
rect 10600 14501 10609 14535
rect 10609 14501 10643 14535
rect 10643 14501 10652 14535
rect 11152 14535 11204 14544
rect 10600 14492 10652 14501
rect 11152 14501 11161 14535
rect 11161 14501 11195 14535
rect 11195 14501 11204 14535
rect 11152 14492 11204 14501
rect 14832 14569 14841 14603
rect 14841 14569 14875 14603
rect 14875 14569 14884 14603
rect 14832 14560 14884 14569
rect 15844 14603 15896 14612
rect 15844 14569 15853 14603
rect 15853 14569 15887 14603
rect 15887 14569 15896 14603
rect 15844 14560 15896 14569
rect 16396 14603 16448 14612
rect 16396 14569 16405 14603
rect 16405 14569 16439 14603
rect 16439 14569 16448 14603
rect 16396 14560 16448 14569
rect 18328 14560 18380 14612
rect 23020 14560 23072 14612
rect 23296 14560 23348 14612
rect 24216 14603 24268 14612
rect 24216 14569 24225 14603
rect 24225 14569 24259 14603
rect 24259 14569 24268 14603
rect 24216 14560 24268 14569
rect 25228 14560 25280 14612
rect 27344 14560 27396 14612
rect 12256 14535 12308 14544
rect 12256 14501 12265 14535
rect 12265 14501 12299 14535
rect 12299 14501 12308 14535
rect 12256 14492 12308 14501
rect 13360 14492 13412 14544
rect 13820 14535 13872 14544
rect 13820 14501 13829 14535
rect 13829 14501 13863 14535
rect 13863 14501 13872 14535
rect 13820 14492 13872 14501
rect 15108 14492 15160 14544
rect 16856 14535 16908 14544
rect 16856 14501 16865 14535
rect 16865 14501 16899 14535
rect 16899 14501 16908 14535
rect 16856 14492 16908 14501
rect 19892 14492 19944 14544
rect 20812 14492 20864 14544
rect 22376 14492 22428 14544
rect 22836 14535 22888 14544
rect 22836 14501 22845 14535
rect 22845 14501 22879 14535
rect 22879 14501 22888 14535
rect 23388 14535 23440 14544
rect 22836 14492 22888 14501
rect 23388 14501 23397 14535
rect 23397 14501 23431 14535
rect 23431 14501 23440 14535
rect 23388 14492 23440 14501
rect 3700 14356 3752 14408
rect 4896 14424 4948 14476
rect 7564 14424 7616 14476
rect 15200 14424 15252 14476
rect 6920 14399 6972 14408
rect 6920 14365 6929 14399
rect 6929 14365 6963 14399
rect 6963 14365 6972 14399
rect 6920 14356 6972 14365
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 13728 14399 13780 14408
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 13820 14356 13872 14408
rect 17224 14467 17276 14476
rect 17224 14433 17233 14467
rect 17233 14433 17267 14467
rect 17267 14433 17276 14467
rect 17224 14424 17276 14433
rect 18788 14424 18840 14476
rect 20168 14424 20220 14476
rect 24952 14467 25004 14476
rect 24952 14433 24970 14467
rect 24970 14433 25004 14467
rect 26424 14467 26476 14476
rect 24952 14424 25004 14433
rect 20352 14356 20404 14408
rect 7472 14331 7524 14340
rect 7472 14297 7481 14331
rect 7481 14297 7515 14331
rect 7515 14297 7524 14331
rect 7472 14288 7524 14297
rect 10140 14288 10192 14340
rect 21548 14331 21600 14340
rect 21548 14297 21557 14331
rect 21557 14297 21591 14331
rect 21591 14297 21600 14331
rect 21548 14288 21600 14297
rect 26424 14433 26433 14467
rect 26433 14433 26467 14467
rect 26467 14433 26476 14467
rect 26424 14424 26476 14433
rect 26792 14424 26844 14476
rect 39120 14603 39172 14612
rect 28264 14535 28316 14544
rect 28264 14501 28273 14535
rect 28273 14501 28307 14535
rect 28307 14501 28316 14535
rect 28264 14492 28316 14501
rect 29276 14535 29328 14544
rect 29276 14501 29285 14535
rect 29285 14501 29319 14535
rect 29319 14501 29328 14535
rect 29276 14492 29328 14501
rect 30196 14492 30248 14544
rect 31484 14535 31536 14544
rect 31484 14501 31493 14535
rect 31493 14501 31527 14535
rect 31527 14501 31536 14535
rect 31484 14492 31536 14501
rect 31760 14492 31812 14544
rect 32404 14492 32456 14544
rect 39120 14569 39129 14603
rect 39129 14569 39163 14603
rect 39163 14569 39172 14603
rect 39120 14560 39172 14569
rect 34428 14535 34480 14544
rect 34428 14501 34437 14535
rect 34437 14501 34471 14535
rect 34471 14501 34480 14535
rect 34428 14492 34480 14501
rect 35256 14492 35308 14544
rect 36268 14535 36320 14544
rect 36268 14501 36277 14535
rect 36277 14501 36311 14535
rect 36311 14501 36320 14535
rect 36268 14492 36320 14501
rect 36820 14535 36872 14544
rect 36820 14501 36829 14535
rect 36829 14501 36863 14535
rect 36863 14501 36872 14535
rect 36820 14492 36872 14501
rect 39672 14492 39724 14544
rect 42616 14560 42668 14612
rect 43536 14560 43588 14612
rect 44916 14560 44968 14612
rect 41420 14492 41472 14544
rect 42248 14535 42300 14544
rect 42248 14501 42257 14535
rect 42257 14501 42291 14535
rect 42291 14501 42300 14535
rect 42248 14492 42300 14501
rect 28080 14467 28132 14476
rect 28080 14433 28089 14467
rect 28089 14433 28123 14467
rect 28123 14433 28132 14467
rect 28080 14424 28132 14433
rect 29000 14424 29052 14476
rect 31300 14424 31352 14476
rect 31944 14467 31996 14476
rect 31944 14433 31953 14467
rect 31953 14433 31987 14467
rect 31987 14433 31996 14467
rect 31944 14424 31996 14433
rect 40960 14424 41012 14476
rect 43536 14424 43588 14476
rect 29184 14399 29236 14408
rect 29184 14365 29193 14399
rect 29193 14365 29227 14399
rect 29227 14365 29236 14399
rect 29184 14356 29236 14365
rect 31852 14356 31904 14408
rect 32496 14399 32548 14408
rect 32496 14365 32505 14399
rect 32505 14365 32539 14399
rect 32539 14365 32548 14399
rect 32496 14356 32548 14365
rect 32680 14356 32732 14408
rect 30840 14288 30892 14340
rect 34980 14356 35032 14408
rect 39580 14399 39632 14408
rect 39580 14365 39589 14399
rect 39589 14365 39623 14399
rect 39623 14365 39632 14399
rect 39580 14356 39632 14365
rect 37648 14288 37700 14340
rect 5540 14220 5592 14272
rect 8668 14220 8720 14272
rect 25320 14263 25372 14272
rect 25320 14229 25329 14263
rect 25329 14229 25363 14263
rect 25363 14229 25372 14263
rect 25320 14220 25372 14229
rect 26976 14263 27028 14272
rect 26976 14229 26985 14263
rect 26985 14229 27019 14263
rect 27019 14229 27028 14263
rect 26976 14220 27028 14229
rect 31300 14220 31352 14272
rect 32864 14220 32916 14272
rect 39212 14220 39264 14272
rect 40500 14263 40552 14272
rect 40500 14229 40509 14263
rect 40509 14229 40543 14263
rect 40543 14229 40552 14263
rect 40500 14220 40552 14229
rect 41328 14263 41380 14272
rect 41328 14229 41337 14263
rect 41337 14229 41371 14263
rect 41371 14229 41380 14263
rect 41328 14220 41380 14229
rect 42984 14220 43036 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 3700 14059 3752 14068
rect 3700 14025 3709 14059
rect 3709 14025 3743 14059
rect 3743 14025 3752 14059
rect 3700 14016 3752 14025
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 6920 14016 6972 14068
rect 10600 14016 10652 14068
rect 12256 14016 12308 14068
rect 12532 14016 12584 14068
rect 13728 14016 13780 14068
rect 13820 14016 13872 14068
rect 14004 14016 14056 14068
rect 15200 14016 15252 14068
rect 6828 13948 6880 14000
rect 7472 13991 7524 14000
rect 7104 13880 7156 13932
rect 7472 13957 7481 13991
rect 7481 13957 7515 13991
rect 7515 13957 7524 13991
rect 7472 13948 7524 13957
rect 12072 13948 12124 14000
rect 4620 13812 4672 13864
rect 4988 13812 5040 13864
rect 6736 13744 6788 13796
rect 7012 13787 7064 13796
rect 7012 13753 7021 13787
rect 7021 13753 7055 13787
rect 7055 13753 7064 13787
rect 8668 13880 8720 13932
rect 10140 13923 10192 13932
rect 10140 13889 10149 13923
rect 10149 13889 10183 13923
rect 10183 13889 10192 13923
rect 10140 13880 10192 13889
rect 12716 13812 12768 13864
rect 15108 13880 15160 13932
rect 15936 13812 15988 13864
rect 17500 13812 17552 13864
rect 7012 13744 7064 13753
rect 8484 13744 8536 13796
rect 9128 13787 9180 13796
rect 9128 13753 9137 13787
rect 9137 13753 9171 13787
rect 9171 13753 9180 13787
rect 9128 13744 9180 13753
rect 5448 13719 5500 13728
rect 5448 13685 5457 13719
rect 5457 13685 5491 13719
rect 5491 13685 5500 13719
rect 5448 13676 5500 13685
rect 6828 13676 6880 13728
rect 9956 13719 10008 13728
rect 9956 13685 9965 13719
rect 9965 13685 9999 13719
rect 9999 13685 10008 13719
rect 12992 13744 13044 13796
rect 15292 13744 15344 13796
rect 15568 13787 15620 13796
rect 15568 13753 15577 13787
rect 15577 13753 15611 13787
rect 15611 13753 15620 13787
rect 15568 13744 15620 13753
rect 18696 13744 18748 13796
rect 19432 13812 19484 13864
rect 20168 14016 20220 14068
rect 20812 14016 20864 14068
rect 22376 14059 22428 14068
rect 22376 14025 22385 14059
rect 22385 14025 22419 14059
rect 22419 14025 22428 14059
rect 22376 14016 22428 14025
rect 23112 14059 23164 14068
rect 23112 14025 23121 14059
rect 23121 14025 23155 14059
rect 23155 14025 23164 14059
rect 23112 14016 23164 14025
rect 20904 13948 20956 14000
rect 21088 13991 21140 14000
rect 21088 13957 21097 13991
rect 21097 13957 21131 13991
rect 21131 13957 21140 13991
rect 21088 13948 21140 13957
rect 22836 13948 22888 14000
rect 23848 14016 23900 14068
rect 24952 14059 25004 14068
rect 24952 14025 24961 14059
rect 24961 14025 24995 14059
rect 24995 14025 25004 14059
rect 24952 14016 25004 14025
rect 26424 14059 26476 14068
rect 26424 14025 26433 14059
rect 26433 14025 26467 14059
rect 26467 14025 26476 14059
rect 26424 14016 26476 14025
rect 27344 14016 27396 14068
rect 28080 14059 28132 14068
rect 28080 14025 28089 14059
rect 28089 14025 28123 14059
rect 28123 14025 28132 14059
rect 28080 14016 28132 14025
rect 29184 14016 29236 14068
rect 29092 13991 29144 14000
rect 21456 13812 21508 13864
rect 25320 13880 25372 13932
rect 25872 13880 25924 13932
rect 23112 13812 23164 13864
rect 27344 13880 27396 13932
rect 20260 13744 20312 13796
rect 26976 13812 27028 13864
rect 29092 13957 29101 13991
rect 29101 13957 29135 13991
rect 29135 13957 29144 13991
rect 29092 13948 29144 13957
rect 29276 13948 29328 14000
rect 29828 13948 29880 14000
rect 32312 14016 32364 14068
rect 32404 14016 32456 14068
rect 33324 14016 33376 14068
rect 34428 14016 34480 14068
rect 36268 14016 36320 14068
rect 37648 14059 37700 14068
rect 37648 14025 37657 14059
rect 37657 14025 37691 14059
rect 37691 14025 37700 14059
rect 37648 14016 37700 14025
rect 31300 13948 31352 14000
rect 31484 13948 31536 14000
rect 34520 13948 34572 14000
rect 38384 14016 38436 14068
rect 39212 14059 39264 14068
rect 39212 14025 39221 14059
rect 39221 14025 39255 14059
rect 39255 14025 39264 14059
rect 39212 14016 39264 14025
rect 39580 14016 39632 14068
rect 41328 14016 41380 14068
rect 42984 14059 43036 14068
rect 31852 13923 31904 13932
rect 31852 13889 31861 13923
rect 31861 13889 31895 13923
rect 31895 13889 31904 13923
rect 31852 13880 31904 13889
rect 32956 13880 33008 13932
rect 34152 13880 34204 13932
rect 35900 13880 35952 13932
rect 36820 13880 36872 13932
rect 37188 13923 37240 13932
rect 37188 13889 37197 13923
rect 37197 13889 37231 13923
rect 37231 13889 37240 13923
rect 37188 13880 37240 13889
rect 28816 13812 28868 13864
rect 34888 13855 34940 13864
rect 34888 13821 34897 13855
rect 34897 13821 34931 13855
rect 34931 13821 34940 13855
rect 34888 13812 34940 13821
rect 24952 13744 25004 13796
rect 25228 13787 25280 13796
rect 25228 13753 25237 13787
rect 25237 13753 25271 13787
rect 25271 13753 25280 13787
rect 25228 13744 25280 13753
rect 29092 13744 29144 13796
rect 29460 13787 29512 13796
rect 29460 13753 29469 13787
rect 29469 13753 29503 13787
rect 29503 13753 29512 13787
rect 29460 13744 29512 13753
rect 31576 13744 31628 13796
rect 32036 13744 32088 13796
rect 32404 13744 32456 13796
rect 33324 13744 33376 13796
rect 34520 13744 34572 13796
rect 36728 13787 36780 13796
rect 36728 13753 36737 13787
rect 36737 13753 36771 13787
rect 36771 13753 36780 13787
rect 36728 13744 36780 13753
rect 38200 13948 38252 14000
rect 39672 13991 39724 14000
rect 39672 13957 39681 13991
rect 39681 13957 39715 13991
rect 39715 13957 39724 13991
rect 39672 13948 39724 13957
rect 40500 13948 40552 14000
rect 41420 13991 41472 14000
rect 38476 13880 38528 13932
rect 40960 13923 41012 13932
rect 40960 13889 40969 13923
rect 40969 13889 41003 13923
rect 41003 13889 41012 13923
rect 40960 13880 41012 13889
rect 9956 13676 10008 13685
rect 17224 13676 17276 13728
rect 20352 13719 20404 13728
rect 20352 13685 20361 13719
rect 20361 13685 20395 13719
rect 20395 13685 20404 13719
rect 20352 13676 20404 13685
rect 22376 13676 22428 13728
rect 23112 13676 23164 13728
rect 24400 13676 24452 13728
rect 26700 13719 26752 13728
rect 26700 13685 26709 13719
rect 26709 13685 26743 13719
rect 26743 13685 26752 13719
rect 26700 13676 26752 13685
rect 32772 13676 32824 13728
rect 32956 13676 33008 13728
rect 36268 13676 36320 13728
rect 38384 13787 38436 13796
rect 38384 13753 38393 13787
rect 38393 13753 38427 13787
rect 38427 13753 38436 13787
rect 41420 13957 41429 13991
rect 41429 13957 41463 13991
rect 41463 13957 41472 13991
rect 41420 13948 41472 13957
rect 42156 13991 42208 14000
rect 42156 13957 42165 13991
rect 42165 13957 42199 13991
rect 42199 13957 42208 13991
rect 42156 13948 42208 13957
rect 42984 14025 42993 14059
rect 42993 14025 43027 14059
rect 43027 14025 43036 14059
rect 42984 14016 43036 14025
rect 43904 13923 43956 13932
rect 43904 13889 43913 13923
rect 43913 13889 43947 13923
rect 43947 13889 43956 13923
rect 43904 13880 43956 13889
rect 38384 13744 38436 13753
rect 41604 13744 41656 13796
rect 42616 13676 42668 13728
rect 43536 13719 43588 13728
rect 43536 13685 43545 13719
rect 43545 13685 43579 13719
rect 43579 13685 43588 13719
rect 43536 13676 43588 13685
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 10508 13515 10560 13524
rect 7104 13447 7156 13456
rect 7104 13413 7113 13447
rect 7113 13413 7147 13447
rect 7147 13413 7156 13447
rect 7104 13404 7156 13413
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 10508 13481 10517 13515
rect 10517 13481 10551 13515
rect 10551 13481 10560 13515
rect 10508 13472 10560 13481
rect 12716 13472 12768 13524
rect 15108 13472 15160 13524
rect 16764 13472 16816 13524
rect 18328 13472 18380 13524
rect 21456 13472 21508 13524
rect 23112 13472 23164 13524
rect 23756 13472 23808 13524
rect 25320 13472 25372 13524
rect 29184 13472 29236 13524
rect 29460 13472 29512 13524
rect 31576 13515 31628 13524
rect 31576 13481 31585 13515
rect 31585 13481 31619 13515
rect 31619 13481 31628 13515
rect 31576 13472 31628 13481
rect 31760 13472 31812 13524
rect 36728 13472 36780 13524
rect 11244 13447 11296 13456
rect 11244 13413 11253 13447
rect 11253 13413 11287 13447
rect 11287 13413 11296 13447
rect 11244 13404 11296 13413
rect 15844 13404 15896 13456
rect 18788 13404 18840 13456
rect 21180 13447 21232 13456
rect 21180 13413 21189 13447
rect 21189 13413 21223 13447
rect 21223 13413 21232 13447
rect 21180 13404 21232 13413
rect 23480 13404 23532 13456
rect 25228 13404 25280 13456
rect 26332 13404 26384 13456
rect 32496 13404 32548 13456
rect 32864 13447 32916 13456
rect 32864 13413 32873 13447
rect 32873 13413 32907 13447
rect 32907 13413 32916 13447
rect 32864 13404 32916 13413
rect 34888 13404 34940 13456
rect 36268 13447 36320 13456
rect 36268 13413 36277 13447
rect 36277 13413 36311 13447
rect 36311 13413 36320 13447
rect 36268 13404 36320 13413
rect 39672 13404 39724 13456
rect 41604 13447 41656 13456
rect 41604 13413 41613 13447
rect 41613 13413 41647 13447
rect 41647 13413 41656 13447
rect 41604 13404 41656 13413
rect 9220 13336 9272 13388
rect 14188 13379 14240 13388
rect 14188 13345 14197 13379
rect 14197 13345 14231 13379
rect 14231 13345 14240 13379
rect 14188 13336 14240 13345
rect 18604 13336 18656 13388
rect 19248 13379 19300 13388
rect 19248 13345 19257 13379
rect 19257 13345 19291 13379
rect 19291 13345 19300 13379
rect 19248 13336 19300 13345
rect 19432 13336 19484 13388
rect 24860 13336 24912 13388
rect 26700 13336 26752 13388
rect 28816 13336 28868 13388
rect 7656 13311 7708 13320
rect 6828 13200 6880 13252
rect 7656 13277 7665 13311
rect 7665 13277 7699 13311
rect 7699 13277 7708 13311
rect 7656 13268 7708 13277
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 11152 13268 11204 13277
rect 11428 13268 11480 13320
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 11888 13268 11940 13320
rect 12440 13268 12492 13320
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 15108 13268 15160 13320
rect 15384 13311 15436 13320
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 15384 13268 15436 13277
rect 17040 13311 17092 13320
rect 14004 13200 14056 13252
rect 15568 13200 15620 13252
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 20168 13268 20220 13320
rect 21364 13268 21416 13320
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 22376 13268 22428 13320
rect 23572 13311 23624 13320
rect 23572 13277 23581 13311
rect 23581 13277 23615 13311
rect 23615 13277 23624 13311
rect 23572 13268 23624 13277
rect 24124 13268 24176 13320
rect 30564 13336 30616 13388
rect 31300 13336 31352 13388
rect 33876 13379 33928 13388
rect 33876 13345 33885 13379
rect 33885 13345 33919 13379
rect 33919 13345 33928 13379
rect 33876 13336 33928 13345
rect 33968 13336 34020 13388
rect 34520 13336 34572 13388
rect 37832 13336 37884 13388
rect 43260 13379 43312 13388
rect 43260 13345 43269 13379
rect 43269 13345 43303 13379
rect 43303 13345 43312 13379
rect 43260 13336 43312 13345
rect 32864 13268 32916 13320
rect 34796 13268 34848 13320
rect 36176 13311 36228 13320
rect 36176 13277 36185 13311
rect 36185 13277 36219 13311
rect 36219 13277 36228 13311
rect 36176 13268 36228 13277
rect 36636 13268 36688 13320
rect 37188 13268 37240 13320
rect 39580 13311 39632 13320
rect 39580 13277 39589 13311
rect 39589 13277 39623 13311
rect 39623 13277 39632 13311
rect 39580 13268 39632 13277
rect 42616 13268 42668 13320
rect 26884 13200 26936 13252
rect 31392 13200 31444 13252
rect 34336 13200 34388 13252
rect 38292 13200 38344 13252
rect 40868 13200 40920 13252
rect 41696 13200 41748 13252
rect 44180 13200 44232 13252
rect 6736 13175 6788 13184
rect 6736 13141 6745 13175
rect 6745 13141 6779 13175
rect 6779 13141 6788 13175
rect 6736 13132 6788 13141
rect 10048 13132 10100 13184
rect 14372 13175 14424 13184
rect 14372 13141 14381 13175
rect 14381 13141 14415 13175
rect 14415 13141 14424 13175
rect 14372 13132 14424 13141
rect 18052 13132 18104 13184
rect 18604 13175 18656 13184
rect 18604 13141 18613 13175
rect 18613 13141 18647 13175
rect 18647 13141 18656 13175
rect 18604 13132 18656 13141
rect 23756 13132 23808 13184
rect 25228 13132 25280 13184
rect 29736 13132 29788 13184
rect 32404 13132 32456 13184
rect 38200 13175 38252 13184
rect 38200 13141 38209 13175
rect 38209 13141 38243 13175
rect 38243 13141 38252 13175
rect 38200 13132 38252 13141
rect 40960 13132 41012 13184
rect 43168 13132 43220 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 4712 12928 4764 12980
rect 5356 12971 5408 12980
rect 5356 12937 5365 12971
rect 5365 12937 5399 12971
rect 5399 12937 5408 12971
rect 5356 12928 5408 12937
rect 6736 12928 6788 12980
rect 9220 12928 9272 12980
rect 11428 12971 11480 12980
rect 11428 12937 11437 12971
rect 11437 12937 11471 12971
rect 11471 12937 11480 12971
rect 11428 12928 11480 12937
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 15292 12971 15344 12980
rect 9128 12860 9180 12912
rect 9864 12860 9916 12912
rect 11244 12860 11296 12912
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 15844 12971 15896 12980
rect 15844 12937 15853 12971
rect 15853 12937 15887 12971
rect 15887 12937 15896 12971
rect 15844 12928 15896 12937
rect 19432 12928 19484 12980
rect 20076 12971 20128 12980
rect 20076 12937 20085 12971
rect 20085 12937 20119 12971
rect 20119 12937 20128 12971
rect 20076 12928 20128 12937
rect 21364 12971 21416 12980
rect 21364 12937 21373 12971
rect 21373 12937 21407 12971
rect 21407 12937 21416 12971
rect 21364 12928 21416 12937
rect 22376 12971 22428 12980
rect 22376 12937 22385 12971
rect 22385 12937 22419 12971
rect 22419 12937 22428 12971
rect 22376 12928 22428 12937
rect 23480 12971 23532 12980
rect 23480 12937 23489 12971
rect 23489 12937 23523 12971
rect 23523 12937 23532 12971
rect 23480 12928 23532 12937
rect 27620 12928 27672 12980
rect 30564 12971 30616 12980
rect 30564 12937 30573 12971
rect 30573 12937 30607 12971
rect 30607 12937 30616 12971
rect 30564 12928 30616 12937
rect 31300 12928 31352 12980
rect 32496 12971 32548 12980
rect 32496 12937 32505 12971
rect 32505 12937 32539 12971
rect 32539 12937 32548 12971
rect 32496 12928 32548 12937
rect 32864 12971 32916 12980
rect 32864 12937 32873 12971
rect 32873 12937 32907 12971
rect 32907 12937 32916 12971
rect 32864 12928 32916 12937
rect 33876 12928 33928 12980
rect 34336 12971 34388 12980
rect 34336 12937 34345 12971
rect 34345 12937 34379 12971
rect 34379 12937 34388 12971
rect 34336 12928 34388 12937
rect 34520 12928 34572 12980
rect 35348 12928 35400 12980
rect 36268 12928 36320 12980
rect 37832 12971 37884 12980
rect 37832 12937 37841 12971
rect 37841 12937 37875 12971
rect 37875 12937 37884 12971
rect 37832 12928 37884 12937
rect 39672 12928 39724 12980
rect 41604 12928 41656 12980
rect 42616 12928 42668 12980
rect 43260 12928 43312 12980
rect 4620 12792 4672 12844
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 11612 12792 11664 12844
rect 5356 12724 5408 12776
rect 7104 12699 7156 12708
rect 7104 12665 7113 12699
rect 7113 12665 7147 12699
rect 7147 12665 7156 12699
rect 7104 12656 7156 12665
rect 7748 12656 7800 12708
rect 9220 12699 9272 12708
rect 9220 12665 9229 12699
rect 9229 12665 9263 12699
rect 9263 12665 9272 12699
rect 9220 12656 9272 12665
rect 10140 12699 10192 12708
rect 10140 12665 10149 12699
rect 10149 12665 10183 12699
rect 10183 12665 10192 12699
rect 10140 12656 10192 12665
rect 21180 12860 21232 12912
rect 30472 12860 30524 12912
rect 32680 12860 32732 12912
rect 34704 12860 34756 12912
rect 12992 12792 13044 12844
rect 18420 12792 18472 12844
rect 20168 12835 20220 12844
rect 20168 12801 20177 12835
rect 20177 12801 20211 12835
rect 20211 12801 20220 12835
rect 20168 12792 20220 12801
rect 23756 12835 23808 12844
rect 23756 12801 23765 12835
rect 23765 12801 23799 12835
rect 23799 12801 23808 12835
rect 23756 12792 23808 12801
rect 24584 12792 24636 12844
rect 24860 12835 24912 12844
rect 24860 12801 24869 12835
rect 24869 12801 24903 12835
rect 24903 12801 24912 12835
rect 28816 12835 28868 12844
rect 24860 12792 24912 12801
rect 28816 12801 28825 12835
rect 28825 12801 28859 12835
rect 28859 12801 28868 12835
rect 28816 12792 28868 12801
rect 29920 12792 29972 12844
rect 32588 12792 32640 12844
rect 34428 12792 34480 12844
rect 15752 12724 15804 12776
rect 16948 12767 17000 12776
rect 9956 12631 10008 12640
rect 9956 12597 9965 12631
rect 9965 12597 9999 12631
rect 9999 12597 10008 12631
rect 13176 12656 13228 12708
rect 13636 12656 13688 12708
rect 13820 12656 13872 12708
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 19248 12767 19300 12776
rect 19248 12733 19257 12767
rect 19257 12733 19291 12767
rect 19291 12733 19300 12767
rect 19248 12724 19300 12733
rect 25780 12767 25832 12776
rect 18236 12656 18288 12708
rect 20076 12656 20128 12708
rect 25780 12733 25789 12767
rect 25789 12733 25823 12767
rect 25823 12733 25832 12767
rect 25780 12724 25832 12733
rect 27620 12767 27672 12776
rect 27620 12733 27629 12767
rect 27629 12733 27663 12767
rect 27663 12733 27672 12767
rect 27620 12724 27672 12733
rect 28080 12767 28132 12776
rect 28080 12733 28089 12767
rect 28089 12733 28123 12767
rect 28123 12733 28132 12767
rect 28080 12724 28132 12733
rect 33784 12724 33836 12776
rect 34336 12724 34388 12776
rect 34704 12724 34756 12776
rect 35348 12767 35400 12776
rect 35348 12733 35357 12767
rect 35357 12733 35391 12767
rect 35391 12733 35400 12767
rect 35348 12724 35400 12733
rect 23480 12656 23532 12708
rect 23940 12656 23992 12708
rect 9956 12588 10008 12597
rect 11244 12588 11296 12640
rect 14188 12631 14240 12640
rect 14188 12597 14197 12631
rect 14197 12597 14231 12631
rect 14231 12597 14240 12631
rect 14188 12588 14240 12597
rect 16764 12588 16816 12640
rect 18420 12631 18472 12640
rect 18420 12597 18429 12631
rect 18429 12597 18463 12631
rect 18463 12597 18472 12631
rect 18420 12588 18472 12597
rect 18972 12631 19024 12640
rect 18972 12597 18981 12631
rect 18981 12597 19015 12631
rect 19015 12597 19024 12631
rect 18972 12588 19024 12597
rect 22836 12588 22888 12640
rect 23112 12631 23164 12640
rect 23112 12597 23121 12631
rect 23121 12597 23155 12631
rect 23155 12597 23164 12631
rect 23112 12588 23164 12597
rect 25412 12588 25464 12640
rect 26332 12656 26384 12708
rect 28632 12656 28684 12708
rect 29736 12699 29788 12708
rect 29736 12665 29745 12699
rect 29745 12665 29779 12699
rect 29779 12665 29788 12699
rect 29736 12656 29788 12665
rect 31300 12656 31352 12708
rect 31576 12699 31628 12708
rect 31576 12665 31585 12699
rect 31585 12665 31619 12699
rect 31619 12665 31628 12699
rect 31576 12656 31628 12665
rect 31668 12699 31720 12708
rect 31668 12665 31677 12699
rect 31677 12665 31711 12699
rect 31711 12665 31720 12699
rect 31668 12656 31720 12665
rect 36544 12656 36596 12708
rect 37096 12792 37148 12844
rect 37188 12835 37240 12844
rect 37188 12801 37197 12835
rect 37197 12801 37231 12835
rect 37231 12801 37240 12835
rect 37188 12792 37240 12801
rect 41512 12860 41564 12912
rect 39580 12835 39632 12844
rect 39580 12801 39589 12835
rect 39589 12801 39623 12835
rect 39623 12801 39632 12835
rect 39580 12792 39632 12801
rect 42248 12792 42300 12844
rect 43168 12835 43220 12844
rect 43168 12801 43177 12835
rect 43177 12801 43211 12835
rect 43211 12801 43220 12835
rect 43168 12792 43220 12801
rect 39120 12724 39172 12776
rect 43996 12724 44048 12776
rect 37004 12699 37056 12708
rect 37004 12665 37013 12699
rect 37013 12665 37047 12699
rect 37047 12665 37056 12699
rect 37004 12656 37056 12665
rect 40868 12699 40920 12708
rect 40868 12665 40877 12699
rect 40877 12665 40911 12699
rect 40911 12665 40920 12699
rect 40868 12656 40920 12665
rect 40960 12699 41012 12708
rect 40960 12665 40969 12699
rect 40969 12665 41003 12699
rect 41003 12665 41012 12699
rect 40960 12656 41012 12665
rect 41880 12656 41932 12708
rect 25688 12588 25740 12640
rect 35256 12588 35308 12640
rect 43536 12588 43588 12640
rect 44456 12588 44508 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 7012 12384 7064 12436
rect 8852 12384 8904 12436
rect 10140 12384 10192 12436
rect 15108 12427 15160 12436
rect 15108 12393 15117 12427
rect 15117 12393 15151 12427
rect 15151 12393 15160 12427
rect 15108 12384 15160 12393
rect 15844 12427 15896 12436
rect 15844 12393 15853 12427
rect 15853 12393 15887 12427
rect 15887 12393 15896 12427
rect 15844 12384 15896 12393
rect 15936 12384 15988 12436
rect 16948 12384 17000 12436
rect 20352 12384 20404 12436
rect 22928 12384 22980 12436
rect 6828 12359 6880 12368
rect 6828 12325 6837 12359
rect 6837 12325 6871 12359
rect 6871 12325 6880 12359
rect 6828 12316 6880 12325
rect 7104 12359 7156 12368
rect 7104 12325 7113 12359
rect 7113 12325 7147 12359
rect 7147 12325 7156 12359
rect 7104 12316 7156 12325
rect 7656 12359 7708 12368
rect 7656 12325 7665 12359
rect 7665 12325 7699 12359
rect 7699 12325 7708 12359
rect 7656 12316 7708 12325
rect 9128 12316 9180 12368
rect 9772 12359 9824 12368
rect 9772 12325 9781 12359
rect 9781 12325 9815 12359
rect 9815 12325 9824 12359
rect 9772 12316 9824 12325
rect 9864 12359 9916 12368
rect 9864 12325 9873 12359
rect 9873 12325 9907 12359
rect 9907 12325 9916 12359
rect 9864 12316 9916 12325
rect 11612 12316 11664 12368
rect 12808 12359 12860 12368
rect 12808 12325 12817 12359
rect 12817 12325 12851 12359
rect 12851 12325 12860 12359
rect 12808 12316 12860 12325
rect 13176 12316 13228 12368
rect 17040 12316 17092 12368
rect 17868 12359 17920 12368
rect 17868 12325 17877 12359
rect 17877 12325 17911 12359
rect 17911 12325 17920 12359
rect 17868 12316 17920 12325
rect 17960 12359 18012 12368
rect 17960 12325 17969 12359
rect 17969 12325 18003 12359
rect 18003 12325 18012 12359
rect 17960 12316 18012 12325
rect 18972 12316 19024 12368
rect 20260 12359 20312 12368
rect 20260 12325 20269 12359
rect 20269 12325 20303 12359
rect 20303 12325 20312 12359
rect 20260 12316 20312 12325
rect 21088 12359 21140 12368
rect 21088 12325 21097 12359
rect 21097 12325 21131 12359
rect 21131 12325 21140 12359
rect 21088 12316 21140 12325
rect 22836 12316 22888 12368
rect 24032 12384 24084 12436
rect 24584 12384 24636 12436
rect 26700 12384 26752 12436
rect 28080 12384 28132 12436
rect 28908 12384 28960 12436
rect 29736 12384 29788 12436
rect 29920 12427 29972 12436
rect 29920 12393 29929 12427
rect 29929 12393 29963 12427
rect 29963 12393 29972 12427
rect 29920 12384 29972 12393
rect 31668 12384 31720 12436
rect 34704 12384 34756 12436
rect 36176 12427 36228 12436
rect 36176 12393 36185 12427
rect 36185 12393 36219 12427
rect 36219 12393 36228 12427
rect 36176 12384 36228 12393
rect 38200 12384 38252 12436
rect 39120 12384 39172 12436
rect 43168 12427 43220 12436
rect 23940 12359 23992 12368
rect 23940 12325 23949 12359
rect 23949 12325 23983 12359
rect 23983 12325 23992 12359
rect 23940 12316 23992 12325
rect 24400 12316 24452 12368
rect 25228 12316 25280 12368
rect 25872 12316 25924 12368
rect 5448 12248 5500 12300
rect 6092 12248 6144 12300
rect 8576 12248 8628 12300
rect 15384 12248 15436 12300
rect 18880 12248 18932 12300
rect 19156 12248 19208 12300
rect 26608 12248 26660 12300
rect 27620 12316 27672 12368
rect 30564 12359 30616 12368
rect 30564 12325 30573 12359
rect 30573 12325 30607 12359
rect 30607 12325 30616 12359
rect 30564 12316 30616 12325
rect 32036 12316 32088 12368
rect 34428 12359 34480 12368
rect 34428 12325 34437 12359
rect 34437 12325 34471 12359
rect 34471 12325 34480 12359
rect 34428 12316 34480 12325
rect 34796 12316 34848 12368
rect 35164 12316 35216 12368
rect 39672 12316 39724 12368
rect 39948 12316 40000 12368
rect 40868 12359 40920 12368
rect 40868 12325 40877 12359
rect 40877 12325 40911 12359
rect 40911 12325 40920 12359
rect 40868 12316 40920 12325
rect 43168 12393 43177 12427
rect 43177 12393 43211 12427
rect 43211 12393 43220 12427
rect 43168 12384 43220 12393
rect 42248 12316 42300 12368
rect 43536 12359 43588 12368
rect 43536 12325 43545 12359
rect 43545 12325 43579 12359
rect 43579 12325 43588 12359
rect 43536 12316 43588 12325
rect 44180 12316 44232 12368
rect 26976 12291 27028 12300
rect 26976 12257 26985 12291
rect 26985 12257 27019 12291
rect 27019 12257 27028 12291
rect 26976 12248 27028 12257
rect 31300 12248 31352 12300
rect 36084 12248 36136 12300
rect 36728 12248 36780 12300
rect 38016 12248 38068 12300
rect 7012 12223 7064 12232
rect 7012 12189 7021 12223
rect 7021 12189 7055 12223
rect 7055 12189 7064 12223
rect 7012 12180 7064 12189
rect 9220 12180 9272 12232
rect 12164 12180 12216 12232
rect 14280 12180 14332 12232
rect 20996 12223 21048 12232
rect 20996 12189 21005 12223
rect 21005 12189 21039 12223
rect 21039 12189 21048 12223
rect 20996 12180 21048 12189
rect 25780 12180 25832 12232
rect 28632 12223 28684 12232
rect 28632 12189 28641 12223
rect 28641 12189 28675 12223
rect 28675 12189 28684 12223
rect 28632 12180 28684 12189
rect 30472 12223 30524 12232
rect 30472 12189 30481 12223
rect 30481 12189 30515 12223
rect 30515 12189 30524 12223
rect 30472 12180 30524 12189
rect 32220 12223 32272 12232
rect 32220 12189 32229 12223
rect 32229 12189 32263 12223
rect 32263 12189 32272 12223
rect 32220 12180 32272 12189
rect 32588 12223 32640 12232
rect 32588 12189 32597 12223
rect 32597 12189 32631 12223
rect 32631 12189 32640 12223
rect 32588 12180 32640 12189
rect 39672 12223 39724 12232
rect 18420 12155 18472 12164
rect 18420 12121 18429 12155
rect 18429 12121 18463 12155
rect 18463 12121 18472 12155
rect 18420 12112 18472 12121
rect 21548 12155 21600 12164
rect 21548 12121 21557 12155
rect 21557 12121 21591 12155
rect 21591 12121 21600 12155
rect 21548 12112 21600 12121
rect 34244 12112 34296 12164
rect 39672 12189 39681 12223
rect 39681 12189 39715 12223
rect 39715 12189 39724 12223
rect 39672 12180 39724 12189
rect 40776 12180 40828 12232
rect 41512 12223 41564 12232
rect 41512 12189 41521 12223
rect 41521 12189 41555 12223
rect 41555 12189 41564 12223
rect 41512 12180 41564 12189
rect 41880 12223 41932 12232
rect 41880 12189 41889 12223
rect 41889 12189 41923 12223
rect 41923 12189 41932 12223
rect 41880 12180 41932 12189
rect 44456 12180 44508 12232
rect 41328 12155 41380 12164
rect 41328 12121 41337 12155
rect 41337 12121 41371 12155
rect 41371 12121 41380 12155
rect 41328 12112 41380 12121
rect 42156 12112 42208 12164
rect 43352 12112 43404 12164
rect 11612 12087 11664 12096
rect 11612 12053 11621 12087
rect 11621 12053 11655 12087
rect 11655 12053 11664 12087
rect 11612 12044 11664 12053
rect 13268 12044 13320 12096
rect 14096 12044 14148 12096
rect 23204 12044 23256 12096
rect 31576 12044 31628 12096
rect 33784 12044 33836 12096
rect 36912 12044 36964 12096
rect 37096 12087 37148 12096
rect 37096 12053 37105 12087
rect 37105 12053 37139 12087
rect 37139 12053 37148 12087
rect 37096 12044 37148 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 7012 11840 7064 11892
rect 8576 11883 8628 11892
rect 8576 11849 8585 11883
rect 8585 11849 8619 11883
rect 8619 11849 8628 11883
rect 8576 11840 8628 11849
rect 9772 11840 9824 11892
rect 6092 11815 6144 11824
rect 6092 11781 6101 11815
rect 6101 11781 6135 11815
rect 6135 11781 6144 11815
rect 6092 11772 6144 11781
rect 7104 11815 7156 11824
rect 7104 11781 7113 11815
rect 7113 11781 7147 11815
rect 7147 11781 7156 11815
rect 7104 11772 7156 11781
rect 9864 11704 9916 11756
rect 5540 11636 5592 11688
rect 11520 11840 11572 11892
rect 12808 11840 12860 11892
rect 14188 11840 14240 11892
rect 14372 11840 14424 11892
rect 17868 11883 17920 11892
rect 11612 11772 11664 11824
rect 14832 11772 14884 11824
rect 14096 11704 14148 11756
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 18328 11840 18380 11892
rect 19340 11840 19392 11892
rect 20076 11840 20128 11892
rect 21088 11840 21140 11892
rect 24124 11840 24176 11892
rect 26608 11883 26660 11892
rect 26608 11849 26617 11883
rect 26617 11849 26651 11883
rect 26651 11849 26660 11883
rect 26608 11840 26660 11849
rect 30564 11883 30616 11892
rect 30564 11849 30573 11883
rect 30573 11849 30607 11883
rect 30607 11849 30616 11883
rect 30564 11840 30616 11849
rect 32036 11840 32088 11892
rect 34428 11840 34480 11892
rect 38016 11883 38068 11892
rect 38016 11849 38025 11883
rect 38025 11849 38059 11883
rect 38059 11849 38068 11883
rect 38016 11840 38068 11849
rect 38660 11883 38712 11892
rect 38660 11849 38669 11883
rect 38669 11849 38703 11883
rect 38703 11849 38712 11883
rect 38660 11840 38712 11849
rect 39948 11883 40000 11892
rect 39948 11849 39957 11883
rect 39957 11849 39991 11883
rect 39991 11849 40000 11883
rect 39948 11840 40000 11849
rect 40776 11883 40828 11892
rect 40776 11849 40785 11883
rect 40785 11849 40819 11883
rect 40819 11849 40828 11883
rect 40776 11840 40828 11849
rect 42248 11883 42300 11892
rect 42248 11849 42257 11883
rect 42257 11849 42291 11883
rect 42291 11849 42300 11883
rect 42248 11840 42300 11849
rect 43076 11840 43128 11892
rect 44456 11883 44508 11892
rect 17960 11772 18012 11824
rect 23572 11772 23624 11824
rect 20260 11704 20312 11756
rect 21364 11704 21416 11756
rect 24032 11747 24084 11756
rect 24032 11713 24041 11747
rect 24041 11713 24075 11747
rect 24075 11713 24084 11747
rect 24032 11704 24084 11713
rect 25504 11772 25556 11824
rect 30472 11772 30524 11824
rect 36728 11815 36780 11824
rect 36728 11781 36737 11815
rect 36737 11781 36771 11815
rect 36771 11781 36780 11815
rect 41880 11815 41932 11824
rect 36728 11772 36780 11781
rect 41880 11781 41889 11815
rect 41889 11781 41923 11815
rect 41923 11781 41932 11815
rect 41880 11772 41932 11781
rect 44456 11849 44465 11883
rect 44465 11849 44499 11883
rect 44499 11849 44508 11883
rect 44456 11840 44508 11849
rect 25872 11704 25924 11756
rect 32220 11704 32272 11756
rect 35256 11747 35308 11756
rect 35256 11713 35265 11747
rect 35265 11713 35299 11747
rect 35299 11713 35308 11747
rect 35256 11704 35308 11713
rect 36544 11704 36596 11756
rect 37464 11704 37516 11756
rect 37924 11704 37976 11756
rect 38476 11704 38528 11756
rect 39672 11704 39724 11756
rect 41328 11747 41380 11756
rect 41328 11713 41337 11747
rect 41337 11713 41371 11747
rect 41371 11713 41380 11747
rect 41328 11704 41380 11713
rect 41696 11704 41748 11756
rect 43076 11747 43128 11756
rect 43076 11713 43085 11747
rect 43085 11713 43119 11747
rect 43119 11713 43128 11747
rect 43076 11704 43128 11713
rect 43352 11747 43404 11756
rect 43352 11713 43361 11747
rect 43361 11713 43395 11747
rect 43395 11713 43404 11747
rect 43352 11704 43404 11713
rect 17684 11636 17736 11688
rect 18420 11636 18472 11688
rect 21548 11636 21600 11688
rect 27528 11679 27580 11688
rect 27528 11645 27537 11679
rect 27537 11645 27571 11679
rect 27571 11645 27580 11679
rect 27804 11679 27856 11688
rect 27528 11636 27580 11645
rect 27804 11645 27813 11679
rect 27813 11645 27847 11679
rect 27847 11645 27856 11679
rect 27804 11636 27856 11645
rect 28080 11679 28132 11688
rect 28080 11645 28089 11679
rect 28089 11645 28123 11679
rect 28123 11645 28132 11679
rect 28080 11636 28132 11645
rect 29276 11679 29328 11688
rect 29276 11645 29285 11679
rect 29285 11645 29319 11679
rect 29319 11645 29328 11679
rect 29276 11636 29328 11645
rect 31208 11636 31260 11688
rect 31760 11679 31812 11688
rect 31760 11645 31769 11679
rect 31769 11645 31803 11679
rect 31803 11645 31812 11679
rect 31760 11636 31812 11645
rect 33232 11679 33284 11688
rect 33232 11645 33241 11679
rect 33241 11645 33275 11679
rect 33275 11645 33284 11679
rect 33232 11636 33284 11645
rect 14004 11611 14056 11620
rect 14004 11577 14013 11611
rect 14013 11577 14047 11611
rect 14047 11577 14056 11611
rect 14004 11568 14056 11577
rect 10232 11500 10284 11552
rect 12256 11543 12308 11552
rect 12256 11509 12265 11543
rect 12265 11509 12299 11543
rect 12299 11509 12308 11543
rect 12256 11500 12308 11509
rect 13176 11500 13228 11552
rect 13360 11500 13412 11552
rect 24124 11611 24176 11620
rect 24124 11577 24133 11611
rect 24133 11577 24167 11611
rect 24167 11577 24176 11611
rect 24124 11568 24176 11577
rect 25688 11611 25740 11620
rect 25688 11577 25697 11611
rect 25697 11577 25731 11611
rect 25731 11577 25740 11611
rect 25688 11568 25740 11577
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 18880 11500 18932 11552
rect 20076 11543 20128 11552
rect 20076 11509 20085 11543
rect 20085 11509 20119 11543
rect 20119 11509 20128 11543
rect 20076 11500 20128 11509
rect 20444 11500 20496 11552
rect 20996 11500 21048 11552
rect 22928 11500 22980 11552
rect 25228 11500 25280 11552
rect 26700 11500 26752 11552
rect 28908 11500 28960 11552
rect 33968 11636 34020 11688
rect 38660 11636 38712 11688
rect 39120 11636 39172 11688
rect 33508 11543 33560 11552
rect 33508 11509 33517 11543
rect 33517 11509 33551 11543
rect 33551 11509 33560 11543
rect 33508 11500 33560 11509
rect 34244 11543 34296 11552
rect 34244 11509 34253 11543
rect 34253 11509 34287 11543
rect 34287 11509 34296 11543
rect 34244 11500 34296 11509
rect 35072 11543 35124 11552
rect 35072 11509 35081 11543
rect 35081 11509 35115 11543
rect 35115 11509 35124 11543
rect 35072 11500 35124 11509
rect 36176 11543 36228 11552
rect 36176 11509 36185 11543
rect 36185 11509 36219 11543
rect 36219 11509 36228 11543
rect 36176 11500 36228 11509
rect 37004 11500 37056 11552
rect 37740 11500 37792 11552
rect 41512 11568 41564 11620
rect 42892 11543 42944 11552
rect 42892 11509 42901 11543
rect 42901 11509 42935 11543
rect 42935 11509 42944 11543
rect 42892 11500 42944 11509
rect 43536 11500 43588 11552
rect 44180 11500 44232 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 9864 11160 9916 11212
rect 10048 11296 10100 11348
rect 13820 11296 13872 11348
rect 14004 11339 14056 11348
rect 14004 11305 14013 11339
rect 14013 11305 14047 11339
rect 14047 11305 14056 11339
rect 14004 11296 14056 11305
rect 19064 11339 19116 11348
rect 19064 11305 19073 11339
rect 19073 11305 19107 11339
rect 19107 11305 19116 11339
rect 19064 11296 19116 11305
rect 22836 11296 22888 11348
rect 24400 11296 24452 11348
rect 25872 11339 25924 11348
rect 11428 11271 11480 11280
rect 11428 11237 11437 11271
rect 11437 11237 11471 11271
rect 11471 11237 11480 11271
rect 11428 11228 11480 11237
rect 12164 11228 12216 11280
rect 13360 11228 13412 11280
rect 13636 11271 13688 11280
rect 13636 11237 13645 11271
rect 13645 11237 13679 11271
rect 13679 11237 13688 11271
rect 13636 11228 13688 11237
rect 17132 11271 17184 11280
rect 17132 11237 17141 11271
rect 17141 11237 17175 11271
rect 17175 11237 17184 11271
rect 17132 11228 17184 11237
rect 19156 11228 19208 11280
rect 23388 11271 23440 11280
rect 10232 11203 10284 11212
rect 10232 11169 10241 11203
rect 10241 11169 10275 11203
rect 10275 11169 10284 11203
rect 10232 11160 10284 11169
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 15936 11203 15988 11212
rect 15936 11169 15945 11203
rect 15945 11169 15979 11203
rect 15979 11169 15988 11203
rect 15936 11160 15988 11169
rect 18788 11160 18840 11212
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 23388 11237 23397 11271
rect 23397 11237 23431 11271
rect 23431 11237 23440 11271
rect 23388 11228 23440 11237
rect 23572 11228 23624 11280
rect 25872 11305 25881 11339
rect 25881 11305 25915 11339
rect 25915 11305 25924 11339
rect 25872 11296 25924 11305
rect 26976 11296 27028 11348
rect 28632 11296 28684 11348
rect 29276 11296 29328 11348
rect 30748 11296 30800 11348
rect 32772 11296 32824 11348
rect 34428 11296 34480 11348
rect 35256 11339 35308 11348
rect 35256 11305 35265 11339
rect 35265 11305 35299 11339
rect 35299 11305 35308 11339
rect 35256 11296 35308 11305
rect 37004 11296 37056 11348
rect 37464 11339 37516 11348
rect 37464 11305 37473 11339
rect 37473 11305 37507 11339
rect 37507 11305 37516 11339
rect 37464 11296 37516 11305
rect 37740 11296 37792 11348
rect 26700 11228 26752 11280
rect 29920 11271 29972 11280
rect 29920 11237 29929 11271
rect 29929 11237 29963 11271
rect 29963 11237 29972 11271
rect 29920 11228 29972 11237
rect 32036 11228 32088 11280
rect 33600 11228 33652 11280
rect 35072 11228 35124 11280
rect 36176 11228 36228 11280
rect 36912 11228 36964 11280
rect 37832 11271 37884 11280
rect 37832 11237 37841 11271
rect 37841 11237 37875 11271
rect 37875 11237 37884 11271
rect 37832 11228 37884 11237
rect 39120 11296 39172 11348
rect 43076 11339 43128 11348
rect 43076 11305 43085 11339
rect 43085 11305 43119 11339
rect 43119 11305 43128 11339
rect 43076 11296 43128 11305
rect 41420 11271 41472 11280
rect 21456 11160 21508 11212
rect 22928 11160 22980 11212
rect 27160 11160 27212 11212
rect 28724 11160 28776 11212
rect 33508 11160 33560 11212
rect 39304 11203 39356 11212
rect 39304 11169 39313 11203
rect 39313 11169 39347 11203
rect 39347 11169 39356 11203
rect 39304 11160 39356 11169
rect 41420 11237 41429 11271
rect 41429 11237 41463 11271
rect 41463 11237 41472 11271
rect 41420 11228 41472 11237
rect 44180 11228 44232 11280
rect 10324 11092 10376 11144
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 16120 11135 16172 11144
rect 10140 11024 10192 11076
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 16672 11092 16724 11144
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 22284 11135 22336 11144
rect 22284 11101 22293 11135
rect 22293 11101 22327 11135
rect 22327 11101 22336 11135
rect 22284 11092 22336 11101
rect 23480 11092 23532 11144
rect 26516 11135 26568 11144
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 29828 11135 29880 11144
rect 29828 11101 29837 11135
rect 29837 11101 29871 11135
rect 29871 11101 29880 11135
rect 29828 11092 29880 11101
rect 12256 11024 12308 11076
rect 13084 11024 13136 11076
rect 24124 11024 24176 11076
rect 28724 11024 28776 11076
rect 31944 11092 31996 11144
rect 32312 11092 32364 11144
rect 36912 11092 36964 11144
rect 37188 11092 37240 11144
rect 40040 11135 40092 11144
rect 31300 11024 31352 11076
rect 36728 11067 36780 11076
rect 36728 11033 36737 11067
rect 36737 11033 36771 11067
rect 36771 11033 36780 11067
rect 36728 11024 36780 11033
rect 36820 11024 36872 11076
rect 40040 11101 40049 11135
rect 40049 11101 40083 11135
rect 40083 11101 40092 11135
rect 40040 11092 40092 11101
rect 41328 11135 41380 11144
rect 41328 11101 41337 11135
rect 41337 11101 41371 11135
rect 41371 11101 41380 11135
rect 43444 11135 43496 11144
rect 41328 11092 41380 11101
rect 41880 11067 41932 11076
rect 41880 11033 41889 11067
rect 41889 11033 41923 11067
rect 41923 11033 41932 11067
rect 41880 11024 41932 11033
rect 43444 11101 43453 11135
rect 43453 11101 43487 11135
rect 43487 11101 43496 11135
rect 43444 11092 43496 11101
rect 43720 11135 43772 11144
rect 43720 11101 43729 11135
rect 43729 11101 43763 11135
rect 43763 11101 43772 11135
rect 43720 11092 43772 11101
rect 19984 10999 20036 11008
rect 19984 10965 19993 10999
rect 19993 10965 20027 10999
rect 20027 10965 20036 10999
rect 19984 10956 20036 10965
rect 25136 10999 25188 11008
rect 25136 10965 25145 10999
rect 25145 10965 25179 10999
rect 25179 10965 25188 10999
rect 25136 10956 25188 10965
rect 26332 10956 26384 11008
rect 33232 10999 33284 11008
rect 33232 10965 33241 10999
rect 33241 10965 33275 10999
rect 33275 10965 33284 10999
rect 33232 10956 33284 10965
rect 38660 10956 38712 11008
rect 39028 10956 39080 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 9864 10795 9916 10804
rect 9864 10761 9873 10795
rect 9873 10761 9907 10795
rect 9907 10761 9916 10795
rect 9864 10752 9916 10761
rect 11428 10752 11480 10804
rect 12164 10795 12216 10804
rect 12164 10761 12173 10795
rect 12173 10761 12207 10795
rect 12207 10761 12216 10795
rect 12164 10752 12216 10761
rect 13360 10752 13412 10804
rect 15016 10752 15068 10804
rect 16672 10752 16724 10804
rect 17132 10795 17184 10804
rect 17132 10761 17141 10795
rect 17141 10761 17175 10795
rect 17175 10761 17184 10795
rect 17132 10752 17184 10761
rect 17500 10752 17552 10804
rect 18788 10752 18840 10804
rect 21456 10795 21508 10804
rect 21456 10761 21465 10795
rect 21465 10761 21499 10795
rect 21499 10761 21508 10795
rect 21456 10752 21508 10761
rect 25228 10752 25280 10804
rect 26516 10752 26568 10804
rect 27620 10752 27672 10804
rect 28724 10795 28776 10804
rect 28724 10761 28733 10795
rect 28733 10761 28767 10795
rect 28767 10761 28776 10795
rect 28724 10752 28776 10761
rect 29828 10752 29880 10804
rect 29920 10752 29972 10804
rect 32036 10752 32088 10804
rect 33508 10752 33560 10804
rect 33784 10752 33836 10804
rect 34336 10795 34388 10804
rect 34336 10761 34345 10795
rect 34345 10761 34379 10795
rect 34379 10761 34388 10795
rect 34336 10752 34388 10761
rect 36176 10795 36228 10804
rect 36176 10761 36185 10795
rect 36185 10761 36219 10795
rect 36219 10761 36228 10795
rect 36176 10752 36228 10761
rect 37740 10795 37792 10804
rect 37740 10761 37749 10795
rect 37749 10761 37783 10795
rect 37783 10761 37792 10795
rect 37740 10752 37792 10761
rect 37832 10752 37884 10804
rect 38660 10795 38712 10804
rect 38660 10761 38669 10795
rect 38669 10761 38703 10795
rect 38703 10761 38712 10795
rect 38660 10752 38712 10761
rect 39304 10752 39356 10804
rect 41420 10752 41472 10804
rect 42892 10795 42944 10804
rect 42892 10761 42901 10795
rect 42901 10761 42935 10795
rect 42935 10761 42944 10795
rect 42892 10752 42944 10761
rect 43444 10795 43496 10804
rect 43444 10761 43453 10795
rect 43453 10761 43487 10795
rect 43487 10761 43496 10795
rect 44180 10795 44232 10804
rect 43444 10752 43496 10761
rect 15936 10684 15988 10736
rect 10324 10659 10376 10668
rect 10324 10625 10333 10659
rect 10333 10625 10367 10659
rect 10367 10625 10376 10659
rect 10324 10616 10376 10625
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 16120 10616 16172 10668
rect 11336 10548 11388 10600
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 15016 10548 15068 10600
rect 15660 10548 15712 10600
rect 23388 10684 23440 10736
rect 31300 10727 31352 10736
rect 31300 10693 31309 10727
rect 31309 10693 31343 10727
rect 31343 10693 31352 10727
rect 31300 10684 31352 10693
rect 33692 10684 33744 10736
rect 18236 10616 18288 10668
rect 18052 10548 18104 10600
rect 22284 10616 22336 10668
rect 19432 10548 19484 10600
rect 19984 10548 20036 10600
rect 23572 10548 23624 10600
rect 23756 10591 23808 10600
rect 23756 10557 23774 10591
rect 23774 10557 23808 10591
rect 23756 10548 23808 10557
rect 25136 10548 25188 10600
rect 26148 10548 26200 10600
rect 26884 10591 26936 10600
rect 26884 10557 26893 10591
rect 26893 10557 26927 10591
rect 26927 10557 26936 10591
rect 26884 10548 26936 10557
rect 26976 10548 27028 10600
rect 27252 10591 27304 10600
rect 27252 10557 27261 10591
rect 27261 10557 27295 10591
rect 27295 10557 27304 10591
rect 27252 10548 27304 10557
rect 31944 10616 31996 10668
rect 32772 10659 32824 10668
rect 32772 10625 32781 10659
rect 32781 10625 32815 10659
rect 32815 10625 32824 10659
rect 32772 10616 32824 10625
rect 34796 10616 34848 10668
rect 36728 10684 36780 10736
rect 36820 10659 36872 10668
rect 36820 10625 36829 10659
rect 36829 10625 36863 10659
rect 36863 10625 36872 10659
rect 36820 10616 36872 10625
rect 39948 10684 40000 10736
rect 38108 10616 38160 10668
rect 40040 10616 40092 10668
rect 41972 10659 42024 10668
rect 41972 10625 41981 10659
rect 41981 10625 42015 10659
rect 42015 10625 42024 10659
rect 41972 10616 42024 10625
rect 30196 10591 30248 10600
rect 30196 10557 30205 10591
rect 30205 10557 30239 10591
rect 30239 10557 30248 10591
rect 30196 10548 30248 10557
rect 34336 10548 34388 10600
rect 38660 10548 38712 10600
rect 39120 10548 39172 10600
rect 41880 10548 41932 10600
rect 10232 10480 10284 10532
rect 10508 10480 10560 10532
rect 13544 10480 13596 10532
rect 16672 10480 16724 10532
rect 20076 10523 20128 10532
rect 20076 10489 20085 10523
rect 20085 10489 20119 10523
rect 20119 10489 20128 10523
rect 20076 10480 20128 10489
rect 22928 10480 22980 10532
rect 23480 10480 23532 10532
rect 30748 10523 30800 10532
rect 30748 10489 30757 10523
rect 30757 10489 30791 10523
rect 30791 10489 30800 10523
rect 30748 10480 30800 10489
rect 30840 10523 30892 10532
rect 30840 10489 30849 10523
rect 30849 10489 30883 10523
rect 30883 10489 30892 10523
rect 32128 10523 32180 10532
rect 30840 10480 30892 10489
rect 32128 10489 32137 10523
rect 32137 10489 32171 10523
rect 32171 10489 32180 10523
rect 32128 10480 32180 10489
rect 39580 10523 39632 10532
rect 20996 10455 21048 10464
rect 20996 10421 21005 10455
rect 21005 10421 21039 10455
rect 21039 10421 21048 10455
rect 20996 10412 21048 10421
rect 23388 10412 23440 10464
rect 24676 10412 24728 10464
rect 25412 10455 25464 10464
rect 25412 10421 25421 10455
rect 25421 10421 25455 10455
rect 25455 10421 25464 10455
rect 25412 10412 25464 10421
rect 26700 10412 26752 10464
rect 26884 10455 26936 10464
rect 26884 10421 26893 10455
rect 26893 10421 26927 10455
rect 26927 10421 26936 10455
rect 26884 10412 26936 10421
rect 32036 10412 32088 10464
rect 32588 10412 32640 10464
rect 33140 10412 33192 10464
rect 33600 10455 33652 10464
rect 33600 10421 33609 10455
rect 33609 10421 33643 10455
rect 33643 10421 33652 10455
rect 33600 10412 33652 10421
rect 34612 10455 34664 10464
rect 34612 10421 34621 10455
rect 34621 10421 34655 10455
rect 34655 10421 34664 10455
rect 34612 10412 34664 10421
rect 36728 10412 36780 10464
rect 39580 10489 39589 10523
rect 39589 10489 39623 10523
rect 39623 10489 39632 10523
rect 39580 10480 39632 10489
rect 44180 10761 44189 10795
rect 44189 10761 44223 10795
rect 44223 10761 44232 10795
rect 44180 10752 44232 10761
rect 40500 10412 40552 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 11428 10208 11480 10260
rect 11796 10251 11848 10260
rect 11796 10217 11805 10251
rect 11805 10217 11839 10251
rect 11839 10217 11848 10251
rect 11796 10208 11848 10217
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 13636 10208 13688 10260
rect 15384 10208 15436 10260
rect 16120 10208 16172 10260
rect 18052 10251 18104 10260
rect 18052 10217 18061 10251
rect 18061 10217 18095 10251
rect 18095 10217 18104 10251
rect 18052 10208 18104 10217
rect 19064 10208 19116 10260
rect 23572 10208 23624 10260
rect 27160 10251 27212 10260
rect 27160 10217 27169 10251
rect 27169 10217 27203 10251
rect 27203 10217 27212 10251
rect 27160 10208 27212 10217
rect 27252 10208 27304 10260
rect 28908 10208 28960 10260
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 10232 10072 10284 10124
rect 13820 10183 13872 10192
rect 13820 10149 13829 10183
rect 13829 10149 13863 10183
rect 13863 10149 13872 10183
rect 13820 10140 13872 10149
rect 16672 10140 16724 10192
rect 11704 10115 11756 10124
rect 11704 10081 11713 10115
rect 11713 10081 11747 10115
rect 11747 10081 11756 10115
rect 11704 10072 11756 10081
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 19156 10140 19208 10192
rect 19340 10140 19392 10192
rect 19984 10140 20036 10192
rect 22928 10140 22980 10192
rect 24676 10140 24728 10192
rect 24952 10183 25004 10192
rect 24952 10149 24961 10183
rect 24961 10149 24995 10183
rect 24995 10149 25004 10183
rect 24952 10140 25004 10149
rect 25504 10183 25556 10192
rect 25504 10149 25513 10183
rect 25513 10149 25547 10183
rect 25547 10149 25556 10183
rect 25504 10140 25556 10149
rect 26792 10183 26844 10192
rect 26792 10149 26801 10183
rect 26801 10149 26835 10183
rect 26835 10149 26844 10183
rect 26792 10140 26844 10149
rect 30840 10251 30892 10260
rect 30840 10217 30849 10251
rect 30849 10217 30883 10251
rect 30883 10217 30892 10251
rect 30840 10208 30892 10217
rect 32128 10251 32180 10260
rect 32128 10217 32137 10251
rect 32137 10217 32171 10251
rect 32171 10217 32180 10251
rect 32128 10208 32180 10217
rect 32588 10251 32640 10260
rect 32588 10217 32597 10251
rect 32597 10217 32631 10251
rect 32631 10217 32640 10251
rect 32588 10208 32640 10217
rect 34612 10208 34664 10260
rect 34796 10208 34848 10260
rect 36084 10251 36136 10260
rect 36084 10217 36093 10251
rect 36093 10217 36127 10251
rect 36127 10217 36136 10251
rect 36084 10208 36136 10217
rect 37740 10208 37792 10260
rect 31944 10140 31996 10192
rect 33140 10140 33192 10192
rect 36912 10183 36964 10192
rect 36912 10149 36921 10183
rect 36921 10149 36955 10183
rect 36955 10149 36964 10183
rect 36912 10140 36964 10149
rect 39120 10208 39172 10260
rect 41420 10208 41472 10260
rect 41972 10251 42024 10260
rect 41972 10217 41981 10251
rect 41981 10217 42015 10251
rect 42015 10217 42024 10251
rect 41972 10208 42024 10217
rect 39948 10140 40000 10192
rect 41328 10183 41380 10192
rect 41328 10149 41337 10183
rect 41337 10149 41371 10183
rect 41371 10149 41380 10183
rect 41328 10140 41380 10149
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 27068 10072 27120 10124
rect 15844 10004 15896 10056
rect 16488 10004 16540 10056
rect 20076 10004 20128 10056
rect 22468 10004 22520 10056
rect 23020 10047 23072 10056
rect 23020 10013 23029 10047
rect 23029 10013 23063 10047
rect 23063 10013 23072 10047
rect 23020 10004 23072 10013
rect 23664 10004 23716 10056
rect 24860 10047 24912 10056
rect 24860 10013 24869 10047
rect 24869 10013 24903 10047
rect 24903 10013 24912 10047
rect 24860 10004 24912 10013
rect 11704 9936 11756 9988
rect 13912 9936 13964 9988
rect 14280 9979 14332 9988
rect 14280 9945 14289 9979
rect 14289 9945 14323 9979
rect 14323 9945 14332 9979
rect 14280 9936 14332 9945
rect 17592 9911 17644 9920
rect 17592 9877 17601 9911
rect 17601 9877 17635 9911
rect 17635 9877 17644 9911
rect 17592 9868 17644 9877
rect 21272 9868 21324 9920
rect 21364 9868 21416 9920
rect 23020 9868 23072 9920
rect 26884 9936 26936 9988
rect 28080 10072 28132 10124
rect 28448 10115 28500 10124
rect 28448 10081 28457 10115
rect 28457 10081 28491 10115
rect 28491 10081 28500 10115
rect 28448 10072 28500 10081
rect 31760 10072 31812 10124
rect 36544 10072 36596 10124
rect 36820 10072 36872 10124
rect 39580 10072 39632 10124
rect 40132 10115 40184 10124
rect 40132 10081 40141 10115
rect 40141 10081 40175 10115
rect 40175 10081 40184 10115
rect 40132 10072 40184 10081
rect 28724 10047 28776 10056
rect 28724 10013 28733 10047
rect 28733 10013 28767 10047
rect 28767 10013 28776 10047
rect 28724 10004 28776 10013
rect 29552 10047 29604 10056
rect 29552 10013 29561 10047
rect 29561 10013 29595 10047
rect 29595 10013 29604 10047
rect 29552 10004 29604 10013
rect 33784 10004 33836 10056
rect 35716 10047 35768 10056
rect 35716 10013 35725 10047
rect 35725 10013 35759 10047
rect 35759 10013 35768 10047
rect 35716 10004 35768 10013
rect 37924 10004 37976 10056
rect 38108 10047 38160 10056
rect 38108 10013 38117 10047
rect 38117 10013 38151 10047
rect 38151 10013 38160 10047
rect 38108 10004 38160 10013
rect 28172 9936 28224 9988
rect 32956 9936 33008 9988
rect 34704 9936 34756 9988
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 10232 9664 10284 9716
rect 10508 9707 10560 9716
rect 10508 9673 10517 9707
rect 10517 9673 10551 9707
rect 10551 9673 10560 9707
rect 10508 9664 10560 9673
rect 11704 9664 11756 9716
rect 12164 9707 12216 9716
rect 12164 9673 12173 9707
rect 12173 9673 12207 9707
rect 12207 9673 12216 9707
rect 12164 9664 12216 9673
rect 13912 9664 13964 9716
rect 10140 9639 10192 9648
rect 10140 9605 10149 9639
rect 10149 9605 10183 9639
rect 10183 9605 10192 9639
rect 10140 9596 10192 9605
rect 10692 9528 10744 9580
rect 14188 9596 14240 9648
rect 15844 9664 15896 9716
rect 16672 9707 16724 9716
rect 16672 9673 16681 9707
rect 16681 9673 16715 9707
rect 16715 9673 16724 9707
rect 16672 9664 16724 9673
rect 18512 9707 18564 9716
rect 18512 9673 18521 9707
rect 18521 9673 18555 9707
rect 18555 9673 18564 9707
rect 18512 9664 18564 9673
rect 19156 9707 19208 9716
rect 19156 9673 19165 9707
rect 19165 9673 19199 9707
rect 19199 9673 19208 9707
rect 19156 9664 19208 9673
rect 21272 9707 21324 9716
rect 21272 9673 21281 9707
rect 21281 9673 21315 9707
rect 21315 9673 21324 9707
rect 21272 9664 21324 9673
rect 22468 9707 22520 9716
rect 22468 9673 22477 9707
rect 22477 9673 22511 9707
rect 22511 9673 22520 9707
rect 22468 9664 22520 9673
rect 22928 9664 22980 9716
rect 24676 9664 24728 9716
rect 25412 9664 25464 9716
rect 27068 9664 27120 9716
rect 28172 9707 28224 9716
rect 28172 9673 28181 9707
rect 28181 9673 28215 9707
rect 28215 9673 28224 9707
rect 28172 9664 28224 9673
rect 28448 9707 28500 9716
rect 28448 9673 28457 9707
rect 28457 9673 28491 9707
rect 28491 9673 28500 9707
rect 28448 9664 28500 9673
rect 28908 9664 28960 9716
rect 29920 9664 29972 9716
rect 32036 9664 32088 9716
rect 36728 9707 36780 9716
rect 36728 9673 36737 9707
rect 36737 9673 36771 9707
rect 36771 9673 36780 9707
rect 36728 9664 36780 9673
rect 37740 9707 37792 9716
rect 37740 9673 37749 9707
rect 37749 9673 37783 9707
rect 37783 9673 37792 9707
rect 37740 9664 37792 9673
rect 37924 9664 37976 9716
rect 39948 9664 40000 9716
rect 41512 9664 41564 9716
rect 16580 9596 16632 9648
rect 23664 9596 23716 9648
rect 14280 9571 14332 9580
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 21548 9571 21600 9580
rect 21548 9537 21557 9571
rect 21557 9537 21591 9571
rect 21591 9537 21600 9571
rect 21548 9528 21600 9537
rect 21824 9571 21876 9580
rect 21824 9537 21833 9571
rect 21833 9537 21867 9571
rect 21867 9537 21876 9571
rect 21824 9528 21876 9537
rect 23388 9528 23440 9580
rect 24952 9596 25004 9648
rect 28816 9596 28868 9648
rect 27620 9571 27672 9580
rect 27620 9537 27629 9571
rect 27629 9537 27663 9571
rect 27663 9537 27672 9571
rect 27620 9528 27672 9537
rect 28724 9528 28776 9580
rect 29276 9571 29328 9580
rect 29276 9537 29285 9571
rect 29285 9537 29319 9571
rect 29319 9537 29328 9571
rect 29276 9528 29328 9537
rect 29552 9528 29604 9580
rect 14924 9503 14976 9512
rect 10508 9392 10560 9444
rect 11244 9392 11296 9444
rect 14924 9469 14933 9503
rect 14933 9469 14967 9503
rect 14967 9469 14976 9503
rect 14924 9460 14976 9469
rect 13544 9392 13596 9444
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 12440 9324 12492 9376
rect 13636 9324 13688 9376
rect 13820 9324 13872 9376
rect 18512 9460 18564 9512
rect 19892 9460 19944 9512
rect 23572 9460 23624 9512
rect 25320 9503 25372 9512
rect 25320 9469 25329 9503
rect 25329 9469 25363 9503
rect 25363 9469 25372 9503
rect 25320 9460 25372 9469
rect 18512 9324 18564 9376
rect 19984 9324 20036 9376
rect 27252 9460 27304 9512
rect 31024 9503 31076 9512
rect 31024 9469 31033 9503
rect 31033 9469 31067 9503
rect 31067 9469 31076 9503
rect 31024 9460 31076 9469
rect 34520 9596 34572 9648
rect 38568 9596 38620 9648
rect 33784 9571 33836 9580
rect 33784 9537 33793 9571
rect 33793 9537 33827 9571
rect 33827 9537 33836 9571
rect 33784 9528 33836 9537
rect 34704 9528 34756 9580
rect 33968 9460 34020 9512
rect 35808 9503 35860 9512
rect 35808 9469 35817 9503
rect 35817 9469 35851 9503
rect 35851 9469 35860 9503
rect 35808 9460 35860 9469
rect 39120 9460 39172 9512
rect 40500 9503 40552 9512
rect 40500 9469 40509 9503
rect 40509 9469 40543 9503
rect 40543 9469 40552 9503
rect 40500 9460 40552 9469
rect 20628 9367 20680 9376
rect 20628 9333 20637 9367
rect 20637 9333 20671 9367
rect 20671 9333 20680 9367
rect 20628 9324 20680 9333
rect 21272 9324 21324 9376
rect 27804 9392 27856 9444
rect 28908 9392 28960 9444
rect 33140 9392 33192 9444
rect 36084 9392 36136 9444
rect 39948 9392 40000 9444
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 10692 9163 10744 9172
rect 10692 9129 10701 9163
rect 10701 9129 10735 9163
rect 10735 9129 10744 9163
rect 10692 9120 10744 9129
rect 11244 9163 11296 9172
rect 11244 9129 11253 9163
rect 11253 9129 11287 9163
rect 11287 9129 11296 9163
rect 11244 9120 11296 9129
rect 12440 9163 12492 9172
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 12440 9120 12492 9129
rect 14188 9120 14240 9172
rect 21548 9120 21600 9172
rect 23204 9120 23256 9172
rect 23388 9120 23440 9172
rect 24860 9163 24912 9172
rect 24860 9129 24869 9163
rect 24869 9129 24903 9163
rect 24903 9129 24912 9163
rect 24860 9120 24912 9129
rect 25320 9120 25372 9172
rect 29276 9120 29328 9172
rect 33968 9120 34020 9172
rect 35716 9163 35768 9172
rect 35716 9129 35725 9163
rect 35725 9129 35759 9163
rect 35759 9129 35768 9163
rect 35716 9120 35768 9129
rect 37096 9120 37148 9172
rect 39120 9120 39172 9172
rect 40132 9163 40184 9172
rect 40132 9129 40141 9163
rect 40141 9129 40175 9163
rect 40175 9129 40184 9163
rect 40132 9120 40184 9129
rect 40500 9120 40552 9172
rect 11704 8984 11756 9036
rect 13452 9052 13504 9104
rect 13544 9052 13596 9104
rect 17592 9052 17644 9104
rect 19892 9052 19944 9104
rect 20628 9052 20680 9104
rect 21824 9052 21876 9104
rect 23020 9095 23072 9104
rect 14188 9027 14240 9036
rect 14188 8993 14197 9027
rect 14197 8993 14231 9027
rect 14231 8993 14240 9027
rect 14188 8984 14240 8993
rect 14280 8984 14332 9036
rect 18696 8984 18748 9036
rect 19432 9027 19484 9036
rect 19432 8993 19441 9027
rect 19441 8993 19475 9027
rect 19475 8993 19484 9027
rect 19432 8984 19484 8993
rect 23020 9061 23029 9095
rect 23029 9061 23063 9095
rect 23063 9061 23072 9095
rect 23020 9052 23072 9061
rect 26792 9052 26844 9104
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 17500 8916 17552 8968
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 21180 8916 21232 8968
rect 27252 8984 27304 9036
rect 28448 9052 28500 9104
rect 28724 9027 28776 9036
rect 28724 8993 28733 9027
rect 28733 8993 28767 9027
rect 28767 8993 28776 9027
rect 28724 8984 28776 8993
rect 29552 9052 29604 9104
rect 29736 8984 29788 9036
rect 33600 9027 33652 9036
rect 33600 8993 33609 9027
rect 33609 8993 33643 9027
rect 33643 8993 33652 9027
rect 33600 8984 33652 8993
rect 34704 9027 34756 9036
rect 34704 8993 34713 9027
rect 34713 8993 34747 9027
rect 34747 8993 34756 9027
rect 34704 8984 34756 8993
rect 35808 9052 35860 9104
rect 36544 9027 36596 9036
rect 36544 8993 36553 9027
rect 36553 8993 36587 9027
rect 36587 8993 36596 9027
rect 36544 8984 36596 8993
rect 39948 8984 40000 9036
rect 27160 8916 27212 8968
rect 28172 8916 28224 8968
rect 14372 8823 14424 8832
rect 14372 8789 14381 8823
rect 14381 8789 14415 8823
rect 14415 8789 14424 8823
rect 14372 8780 14424 8789
rect 16488 8780 16540 8832
rect 30012 8780 30064 8832
rect 31024 8823 31076 8832
rect 31024 8789 31033 8823
rect 31033 8789 31067 8823
rect 31067 8789 31076 8823
rect 31024 8780 31076 8789
rect 33416 8780 33468 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 11244 8576 11296 8628
rect 11520 8576 11572 8628
rect 13452 8619 13504 8628
rect 11796 8508 11848 8560
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 17592 8576 17644 8628
rect 18696 8576 18748 8628
rect 19432 8619 19484 8628
rect 19432 8585 19441 8619
rect 19441 8585 19475 8619
rect 19475 8585 19484 8619
rect 19432 8576 19484 8585
rect 20444 8576 20496 8628
rect 20628 8619 20680 8628
rect 20628 8585 20637 8619
rect 20637 8585 20671 8619
rect 20671 8585 20680 8619
rect 20628 8576 20680 8585
rect 20996 8619 21048 8628
rect 20996 8585 21005 8619
rect 21005 8585 21039 8619
rect 21039 8585 21048 8619
rect 20996 8576 21048 8585
rect 27160 8619 27212 8628
rect 27160 8585 27169 8619
rect 27169 8585 27203 8619
rect 27203 8585 27212 8619
rect 27160 8576 27212 8585
rect 28448 8619 28500 8628
rect 28448 8585 28457 8619
rect 28457 8585 28491 8619
rect 28491 8585 28500 8619
rect 28448 8576 28500 8585
rect 28724 8619 28776 8628
rect 28724 8585 28733 8619
rect 28733 8585 28767 8619
rect 28767 8585 28776 8619
rect 28724 8576 28776 8585
rect 33600 8619 33652 8628
rect 33600 8585 33609 8619
rect 33609 8585 33643 8619
rect 33643 8585 33652 8619
rect 33600 8576 33652 8585
rect 33968 8576 34020 8628
rect 36544 8619 36596 8628
rect 12440 8508 12492 8560
rect 13084 8551 13136 8560
rect 13084 8517 13093 8551
rect 13093 8517 13127 8551
rect 13127 8517 13136 8551
rect 13084 8508 13136 8517
rect 16580 8508 16632 8560
rect 13636 8440 13688 8492
rect 21824 8508 21876 8560
rect 30012 8483 30064 8492
rect 30012 8449 30021 8483
rect 30021 8449 30055 8483
rect 30055 8449 30064 8483
rect 30012 8440 30064 8449
rect 34244 8440 34296 8492
rect 36544 8585 36553 8619
rect 36553 8585 36587 8619
rect 36587 8585 36596 8619
rect 36544 8576 36596 8585
rect 14372 8415 14424 8424
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 17776 8372 17828 8424
rect 17868 8372 17920 8424
rect 20352 8372 20404 8424
rect 14096 8304 14148 8356
rect 17500 8304 17552 8356
rect 21364 8347 21416 8356
rect 21364 8313 21373 8347
rect 21373 8313 21407 8347
rect 21407 8313 21416 8347
rect 21364 8304 21416 8313
rect 26424 8372 26476 8424
rect 27252 8372 27304 8424
rect 29736 8415 29788 8424
rect 29368 8304 29420 8356
rect 29736 8381 29745 8415
rect 29745 8381 29779 8415
rect 29779 8381 29788 8415
rect 29736 8372 29788 8381
rect 34520 8372 34572 8424
rect 35072 8372 35124 8424
rect 35716 8440 35768 8492
rect 33232 8304 33284 8356
rect 15108 8279 15160 8288
rect 15108 8245 15117 8279
rect 15117 8245 15151 8279
rect 15151 8245 15160 8279
rect 15108 8236 15160 8245
rect 21180 8236 21232 8288
rect 26148 8279 26200 8288
rect 26148 8245 26157 8279
rect 26157 8245 26191 8279
rect 26191 8245 26200 8279
rect 26148 8236 26200 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 12716 8075 12768 8084
rect 12716 8041 12725 8075
rect 12725 8041 12759 8075
rect 12759 8041 12768 8075
rect 12716 8032 12768 8041
rect 14924 8032 14976 8084
rect 15752 8075 15804 8084
rect 15752 8041 15761 8075
rect 15761 8041 15795 8075
rect 15795 8041 15804 8075
rect 15752 8032 15804 8041
rect 15844 8032 15896 8084
rect 16488 8075 16540 8084
rect 16488 8041 16497 8075
rect 16497 8041 16531 8075
rect 16531 8041 16540 8075
rect 16488 8032 16540 8041
rect 17224 8075 17276 8084
rect 17224 8041 17233 8075
rect 17233 8041 17267 8075
rect 17267 8041 17276 8075
rect 17224 8032 17276 8041
rect 17500 8075 17552 8084
rect 17500 8041 17509 8075
rect 17509 8041 17543 8075
rect 17543 8041 17552 8075
rect 17500 8032 17552 8041
rect 21180 8075 21232 8084
rect 14188 7964 14240 8016
rect 15108 7964 15160 8016
rect 13084 7939 13136 7948
rect 13084 7905 13093 7939
rect 13093 7905 13127 7939
rect 13127 7905 13136 7939
rect 13084 7896 13136 7905
rect 15936 7964 15988 8016
rect 16580 7896 16632 7948
rect 18788 7964 18840 8016
rect 21180 8041 21189 8075
rect 21189 8041 21223 8075
rect 21223 8041 21232 8075
rect 21180 8032 21232 8041
rect 21364 8075 21416 8084
rect 21364 8041 21373 8075
rect 21373 8041 21407 8075
rect 21407 8041 21416 8075
rect 21364 8032 21416 8041
rect 26424 8032 26476 8084
rect 29368 8075 29420 8084
rect 29368 8041 29377 8075
rect 29377 8041 29411 8075
rect 29411 8041 29420 8075
rect 29368 8032 29420 8041
rect 29736 8075 29788 8084
rect 29736 8041 29745 8075
rect 29745 8041 29779 8075
rect 29779 8041 29788 8075
rect 29736 8032 29788 8041
rect 34704 8075 34756 8084
rect 34704 8041 34713 8075
rect 34713 8041 34747 8075
rect 34747 8041 34756 8075
rect 34704 8032 34756 8041
rect 35072 8075 35124 8084
rect 35072 8041 35081 8075
rect 35081 8041 35115 8075
rect 35115 8041 35124 8075
rect 35072 8032 35124 8041
rect 17132 7896 17184 7948
rect 17960 7896 18012 7948
rect 19616 7896 19668 7948
rect 20904 7939 20956 7948
rect 20904 7905 20948 7939
rect 20948 7905 20956 7939
rect 20904 7896 20956 7905
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 18512 7828 18564 7880
rect 13176 7692 13228 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 13084 7488 13136 7540
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 16580 7488 16632 7540
rect 20352 7531 20404 7540
rect 20352 7497 20361 7531
rect 20361 7497 20395 7531
rect 20395 7497 20404 7531
rect 20352 7488 20404 7497
rect 20904 7531 20956 7540
rect 20904 7497 20913 7531
rect 20913 7497 20947 7531
rect 20947 7497 20956 7531
rect 20904 7488 20956 7497
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 18880 7352 18932 7404
rect 13544 7327 13596 7336
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 8576 7216 8628 7268
rect 14648 7216 14700 7268
rect 17776 7284 17828 7336
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 17408 7216 17460 7268
rect 15568 7148 15620 7200
rect 17040 7148 17092 7200
rect 17684 7191 17736 7200
rect 17684 7157 17693 7191
rect 17693 7157 17727 7191
rect 17727 7157 17736 7191
rect 17684 7148 17736 7157
rect 18052 7148 18104 7200
rect 18788 7216 18840 7268
rect 19616 7216 19668 7268
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 13176 6944 13228 6996
rect 15108 6944 15160 6996
rect 17868 6987 17920 6996
rect 17868 6953 17877 6987
rect 17877 6953 17911 6987
rect 17911 6953 17920 6987
rect 17868 6944 17920 6953
rect 18512 6987 18564 6996
rect 18512 6953 18521 6987
rect 18521 6953 18555 6987
rect 18555 6953 18564 6987
rect 18512 6944 18564 6953
rect 18880 6987 18932 6996
rect 18880 6953 18889 6987
rect 18889 6953 18923 6987
rect 18923 6953 18932 6987
rect 18880 6944 18932 6953
rect 17040 6876 17092 6928
rect 18788 6876 18840 6928
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 15016 6808 15068 6860
rect 15936 6851 15988 6860
rect 15936 6817 15945 6851
rect 15945 6817 15979 6851
rect 15979 6817 15988 6851
rect 15936 6808 15988 6817
rect 17408 6851 17460 6860
rect 17408 6817 17417 6851
rect 17417 6817 17451 6851
rect 17451 6817 17460 6851
rect 17408 6808 17460 6817
rect 15200 6740 15252 6792
rect 14648 6672 14700 6724
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 15200 6443 15252 6452
rect 15200 6409 15209 6443
rect 15209 6409 15243 6443
rect 15243 6409 15252 6443
rect 15200 6400 15252 6409
rect 15568 6443 15620 6452
rect 15568 6409 15577 6443
rect 15577 6409 15611 6443
rect 15611 6409 15620 6443
rect 15568 6400 15620 6409
rect 15936 6400 15988 6452
rect 17132 6443 17184 6452
rect 17132 6409 17141 6443
rect 17141 6409 17175 6443
rect 17175 6409 17184 6443
rect 17132 6400 17184 6409
rect 18052 6400 18104 6452
rect 13728 6332 13780 6384
rect 17776 6332 17828 6384
rect 14648 6264 14700 6316
rect 17040 6264 17092 6316
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 28540 76 28592 128
rect 30472 76 30524 128
<< metal2 >>
rect 2778 49586 2834 50000
rect 2778 49558 2912 49586
rect 2778 49520 2834 49558
rect 110 46472 166 46481
rect 110 46407 166 46416
rect 124 39817 152 46407
rect 2884 42794 2912 49558
rect 8298 49520 8354 50000
rect 13818 49586 13874 50000
rect 19430 49586 19486 50000
rect 13818 49558 14044 49586
rect 13818 49520 13874 49558
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 2792 42766 2912 42794
rect 110 39808 166 39817
rect 110 39743 166 39752
rect 2792 39409 2820 42766
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 12808 39840 12860 39846
rect 12808 39782 12860 39788
rect 12992 39840 13044 39846
rect 12992 39782 13044 39788
rect 11980 39500 12032 39506
rect 11980 39442 12032 39448
rect 10968 39432 11020 39438
rect 2778 39400 2834 39409
rect 10968 39374 11020 39380
rect 2778 39335 2834 39344
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 8300 38956 8352 38962
rect 8300 38898 8352 38904
rect 2594 38720 2650 38729
rect 2594 38655 2650 38664
rect 2228 25356 2280 25362
rect 2228 25298 2280 25304
rect 2136 25152 2188 25158
rect 2136 25094 2188 25100
rect 110 24984 166 24993
rect 110 24919 166 24928
rect 124 24886 152 24919
rect 112 24880 164 24886
rect 112 24822 164 24828
rect 2148 24274 2176 25094
rect 2240 24818 2268 25298
rect 2228 24812 2280 24818
rect 2228 24754 2280 24760
rect 2240 24410 2268 24754
rect 2412 24676 2464 24682
rect 2412 24618 2464 24624
rect 2228 24404 2280 24410
rect 2228 24346 2280 24352
rect 1492 24268 1544 24274
rect 1492 24210 1544 24216
rect 2136 24268 2188 24274
rect 2136 24210 2188 24216
rect 1504 23526 1532 24210
rect 2424 23866 2452 24618
rect 2504 24132 2556 24138
rect 2504 24074 2556 24080
rect 2412 23860 2464 23866
rect 2412 23802 2464 23808
rect 1492 23520 1544 23526
rect 1492 23462 1544 23468
rect 2320 23520 2372 23526
rect 2372 23480 2452 23508
rect 2320 23462 2372 23468
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1412 4185 1440 21286
rect 1504 11257 1532 23462
rect 2424 23186 2452 23480
rect 2516 23322 2544 24074
rect 2504 23316 2556 23322
rect 2504 23258 2556 23264
rect 2320 23180 2372 23186
rect 2320 23122 2372 23128
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 2332 22574 2360 23122
rect 2320 22568 2372 22574
rect 2320 22510 2372 22516
rect 1952 22432 2004 22438
rect 1952 22374 2004 22380
rect 1964 18465 1992 22374
rect 2136 22092 2188 22098
rect 2136 22034 2188 22040
rect 2148 21486 2176 22034
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 2608 18873 2636 38655
rect 7196 38276 7248 38282
rect 7196 38218 7248 38224
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 7104 37392 7156 37398
rect 7104 37334 7156 37340
rect 6920 37256 6972 37262
rect 6920 37198 6972 37204
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 6932 36922 6960 37198
rect 6920 36916 6972 36922
rect 6920 36858 6972 36864
rect 7116 36582 7144 37334
rect 7208 37262 7236 38218
rect 7656 38208 7708 38214
rect 7656 38150 7708 38156
rect 7668 37738 7696 38150
rect 8312 37874 8340 38898
rect 10980 38826 11008 39374
rect 11152 38956 11204 38962
rect 11152 38898 11204 38904
rect 10876 38820 10928 38826
rect 10876 38762 10928 38768
rect 10968 38820 11020 38826
rect 10968 38762 11020 38768
rect 10232 38480 10284 38486
rect 10232 38422 10284 38428
rect 10048 38344 10100 38350
rect 10048 38286 10100 38292
rect 10060 37874 10088 38286
rect 10244 37942 10272 38422
rect 10888 38350 10916 38762
rect 10876 38344 10928 38350
rect 10876 38286 10928 38292
rect 11164 38282 11192 38898
rect 11992 38894 12020 39442
rect 12820 38894 12848 39782
rect 13004 39545 13032 39782
rect 12990 39536 13046 39545
rect 12990 39471 13046 39480
rect 12992 39432 13044 39438
rect 12992 39374 13044 39380
rect 11980 38888 12032 38894
rect 11980 38830 12032 38836
rect 12808 38888 12860 38894
rect 12808 38830 12860 38836
rect 11888 38752 11940 38758
rect 11888 38694 11940 38700
rect 11900 38418 11928 38694
rect 11888 38412 11940 38418
rect 11888 38354 11940 38360
rect 11244 38344 11296 38350
rect 11244 38286 11296 38292
rect 11152 38276 11204 38282
rect 11152 38218 11204 38224
rect 10232 37936 10284 37942
rect 10232 37878 10284 37884
rect 8300 37868 8352 37874
rect 8300 37810 8352 37816
rect 9496 37868 9548 37874
rect 9496 37810 9548 37816
rect 10048 37868 10100 37874
rect 10048 37810 10100 37816
rect 9508 37738 9536 37810
rect 7656 37732 7708 37738
rect 7656 37674 7708 37680
rect 9036 37732 9088 37738
rect 9036 37674 9088 37680
rect 9220 37732 9272 37738
rect 9220 37674 9272 37680
rect 9496 37732 9548 37738
rect 9496 37674 9548 37680
rect 7196 37256 7248 37262
rect 7196 37198 7248 37204
rect 5540 36576 5592 36582
rect 5540 36518 5592 36524
rect 6184 36576 6236 36582
rect 6184 36518 6236 36524
rect 7104 36576 7156 36582
rect 7104 36518 7156 36524
rect 5264 36236 5316 36242
rect 5264 36178 5316 36184
rect 4620 36032 4672 36038
rect 4620 35974 4672 35980
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4632 35630 4660 35974
rect 4620 35624 4672 35630
rect 4620 35566 4672 35572
rect 4160 35488 4212 35494
rect 4160 35430 4212 35436
rect 4172 35154 4200 35430
rect 4160 35148 4212 35154
rect 4160 35090 4212 35096
rect 4068 35080 4120 35086
rect 4068 35022 4120 35028
rect 3332 34536 3384 34542
rect 3332 34478 3384 34484
rect 3344 33658 3372 34478
rect 4080 33862 4108 35022
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4068 33856 4120 33862
rect 4068 33798 4120 33804
rect 3332 33652 3384 33658
rect 3332 33594 3384 33600
rect 3700 33448 3752 33454
rect 3700 33390 3752 33396
rect 3976 33448 4028 33454
rect 3976 33390 4028 33396
rect 3516 32972 3568 32978
rect 3516 32914 3568 32920
rect 3240 32768 3292 32774
rect 3240 32710 3292 32716
rect 3252 32570 3280 32710
rect 3240 32564 3292 32570
rect 3240 32506 3292 32512
rect 3240 32360 3292 32366
rect 3240 32302 3292 32308
rect 3056 30320 3108 30326
rect 3056 30262 3108 30268
rect 2964 30048 3016 30054
rect 2964 29990 3016 29996
rect 2976 29102 3004 29990
rect 2964 29096 3016 29102
rect 2964 29038 3016 29044
rect 2976 28014 3004 29038
rect 2964 28008 3016 28014
rect 2964 27950 3016 27956
rect 3068 25702 3096 30262
rect 3148 30116 3200 30122
rect 3148 30058 3200 30064
rect 3160 29510 3188 30058
rect 3148 29504 3200 29510
rect 3148 29446 3200 29452
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 2964 25356 3016 25362
rect 2964 25298 3016 25304
rect 2976 24410 3004 25298
rect 2964 24404 3016 24410
rect 2964 24346 3016 24352
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2976 23662 3004 24210
rect 2964 23656 3016 23662
rect 2884 23616 2964 23644
rect 2884 23322 2912 23616
rect 2964 23598 3016 23604
rect 3068 23474 3096 25638
rect 3160 25140 3188 29446
rect 3252 29102 3280 32302
rect 3528 32230 3556 32914
rect 3516 32224 3568 32230
rect 3516 32166 3568 32172
rect 3330 31648 3386 31657
rect 3330 31583 3386 31592
rect 3240 29096 3292 29102
rect 3240 29038 3292 29044
rect 3252 28422 3280 29038
rect 3240 28416 3292 28422
rect 3240 28358 3292 28364
rect 3240 25152 3292 25158
rect 3160 25112 3240 25140
rect 3240 25094 3292 25100
rect 3148 23792 3200 23798
rect 3148 23734 3200 23740
rect 2976 23446 3096 23474
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2884 22642 2912 22918
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2688 21888 2740 21894
rect 2688 21830 2740 21836
rect 2594 18864 2650 18873
rect 2594 18799 2650 18808
rect 1950 18456 2006 18465
rect 1950 18391 2006 18400
rect 2700 16658 2728 21830
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2792 20058 2820 20334
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2792 19292 2820 19994
rect 2976 19378 3004 23446
rect 3160 22982 3188 23734
rect 3148 22976 3200 22982
rect 3148 22918 3200 22924
rect 3252 20534 3280 25094
rect 3344 23746 3372 31583
rect 3528 30122 3556 32166
rect 3712 30326 3740 33390
rect 3988 33046 4016 33390
rect 4080 33114 4108 33798
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4068 33108 4120 33114
rect 4068 33050 4120 33056
rect 3976 33040 4028 33046
rect 3976 32982 4028 32988
rect 3988 32774 4016 32982
rect 3976 32768 4028 32774
rect 3976 32710 4028 32716
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4632 32434 4660 35566
rect 4712 35488 4764 35494
rect 4712 35430 4764 35436
rect 4724 35290 4752 35430
rect 5276 35290 5304 36178
rect 5552 35834 5580 36518
rect 6092 36304 6144 36310
rect 6092 36246 6144 36252
rect 6000 36168 6052 36174
rect 6000 36110 6052 36116
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 6012 35290 6040 36110
rect 6104 35834 6132 36246
rect 6092 35828 6144 35834
rect 6092 35770 6144 35776
rect 6196 35766 6224 36518
rect 7116 36038 7144 36518
rect 7208 36310 7236 37198
rect 7668 37194 7696 37674
rect 8944 37256 8996 37262
rect 8944 37198 8996 37204
rect 7656 37188 7708 37194
rect 7656 37130 7708 37136
rect 8956 36922 8984 37198
rect 8944 36916 8996 36922
rect 8944 36858 8996 36864
rect 8208 36780 8260 36786
rect 8208 36722 8260 36728
rect 8220 36310 8248 36722
rect 7196 36304 7248 36310
rect 7196 36246 7248 36252
rect 7840 36304 7892 36310
rect 7840 36246 7892 36252
rect 8208 36304 8260 36310
rect 8208 36246 8260 36252
rect 7104 36032 7156 36038
rect 7104 35974 7156 35980
rect 6184 35760 6236 35766
rect 6184 35702 6236 35708
rect 7116 35562 7144 35974
rect 7196 35692 7248 35698
rect 7196 35634 7248 35640
rect 7104 35556 7156 35562
rect 7104 35498 7156 35504
rect 4712 35284 4764 35290
rect 4712 35226 4764 35232
rect 5264 35284 5316 35290
rect 5264 35226 5316 35232
rect 6000 35284 6052 35290
rect 6000 35226 6052 35232
rect 4724 34406 4752 35226
rect 6092 35216 6144 35222
rect 6092 35158 6144 35164
rect 4896 34536 4948 34542
rect 4896 34478 4948 34484
rect 4712 34400 4764 34406
rect 4712 34342 4764 34348
rect 4712 34060 4764 34066
rect 4712 34002 4764 34008
rect 4724 33318 4752 34002
rect 4712 33312 4764 33318
rect 4712 33254 4764 33260
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 4528 32360 4580 32366
rect 4528 32302 4580 32308
rect 4540 31890 4568 32302
rect 3792 31884 3844 31890
rect 3792 31826 3844 31832
rect 4528 31884 4580 31890
rect 4580 31844 4660 31872
rect 4528 31826 4580 31832
rect 3804 31142 3832 31826
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4632 31482 4660 31844
rect 4620 31476 4672 31482
rect 4620 31418 4672 31424
rect 3792 31136 3844 31142
rect 3792 31078 3844 31084
rect 3700 30320 3752 30326
rect 3700 30262 3752 30268
rect 3516 30116 3568 30122
rect 3516 30058 3568 30064
rect 3804 28404 3832 31078
rect 4620 30932 4672 30938
rect 4620 30874 4672 30880
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 3884 30116 3936 30122
rect 3884 30058 3936 30064
rect 3896 29646 3924 30058
rect 4632 30054 4660 30874
rect 4620 30048 4672 30054
rect 4620 29990 4672 29996
rect 4632 29782 4660 29990
rect 4620 29776 4672 29782
rect 4620 29718 4672 29724
rect 3884 29640 3936 29646
rect 3884 29582 3936 29588
rect 3896 28558 3924 29582
rect 4068 29504 4120 29510
rect 4068 29446 4120 29452
rect 3976 28960 4028 28966
rect 3974 28928 3976 28937
rect 4028 28928 4030 28937
rect 3974 28863 4030 28872
rect 3884 28552 3936 28558
rect 3884 28494 3936 28500
rect 3804 28376 3924 28404
rect 3896 28014 3924 28376
rect 3792 28008 3844 28014
rect 3792 27950 3844 27956
rect 3884 28008 3936 28014
rect 3884 27950 3936 27956
rect 3804 26450 3832 27950
rect 3896 27316 3924 27950
rect 3988 27606 4016 28863
rect 4080 28694 4108 29446
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4528 29028 4580 29034
rect 4632 29016 4660 29718
rect 4580 28988 4660 29016
rect 4528 28970 4580 28976
rect 4540 28937 4568 28970
rect 4526 28928 4582 28937
rect 4526 28863 4582 28872
rect 4068 28688 4120 28694
rect 4068 28630 4120 28636
rect 4620 28620 4672 28626
rect 4620 28562 4672 28568
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4068 28076 4120 28082
rect 4068 28018 4120 28024
rect 3976 27600 4028 27606
rect 3976 27542 4028 27548
rect 4080 27538 4108 28018
rect 4632 27878 4660 28562
rect 4620 27872 4672 27878
rect 4620 27814 4672 27820
rect 4632 27674 4660 27814
rect 4620 27668 4672 27674
rect 4620 27610 4672 27616
rect 4068 27532 4120 27538
rect 4068 27474 4120 27480
rect 3976 27328 4028 27334
rect 3896 27288 3976 27316
rect 3976 27270 4028 27276
rect 3792 26444 3844 26450
rect 3792 26386 3844 26392
rect 3988 25974 4016 27270
rect 4080 26586 4108 27474
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4724 27146 4752 33254
rect 4908 31958 4936 34478
rect 6104 34406 6132 35158
rect 6460 35080 6512 35086
rect 6460 35022 6512 35028
rect 6472 34406 6500 35022
rect 7208 34950 7236 35634
rect 7852 35494 7880 36246
rect 8208 36168 8260 36174
rect 8208 36110 8260 36116
rect 8220 35494 8248 36110
rect 8956 35698 8984 36858
rect 9048 36310 9076 37674
rect 9232 37466 9260 37674
rect 9220 37460 9272 37466
rect 9220 37402 9272 37408
rect 9232 36786 9260 37402
rect 10244 37398 10272 37878
rect 11256 37738 11284 38286
rect 11900 38010 11928 38354
rect 11992 38010 12020 38830
rect 12820 38010 12848 38830
rect 11888 38004 11940 38010
rect 11888 37946 11940 37952
rect 11980 38004 12032 38010
rect 11980 37946 12032 37952
rect 12808 38004 12860 38010
rect 12808 37946 12860 37952
rect 12820 37806 12848 37946
rect 12808 37800 12860 37806
rect 12808 37742 12860 37748
rect 10876 37732 10928 37738
rect 10876 37674 10928 37680
rect 11244 37732 11296 37738
rect 11244 37674 11296 37680
rect 10888 37466 10916 37674
rect 10876 37460 10928 37466
rect 10876 37402 10928 37408
rect 10232 37392 10284 37398
rect 10232 37334 10284 37340
rect 10244 36922 10272 37334
rect 10232 36916 10284 36922
rect 10232 36858 10284 36864
rect 9220 36780 9272 36786
rect 9220 36722 9272 36728
rect 10244 36650 10272 36858
rect 10888 36786 10916 37402
rect 13004 37398 13032 39374
rect 13636 39296 13688 39302
rect 13636 39238 13688 39244
rect 13176 38344 13228 38350
rect 13176 38286 13228 38292
rect 13188 37738 13216 38286
rect 13648 37806 13676 39238
rect 13728 38820 13780 38826
rect 13728 38762 13780 38768
rect 13740 38554 13768 38762
rect 13728 38548 13780 38554
rect 13728 38490 13780 38496
rect 13820 38480 13872 38486
rect 13820 38422 13872 38428
rect 13832 38010 13860 38422
rect 13820 38004 13872 38010
rect 13820 37946 13872 37952
rect 14016 37942 14044 49558
rect 19352 49558 19486 49586
rect 19352 42362 19380 49558
rect 19430 49520 19486 49558
rect 24950 49586 25006 50000
rect 30470 49586 30526 50000
rect 36082 49586 36138 50000
rect 41602 49586 41658 50000
rect 47122 49586 47178 50000
rect 24950 49558 25084 49586
rect 24950 49520 25006 49558
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 23110 43888 23166 43897
rect 25056 43858 25084 49558
rect 30300 49558 30526 49586
rect 30300 43897 30328 49558
rect 30470 49520 30526 49558
rect 35912 49558 36138 49586
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 30748 44328 30800 44334
rect 30748 44270 30800 44276
rect 31852 44328 31904 44334
rect 31852 44270 31904 44276
rect 30286 43888 30342 43897
rect 23110 43823 23112 43832
rect 23164 43823 23166 43832
rect 25044 43852 25096 43858
rect 23112 43794 23164 43800
rect 30286 43823 30342 43832
rect 25044 43794 25096 43800
rect 23124 43450 23152 43794
rect 23572 43648 23624 43654
rect 23572 43590 23624 43596
rect 23848 43648 23900 43654
rect 23848 43590 23900 43596
rect 24032 43648 24084 43654
rect 24032 43590 24084 43596
rect 22376 43444 22428 43450
rect 22376 43386 22428 43392
rect 23112 43444 23164 43450
rect 23112 43386 23164 43392
rect 21640 43104 21692 43110
rect 21640 43046 21692 43052
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 18512 42356 18564 42362
rect 18512 42298 18564 42304
rect 19340 42356 19392 42362
rect 19340 42298 19392 42304
rect 17314 39808 17370 39817
rect 17314 39743 17370 39752
rect 14832 39500 14884 39506
rect 14832 39442 14884 39448
rect 16120 39500 16172 39506
rect 16120 39442 16172 39448
rect 14844 38894 14872 39442
rect 15016 39296 15068 39302
rect 15016 39238 15068 39244
rect 14832 38888 14884 38894
rect 14832 38830 14884 38836
rect 14004 37936 14056 37942
rect 14004 37878 14056 37884
rect 13912 37868 13964 37874
rect 13912 37810 13964 37816
rect 13636 37800 13688 37806
rect 13636 37742 13688 37748
rect 13176 37732 13228 37738
rect 13176 37674 13228 37680
rect 11428 37392 11480 37398
rect 11428 37334 11480 37340
rect 12992 37392 13044 37398
rect 12992 37334 13044 37340
rect 11336 37256 11388 37262
rect 11336 37198 11388 37204
rect 11348 36922 11376 37198
rect 11336 36916 11388 36922
rect 11336 36858 11388 36864
rect 10876 36780 10928 36786
rect 10876 36722 10928 36728
rect 9864 36644 9916 36650
rect 9864 36586 9916 36592
rect 10232 36644 10284 36650
rect 10232 36586 10284 36592
rect 9036 36304 9088 36310
rect 9036 36246 9088 36252
rect 9876 36038 9904 36586
rect 10888 36310 10916 36722
rect 11440 36582 11468 37334
rect 12900 37256 12952 37262
rect 12900 37198 12952 37204
rect 11980 36916 12032 36922
rect 11980 36858 12032 36864
rect 11428 36576 11480 36582
rect 11428 36518 11480 36524
rect 11440 36378 11468 36518
rect 11428 36372 11480 36378
rect 11428 36314 11480 36320
rect 10140 36304 10192 36310
rect 10140 36246 10192 36252
rect 10876 36304 10928 36310
rect 10876 36246 10928 36252
rect 11796 36304 11848 36310
rect 11796 36246 11848 36252
rect 9864 36032 9916 36038
rect 9864 35974 9916 35980
rect 8944 35692 8996 35698
rect 8944 35634 8996 35640
rect 7840 35488 7892 35494
rect 7840 35430 7892 35436
rect 8208 35488 8260 35494
rect 8208 35430 8260 35436
rect 7852 35204 7880 35430
rect 7932 35216 7984 35222
rect 7852 35176 7932 35204
rect 7196 34944 7248 34950
rect 7196 34886 7248 34892
rect 5356 34400 5408 34406
rect 5356 34342 5408 34348
rect 6092 34400 6144 34406
rect 6092 34342 6144 34348
rect 6460 34400 6512 34406
rect 6460 34342 6512 34348
rect 5368 34066 5396 34342
rect 5172 34060 5224 34066
rect 5172 34002 5224 34008
rect 5356 34060 5408 34066
rect 5356 34002 5408 34008
rect 4988 33992 5040 33998
rect 4988 33934 5040 33940
rect 5000 33522 5028 33934
rect 4988 33516 5040 33522
rect 4988 33458 5040 33464
rect 5000 33114 5028 33458
rect 4988 33108 5040 33114
rect 4988 33050 5040 33056
rect 5184 32978 5212 34002
rect 6104 33386 6132 34342
rect 6184 34060 6236 34066
rect 6184 34002 6236 34008
rect 6196 33658 6224 34002
rect 6184 33652 6236 33658
rect 6184 33594 6236 33600
rect 6472 33454 6500 34342
rect 7208 34202 7236 34886
rect 7288 34536 7340 34542
rect 7288 34478 7340 34484
rect 7196 34196 7248 34202
rect 7196 34138 7248 34144
rect 7300 33862 7328 34478
rect 7852 34406 7880 35176
rect 7932 35158 7984 35164
rect 7932 35080 7984 35086
rect 7932 35022 7984 35028
rect 7944 34610 7972 35022
rect 8220 34746 8248 35430
rect 8956 35222 8984 35634
rect 9312 35556 9364 35562
rect 9312 35498 9364 35504
rect 9324 35222 9352 35498
rect 8944 35216 8996 35222
rect 8944 35158 8996 35164
rect 9312 35216 9364 35222
rect 9312 35158 9364 35164
rect 8576 35080 8628 35086
rect 8576 35022 8628 35028
rect 8208 34740 8260 34746
rect 8208 34682 8260 34688
rect 7932 34604 7984 34610
rect 7932 34546 7984 34552
rect 7840 34400 7892 34406
rect 7840 34342 7892 34348
rect 8300 34400 8352 34406
rect 8300 34342 8352 34348
rect 8312 34134 8340 34342
rect 8588 34202 8616 35022
rect 8852 34944 8904 34950
rect 8852 34886 8904 34892
rect 8760 34604 8812 34610
rect 8864 34592 8892 34886
rect 9324 34746 9352 35158
rect 9312 34740 9364 34746
rect 9312 34682 9364 34688
rect 8812 34564 8892 34592
rect 8760 34546 8812 34552
rect 8864 34202 8892 34564
rect 8576 34196 8628 34202
rect 8576 34138 8628 34144
rect 8852 34196 8904 34202
rect 8852 34138 8904 34144
rect 9324 34134 9352 34682
rect 9496 34604 9548 34610
rect 9496 34546 9548 34552
rect 8300 34128 8352 34134
rect 8300 34070 8352 34076
rect 9312 34128 9364 34134
rect 9312 34070 9364 34076
rect 8024 34060 8076 34066
rect 8024 34002 8076 34008
rect 8484 34060 8536 34066
rect 8484 34002 8536 34008
rect 7288 33856 7340 33862
rect 7288 33798 7340 33804
rect 7300 33658 7328 33798
rect 8036 33658 8064 34002
rect 7288 33652 7340 33658
rect 7288 33594 7340 33600
rect 8024 33652 8076 33658
rect 8024 33594 8076 33600
rect 8392 33652 8444 33658
rect 8392 33594 8444 33600
rect 6460 33448 6512 33454
rect 6460 33390 6512 33396
rect 6828 33448 6880 33454
rect 6828 33390 6880 33396
rect 6092 33380 6144 33386
rect 6092 33322 6144 33328
rect 6840 32978 6868 33390
rect 7840 33380 7892 33386
rect 7840 33322 7892 33328
rect 7852 33114 7880 33322
rect 7840 33108 7892 33114
rect 7840 33050 7892 33056
rect 5172 32972 5224 32978
rect 5172 32914 5224 32920
rect 6368 32972 6420 32978
rect 6368 32914 6420 32920
rect 6828 32972 6880 32978
rect 6828 32914 6880 32920
rect 5184 32774 5212 32914
rect 6276 32904 6328 32910
rect 6276 32846 6328 32852
rect 5172 32768 5224 32774
rect 5172 32710 5224 32716
rect 5184 32570 5212 32710
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 5184 32366 5212 32506
rect 5172 32360 5224 32366
rect 5172 32302 5224 32308
rect 6184 32360 6236 32366
rect 6184 32302 6236 32308
rect 6092 32224 6144 32230
rect 6092 32166 6144 32172
rect 4896 31952 4948 31958
rect 4896 31894 4948 31900
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 5172 31680 5224 31686
rect 5172 31622 5224 31628
rect 5184 31278 5212 31622
rect 5172 31272 5224 31278
rect 5172 31214 5224 31220
rect 4988 31136 5040 31142
rect 4988 31078 5040 31084
rect 4896 30728 4948 30734
rect 4896 30670 4948 30676
rect 4908 30054 4936 30670
rect 5000 30161 5028 31078
rect 5080 30184 5132 30190
rect 4986 30152 5042 30161
rect 5080 30126 5132 30132
rect 4986 30087 5042 30096
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4908 29850 4936 29990
rect 4896 29844 4948 29850
rect 4896 29786 4948 29792
rect 5092 29714 5120 30126
rect 5080 29708 5132 29714
rect 5080 29650 5132 29656
rect 5184 29306 5212 31214
rect 5356 31136 5408 31142
rect 5356 31078 5408 31084
rect 5264 30184 5316 30190
rect 5264 30126 5316 30132
rect 5276 29850 5304 30126
rect 5264 29844 5316 29850
rect 5264 29786 5316 29792
rect 5368 29617 5396 31078
rect 5828 30938 5856 31826
rect 5816 30932 5868 30938
rect 5816 30874 5868 30880
rect 5908 30864 5960 30870
rect 5908 30806 5960 30812
rect 5920 30122 5948 30806
rect 6104 30802 6132 32166
rect 6196 31686 6224 32302
rect 6288 32230 6316 32846
rect 6380 32570 6408 32914
rect 7472 32904 7524 32910
rect 7472 32846 7524 32852
rect 6368 32564 6420 32570
rect 6368 32506 6420 32512
rect 7380 32360 7432 32366
rect 7380 32302 7432 32308
rect 6276 32224 6328 32230
rect 6276 32166 6328 32172
rect 6184 31680 6236 31686
rect 6184 31622 6236 31628
rect 6196 30938 6224 31622
rect 6184 30932 6236 30938
rect 6184 30874 6236 30880
rect 6092 30796 6144 30802
rect 6092 30738 6144 30744
rect 6000 30728 6052 30734
rect 6000 30670 6052 30676
rect 6012 30394 6040 30670
rect 6000 30388 6052 30394
rect 6000 30330 6052 30336
rect 5908 30116 5960 30122
rect 5908 30058 5960 30064
rect 6012 29850 6040 30330
rect 6000 29844 6052 29850
rect 6000 29786 6052 29792
rect 6288 29714 6316 32166
rect 7392 31890 7420 32302
rect 6368 31884 6420 31890
rect 6368 31826 6420 31832
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 6380 31142 6408 31826
rect 7012 31340 7064 31346
rect 7012 31282 7064 31288
rect 7024 31210 7052 31282
rect 7012 31204 7064 31210
rect 7012 31146 7064 31152
rect 6368 31136 6420 31142
rect 6368 31078 6420 31084
rect 5908 29708 5960 29714
rect 5908 29650 5960 29656
rect 6276 29708 6328 29714
rect 6276 29650 6328 29656
rect 5354 29608 5410 29617
rect 5354 29543 5410 29552
rect 5172 29300 5224 29306
rect 5172 29242 5224 29248
rect 5920 28966 5948 29650
rect 5816 28960 5868 28966
rect 5816 28902 5868 28908
rect 5908 28960 5960 28966
rect 5908 28902 5960 28908
rect 5172 28688 5224 28694
rect 5172 28630 5224 28636
rect 5184 28218 5212 28630
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 5172 28212 5224 28218
rect 5172 28154 5224 28160
rect 5172 28008 5224 28014
rect 5172 27950 5224 27956
rect 4804 27600 4856 27606
rect 4804 27542 4856 27548
rect 4632 27118 4752 27146
rect 4252 26920 4304 26926
rect 4252 26862 4304 26868
rect 4264 26586 4292 26862
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 4252 26580 4304 26586
rect 4252 26522 4304 26528
rect 4632 26450 4660 27118
rect 4816 26858 4844 27542
rect 5184 27130 5212 27950
rect 5172 27124 5224 27130
rect 5172 27066 5224 27072
rect 4804 26852 4856 26858
rect 4804 26794 4856 26800
rect 4712 26512 4764 26518
rect 4712 26454 4764 26460
rect 4620 26444 4672 26450
rect 4620 26386 4672 26392
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 3976 25968 4028 25974
rect 3976 25910 4028 25916
rect 3700 25696 3752 25702
rect 3700 25638 3752 25644
rect 3608 24744 3660 24750
rect 3608 24686 3660 24692
rect 3424 24404 3476 24410
rect 3424 24346 3476 24352
rect 3436 23866 3464 24346
rect 3424 23860 3476 23866
rect 3424 23802 3476 23808
rect 3344 23718 3464 23746
rect 3332 23588 3384 23594
rect 3332 23530 3384 23536
rect 3344 22982 3372 23530
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 3344 21690 3372 22918
rect 3332 21684 3384 21690
rect 3332 21626 3384 21632
rect 3240 20528 3292 20534
rect 3240 20470 3292 20476
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 2872 19304 2924 19310
rect 2792 19264 2872 19292
rect 2872 19246 2924 19252
rect 2884 18970 2912 19246
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2884 17882 2912 18906
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2976 17338 3004 19314
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 3252 17082 3280 20470
rect 3436 19961 3464 23718
rect 3620 22710 3648 24686
rect 3712 24410 3740 25638
rect 3884 25424 3936 25430
rect 3884 25366 3936 25372
rect 3896 24954 3924 25366
rect 3884 24948 3936 24954
rect 3884 24890 3936 24896
rect 3988 24834 4016 25910
rect 4344 25832 4396 25838
rect 4344 25774 4396 25780
rect 4356 25498 4384 25774
rect 4632 25702 4660 26386
rect 4724 26042 4752 26454
rect 5368 26042 5396 28358
rect 5632 27532 5684 27538
rect 5632 27474 5684 27480
rect 5448 26852 5500 26858
rect 5448 26794 5500 26800
rect 4712 26036 4764 26042
rect 4712 25978 4764 25984
rect 4804 26036 4856 26042
rect 4804 25978 4856 25984
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 4620 25696 4672 25702
rect 4672 25656 4752 25684
rect 4620 25638 4672 25644
rect 4344 25492 4396 25498
rect 4344 25434 4396 25440
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 3896 24806 4016 24834
rect 3792 24744 3844 24750
rect 3792 24686 3844 24692
rect 3700 24404 3752 24410
rect 3700 24346 3752 24352
rect 3804 22982 3832 24686
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3608 22704 3660 22710
rect 3608 22646 3660 22652
rect 3804 22166 3832 22918
rect 3792 22160 3844 22166
rect 3792 22102 3844 22108
rect 3516 21956 3568 21962
rect 3516 21898 3568 21904
rect 3528 21690 3556 21898
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3528 21486 3556 21626
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3896 21010 3924 24806
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 3976 24336 4028 24342
rect 3976 24278 4028 24284
rect 3988 23866 4016 24278
rect 4172 24206 4200 24686
rect 4528 24676 4580 24682
rect 4528 24618 4580 24624
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4540 24138 4568 24618
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4528 24132 4580 24138
rect 4528 24074 4580 24080
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 4080 23798 4108 24006
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 4632 23730 4660 24142
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4252 23588 4304 23594
rect 4252 23530 4304 23536
rect 4264 23254 4292 23530
rect 4724 23474 4752 25656
rect 4632 23446 4752 23474
rect 3976 23248 4028 23254
rect 3976 23190 4028 23196
rect 4252 23248 4304 23254
rect 4252 23190 4304 23196
rect 3988 22778 4016 23190
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 3976 22772 4028 22778
rect 3976 22714 4028 22720
rect 3976 22500 4028 22506
rect 3976 22442 4028 22448
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 3896 20602 3924 20946
rect 3884 20596 3936 20602
rect 3884 20538 3936 20544
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3804 20058 3832 20334
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3422 19952 3478 19961
rect 3422 19887 3478 19896
rect 3792 19916 3844 19922
rect 3792 19858 3844 19864
rect 3804 19514 3832 19858
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3792 17740 3844 17746
rect 3792 17682 3844 17688
rect 3804 17338 3832 17682
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3252 17054 3372 17082
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3252 16658 3280 16934
rect 3344 16658 3372 17054
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 2700 16250 2728 16594
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 3160 16114 3188 16526
rect 3252 16250 3280 16594
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3712 15638 3740 16186
rect 3700 15632 3752 15638
rect 3700 15574 3752 15580
rect 3712 15162 3740 15574
rect 3896 15570 3924 20538
rect 3988 20466 4016 22442
rect 4080 22098 4108 22918
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4632 22642 4660 23446
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4724 22778 4752 23122
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4632 22234 4660 22578
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 4080 21690 4108 22034
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 4712 21412 4764 21418
rect 4712 21354 4764 21360
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4632 20466 4660 20946
rect 4724 20602 4752 21354
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 4724 20330 4752 20538
rect 4712 20324 4764 20330
rect 4712 20266 4764 20272
rect 4724 20058 4752 20266
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4080 18222 4108 19654
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4356 18970 4384 19246
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4632 18290 4660 19790
rect 4724 19446 4752 19994
rect 4816 19718 4844 25978
rect 4988 25152 5040 25158
rect 4988 25094 5040 25100
rect 5000 24818 5028 25094
rect 4988 24812 5040 24818
rect 4988 24754 5040 24760
rect 5264 24744 5316 24750
rect 5264 24686 5316 24692
rect 5080 24064 5132 24070
rect 5080 24006 5132 24012
rect 5092 23662 5120 24006
rect 5172 23792 5224 23798
rect 5172 23734 5224 23740
rect 5080 23656 5132 23662
rect 4894 23624 4950 23633
rect 4894 23559 4950 23568
rect 5000 23616 5080 23644
rect 4908 23526 4936 23559
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 5000 23118 5028 23616
rect 5080 23598 5132 23604
rect 5080 23520 5132 23526
rect 5080 23462 5132 23468
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5000 21554 5028 21830
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 5000 21078 5028 21490
rect 4988 21072 5040 21078
rect 4988 21014 5040 21020
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 4724 19174 4752 19382
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4724 18834 4752 19110
rect 5092 18834 5120 23462
rect 5184 23322 5212 23734
rect 5276 23662 5304 24686
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 5172 23316 5224 23322
rect 5172 23258 5224 23264
rect 5184 23050 5212 23258
rect 5276 23254 5304 23598
rect 5264 23248 5316 23254
rect 5264 23190 5316 23196
rect 5172 23044 5224 23050
rect 5172 22986 5224 22992
rect 5172 22500 5224 22506
rect 5172 22442 5224 22448
rect 5184 22030 5212 22442
rect 5460 22234 5488 26794
rect 5644 26790 5672 27474
rect 5632 26784 5684 26790
rect 5632 26726 5684 26732
rect 5644 26450 5672 26726
rect 5828 26586 5856 28902
rect 5816 26580 5868 26586
rect 5816 26522 5868 26528
rect 5632 26444 5684 26450
rect 5632 26386 5684 26392
rect 5644 25906 5672 26386
rect 5632 25900 5684 25906
rect 5632 25842 5684 25848
rect 5540 25356 5592 25362
rect 5540 25298 5592 25304
rect 5552 24614 5580 25298
rect 5920 24614 5948 28902
rect 6380 27538 6408 31078
rect 7024 30938 7052 31146
rect 7012 30932 7064 30938
rect 7012 30874 7064 30880
rect 7392 30598 7420 31826
rect 7484 31822 7512 32846
rect 7852 32298 7880 33050
rect 8404 32502 8432 33594
rect 8496 33318 8524 34002
rect 9508 33590 9536 34546
rect 9876 34474 9904 35974
rect 10152 35834 10180 36246
rect 10416 36168 10468 36174
rect 10416 36110 10468 36116
rect 11704 36168 11756 36174
rect 11704 36110 11756 36116
rect 10140 35828 10192 35834
rect 10140 35770 10192 35776
rect 10428 35562 10456 36110
rect 11716 35834 11744 36110
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 10416 35556 10468 35562
rect 10416 35498 10468 35504
rect 10876 35556 10928 35562
rect 10876 35498 10928 35504
rect 10428 35086 10456 35498
rect 10692 35488 10744 35494
rect 10692 35430 10744 35436
rect 10704 35222 10732 35430
rect 10692 35216 10744 35222
rect 10692 35158 10744 35164
rect 10416 35080 10468 35086
rect 10416 35022 10468 35028
rect 10428 34678 10456 35022
rect 10888 34950 10916 35498
rect 11716 35222 11744 35770
rect 11808 35766 11836 36246
rect 11992 36174 12020 36858
rect 12912 36378 12940 37198
rect 13004 36922 13032 37334
rect 13188 37262 13216 37674
rect 13648 37466 13676 37742
rect 13636 37460 13688 37466
rect 13636 37402 13688 37408
rect 13176 37256 13228 37262
rect 13176 37198 13228 37204
rect 13924 36922 13952 37810
rect 12992 36916 13044 36922
rect 12992 36858 13044 36864
rect 13912 36916 13964 36922
rect 13912 36858 13964 36864
rect 13924 36632 13952 36858
rect 14280 36780 14332 36786
rect 14280 36722 14332 36728
rect 14648 36780 14700 36786
rect 14648 36722 14700 36728
rect 14004 36644 14056 36650
rect 13924 36604 14004 36632
rect 14004 36586 14056 36592
rect 12900 36372 12952 36378
rect 12900 36314 12952 36320
rect 14004 36236 14056 36242
rect 14004 36178 14056 36184
rect 11980 36168 12032 36174
rect 11980 36110 12032 36116
rect 11796 35760 11848 35766
rect 11796 35702 11848 35708
rect 11704 35216 11756 35222
rect 11704 35158 11756 35164
rect 11152 35012 11204 35018
rect 11152 34954 11204 34960
rect 10876 34944 10928 34950
rect 10876 34886 10928 34892
rect 10888 34746 10916 34886
rect 10876 34740 10928 34746
rect 10876 34682 10928 34688
rect 11164 34678 11192 34954
rect 10416 34672 10468 34678
rect 10416 34614 10468 34620
rect 11152 34672 11204 34678
rect 11152 34614 11204 34620
rect 11808 34474 11836 35702
rect 11992 35698 12020 36110
rect 13636 36032 13688 36038
rect 13636 35974 13688 35980
rect 13648 35698 13676 35974
rect 11980 35692 12032 35698
rect 11980 35634 12032 35640
rect 13636 35692 13688 35698
rect 13636 35634 13688 35640
rect 13452 35556 13504 35562
rect 13452 35498 13504 35504
rect 13728 35556 13780 35562
rect 13728 35498 13780 35504
rect 12900 35488 12952 35494
rect 12900 35430 12952 35436
rect 11888 35148 11940 35154
rect 11888 35090 11940 35096
rect 9864 34468 9916 34474
rect 9864 34410 9916 34416
rect 11796 34468 11848 34474
rect 11796 34410 11848 34416
rect 9588 34128 9640 34134
rect 9588 34070 9640 34076
rect 9600 33590 9628 34070
rect 9876 33998 9904 34410
rect 11900 34406 11928 35090
rect 12716 35080 12768 35086
rect 12716 35022 12768 35028
rect 12256 34536 12308 34542
rect 12256 34478 12308 34484
rect 11888 34400 11940 34406
rect 11888 34342 11940 34348
rect 12268 34202 12296 34478
rect 12348 34400 12400 34406
rect 12348 34342 12400 34348
rect 12256 34196 12308 34202
rect 12256 34138 12308 34144
rect 11888 34128 11940 34134
rect 11888 34070 11940 34076
rect 9772 33992 9824 33998
rect 9772 33934 9824 33940
rect 9864 33992 9916 33998
rect 9864 33934 9916 33940
rect 11336 33992 11388 33998
rect 11336 33934 11388 33940
rect 9784 33658 9812 33934
rect 11348 33658 11376 33934
rect 9772 33652 9824 33658
rect 9772 33594 9824 33600
rect 11336 33652 11388 33658
rect 11336 33594 11388 33600
rect 9496 33584 9548 33590
rect 9496 33526 9548 33532
rect 9588 33584 9640 33590
rect 9588 33526 9640 33532
rect 9588 33448 9640 33454
rect 9588 33390 9640 33396
rect 8852 33380 8904 33386
rect 8852 33322 8904 33328
rect 8484 33312 8536 33318
rect 8484 33254 8536 33260
rect 8496 33114 8524 33254
rect 8484 33108 8536 33114
rect 8484 33050 8536 33056
rect 8864 32570 8892 33322
rect 9600 33114 9628 33390
rect 11348 33134 11376 33594
rect 11520 33448 11572 33454
rect 11520 33390 11572 33396
rect 9588 33108 9640 33114
rect 9588 33050 9640 33056
rect 11256 33106 11376 33134
rect 10416 32904 10468 32910
rect 10416 32846 10468 32852
rect 8852 32564 8904 32570
rect 8852 32506 8904 32512
rect 8392 32496 8444 32502
rect 8392 32438 8444 32444
rect 8300 32428 8352 32434
rect 8300 32370 8352 32376
rect 7840 32292 7892 32298
rect 7840 32234 7892 32240
rect 7472 31816 7524 31822
rect 7472 31758 7524 31764
rect 7840 31748 7892 31754
rect 7840 31690 7892 31696
rect 7852 30870 7880 31690
rect 8312 31686 8340 32370
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 9692 32026 9720 32302
rect 10428 32230 10456 32846
rect 11152 32360 11204 32366
rect 11152 32302 11204 32308
rect 10416 32224 10468 32230
rect 10416 32166 10468 32172
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 8392 31884 8444 31890
rect 8392 31826 8444 31832
rect 9588 31884 9640 31890
rect 9588 31826 9640 31832
rect 10140 31884 10192 31890
rect 10140 31826 10192 31832
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 7840 30864 7892 30870
rect 7840 30806 7892 30812
rect 7472 30796 7524 30802
rect 7472 30738 7524 30744
rect 6736 30592 6788 30598
rect 6736 30534 6788 30540
rect 7380 30592 7432 30598
rect 7380 30534 7432 30540
rect 6460 29640 6512 29646
rect 6460 29582 6512 29588
rect 6472 28694 6500 29582
rect 6460 28688 6512 28694
rect 6460 28630 6512 28636
rect 6552 28688 6604 28694
rect 6552 28630 6604 28636
rect 6460 28552 6512 28558
rect 6460 28494 6512 28500
rect 6472 28150 6500 28494
rect 6564 28218 6592 28630
rect 6552 28212 6604 28218
rect 6552 28154 6604 28160
rect 6460 28144 6512 28150
rect 6460 28086 6512 28092
rect 6472 27674 6500 28086
rect 6460 27668 6512 27674
rect 6460 27610 6512 27616
rect 6368 27532 6420 27538
rect 6368 27474 6420 27480
rect 6000 25696 6052 25702
rect 6000 25638 6052 25644
rect 6012 25430 6040 25638
rect 6000 25424 6052 25430
rect 6000 25366 6052 25372
rect 6368 25356 6420 25362
rect 6368 25298 6420 25304
rect 6380 24886 6408 25298
rect 6748 25294 6776 30534
rect 7484 30258 7512 30738
rect 7472 30252 7524 30258
rect 7472 30194 7524 30200
rect 7564 30116 7616 30122
rect 7564 30058 7616 30064
rect 7576 29782 7604 30058
rect 7852 29850 7880 30806
rect 8116 30728 8168 30734
rect 8116 30670 8168 30676
rect 8128 30258 8156 30670
rect 8116 30252 8168 30258
rect 8116 30194 8168 30200
rect 7840 29844 7892 29850
rect 7840 29786 7892 29792
rect 7564 29776 7616 29782
rect 7564 29718 7616 29724
rect 7932 29776 7984 29782
rect 7932 29718 7984 29724
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6932 29034 6960 29446
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 6920 29028 6972 29034
rect 6920 28970 6972 28976
rect 6932 28762 6960 28970
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 7208 28694 7236 29106
rect 7944 28966 7972 29718
rect 8208 29640 8260 29646
rect 8208 29582 8260 29588
rect 8220 29306 8248 29582
rect 8208 29300 8260 29306
rect 8208 29242 8260 29248
rect 7932 28960 7984 28966
rect 7932 28902 7984 28908
rect 7944 28762 7972 28902
rect 7932 28756 7984 28762
rect 7932 28698 7984 28704
rect 7196 28688 7248 28694
rect 7196 28630 7248 28636
rect 7656 28620 7708 28626
rect 7656 28562 7708 28568
rect 7668 28218 7696 28562
rect 7656 28212 7708 28218
rect 7656 28154 7708 28160
rect 7564 28008 7616 28014
rect 7564 27950 7616 27956
rect 7012 27532 7064 27538
rect 7012 27474 7064 27480
rect 6828 27464 6880 27470
rect 6828 27406 6880 27412
rect 6840 26994 6868 27406
rect 7024 27130 7052 27474
rect 7576 27334 7604 27950
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 7012 27124 7064 27130
rect 7012 27066 7064 27072
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6920 26852 6972 26858
rect 6920 26794 6972 26800
rect 6932 26586 6960 26794
rect 6920 26580 6972 26586
rect 6840 26540 6920 26568
rect 6840 26042 6868 26540
rect 6920 26522 6972 26528
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 6828 25764 6880 25770
rect 6828 25706 6880 25712
rect 6840 25430 6868 25706
rect 6932 25702 6960 26318
rect 6920 25696 6972 25702
rect 6920 25638 6972 25644
rect 6932 25498 6960 25638
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 6828 25424 6880 25430
rect 6828 25366 6880 25372
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6368 24880 6420 24886
rect 6368 24822 6420 24828
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5908 24608 5960 24614
rect 5908 24550 5960 24556
rect 5552 23662 5580 24550
rect 5816 24268 5868 24274
rect 5816 24210 5868 24216
rect 5724 24132 5776 24138
rect 5724 24074 5776 24080
rect 5736 23798 5764 24074
rect 5724 23792 5776 23798
rect 5724 23734 5776 23740
rect 5632 23724 5684 23730
rect 5632 23666 5684 23672
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5552 23186 5580 23598
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 5644 22982 5672 23666
rect 5828 23322 5856 24210
rect 5920 23526 5948 24550
rect 6380 24342 6408 24822
rect 6644 24608 6696 24614
rect 6644 24550 6696 24556
rect 6656 24410 6684 24550
rect 6644 24404 6696 24410
rect 6644 24346 6696 24352
rect 6748 24342 6776 25230
rect 6368 24336 6420 24342
rect 6368 24278 6420 24284
rect 6736 24336 6788 24342
rect 6736 24278 6788 24284
rect 6000 24268 6052 24274
rect 6000 24210 6052 24216
rect 6012 23633 6040 24210
rect 6644 23656 6696 23662
rect 5998 23624 6054 23633
rect 6644 23598 6696 23604
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 5998 23559 6054 23568
rect 6012 23526 6040 23559
rect 6656 23526 6684 23598
rect 5908 23520 5960 23526
rect 5908 23462 5960 23468
rect 6000 23520 6052 23526
rect 6000 23462 6052 23468
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 5816 23316 5868 23322
rect 5816 23258 5868 23264
rect 6656 23254 6684 23462
rect 6644 23248 6696 23254
rect 6644 23190 6696 23196
rect 6748 23186 6776 23598
rect 6736 23180 6788 23186
rect 6736 23122 6788 23128
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 5908 22976 5960 22982
rect 5908 22918 5960 22924
rect 5644 22710 5672 22918
rect 5920 22710 5948 22918
rect 6012 22778 6040 23054
rect 6000 22772 6052 22778
rect 6000 22714 6052 22720
rect 5632 22704 5684 22710
rect 5632 22646 5684 22652
rect 5908 22704 5960 22710
rect 5908 22646 5960 22652
rect 6748 22234 6776 23122
rect 6828 22976 6880 22982
rect 6828 22918 6880 22924
rect 6840 22574 6868 22918
rect 7024 22778 7052 27066
rect 7576 26586 7604 27270
rect 7668 27130 7696 28154
rect 7944 27946 7972 28698
rect 8208 28416 8260 28422
rect 8208 28358 8260 28364
rect 8220 28082 8248 28358
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 7932 27940 7984 27946
rect 7932 27882 7984 27888
rect 7840 27872 7892 27878
rect 7840 27814 7892 27820
rect 7852 27606 7880 27814
rect 7840 27600 7892 27606
rect 7840 27542 7892 27548
rect 7852 27130 7880 27542
rect 7656 27124 7708 27130
rect 7656 27066 7708 27072
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7748 26920 7800 26926
rect 7748 26862 7800 26868
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 7656 25832 7708 25838
rect 7656 25774 7708 25780
rect 7472 25492 7524 25498
rect 7472 25434 7524 25440
rect 7484 24750 7512 25434
rect 7668 25362 7696 25774
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 7104 23588 7156 23594
rect 7104 23530 7156 23536
rect 7116 23186 7144 23530
rect 7104 23180 7156 23186
rect 7104 23122 7156 23128
rect 7208 23050 7236 24210
rect 7392 23254 7420 24210
rect 7564 24132 7616 24138
rect 7564 24074 7616 24080
rect 7576 23662 7604 24074
rect 7668 24070 7696 25298
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7380 23248 7432 23254
rect 7380 23190 7432 23196
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 7300 22778 7328 23122
rect 7012 22772 7064 22778
rect 7288 22772 7340 22778
rect 7064 22732 7144 22760
rect 7012 22714 7064 22720
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 6736 22228 6788 22234
rect 6736 22170 6788 22176
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5184 21146 5212 21966
rect 5460 21690 5488 22170
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5460 21418 5488 21626
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 5172 21140 5224 21146
rect 5172 21082 5224 21088
rect 5552 21010 5580 21286
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5552 20602 5580 20946
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 6748 20466 6776 21286
rect 7024 21146 7052 21966
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 7116 21010 7144 22732
rect 7288 22714 7340 22720
rect 7196 22160 7248 22166
rect 7196 22102 7248 22108
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 7012 20800 7064 20806
rect 7208 20788 7236 22102
rect 7564 21956 7616 21962
rect 7564 21898 7616 21904
rect 7576 21418 7604 21898
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7064 20760 7236 20788
rect 7012 20742 7064 20748
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 5724 20324 5776 20330
rect 5724 20266 5776 20272
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 5184 19514 5212 20198
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 5092 18426 5120 18770
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4068 18216 4120 18222
rect 3988 18176 4068 18204
rect 3988 17338 4016 18176
rect 4068 18158 4120 18164
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 3988 17134 4016 17274
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3988 16250 4016 16594
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3896 15162 3924 15506
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3712 14074 3740 14350
rect 4080 14074 4108 17818
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4632 17134 4660 17682
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4632 16658 4660 17070
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4632 15638 4660 16594
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4724 15706 4752 15982
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4620 15632 4672 15638
rect 4620 15574 4672 15580
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4632 15026 4660 15438
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4620 13864 4672 13870
rect 4816 13814 4844 17002
rect 5092 16658 5120 18362
rect 5276 17746 5304 19654
rect 5552 19514 5580 19790
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5460 18222 5488 19110
rect 5736 18834 5764 20266
rect 6748 19990 6776 20402
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6380 19242 6408 19654
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 5736 18358 5764 18770
rect 5724 18352 5776 18358
rect 5724 18294 5776 18300
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 6380 17882 6408 19178
rect 6564 18970 6592 19722
rect 6748 19446 6776 19926
rect 7024 19514 7052 20742
rect 7576 20505 7604 21354
rect 7668 20602 7696 24006
rect 7760 23730 7788 26862
rect 8208 25696 8260 25702
rect 8208 25638 8260 25644
rect 8220 24818 8248 25638
rect 8312 25430 8340 31622
rect 8404 31142 8432 31826
rect 8852 31204 8904 31210
rect 8852 31146 8904 31152
rect 8944 31204 8996 31210
rect 8944 31146 8996 31152
rect 8392 31136 8444 31142
rect 8392 31078 8444 31084
rect 8404 30297 8432 31078
rect 8864 30938 8892 31146
rect 8852 30932 8904 30938
rect 8852 30874 8904 30880
rect 8484 30864 8536 30870
rect 8484 30806 8536 30812
rect 8390 30288 8446 30297
rect 8390 30223 8446 30232
rect 8496 30054 8524 30806
rect 8484 30048 8536 30054
rect 8484 29990 8536 29996
rect 8496 29034 8524 29990
rect 8864 29782 8892 30874
rect 8852 29776 8904 29782
rect 8852 29718 8904 29724
rect 8484 29028 8536 29034
rect 8484 28970 8536 28976
rect 8496 27606 8524 28970
rect 8956 28966 8984 31146
rect 9600 31142 9628 31826
rect 10152 31346 10180 31826
rect 10140 31340 10192 31346
rect 10140 31282 10192 31288
rect 9680 31204 9732 31210
rect 9680 31146 9732 31152
rect 9588 31136 9640 31142
rect 9588 31078 9640 31084
rect 9036 30252 9088 30258
rect 9036 30194 9088 30200
rect 9048 29850 9076 30194
rect 9496 30116 9548 30122
rect 9496 30058 9548 30064
rect 9036 29844 9088 29850
rect 9036 29786 9088 29792
rect 9128 29028 9180 29034
rect 9128 28970 9180 28976
rect 8944 28960 8996 28966
rect 8944 28902 8996 28908
rect 9140 28694 9168 28970
rect 9508 28762 9536 30058
rect 9496 28756 9548 28762
rect 9496 28698 9548 28704
rect 9128 28688 9180 28694
rect 9128 28630 9180 28636
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9324 28218 9352 28494
rect 9312 28212 9364 28218
rect 9312 28154 9364 28160
rect 8760 28144 8812 28150
rect 8760 28086 8812 28092
rect 8772 27606 8800 28086
rect 8484 27600 8536 27606
rect 8484 27542 8536 27548
rect 8760 27600 8812 27606
rect 8760 27542 8812 27548
rect 8496 27062 8524 27542
rect 9600 27470 9628 31078
rect 9692 30122 9720 31146
rect 10152 31142 10180 31282
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 10048 30796 10100 30802
rect 10048 30738 10100 30744
rect 10060 30394 10088 30738
rect 10152 30598 10180 31078
rect 10140 30592 10192 30598
rect 10140 30534 10192 30540
rect 10324 30592 10376 30598
rect 10324 30534 10376 30540
rect 10048 30388 10100 30394
rect 10048 30330 10100 30336
rect 9680 30116 9732 30122
rect 9680 30058 9732 30064
rect 9692 28937 9720 30058
rect 10140 29708 10192 29714
rect 10140 29650 10192 29656
rect 9862 29064 9918 29073
rect 9862 28999 9864 29008
rect 9916 28999 9918 29008
rect 9864 28970 9916 28976
rect 9678 28928 9734 28937
rect 9678 28863 9734 28872
rect 9876 28694 9904 28970
rect 10152 28966 10180 29650
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 9864 28688 9916 28694
rect 9864 28630 9916 28636
rect 9876 28218 9904 28630
rect 9864 28212 9916 28218
rect 9864 28154 9916 28160
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 9956 27872 10008 27878
rect 9956 27814 10008 27820
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 8484 27056 8536 27062
rect 8484 26998 8536 27004
rect 9600 26926 9628 27406
rect 9692 27062 9720 27814
rect 9772 27668 9824 27674
rect 9772 27610 9824 27616
rect 9680 27056 9732 27062
rect 9680 26998 9732 27004
rect 9784 26994 9812 27610
rect 9864 27532 9916 27538
rect 9864 27474 9916 27480
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8588 25906 8616 26386
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 8772 25498 8800 26726
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8300 25424 8352 25430
rect 8300 25366 8352 25372
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 7840 23724 7892 23730
rect 7944 23712 7972 24686
rect 8772 24682 8800 25434
rect 8944 25152 8996 25158
rect 8944 25094 8996 25100
rect 8956 24750 8984 25094
rect 8944 24744 8996 24750
rect 8944 24686 8996 24692
rect 8576 24676 8628 24682
rect 8576 24618 8628 24624
rect 8760 24676 8812 24682
rect 8760 24618 8812 24624
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8128 23866 8156 24550
rect 8588 24274 8616 24618
rect 8576 24268 8628 24274
rect 8576 24210 8628 24216
rect 8588 23866 8616 24210
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 7892 23684 7972 23712
rect 7840 23666 7892 23672
rect 7852 23322 7880 23666
rect 7840 23316 7892 23322
rect 7840 23258 7892 23264
rect 7852 22778 7880 23258
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 7852 22506 7880 22714
rect 8128 22574 8156 23802
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8300 23588 8352 23594
rect 8300 23530 8352 23536
rect 8208 23316 8260 23322
rect 8208 23258 8260 23264
rect 8220 23186 8248 23258
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 8220 22778 8248 23122
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8116 22568 8168 22574
rect 8116 22510 8168 22516
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 8128 21486 8156 22510
rect 8312 22098 8340 23530
rect 8404 23186 8432 23598
rect 8392 23180 8444 23186
rect 8392 23122 8444 23128
rect 8404 22982 8432 23122
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8404 22234 8432 22918
rect 8772 22545 8800 24006
rect 8956 23730 8984 24686
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 8944 23724 8996 23730
rect 8944 23666 8996 23672
rect 8956 23633 8984 23666
rect 9140 23662 9168 24006
rect 9128 23656 9180 23662
rect 8942 23624 8998 23633
rect 9128 23598 9180 23604
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9496 23656 9548 23662
rect 9496 23598 9548 23604
rect 8942 23559 8998 23568
rect 9232 23322 9260 23598
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9508 23254 9536 23598
rect 9496 23248 9548 23254
rect 9496 23190 9548 23196
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 8758 22536 8814 22545
rect 8758 22471 8814 22480
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 8312 21690 8340 22034
rect 8404 21690 8432 22170
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 8404 21418 8432 21626
rect 8392 21412 8444 21418
rect 8392 21354 8444 21360
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7562 20496 7618 20505
rect 7562 20431 7618 20440
rect 7668 20398 7696 20538
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6748 18358 6776 19382
rect 7024 19242 7052 19450
rect 7576 19242 7604 19790
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7576 19009 7604 19178
rect 7562 19000 7618 19009
rect 7104 18964 7156 18970
rect 7562 18935 7618 18944
rect 7104 18906 7156 18912
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 7116 18086 7144 18906
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 18426 7236 18566
rect 7392 18426 7420 18702
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5276 17338 5304 17682
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6104 16658 6132 16934
rect 7116 16726 7144 18022
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7576 17134 7604 17682
rect 7668 17202 7696 20334
rect 7760 20058 7788 20946
rect 8220 20398 8248 20946
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8300 20324 8352 20330
rect 8300 20266 8352 20272
rect 8312 20058 8340 20266
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 7760 17814 7788 19994
rect 8864 19922 8892 20198
rect 9140 19922 9168 22442
rect 7932 19916 7984 19922
rect 7932 19858 7984 19864
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 7944 19514 7972 19858
rect 8864 19718 8892 19858
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 8312 18630 8340 19178
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8496 18290 8524 18566
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8496 17882 8524 18226
rect 8588 17882 8616 18770
rect 8864 18465 8892 19314
rect 8850 18456 8906 18465
rect 8850 18391 8906 18400
rect 8864 18290 8892 18391
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 7748 17808 7800 17814
rect 7800 17768 7880 17796
rect 7748 17750 7800 17756
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7104 16720 7156 16726
rect 7104 16662 7156 16668
rect 7576 16658 7604 17070
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7668 16794 7696 17002
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4908 14482 4936 16526
rect 5920 16250 5948 16594
rect 6104 16250 6132 16594
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5000 14890 5028 15846
rect 5828 14958 5856 15846
rect 6380 15570 6408 16526
rect 7668 16114 7696 16730
rect 7760 16658 7788 17614
rect 7852 17338 7880 17768
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 7760 16250 7788 16594
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 6472 15638 6500 15914
rect 7668 15706 7696 15914
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6276 15156 6328 15162
rect 6380 15144 6408 15506
rect 6328 15116 6408 15144
rect 6276 15098 6328 15104
rect 6472 15026 6500 15574
rect 8496 15570 8524 15846
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 6460 15020 6512 15026
rect 6460 14962 6512 14968
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 5000 14550 5028 14826
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 5000 13870 5028 14486
rect 4620 13806 4672 13812
rect 4632 13530 4660 13806
rect 4724 13786 4844 13814
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4632 12850 4660 13466
rect 4724 13394 4752 13786
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4724 12986 4752 13330
rect 5368 12986 5396 14758
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 5368 12782 5396 12922
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5460 12306 5488 13670
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 5552 11694 5580 14214
rect 6840 14006 6868 14554
rect 6932 14414 6960 14758
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6932 14074 6960 14350
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6748 13190 6776 13738
rect 6840 13734 6868 13942
rect 7116 13938 7144 15030
rect 7576 14482 7604 15302
rect 8496 15162 8524 15506
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7484 14006 7512 14282
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7012 13796 7064 13802
rect 7116 13784 7144 13874
rect 8496 13802 8524 14758
rect 7064 13756 7144 13784
rect 7012 13738 7064 13744
rect 6828 13728 6880 13734
rect 6880 13688 6960 13716
rect 6828 13670 6880 13676
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6748 12986 6776 13126
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6840 12374 6868 13194
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6932 12322 6960 13688
rect 7116 13462 7144 13756
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7024 12442 7052 12786
rect 7116 12714 7144 13398
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7668 12696 7696 13262
rect 7748 12708 7800 12714
rect 7668 12668 7748 12696
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7668 12374 7696 12668
rect 7748 12650 7800 12656
rect 7104 12368 7156 12374
rect 6932 12316 7104 12322
rect 6932 12310 7156 12316
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 6092 12300 6144 12306
rect 6932 12294 7144 12310
rect 8588 12306 8616 16390
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8864 14890 8892 15302
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 13938 8708 14214
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8864 12442 8892 14826
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9140 12918 9168 13738
rect 9232 13394 9260 23122
rect 9508 22778 9536 23190
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9600 22234 9628 26862
rect 9876 26246 9904 27474
rect 9968 26314 9996 27814
rect 10152 26586 10180 28902
rect 10140 26580 10192 26586
rect 10140 26522 10192 26528
rect 10336 26518 10364 30534
rect 10324 26512 10376 26518
rect 10324 26454 10376 26460
rect 10232 26376 10284 26382
rect 10232 26318 10284 26324
rect 9956 26308 10008 26314
rect 9956 26250 10008 26256
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9876 25702 9904 26182
rect 9956 25832 10008 25838
rect 9956 25774 10008 25780
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9968 25362 9996 25774
rect 10244 25770 10272 26318
rect 10232 25764 10284 25770
rect 10232 25706 10284 25712
rect 10244 25498 10272 25706
rect 10232 25492 10284 25498
rect 10232 25434 10284 25440
rect 9956 25356 10008 25362
rect 9956 25298 10008 25304
rect 9968 24954 9996 25298
rect 9956 24948 10008 24954
rect 9956 24890 10008 24896
rect 9968 24410 9996 24890
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 9968 23474 9996 24346
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 10152 23730 10180 24142
rect 10140 23724 10192 23730
rect 10140 23666 10192 23672
rect 9784 23446 9996 23474
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9692 22438 9720 23122
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9404 21616 9456 21622
rect 9404 21558 9456 21564
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9324 20058 9352 20334
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9416 19242 9444 21558
rect 9600 19310 9628 22170
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9692 21554 9720 22034
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9692 19514 9720 19858
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9404 19236 9456 19242
rect 9404 19178 9456 19184
rect 9784 18426 9812 23446
rect 9954 23080 10010 23089
rect 9864 23044 9916 23050
rect 9916 23024 9954 23032
rect 9916 23015 10010 23024
rect 9916 23004 9996 23015
rect 9864 22986 9916 22992
rect 10140 22432 10192 22438
rect 10244 22420 10272 23462
rect 10192 22392 10272 22420
rect 10140 22374 10192 22380
rect 10152 21962 10180 22374
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 10232 21888 10284 21894
rect 10232 21830 10284 21836
rect 10244 19786 10272 21830
rect 10336 19990 10364 26454
rect 10428 25430 10456 32166
rect 11164 31278 11192 32302
rect 11256 32026 11284 33106
rect 11428 33040 11480 33046
rect 11428 32982 11480 32988
rect 11440 32298 11468 32982
rect 11428 32292 11480 32298
rect 11428 32234 11480 32240
rect 11244 32020 11296 32026
rect 11244 31962 11296 31968
rect 11428 31884 11480 31890
rect 11428 31826 11480 31832
rect 10784 31272 10836 31278
rect 10784 31214 10836 31220
rect 11152 31272 11204 31278
rect 11152 31214 11204 31220
rect 10796 30326 10824 31214
rect 10876 31136 10928 31142
rect 10876 31078 10928 31084
rect 10784 30320 10836 30326
rect 10784 30262 10836 30268
rect 10692 30048 10744 30054
rect 10692 29990 10744 29996
rect 10704 27946 10732 29990
rect 10796 29714 10824 30262
rect 10888 30258 10916 31078
rect 10968 30728 11020 30734
rect 10968 30670 11020 30676
rect 10876 30252 10928 30258
rect 10876 30194 10928 30200
rect 10888 29850 10916 30194
rect 10980 29850 11008 30670
rect 11164 30598 11192 31214
rect 11440 31142 11468 31826
rect 11428 31136 11480 31142
rect 11428 31078 11480 31084
rect 11244 30864 11296 30870
rect 11244 30806 11296 30812
rect 11152 30592 11204 30598
rect 11152 30534 11204 30540
rect 11256 30122 11284 30806
rect 11244 30116 11296 30122
rect 11244 30058 11296 30064
rect 10876 29844 10928 29850
rect 10876 29786 10928 29792
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 11440 29714 11468 31078
rect 11532 30394 11560 33390
rect 11900 33386 11928 34070
rect 11888 33380 11940 33386
rect 11888 33322 11940 33328
rect 11900 33046 11928 33322
rect 12360 33114 12388 34342
rect 12728 33862 12756 35022
rect 12912 34746 12940 35430
rect 13084 35284 13136 35290
rect 13084 35226 13136 35232
rect 12900 34740 12952 34746
rect 12900 34682 12952 34688
rect 13096 34474 13124 35226
rect 13084 34468 13136 34474
rect 13084 34410 13136 34416
rect 12716 33856 12768 33862
rect 12716 33798 12768 33804
rect 13268 33856 13320 33862
rect 13268 33798 13320 33804
rect 12440 33312 12492 33318
rect 12440 33254 12492 33260
rect 12348 33108 12400 33114
rect 12348 33050 12400 33056
rect 11888 33040 11940 33046
rect 11888 32982 11940 32988
rect 11888 32904 11940 32910
rect 11888 32846 11940 32852
rect 11900 32298 11928 32846
rect 11888 32292 11940 32298
rect 11888 32234 11940 32240
rect 12072 31952 12124 31958
rect 12072 31894 12124 31900
rect 12084 31793 12112 31894
rect 12256 31884 12308 31890
rect 12256 31826 12308 31832
rect 12070 31784 12126 31793
rect 12070 31719 12126 31728
rect 12268 31686 12296 31826
rect 12256 31680 12308 31686
rect 12256 31622 12308 31628
rect 12268 30870 12296 31622
rect 12256 30864 12308 30870
rect 12256 30806 12308 30812
rect 11520 30388 11572 30394
rect 11520 30330 11572 30336
rect 12256 30320 12308 30326
rect 12256 30262 12308 30268
rect 10784 29708 10836 29714
rect 10784 29650 10836 29656
rect 11428 29708 11480 29714
rect 11428 29650 11480 29656
rect 10796 29306 10824 29650
rect 10784 29300 10836 29306
rect 10784 29242 10836 29248
rect 10784 29096 10836 29102
rect 10784 29038 10836 29044
rect 10692 27940 10744 27946
rect 10692 27882 10744 27888
rect 10796 27130 10824 29038
rect 11440 28966 11468 29650
rect 11520 29504 11572 29510
rect 11520 29446 11572 29452
rect 10876 28960 10928 28966
rect 10876 28902 10928 28908
rect 11428 28960 11480 28966
rect 11428 28902 11480 28908
rect 10888 28082 10916 28902
rect 10876 28076 10928 28082
rect 10876 28018 10928 28024
rect 10888 27674 10916 28018
rect 10876 27668 10928 27674
rect 10876 27610 10928 27616
rect 10784 27124 10836 27130
rect 10784 27066 10836 27072
rect 10600 26852 10652 26858
rect 10600 26794 10652 26800
rect 10612 26518 10640 26794
rect 10600 26512 10652 26518
rect 10600 26454 10652 26460
rect 10612 25974 10640 26454
rect 10600 25968 10652 25974
rect 10600 25910 10652 25916
rect 11152 25900 11204 25906
rect 11152 25842 11204 25848
rect 10416 25424 10468 25430
rect 10416 25366 10468 25372
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10704 24410 10732 24550
rect 11164 24410 11192 25842
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 11256 24342 11284 24550
rect 11244 24336 11296 24342
rect 11244 24278 11296 24284
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10692 24132 10744 24138
rect 10692 24074 10744 24080
rect 10704 23644 10732 24074
rect 11072 23866 11100 24210
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 10784 23656 10836 23662
rect 10704 23616 10784 23644
rect 10704 23322 10732 23616
rect 10784 23598 10836 23604
rect 11072 23474 11100 23802
rect 11256 23662 11284 24278
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 11072 23446 11192 23474
rect 10692 23316 10744 23322
rect 10692 23258 10744 23264
rect 10704 22574 10732 23258
rect 11164 23254 11192 23446
rect 11152 23248 11204 23254
rect 11152 23190 11204 23196
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 10692 22568 10744 22574
rect 10692 22510 10744 22516
rect 10600 22500 10652 22506
rect 10600 22442 10652 22448
rect 10612 21894 10640 22442
rect 10704 22234 10732 22510
rect 11072 22506 11100 23122
rect 11164 22778 11192 23190
rect 11152 22772 11204 22778
rect 11152 22714 11204 22720
rect 11440 22692 11468 28902
rect 11532 28694 11560 29446
rect 11612 29232 11664 29238
rect 11612 29174 11664 29180
rect 11624 28694 11652 29174
rect 12164 28756 12216 28762
rect 12164 28698 12216 28704
rect 11520 28688 11572 28694
rect 11520 28630 11572 28636
rect 11612 28688 11664 28694
rect 11612 28630 11664 28636
rect 11532 28218 11560 28630
rect 11520 28212 11572 28218
rect 11520 28154 11572 28160
rect 11624 28150 11652 28630
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 11612 28144 11664 28150
rect 11612 28086 11664 28092
rect 11992 26994 12020 28494
rect 12176 28082 12204 28698
rect 12164 28076 12216 28082
rect 12164 28018 12216 28024
rect 12176 27130 12204 28018
rect 12268 27538 12296 30262
rect 12452 29646 12480 33254
rect 13280 33114 13308 33798
rect 13360 33448 13412 33454
rect 13360 33390 13412 33396
rect 13268 33108 13320 33114
rect 13268 33050 13320 33056
rect 12992 32768 13044 32774
rect 12992 32710 13044 32716
rect 13004 32366 13032 32710
rect 12992 32360 13044 32366
rect 12992 32302 13044 32308
rect 13004 31686 13032 32302
rect 13268 31884 13320 31890
rect 13268 31826 13320 31832
rect 12992 31680 13044 31686
rect 12992 31622 13044 31628
rect 13280 31346 13308 31826
rect 13268 31340 13320 31346
rect 13268 31282 13320 31288
rect 12532 31204 12584 31210
rect 12532 31146 12584 31152
rect 13176 31204 13228 31210
rect 13176 31146 13228 31152
rect 12544 30938 12572 31146
rect 12900 31136 12952 31142
rect 12900 31078 12952 31084
rect 12532 30932 12584 30938
rect 12532 30874 12584 30880
rect 12716 29776 12768 29782
rect 12716 29718 12768 29724
rect 12440 29640 12492 29646
rect 12440 29582 12492 29588
rect 12532 29640 12584 29646
rect 12532 29582 12584 29588
rect 12452 28626 12480 29582
rect 12544 29034 12572 29582
rect 12728 29238 12756 29718
rect 12716 29232 12768 29238
rect 12716 29174 12768 29180
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 12532 29028 12584 29034
rect 12532 28970 12584 28976
rect 12544 28694 12572 28970
rect 12820 28762 12848 29106
rect 12808 28756 12860 28762
rect 12808 28698 12860 28704
rect 12532 28688 12584 28694
rect 12532 28630 12584 28636
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12544 27946 12572 28494
rect 12808 28008 12860 28014
rect 12808 27950 12860 27956
rect 12532 27940 12584 27946
rect 12532 27882 12584 27888
rect 12256 27532 12308 27538
rect 12256 27474 12308 27480
rect 12164 27124 12216 27130
rect 12164 27066 12216 27072
rect 11980 26988 12032 26994
rect 11980 26930 12032 26936
rect 12268 26926 12296 27474
rect 12256 26920 12308 26926
rect 12256 26862 12308 26868
rect 12268 26586 12296 26862
rect 12544 26858 12572 27882
rect 12820 27606 12848 27950
rect 12912 27878 12940 31078
rect 12992 30048 13044 30054
rect 12992 29990 13044 29996
rect 13004 29306 13032 29990
rect 13188 29782 13216 31146
rect 13372 30802 13400 33390
rect 13464 33114 13492 35498
rect 13740 35222 13768 35498
rect 14016 35290 14044 36178
rect 14292 35698 14320 36722
rect 14660 36378 14688 36722
rect 14648 36372 14700 36378
rect 14648 36314 14700 36320
rect 14280 35692 14332 35698
rect 14280 35634 14332 35640
rect 14556 35488 14608 35494
rect 14556 35430 14608 35436
rect 14004 35284 14056 35290
rect 14004 35226 14056 35232
rect 13728 35216 13780 35222
rect 13728 35158 13780 35164
rect 13636 34604 13688 34610
rect 13636 34546 13688 34552
rect 13648 33862 13676 34546
rect 13728 34468 13780 34474
rect 13728 34410 13780 34416
rect 13636 33856 13688 33862
rect 13636 33798 13688 33804
rect 13648 33522 13676 33798
rect 13636 33516 13688 33522
rect 13636 33458 13688 33464
rect 13544 33448 13596 33454
rect 13544 33390 13596 33396
rect 13452 33108 13504 33114
rect 13452 33050 13504 33056
rect 13452 32972 13504 32978
rect 13452 32914 13504 32920
rect 13464 32230 13492 32914
rect 13556 32910 13584 33390
rect 13740 33386 13768 34410
rect 14188 34400 14240 34406
rect 14188 34342 14240 34348
rect 14200 34066 14228 34342
rect 14568 34202 14596 35430
rect 14556 34196 14608 34202
rect 14556 34138 14608 34144
rect 14188 34060 14240 34066
rect 14188 34002 14240 34008
rect 14200 33658 14228 34002
rect 14188 33652 14240 33658
rect 14188 33594 14240 33600
rect 14648 33448 14700 33454
rect 14648 33390 14700 33396
rect 13728 33380 13780 33386
rect 13728 33322 13780 33328
rect 13544 32904 13596 32910
rect 13544 32846 13596 32852
rect 13452 32224 13504 32230
rect 13452 32166 13504 32172
rect 13268 30796 13320 30802
rect 13268 30738 13320 30744
rect 13360 30796 13412 30802
rect 13360 30738 13412 30744
rect 13280 30326 13308 30738
rect 13268 30320 13320 30326
rect 13268 30262 13320 30268
rect 13176 29776 13228 29782
rect 13176 29718 13228 29724
rect 13372 29510 13400 30738
rect 13176 29504 13228 29510
rect 13176 29446 13228 29452
rect 13360 29504 13412 29510
rect 13360 29446 13412 29452
rect 12992 29300 13044 29306
rect 12992 29242 13044 29248
rect 12900 27872 12952 27878
rect 12900 27814 12952 27820
rect 12808 27600 12860 27606
rect 12808 27542 12860 27548
rect 12716 27532 12768 27538
rect 12716 27474 12768 27480
rect 12728 27334 12756 27474
rect 12808 27396 12860 27402
rect 12808 27338 12860 27344
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12624 27124 12676 27130
rect 12624 27066 12676 27072
rect 12636 26858 12664 27066
rect 12532 26852 12584 26858
rect 12532 26794 12584 26800
rect 12624 26852 12676 26858
rect 12624 26794 12676 26800
rect 12348 26784 12400 26790
rect 12348 26726 12400 26732
rect 12256 26580 12308 26586
rect 12176 26540 12256 26568
rect 12176 26042 12204 26540
rect 12256 26522 12308 26528
rect 12256 26444 12308 26450
rect 12256 26386 12308 26392
rect 12164 26036 12216 26042
rect 12164 25978 12216 25984
rect 12268 25702 12296 26386
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 11900 25498 11928 25638
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 11796 25356 11848 25362
rect 11796 25298 11848 25304
rect 11980 25356 12032 25362
rect 11980 25298 12032 25304
rect 11808 24886 11836 25298
rect 11796 24880 11848 24886
rect 11796 24822 11848 24828
rect 11992 24750 12020 25298
rect 12268 24954 12296 25638
rect 12360 25430 12388 26726
rect 12544 26586 12572 26794
rect 12728 26738 12756 27270
rect 12820 26994 12848 27338
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12636 26710 12756 26738
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12532 26240 12584 26246
rect 12636 26228 12664 26710
rect 12584 26200 12664 26228
rect 12532 26182 12584 26188
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12348 25424 12400 25430
rect 12348 25366 12400 25372
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 12440 24744 12492 24750
rect 12440 24686 12492 24692
rect 12072 24676 12124 24682
rect 12072 24618 12124 24624
rect 12084 23118 12112 24618
rect 12452 24274 12480 24686
rect 12544 24410 12572 25774
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12360 23322 12388 24142
rect 12452 23866 12480 24210
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 11520 22704 11572 22710
rect 11440 22664 11520 22692
rect 11520 22646 11572 22652
rect 11060 22500 11112 22506
rect 11060 22442 11112 22448
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 11808 22098 11836 22374
rect 12636 22098 12664 26200
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12728 25430 12756 26182
rect 13188 25702 13216 29446
rect 13464 27334 13492 32166
rect 13740 30122 13768 33322
rect 14660 33114 14688 33390
rect 14648 33108 14700 33114
rect 14648 33050 14700 33056
rect 14660 32434 14688 33050
rect 14648 32428 14700 32434
rect 14648 32370 14700 32376
rect 14004 32360 14056 32366
rect 14004 32302 14056 32308
rect 13912 31204 13964 31210
rect 13912 31146 13964 31152
rect 13820 30728 13872 30734
rect 13820 30670 13872 30676
rect 13832 30258 13860 30670
rect 13820 30252 13872 30258
rect 13820 30194 13872 30200
rect 13728 30116 13780 30122
rect 13728 30058 13780 30064
rect 13832 29850 13860 30194
rect 13820 29844 13872 29850
rect 13820 29786 13872 29792
rect 13636 29708 13688 29714
rect 13636 29650 13688 29656
rect 13648 28218 13676 29650
rect 13728 29504 13780 29510
rect 13728 29446 13780 29452
rect 13740 28558 13768 29446
rect 13820 29028 13872 29034
rect 13820 28970 13872 28976
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 13636 28212 13688 28218
rect 13636 28154 13688 28160
rect 13832 28082 13860 28970
rect 13924 28694 13952 31146
rect 13912 28688 13964 28694
rect 13912 28630 13964 28636
rect 13924 28218 13952 28630
rect 13912 28212 13964 28218
rect 13912 28154 13964 28160
rect 13820 28076 13872 28082
rect 13820 28018 13872 28024
rect 13728 27532 13780 27538
rect 13728 27474 13780 27480
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 13740 26790 13768 27474
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 13924 26586 13952 28154
rect 13912 26580 13964 26586
rect 13912 26522 13964 26528
rect 14016 26450 14044 32302
rect 14188 32292 14240 32298
rect 14188 32234 14240 32240
rect 14200 32026 14228 32234
rect 14188 32020 14240 32026
rect 14188 31962 14240 31968
rect 14832 32020 14884 32026
rect 14832 31962 14884 31968
rect 14200 31686 14228 31962
rect 14188 31680 14240 31686
rect 14188 31622 14240 31628
rect 14464 31272 14516 31278
rect 14464 31214 14516 31220
rect 14476 30297 14504 31214
rect 14740 30728 14792 30734
rect 14740 30670 14792 30676
rect 14462 30288 14518 30297
rect 14462 30223 14518 30232
rect 14648 30184 14700 30190
rect 14568 30161 14648 30172
rect 14554 30152 14648 30161
rect 14096 30116 14148 30122
rect 14610 30144 14648 30152
rect 14648 30126 14700 30132
rect 14554 30087 14610 30096
rect 14096 30058 14148 30064
rect 14108 27946 14136 30058
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14660 28694 14688 29106
rect 14752 29034 14780 30670
rect 14740 29028 14792 29034
rect 14740 28970 14792 28976
rect 14648 28688 14700 28694
rect 14648 28630 14700 28636
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14384 28218 14412 28494
rect 14372 28212 14424 28218
rect 14372 28154 14424 28160
rect 14096 27940 14148 27946
rect 14096 27882 14148 27888
rect 14108 27130 14136 27882
rect 14188 27328 14240 27334
rect 14188 27270 14240 27276
rect 14096 27124 14148 27130
rect 14096 27066 14148 27072
rect 14108 26858 14136 27066
rect 14200 26994 14228 27270
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14096 26852 14148 26858
rect 14096 26794 14148 26800
rect 13544 26444 13596 26450
rect 13544 26386 13596 26392
rect 14004 26444 14056 26450
rect 14004 26386 14056 26392
rect 13556 26042 13584 26386
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13544 26036 13596 26042
rect 13544 25978 13596 25984
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 12716 25424 12768 25430
rect 12716 25366 12768 25372
rect 13188 23186 13216 25638
rect 13556 25362 13584 25978
rect 13544 25356 13596 25362
rect 13544 25298 13596 25304
rect 13556 24954 13584 25298
rect 13740 25226 13768 26318
rect 14108 26042 14136 26794
rect 14200 26518 14228 26930
rect 14188 26512 14240 26518
rect 14188 26454 14240 26460
rect 14556 26240 14608 26246
rect 14556 26182 14608 26188
rect 14096 26036 14148 26042
rect 14096 25978 14148 25984
rect 14568 25906 14596 26182
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14568 25430 14596 25842
rect 14740 25764 14792 25770
rect 14740 25706 14792 25712
rect 14556 25424 14608 25430
rect 14556 25366 14608 25372
rect 14464 25356 14516 25362
rect 14464 25298 14516 25304
rect 13728 25220 13780 25226
rect 13728 25162 13780 25168
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13648 24342 13676 24754
rect 14476 24750 14504 25298
rect 14556 25152 14608 25158
rect 14556 25094 14608 25100
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14200 24342 14228 24550
rect 13636 24336 13688 24342
rect 13636 24278 13688 24284
rect 14188 24336 14240 24342
rect 14188 24278 14240 24284
rect 13648 23322 13676 24278
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13740 23662 13768 24074
rect 13832 23866 13860 24210
rect 14476 24070 14504 24686
rect 14568 24410 14596 25094
rect 14648 24744 14700 24750
rect 14648 24686 14700 24692
rect 14556 24404 14608 24410
rect 14556 24346 14608 24352
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13636 23316 13688 23322
rect 13636 23258 13688 23264
rect 13176 23180 13228 23186
rect 13176 23122 13228 23128
rect 13452 23180 13504 23186
rect 13452 23122 13504 23128
rect 13636 23180 13688 23186
rect 13740 23168 13768 23598
rect 13820 23588 13872 23594
rect 13820 23530 13872 23536
rect 13688 23140 13768 23168
rect 13636 23122 13688 23128
rect 12900 22704 12952 22710
rect 12900 22646 12952 22652
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 11612 21956 11664 21962
rect 11664 21916 11744 21944
rect 11612 21898 11664 21904
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 10980 21418 11008 21558
rect 10876 21412 10928 21418
rect 10876 21354 10928 21360
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10520 20058 10548 20878
rect 10796 20262 10824 21014
rect 10888 20602 10916 21354
rect 11612 21072 11664 21078
rect 11612 21014 11664 21020
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 11624 20466 11652 21014
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 10324 19984 10376 19990
rect 10324 19926 10376 19932
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9968 18970 9996 19246
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9784 18222 9812 18362
rect 9772 18216 9824 18222
rect 9692 18176 9772 18204
rect 9692 17134 9720 18176
rect 9772 18158 9824 18164
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9416 16794 9444 17002
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9508 15978 9536 16662
rect 9600 16114 9628 16934
rect 9784 16658 9812 17818
rect 9968 17746 9996 18906
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 9968 17338 9996 17682
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 10152 17066 10180 17682
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9784 15706 9812 16594
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9876 15094 9904 15574
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 10060 15026 10088 15438
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 10152 15162 10180 15370
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10060 13814 10088 14962
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10152 13938 10180 14282
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10060 13786 10180 13814
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9232 12986 9260 13330
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9128 12912 9180 12918
rect 9128 12854 9180 12860
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 9140 12374 9168 12854
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 6092 12242 6144 12248
rect 6104 11830 6132 12242
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7024 11898 7052 12174
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7116 11830 7144 12294
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 11898 8616 12242
rect 9232 12238 9260 12650
rect 9876 12374 9904 12854
rect 9968 12646 9996 13670
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9784 11898 9812 12310
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 9876 11762 9904 12310
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 10060 11354 10088 13126
rect 10152 12714 10180 13786
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 10152 12442 10180 12650
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10244 11642 10272 19722
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10520 19310 10548 19654
rect 10796 19334 10824 20198
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10508 19304 10560 19310
rect 10796 19306 10916 19334
rect 10508 19246 10560 19252
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10428 18154 10456 18702
rect 10520 18222 10548 19246
rect 10692 19236 10744 19242
rect 10692 19178 10744 19184
rect 10704 18766 10732 19178
rect 10888 18970 10916 19306
rect 11072 19174 11100 19858
rect 11624 19310 11652 20402
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10336 16726 10364 18022
rect 10428 17882 10456 18090
rect 10888 18086 10916 18906
rect 11072 18834 11100 19110
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11256 18426 11284 18566
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11256 18222 11284 18362
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10796 16794 10824 17070
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10336 15978 10364 16662
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 14550 10548 15846
rect 10888 15706 10916 16934
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10888 15026 10916 15642
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 10600 14884 10652 14890
rect 10600 14826 10652 14832
rect 10612 14550 10640 14826
rect 11164 14550 11192 14962
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 10520 13530 10548 14486
rect 10612 14074 10640 14486
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 11164 13326 11192 14486
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11256 12918 11284 13398
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11440 12986 11468 13262
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 11256 12646 11284 12854
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11532 11898 11560 15370
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12850 11652 13262
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11624 12374 11652 12786
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11624 11830 11652 12038
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 10152 11614 10272 11642
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 1490 11248 1546 11257
rect 1490 11183 1546 11192
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 9876 10810 9904 11154
rect 10152 11082 10180 11614
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10244 11218 10272 11494
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 10152 10130 10180 11018
rect 10244 10538 10272 11154
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 10336 10674 10364 11086
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 11348 10606 11376 11086
rect 11440 10810 11468 11222
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10244 10130 10272 10474
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 10152 9654 10180 10066
rect 10244 9722 10272 10066
rect 10520 9722 10548 10474
rect 11440 10266 11468 10746
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11716 10130 11744 21916
rect 11808 21690 11836 22034
rect 12636 21690 12664 22034
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12072 21412 12124 21418
rect 12072 21354 12124 21360
rect 12084 20874 12112 21354
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12176 21146 12204 21286
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12268 20942 12296 21286
rect 12256 20936 12308 20942
rect 12256 20878 12308 20884
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 12084 20466 12112 20810
rect 12268 20602 12296 20878
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 11900 19446 11928 19858
rect 12360 19514 12388 19858
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12348 19508 12400 19514
rect 12348 19450 12400 19456
rect 11888 19440 11940 19446
rect 11888 19382 11940 19388
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11808 16658 11836 17818
rect 11900 17134 11928 19382
rect 12256 19236 12308 19242
rect 12256 19178 12308 19184
rect 12268 18970 12296 19178
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12268 18290 12296 18906
rect 12452 18698 12480 19654
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12636 18222 12664 21626
rect 12912 21010 12940 22646
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 13372 22166 13400 22510
rect 13464 22506 13492 23122
rect 13452 22500 13504 22506
rect 13452 22442 13504 22448
rect 13360 22160 13412 22166
rect 13360 22102 13412 22108
rect 13358 21992 13414 22001
rect 13084 21956 13136 21962
rect 13358 21927 13414 21936
rect 13084 21898 13136 21904
rect 13096 21350 13124 21898
rect 13372 21894 13400 21927
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 13096 21010 13124 21286
rect 12900 21004 12952 21010
rect 13084 21004 13136 21010
rect 12900 20946 12952 20952
rect 13004 20964 13084 20992
rect 12912 20602 12940 20946
rect 12900 20596 12952 20602
rect 12820 20556 12900 20584
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12728 19378 12756 20198
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 11992 17270 12020 17682
rect 12176 17338 12204 17682
rect 12728 17610 12756 19314
rect 12820 17814 12848 20556
rect 12900 20538 12952 20544
rect 13004 20262 13032 20964
rect 13084 20946 13136 20952
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13372 20398 13400 20742
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 13004 19922 13032 20198
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 13280 19496 13308 19994
rect 13372 19990 13400 20334
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13360 19508 13412 19514
rect 13280 19468 13360 19496
rect 13280 18902 13308 19468
rect 13360 19450 13412 19456
rect 13268 18896 13320 18902
rect 13268 18838 13320 18844
rect 13464 18850 13492 22442
rect 13648 21962 13676 23122
rect 13728 22636 13780 22642
rect 13728 22578 13780 22584
rect 13740 22438 13768 22578
rect 13728 22432 13780 22438
rect 13728 22374 13780 22380
rect 13636 21956 13688 21962
rect 13636 21898 13688 21904
rect 13740 21706 13768 22374
rect 13648 21678 13768 21706
rect 13648 21486 13676 21678
rect 13636 21480 13688 21486
rect 13636 21422 13688 21428
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13556 19922 13584 20878
rect 13648 20602 13676 21422
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13648 20330 13676 20538
rect 13636 20324 13688 20330
rect 13636 20266 13688 20272
rect 13648 20058 13676 20266
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13556 18970 13584 19858
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13464 18822 13584 18850
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13464 18426 13492 18702
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12808 17808 12860 17814
rect 12808 17750 12860 17756
rect 12912 17746 12940 18158
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11808 15706 11836 16594
rect 12176 15978 12204 16730
rect 12544 16114 12572 16934
rect 13004 16794 13032 17070
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 12268 15570 12296 15846
rect 12544 15706 12572 16050
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12084 14618 12112 15302
rect 12268 15162 12296 15506
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12084 14006 12112 14554
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12268 14074 12296 14486
rect 12452 14414 12480 15030
rect 12544 15026 12572 15302
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 12452 13326 12480 14350
rect 12544 14074 12572 14962
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12728 13870 12756 16390
rect 13188 15570 13216 18090
rect 13556 17746 13584 18822
rect 13832 18426 13860 23530
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 13924 22234 13952 23054
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 13912 22228 13964 22234
rect 13912 22170 13964 22176
rect 13924 21554 13952 22170
rect 14292 22098 14320 22374
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 14004 21616 14056 21622
rect 14004 21558 14056 21564
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 14016 19514 14044 21558
rect 14292 21146 14320 22034
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14016 19174 14044 19450
rect 14370 19408 14426 19417
rect 14370 19343 14426 19352
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14016 18902 14044 19110
rect 14108 18970 14136 19178
rect 14384 18970 14412 19343
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 14108 18698 14136 18906
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13832 18222 13860 18362
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 14384 18086 14412 18770
rect 14476 18426 14504 24006
rect 14568 23594 14596 24346
rect 14660 24138 14688 24686
rect 14648 24132 14700 24138
rect 14648 24074 14700 24080
rect 14752 23866 14780 25706
rect 14844 25362 14872 31962
rect 14924 28620 14976 28626
rect 14924 28562 14976 28568
rect 14936 27878 14964 28562
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 14936 26042 14964 27814
rect 14924 26036 14976 26042
rect 14924 25978 14976 25984
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 14924 24744 14976 24750
rect 14924 24686 14976 24692
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14752 23594 14780 23802
rect 14936 23730 14964 24686
rect 14924 23724 14976 23730
rect 14924 23666 14976 23672
rect 14556 23588 14608 23594
rect 14556 23530 14608 23536
rect 14740 23588 14792 23594
rect 14740 23530 14792 23536
rect 14752 22642 14780 23530
rect 14936 23322 14964 23666
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14832 21344 14884 21350
rect 14832 21286 14884 21292
rect 14844 21010 14872 21286
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 13556 17338 13584 17682
rect 14200 17338 14228 17682
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13832 16250 13860 16594
rect 14016 16590 14044 17070
rect 14200 16794 14228 17274
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 14292 16114 14320 17614
rect 14384 17105 14412 18022
rect 14660 17882 14688 18158
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14370 17096 14426 17105
rect 14370 17031 14426 17040
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13556 15638 13584 15914
rect 14292 15706 14320 16050
rect 14568 15978 14596 16934
rect 14660 16658 14688 17478
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13188 15162 13216 15506
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13372 14550 13400 14894
rect 13556 14822 13584 15574
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12728 13530 12756 13806
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 13004 13326 13032 13738
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 11900 12986 11928 13262
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 13004 12850 13032 13262
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13188 12374 13216 12650
rect 12808 12368 12860 12374
rect 12808 12310 12860 12316
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12176 11286 12204 12174
rect 12820 11898 12848 12310
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 13188 11558 13216 12310
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 12176 10810 12204 11222
rect 12268 11082 12296 11494
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10520 9450 10548 9658
rect 10704 9586 10732 9998
rect 11716 9994 11744 10066
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11716 9722 11744 9930
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10704 9178 10732 9522
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 11256 9178 11284 9386
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 11256 8634 11284 9114
rect 11532 8634 11560 9318
rect 11704 9036 11756 9042
rect 11808 9024 11836 10202
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12176 9722 12204 10066
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 9178 12480 9318
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 11756 8996 11836 9024
rect 11704 8978 11756 8984
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11808 8566 11836 8996
rect 12452 8566 12480 9114
rect 13096 8974 13124 11018
rect 13188 10674 13216 11494
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13280 10606 13308 12038
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 11286 13400 11494
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13372 10810 13400 11222
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13280 10266 13308 10542
rect 13556 10538 13584 14758
rect 13832 14550 13860 14826
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13832 14414 13860 14486
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13740 14074 13768 14350
rect 13832 14074 13860 14350
rect 14016 14074 14044 15302
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14844 14618 14872 14826
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 13648 11286 13676 12650
rect 13832 11354 13860 12650
rect 14016 11626 14044 13194
rect 14200 12646 14228 13330
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14108 11762 14136 12038
rect 14200 11898 14228 12582
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14292 11762 14320 12174
rect 14384 11898 14412 13126
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14096 11756 14148 11762
rect 14280 11756 14332 11762
rect 14096 11698 14148 11704
rect 14200 11716 14280 11744
rect 14004 11620 14056 11626
rect 14004 11562 14056 11568
rect 14016 11354 14044 11562
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13648 10266 13676 11222
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13556 9110 13584 9386
rect 13832 9382 13860 10134
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13924 9722 13952 9930
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14200 9654 14228 11716
rect 14280 11698 14332 11704
rect 14844 10577 14872 11766
rect 15028 10810 15056 39238
rect 16132 38758 16160 39442
rect 17328 39370 17356 39743
rect 17316 39364 17368 39370
rect 17316 39306 17368 39312
rect 15844 38752 15896 38758
rect 15844 38694 15896 38700
rect 16120 38752 16172 38758
rect 16120 38694 16172 38700
rect 16304 38752 16356 38758
rect 16304 38694 16356 38700
rect 16856 38752 16908 38758
rect 16856 38694 16908 38700
rect 15476 38480 15528 38486
rect 15476 38422 15528 38428
rect 15384 38344 15436 38350
rect 15384 38286 15436 38292
rect 15396 37466 15424 38286
rect 15488 38010 15516 38422
rect 15476 38004 15528 38010
rect 15476 37946 15528 37952
rect 15856 37777 15884 38694
rect 16132 38350 16160 38694
rect 16120 38344 16172 38350
rect 16120 38286 16172 38292
rect 15842 37768 15898 37777
rect 15842 37703 15898 37712
rect 15384 37460 15436 37466
rect 15384 37402 15436 37408
rect 16316 37330 16344 38694
rect 16868 38282 16896 38694
rect 17774 38448 17830 38457
rect 17774 38383 17776 38392
rect 17828 38383 17830 38392
rect 17776 38354 17828 38360
rect 16856 38276 16908 38282
rect 16856 38218 16908 38224
rect 16868 37806 16896 38218
rect 17788 38010 17816 38354
rect 17776 38004 17828 38010
rect 17776 37946 17828 37952
rect 16856 37800 16908 37806
rect 16856 37742 16908 37748
rect 18328 37664 18380 37670
rect 18328 37606 18380 37612
rect 16304 37324 16356 37330
rect 16304 37266 16356 37272
rect 17868 37324 17920 37330
rect 17868 37266 17920 37272
rect 15752 37256 15804 37262
rect 15752 37198 15804 37204
rect 15764 36650 15792 37198
rect 16316 36922 16344 37266
rect 17880 36922 17908 37266
rect 16304 36916 16356 36922
rect 16304 36858 16356 36864
rect 17868 36916 17920 36922
rect 17868 36858 17920 36864
rect 18340 36786 18368 37606
rect 18420 37392 18472 37398
rect 18420 37334 18472 37340
rect 18432 37126 18460 37334
rect 18524 37330 18552 42298
rect 21364 42016 21416 42022
rect 21364 41958 21416 41964
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 21376 41750 21404 41958
rect 21364 41744 21416 41750
rect 21364 41686 21416 41692
rect 19248 41200 19300 41206
rect 19248 41142 19300 41148
rect 19064 41064 19116 41070
rect 19064 41006 19116 41012
rect 19076 39409 19104 41006
rect 19062 39400 19118 39409
rect 19062 39335 19118 39344
rect 19076 38418 19104 39335
rect 19064 38412 19116 38418
rect 19064 38354 19116 38360
rect 19076 38010 19104 38354
rect 19064 38004 19116 38010
rect 19064 37946 19116 37952
rect 19260 37806 19288 41142
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 21180 40588 21232 40594
rect 21180 40530 21232 40536
rect 21192 39846 21220 40530
rect 21180 39840 21232 39846
rect 21180 39782 21232 39788
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 21192 38962 21220 39782
rect 21456 39432 21508 39438
rect 21456 39374 21508 39380
rect 21180 38956 21232 38962
rect 21180 38898 21232 38904
rect 21192 38865 21220 38898
rect 21178 38856 21234 38865
rect 21178 38791 21234 38800
rect 21468 38758 21496 39374
rect 20996 38752 21048 38758
rect 20996 38694 21048 38700
rect 21456 38752 21508 38758
rect 21456 38694 21508 38700
rect 21548 38752 21600 38758
rect 21548 38694 21600 38700
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 21008 38486 21036 38694
rect 20996 38480 21048 38486
rect 20996 38422 21048 38428
rect 21088 38480 21140 38486
rect 21088 38422 21140 38428
rect 19340 38208 19392 38214
rect 19340 38150 19392 38156
rect 19616 38208 19668 38214
rect 19616 38150 19668 38156
rect 19352 37874 19380 38150
rect 19340 37868 19392 37874
rect 19340 37810 19392 37816
rect 19248 37800 19300 37806
rect 19248 37742 19300 37748
rect 19352 37466 19380 37810
rect 19628 37738 19656 38150
rect 21008 38010 21036 38422
rect 21100 38214 21128 38422
rect 21088 38208 21140 38214
rect 21088 38150 21140 38156
rect 20996 38004 21048 38010
rect 20996 37946 21048 37952
rect 21100 37874 21128 38150
rect 21088 37868 21140 37874
rect 21088 37810 21140 37816
rect 19616 37732 19668 37738
rect 19616 37674 19668 37680
rect 20168 37732 20220 37738
rect 20168 37674 20220 37680
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19340 37460 19392 37466
rect 19340 37402 19392 37408
rect 18512 37324 18564 37330
rect 18512 37266 18564 37272
rect 20180 37262 20208 37674
rect 18972 37256 19024 37262
rect 18972 37198 19024 37204
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 18420 37120 18472 37126
rect 18420 37062 18472 37068
rect 18328 36780 18380 36786
rect 18328 36722 18380 36728
rect 18432 36650 18460 37062
rect 15568 36644 15620 36650
rect 15568 36586 15620 36592
rect 15752 36644 15804 36650
rect 15752 36586 15804 36592
rect 18420 36644 18472 36650
rect 18420 36586 18472 36592
rect 15580 36038 15608 36586
rect 18432 36378 18460 36586
rect 18984 36378 19012 37198
rect 19064 36644 19116 36650
rect 19064 36586 19116 36592
rect 18420 36372 18472 36378
rect 18420 36314 18472 36320
rect 18972 36372 19024 36378
rect 18972 36314 19024 36320
rect 17684 36304 17736 36310
rect 17684 36246 17736 36252
rect 16212 36236 16264 36242
rect 16212 36178 16264 36184
rect 15660 36168 15712 36174
rect 15660 36110 15712 36116
rect 15568 36032 15620 36038
rect 15568 35974 15620 35980
rect 15292 35760 15344 35766
rect 15292 35702 15344 35708
rect 15304 35562 15332 35702
rect 15292 35556 15344 35562
rect 15292 35498 15344 35504
rect 15304 34746 15332 35498
rect 15672 35222 15700 36110
rect 16028 36032 16080 36038
rect 16028 35974 16080 35980
rect 15660 35216 15712 35222
rect 15660 35158 15712 35164
rect 15292 34740 15344 34746
rect 15292 34682 15344 34688
rect 15304 34474 15332 34682
rect 15568 34672 15620 34678
rect 15672 34660 15700 35158
rect 16040 35018 16068 35974
rect 16224 35834 16252 36178
rect 17408 36168 17460 36174
rect 17408 36110 17460 36116
rect 16212 35828 16264 35834
rect 16212 35770 16264 35776
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 17236 35193 17264 35430
rect 17222 35184 17278 35193
rect 17222 35119 17224 35128
rect 17276 35119 17278 35128
rect 17224 35090 17276 35096
rect 16580 35080 16632 35086
rect 16580 35022 16632 35028
rect 16028 35012 16080 35018
rect 16028 34954 16080 34960
rect 15620 34632 15700 34660
rect 15568 34614 15620 34620
rect 16040 34610 16068 34954
rect 16212 34944 16264 34950
rect 16212 34886 16264 34892
rect 16028 34604 16080 34610
rect 16028 34546 16080 34552
rect 15292 34468 15344 34474
rect 15292 34410 15344 34416
rect 15304 34134 15332 34410
rect 15292 34128 15344 34134
rect 15292 34070 15344 34076
rect 16224 34066 16252 34886
rect 16592 34746 16620 35022
rect 17236 34746 17264 35090
rect 17420 34950 17448 36110
rect 17696 35494 17724 36246
rect 19076 36106 19104 36586
rect 19248 36236 19300 36242
rect 19248 36178 19300 36184
rect 19064 36100 19116 36106
rect 19064 36042 19116 36048
rect 17684 35488 17736 35494
rect 17684 35430 17736 35436
rect 17696 35222 17724 35430
rect 17684 35216 17736 35222
rect 17684 35158 17736 35164
rect 18420 35080 18472 35086
rect 18420 35022 18472 35028
rect 17408 34944 17460 34950
rect 17408 34886 17460 34892
rect 16580 34740 16632 34746
rect 16580 34682 16632 34688
rect 17224 34740 17276 34746
rect 17224 34682 17276 34688
rect 16212 34060 16264 34066
rect 16212 34002 16264 34008
rect 16224 33658 16252 34002
rect 16592 33658 16620 34682
rect 17420 34202 17448 34886
rect 18432 34610 18460 35022
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 18420 34604 18472 34610
rect 18420 34546 18472 34552
rect 18236 34536 18288 34542
rect 18236 34478 18288 34484
rect 17408 34196 17460 34202
rect 17408 34138 17460 34144
rect 17132 34060 17184 34066
rect 17132 34002 17184 34008
rect 17684 34060 17736 34066
rect 17684 34002 17736 34008
rect 17144 33658 17172 34002
rect 16212 33652 16264 33658
rect 16212 33594 16264 33600
rect 16580 33652 16632 33658
rect 16580 33594 16632 33600
rect 17132 33652 17184 33658
rect 17132 33594 17184 33600
rect 15476 33380 15528 33386
rect 15476 33322 15528 33328
rect 15488 33046 15516 33322
rect 17144 33134 17172 33594
rect 17696 33386 17724 34002
rect 17684 33380 17736 33386
rect 17684 33322 17736 33328
rect 17144 33106 17264 33134
rect 15476 33040 15528 33046
rect 17236 33017 17264 33106
rect 17408 33040 17460 33046
rect 15476 32982 15528 32988
rect 17222 33008 17278 33017
rect 15292 32904 15344 32910
rect 15292 32846 15344 32852
rect 15304 32434 15332 32846
rect 15488 32570 15516 32982
rect 17408 32982 17460 32988
rect 17222 32943 17278 32952
rect 17316 32768 17368 32774
rect 17316 32710 17368 32716
rect 15476 32564 15528 32570
rect 15476 32506 15528 32512
rect 15292 32428 15344 32434
rect 15292 32370 15344 32376
rect 15660 32360 15712 32366
rect 15660 32302 15712 32308
rect 15672 32026 15700 32302
rect 17328 32026 17356 32710
rect 17420 32570 17448 32982
rect 17408 32564 17460 32570
rect 17408 32506 17460 32512
rect 17868 32292 17920 32298
rect 17868 32234 17920 32240
rect 15660 32020 15712 32026
rect 15660 31962 15712 31968
rect 17316 32020 17368 32026
rect 17316 31962 17368 31968
rect 17880 31890 17908 32234
rect 16488 31884 16540 31890
rect 16488 31826 16540 31832
rect 17316 31884 17368 31890
rect 17316 31826 17368 31832
rect 17868 31884 17920 31890
rect 17868 31826 17920 31832
rect 15474 31784 15530 31793
rect 15292 31748 15344 31754
rect 16500 31754 16528 31826
rect 15474 31719 15530 31728
rect 16488 31748 16540 31754
rect 15292 31690 15344 31696
rect 15304 31278 15332 31690
rect 15292 31272 15344 31278
rect 15292 31214 15344 31220
rect 15488 30802 15516 31719
rect 16488 31690 16540 31696
rect 16500 31482 16528 31690
rect 16488 31476 16540 31482
rect 16488 31418 16540 31424
rect 17328 31210 17356 31826
rect 17880 31686 17908 31826
rect 17868 31680 17920 31686
rect 17868 31622 17920 31628
rect 17316 31204 17368 31210
rect 17316 31146 17368 31152
rect 17776 31204 17828 31210
rect 17776 31146 17828 31152
rect 15476 30796 15528 30802
rect 15476 30738 15528 30744
rect 17132 30796 17184 30802
rect 17132 30738 17184 30744
rect 15488 30394 15516 30738
rect 16948 30728 17000 30734
rect 16948 30670 17000 30676
rect 15476 30388 15528 30394
rect 15476 30330 15528 30336
rect 15660 30116 15712 30122
rect 15660 30058 15712 30064
rect 15476 29776 15528 29782
rect 15476 29718 15528 29724
rect 15384 29640 15436 29646
rect 15384 29582 15436 29588
rect 15396 29170 15424 29582
rect 15488 29306 15516 29718
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 15384 29164 15436 29170
rect 15384 29106 15436 29112
rect 15488 29073 15516 29242
rect 15474 29064 15530 29073
rect 15474 28999 15530 29008
rect 15476 28960 15528 28966
rect 15476 28902 15528 28908
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15304 27674 15332 28358
rect 15292 27668 15344 27674
rect 15292 27610 15344 27616
rect 15304 27130 15332 27610
rect 15488 27606 15516 28902
rect 15672 28218 15700 30058
rect 16960 29782 16988 30670
rect 17144 30054 17172 30738
rect 17788 30666 17816 31146
rect 17880 31142 17908 31622
rect 17868 31136 17920 31142
rect 17868 31078 17920 31084
rect 17776 30660 17828 30666
rect 17776 30602 17828 30608
rect 17684 30184 17736 30190
rect 17684 30126 17736 30132
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 16948 29776 17000 29782
rect 16948 29718 17000 29724
rect 16120 29640 16172 29646
rect 16120 29582 16172 29588
rect 16946 29608 17002 29617
rect 16132 28762 16160 29582
rect 16946 29543 17002 29552
rect 16488 29028 16540 29034
rect 16488 28970 16540 28976
rect 16120 28756 16172 28762
rect 16120 28698 16172 28704
rect 16028 28416 16080 28422
rect 16028 28358 16080 28364
rect 15660 28212 15712 28218
rect 15660 28154 15712 28160
rect 15672 27946 15700 28154
rect 15660 27940 15712 27946
rect 15660 27882 15712 27888
rect 16040 27878 16068 28358
rect 16132 28082 16160 28698
rect 16500 28694 16528 28970
rect 16578 28928 16634 28937
rect 16578 28863 16634 28872
rect 16488 28688 16540 28694
rect 16488 28630 16540 28636
rect 16592 28558 16620 28863
rect 16764 28688 16816 28694
rect 16764 28630 16816 28636
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 16028 27872 16080 27878
rect 16028 27814 16080 27820
rect 15476 27600 15528 27606
rect 15476 27542 15528 27548
rect 15292 27124 15344 27130
rect 15292 27066 15344 27072
rect 15488 26994 15516 27542
rect 16040 27470 16068 27814
rect 16592 27674 16620 28494
rect 16776 28218 16804 28630
rect 16764 28212 16816 28218
rect 16764 28154 16816 28160
rect 16960 28150 16988 29543
rect 17040 28960 17092 28966
rect 17040 28902 17092 28908
rect 16948 28144 17000 28150
rect 16948 28086 17000 28092
rect 17052 28082 17080 28902
rect 17144 28218 17172 29990
rect 17408 29776 17460 29782
rect 17460 29736 17540 29764
rect 17408 29718 17460 29724
rect 17512 29034 17540 29736
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17224 29028 17276 29034
rect 17224 28970 17276 28976
rect 17500 29028 17552 29034
rect 17500 28970 17552 28976
rect 17236 28558 17264 28970
rect 17512 28694 17540 28970
rect 17500 28688 17552 28694
rect 17500 28630 17552 28636
rect 17224 28552 17276 28558
rect 17224 28494 17276 28500
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 16580 27668 16632 27674
rect 16580 27610 16632 27616
rect 17052 27606 17080 28018
rect 17040 27600 17092 27606
rect 17040 27542 17092 27548
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 15476 26512 15528 26518
rect 15476 26454 15528 26460
rect 15488 26042 15516 26454
rect 15844 26376 15896 26382
rect 15948 26364 15976 26726
rect 16040 26518 16068 27406
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16868 26586 16896 27338
rect 17052 27130 17080 27542
rect 17040 27124 17092 27130
rect 17040 27066 17092 27072
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 16028 26512 16080 26518
rect 16028 26454 16080 26460
rect 17236 26382 17264 28494
rect 17604 27606 17632 29582
rect 17696 28558 17724 30126
rect 17684 28552 17736 28558
rect 17684 28494 17736 28500
rect 17592 27600 17644 27606
rect 17592 27542 17644 27548
rect 17604 26994 17632 27542
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17316 26784 17368 26790
rect 17316 26726 17368 26732
rect 15896 26336 15976 26364
rect 15844 26318 15896 26324
rect 15948 26042 15976 26336
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 17236 26042 17264 26318
rect 15476 26036 15528 26042
rect 15476 25978 15528 25984
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 17224 26036 17276 26042
rect 17224 25978 17276 25984
rect 17328 25838 17356 26726
rect 17500 26512 17552 26518
rect 17500 26454 17552 26460
rect 17512 26042 17540 26454
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17316 25832 17368 25838
rect 17316 25774 17368 25780
rect 17132 25696 17184 25702
rect 17132 25638 17184 25644
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 15304 24614 15332 25298
rect 16500 24682 16528 25298
rect 17144 25294 17172 25638
rect 17696 25498 17724 28494
rect 17788 27928 17816 30602
rect 17880 30258 17908 31078
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17880 29306 17908 30194
rect 18248 29578 18276 34478
rect 18432 34202 18460 34546
rect 18524 34542 18552 34886
rect 18512 34536 18564 34542
rect 18512 34478 18564 34484
rect 18420 34196 18472 34202
rect 18420 34138 18472 34144
rect 18524 33386 18552 34478
rect 18604 33448 18656 33454
rect 18604 33390 18656 33396
rect 18512 33380 18564 33386
rect 18512 33322 18564 33328
rect 18524 32366 18552 33322
rect 18616 33114 18644 33390
rect 18696 33380 18748 33386
rect 18696 33322 18748 33328
rect 18604 33108 18656 33114
rect 18604 33050 18656 33056
rect 18616 32434 18644 33050
rect 18708 33046 18736 33322
rect 19076 33114 19104 36042
rect 19260 35834 19288 36178
rect 19248 35828 19300 35834
rect 19248 35770 19300 35776
rect 19156 35216 19208 35222
rect 19156 35158 19208 35164
rect 19168 34678 19196 35158
rect 19156 34672 19208 34678
rect 19156 34614 19208 34620
rect 19168 33386 19196 34614
rect 19352 33998 19380 37198
rect 19892 36644 19944 36650
rect 19892 36586 19944 36592
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19904 36310 19932 36586
rect 20260 36372 20312 36378
rect 20260 36314 20312 36320
rect 19892 36304 19944 36310
rect 19892 36246 19944 36252
rect 19892 35556 19944 35562
rect 19892 35498 19944 35504
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19904 35222 19932 35498
rect 19892 35216 19944 35222
rect 19892 35158 19944 35164
rect 20272 34746 20300 36314
rect 21100 36310 21128 37810
rect 21468 36922 21496 38694
rect 21560 37398 21588 38694
rect 21548 37392 21600 37398
rect 21548 37334 21600 37340
rect 21652 37244 21680 43046
rect 22100 42560 22152 42566
rect 22100 42502 22152 42508
rect 22112 42226 22140 42502
rect 22100 42220 22152 42226
rect 22100 42162 22152 42168
rect 22112 41818 22140 42162
rect 22100 41812 22152 41818
rect 22100 41754 22152 41760
rect 22100 41676 22152 41682
rect 22100 41618 22152 41624
rect 22112 40934 22140 41618
rect 22100 40928 22152 40934
rect 22100 40870 22152 40876
rect 22112 38894 22140 40870
rect 22284 39840 22336 39846
rect 22284 39782 22336 39788
rect 22192 39636 22244 39642
rect 22192 39578 22244 39584
rect 22204 39098 22232 39578
rect 22192 39092 22244 39098
rect 22192 39034 22244 39040
rect 22204 39001 22232 39034
rect 22190 38992 22246 39001
rect 22190 38927 22246 38936
rect 22100 38888 22152 38894
rect 22100 38830 22152 38836
rect 22296 38486 22324 39782
rect 22284 38480 22336 38486
rect 22284 38422 22336 38428
rect 21916 38344 21968 38350
rect 21916 38286 21968 38292
rect 21732 38208 21784 38214
rect 21732 38150 21784 38156
rect 21744 37874 21772 38150
rect 21928 37874 21956 38286
rect 21732 37868 21784 37874
rect 21732 37810 21784 37816
rect 21916 37868 21968 37874
rect 21916 37810 21968 37816
rect 21744 37466 21772 37810
rect 21824 37664 21876 37670
rect 21824 37606 21876 37612
rect 21732 37460 21784 37466
rect 21732 37402 21784 37408
rect 21836 37398 21864 37606
rect 21824 37392 21876 37398
rect 21824 37334 21876 37340
rect 21560 37216 21680 37244
rect 21456 36916 21508 36922
rect 21456 36858 21508 36864
rect 21364 36576 21416 36582
rect 21364 36518 21416 36524
rect 21088 36304 21140 36310
rect 21088 36246 21140 36252
rect 20720 36168 20772 36174
rect 20720 36110 20772 36116
rect 20732 35290 20760 36110
rect 21100 35834 21128 36246
rect 21088 35828 21140 35834
rect 21088 35770 21140 35776
rect 21376 35562 21404 36518
rect 21364 35556 21416 35562
rect 21364 35498 21416 35504
rect 21376 35290 21404 35498
rect 20720 35284 20772 35290
rect 20720 35226 20772 35232
rect 21272 35284 21324 35290
rect 21272 35226 21324 35232
rect 21364 35284 21416 35290
rect 21364 35226 21416 35232
rect 20536 35080 20588 35086
rect 20536 35022 20588 35028
rect 20260 34740 20312 34746
rect 20260 34682 20312 34688
rect 20272 34542 20300 34682
rect 20260 34536 20312 34542
rect 20260 34478 20312 34484
rect 20548 34474 20576 35022
rect 21284 34746 21312 35226
rect 21272 34740 21324 34746
rect 21272 34682 21324 34688
rect 21178 34640 21234 34649
rect 21178 34575 21234 34584
rect 20076 34468 20128 34474
rect 20076 34410 20128 34416
rect 20536 34468 20588 34474
rect 20536 34410 20588 34416
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19432 34128 19484 34134
rect 19432 34070 19484 34076
rect 19340 33992 19392 33998
rect 19340 33934 19392 33940
rect 19352 33590 19380 33934
rect 19444 33658 19472 34070
rect 19892 33924 19944 33930
rect 19892 33866 19944 33872
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 19340 33584 19392 33590
rect 19340 33526 19392 33532
rect 19156 33380 19208 33386
rect 19156 33322 19208 33328
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19064 33108 19116 33114
rect 19064 33050 19116 33056
rect 18696 33040 18748 33046
rect 18696 32982 18748 32988
rect 19340 33040 19392 33046
rect 19340 32982 19392 32988
rect 18604 32428 18656 32434
rect 18604 32370 18656 32376
rect 18512 32360 18564 32366
rect 18512 32302 18564 32308
rect 18708 31414 18736 32982
rect 19352 32842 19380 32982
rect 19904 32910 19932 33866
rect 19892 32904 19944 32910
rect 19892 32846 19944 32852
rect 19340 32836 19392 32842
rect 19340 32778 19392 32784
rect 19352 32570 19380 32778
rect 19340 32564 19392 32570
rect 19340 32506 19392 32512
rect 19892 32292 19944 32298
rect 19892 32234 19944 32240
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19432 31952 19484 31958
rect 19432 31894 19484 31900
rect 19340 31816 19392 31822
rect 19340 31758 19392 31764
rect 18972 31680 19024 31686
rect 18972 31622 19024 31628
rect 18696 31408 18748 31414
rect 18696 31350 18748 31356
rect 18984 31278 19012 31622
rect 19352 31414 19380 31758
rect 19444 31482 19472 31894
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 19340 31408 19392 31414
rect 19340 31350 19392 31356
rect 18972 31272 19024 31278
rect 18972 31214 19024 31220
rect 18880 30728 18932 30734
rect 18880 30670 18932 30676
rect 18328 30592 18380 30598
rect 18328 30534 18380 30540
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 18340 30190 18368 30534
rect 18800 30190 18828 30534
rect 18892 30258 18920 30670
rect 18880 30252 18932 30258
rect 18880 30194 18932 30200
rect 18328 30184 18380 30190
rect 18328 30126 18380 30132
rect 18788 30184 18840 30190
rect 18788 30126 18840 30132
rect 18800 29714 18828 30126
rect 18880 29844 18932 29850
rect 18880 29786 18932 29792
rect 18696 29708 18748 29714
rect 18696 29650 18748 29656
rect 18788 29708 18840 29714
rect 18788 29650 18840 29656
rect 18236 29572 18288 29578
rect 18236 29514 18288 29520
rect 17868 29300 17920 29306
rect 17868 29242 17920 29248
rect 18708 28966 18736 29650
rect 18892 29102 18920 29786
rect 18984 29646 19012 31214
rect 19248 31204 19300 31210
rect 19248 31146 19300 31152
rect 19260 30938 19288 31146
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19260 30394 19288 30874
rect 19904 30802 19932 32234
rect 19892 30796 19944 30802
rect 19892 30738 19944 30744
rect 19248 30388 19300 30394
rect 19248 30330 19300 30336
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 18880 29096 18932 29102
rect 18880 29038 18932 29044
rect 18696 28960 18748 28966
rect 18696 28902 18748 28908
rect 19432 28960 19484 28966
rect 19432 28902 19484 28908
rect 18144 28620 18196 28626
rect 18144 28562 18196 28568
rect 18972 28620 19024 28626
rect 18972 28562 19024 28568
rect 19340 28620 19392 28626
rect 19340 28562 19392 28568
rect 18156 28218 18184 28562
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 18144 28212 18196 28218
rect 18144 28154 18196 28160
rect 18248 28014 18276 28358
rect 18984 28121 19012 28562
rect 18970 28112 19026 28121
rect 18970 28047 19026 28056
rect 19064 28076 19116 28082
rect 18236 28008 18288 28014
rect 18236 27950 18288 27956
rect 17868 27940 17920 27946
rect 17788 27900 17868 27928
rect 17868 27882 17920 27888
rect 17684 25492 17736 25498
rect 17684 25434 17736 25440
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17132 25288 17184 25294
rect 17132 25230 17184 25236
rect 17512 24886 17540 25298
rect 17880 24954 17908 27882
rect 18248 27674 18276 27950
rect 18984 27878 19012 28047
rect 19064 28018 19116 28024
rect 18972 27872 19024 27878
rect 18972 27814 19024 27820
rect 18236 27668 18288 27674
rect 18236 27610 18288 27616
rect 17960 27328 18012 27334
rect 17960 27270 18012 27276
rect 17972 26926 18000 27270
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 18420 26988 18472 26994
rect 18420 26930 18472 26936
rect 17960 26920 18012 26926
rect 17960 26862 18012 26868
rect 18156 26586 18184 26930
rect 18236 26852 18288 26858
rect 18236 26794 18288 26800
rect 18144 26580 18196 26586
rect 18144 26522 18196 26528
rect 18248 26042 18276 26794
rect 18432 26382 18460 26930
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18236 26036 18288 26042
rect 18236 25978 18288 25984
rect 18052 25832 18104 25838
rect 18052 25774 18104 25780
rect 18064 25498 18092 25774
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17132 24744 17184 24750
rect 17132 24686 17184 24692
rect 17776 24744 17828 24750
rect 17776 24686 17828 24692
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 15292 24608 15344 24614
rect 15292 24550 15344 24556
rect 17144 24342 17172 24686
rect 17684 24676 17736 24682
rect 17684 24618 17736 24624
rect 17408 24608 17460 24614
rect 17408 24550 17460 24556
rect 15660 24336 15712 24342
rect 15660 24278 15712 24284
rect 17132 24336 17184 24342
rect 17132 24278 17184 24284
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15304 23866 15332 24142
rect 15292 23860 15344 23866
rect 15292 23802 15344 23808
rect 15672 23594 15700 24278
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 16212 24064 16264 24070
rect 16212 24006 16264 24012
rect 15660 23588 15712 23594
rect 15660 23530 15712 23536
rect 15108 23248 15160 23254
rect 15108 23190 15160 23196
rect 15120 22574 15148 23190
rect 16224 23186 16252 24006
rect 17328 23254 17356 24142
rect 17420 23866 17448 24550
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 17408 23520 17460 23526
rect 17460 23497 17540 23508
rect 17460 23488 17554 23497
rect 17460 23480 17498 23488
rect 17408 23462 17460 23468
rect 17498 23423 17554 23432
rect 17316 23248 17368 23254
rect 17316 23190 17368 23196
rect 16212 23180 16264 23186
rect 16212 23122 16264 23128
rect 16224 22778 16252 23122
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16776 22778 16804 22986
rect 17328 22778 17356 23190
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 17316 22772 17368 22778
rect 17316 22714 17368 22720
rect 15108 22568 15160 22574
rect 15108 22510 15160 22516
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 15212 21690 15240 22102
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15580 21350 15608 22374
rect 17328 22166 17356 22714
rect 17316 22160 17368 22166
rect 17316 22102 17368 22108
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16028 21956 16080 21962
rect 16028 21898 16080 21904
rect 16040 21554 16068 21898
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 15304 20602 15332 20946
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 19990 15516 20198
rect 15580 19990 15608 21286
rect 15764 21146 15792 21354
rect 16132 21146 16160 21966
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 17316 21072 17368 21078
rect 17316 21014 17368 21020
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16960 20505 16988 20878
rect 16946 20496 17002 20505
rect 16946 20431 17002 20440
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16408 20058 16436 20198
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 15476 19984 15528 19990
rect 15476 19926 15528 19932
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15488 19514 15516 19926
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15580 19446 15608 19926
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16132 19446 16160 19790
rect 16592 19514 16620 20198
rect 16960 20058 16988 20431
rect 17328 20262 17356 21014
rect 17316 20256 17368 20262
rect 17316 20198 17368 20204
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15764 18902 15792 19178
rect 15752 18896 15804 18902
rect 15752 18838 15804 18844
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15948 18222 15976 18362
rect 16040 18222 16068 18566
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15292 18148 15344 18154
rect 15292 18090 15344 18096
rect 15304 17678 15332 18090
rect 16776 18086 16804 18770
rect 16960 18630 16988 19790
rect 17222 19000 17278 19009
rect 17222 18935 17278 18944
rect 17236 18902 17264 18935
rect 17328 18902 17356 20198
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17316 18896 17368 18902
rect 17316 18838 17368 18844
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16960 18465 16988 18566
rect 16946 18456 17002 18465
rect 16946 18391 17002 18400
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15304 16794 15332 17614
rect 15672 17066 15700 17818
rect 16224 17338 16252 18022
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 16132 16658 16160 16934
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15120 14550 15148 14962
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15120 13938 15148 14486
rect 15212 14482 15240 15846
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15212 14074 15240 14418
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15120 13530 15148 13874
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15120 12442 15148 13262
rect 15304 12986 15332 13738
rect 15396 13326 15424 15438
rect 15488 15026 15516 16390
rect 15580 16250 15608 16594
rect 16224 16590 16252 16934
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15856 15638 15884 16390
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15856 14618 15884 15574
rect 15948 14822 15976 15574
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16684 15026 16712 15438
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15948 13870 15976 14758
rect 16408 14618 16436 14962
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15580 13258 15608 13738
rect 16776 13530 16804 18022
rect 17236 17882 17264 18838
rect 17328 18426 17356 18838
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17696 17882 17724 24618
rect 17788 24274 17816 24686
rect 17776 24268 17828 24274
rect 17776 24210 17828 24216
rect 17960 24268 18012 24274
rect 17960 24210 18012 24216
rect 17972 23866 18000 24210
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 17972 23526 18000 23802
rect 18236 23588 18288 23594
rect 18236 23530 18288 23536
rect 17960 23520 18012 23526
rect 17960 23462 18012 23468
rect 18248 23118 18276 23530
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17880 22166 17908 22986
rect 18328 22704 18380 22710
rect 18328 22646 18380 22652
rect 18052 22500 18104 22506
rect 18052 22442 18104 22448
rect 18064 22166 18092 22442
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 18052 22160 18104 22166
rect 18052 22102 18104 22108
rect 17880 21690 17908 22102
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 18064 21622 18092 22102
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 17960 20868 18012 20874
rect 17960 20810 18012 20816
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17880 18902 17908 19722
rect 17972 18970 18000 20810
rect 18064 19990 18092 21558
rect 18236 21412 18288 21418
rect 18236 21354 18288 21360
rect 18248 20806 18276 21354
rect 18340 21010 18368 22646
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18156 20058 18184 20402
rect 18248 20330 18276 20742
rect 18236 20324 18288 20330
rect 18236 20266 18288 20272
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18052 19984 18104 19990
rect 18052 19926 18104 19932
rect 18064 19514 18092 19926
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18248 19242 18276 19450
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18236 19236 18288 19242
rect 18236 19178 18288 19184
rect 18156 18970 18184 19178
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 17880 17746 17908 18022
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 16868 17338 16896 17682
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17868 16992 17920 16998
rect 17972 16980 18000 17682
rect 18248 17610 18276 18090
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18050 17368 18106 17377
rect 18050 17303 18106 17312
rect 17920 16952 18000 16980
rect 17868 16934 17920 16940
rect 17512 16726 17540 16934
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17880 15978 17908 16934
rect 18064 16590 18092 17303
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 18064 16182 18092 16526
rect 18052 16176 18104 16182
rect 18052 16118 18104 16124
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 18064 15638 18092 16118
rect 18156 16046 18184 17478
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18248 16794 18276 17070
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18248 16046 18276 16730
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 18064 15162 18092 15574
rect 18248 15570 18276 15982
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16868 14550 16896 14826
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 15844 13456 15896 13462
rect 15844 13398 15896 13404
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15856 12986 15884 13398
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15396 11558 15424 12242
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15028 10606 15056 10746
rect 15016 10600 15068 10606
rect 14830 10568 14886 10577
rect 15016 10542 15068 10548
rect 14830 10503 14886 10512
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12728 8090 12756 8910
rect 13096 8566 13124 8910
rect 13464 8634 13492 9046
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 13096 7546 13124 7890
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13188 7410 13216 7686
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 1398 4176 1454 4185
rect 1398 4111 1454 4120
rect 3054 4176 3110 4185
rect 3054 4111 3110 4120
rect 2778 82 2834 480
rect 3068 82 3096 4111
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 2778 54 3096 82
rect 8298 82 8354 480
rect 8588 82 8616 7210
rect 13188 7002 13216 7346
rect 13556 7342 13584 9046
rect 13648 8498 13676 9318
rect 14200 9178 14228 9590
rect 14292 9586 14320 9930
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14292 9042 14320 9522
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13188 4185 13216 6598
rect 13740 6390 13768 6802
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13174 4176 13230 4185
rect 13174 4111 13230 4120
rect 8298 54 8616 82
rect 13818 82 13874 480
rect 14108 82 14136 8298
rect 14200 8022 14228 8978
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14384 8430 14412 8774
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14936 8090 14964 9454
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14188 8016 14240 8022
rect 14188 7958 14240 7964
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14660 6730 14688 7210
rect 15028 6866 15056 10542
rect 15396 10266 15424 11494
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15672 10606 15700 11154
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15120 8022 15148 8230
rect 15764 8090 15792 12718
rect 15856 12442 15884 12922
rect 16960 12782 16988 15030
rect 18340 14958 18368 16934
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18340 14618 18368 14894
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 17236 13734 17264 14418
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 18432 13814 18460 26318
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18788 24336 18840 24342
rect 18788 24278 18840 24284
rect 18800 23662 18828 24278
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18616 23254 18644 23462
rect 18604 23248 18656 23254
rect 18604 23190 18656 23196
rect 18616 22438 18644 23190
rect 18788 23112 18840 23118
rect 18788 23054 18840 23060
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 18708 22574 18736 22918
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 18708 22234 18736 22510
rect 18696 22228 18748 22234
rect 18696 22170 18748 22176
rect 18800 22166 18828 23054
rect 18788 22160 18840 22166
rect 18788 22102 18840 22108
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18616 21554 18644 21966
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18524 21146 18552 21490
rect 18512 21140 18564 21146
rect 18512 21082 18564 21088
rect 18616 20466 18644 21490
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18616 18970 18644 19790
rect 18800 19378 18828 20266
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18524 17746 18552 18022
rect 18892 17814 18920 25638
rect 18984 23497 19012 27814
rect 19076 27538 19104 28018
rect 19352 27674 19380 28562
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19064 27532 19116 27538
rect 19064 27474 19116 27480
rect 19076 27130 19104 27474
rect 19064 27124 19116 27130
rect 19064 27066 19116 27072
rect 19064 26444 19116 26450
rect 19064 26386 19116 26392
rect 19076 26042 19104 26386
rect 19064 26036 19116 26042
rect 19064 25978 19116 25984
rect 19444 25362 19472 28902
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 20088 28694 20116 34410
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 20996 33992 21048 33998
rect 20996 33934 21048 33940
rect 21008 33658 21036 33934
rect 20996 33652 21048 33658
rect 20996 33594 21048 33600
rect 21100 33522 21128 34342
rect 21088 33516 21140 33522
rect 21088 33458 21140 33464
rect 20904 33448 20956 33454
rect 20902 33416 20904 33425
rect 20956 33416 20958 33425
rect 20902 33351 20958 33360
rect 20916 33318 20944 33351
rect 20904 33312 20956 33318
rect 20904 33254 20956 33260
rect 21192 33134 21220 34575
rect 21272 34128 21324 34134
rect 21272 34070 21324 34076
rect 21284 33658 21312 34070
rect 21272 33652 21324 33658
rect 21272 33594 21324 33600
rect 21284 33318 21312 33594
rect 21272 33312 21324 33318
rect 21324 33272 21496 33300
rect 21272 33254 21324 33260
rect 20260 33108 20312 33114
rect 21192 33106 21312 33134
rect 20260 33050 20312 33056
rect 20272 32434 20300 33050
rect 20444 32904 20496 32910
rect 20444 32846 20496 32852
rect 20260 32428 20312 32434
rect 20260 32370 20312 32376
rect 20456 32298 20484 32846
rect 20444 32292 20496 32298
rect 20444 32234 20496 32240
rect 21180 32292 21232 32298
rect 21180 32234 21232 32240
rect 20456 31822 20484 32234
rect 21192 31958 21220 32234
rect 21180 31952 21232 31958
rect 21180 31894 21232 31900
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 20444 30184 20496 30190
rect 20444 30126 20496 30132
rect 20456 29510 20484 30126
rect 20916 29850 20944 31078
rect 20996 30116 21048 30122
rect 20996 30058 21048 30064
rect 20904 29844 20956 29850
rect 20904 29786 20956 29792
rect 20260 29504 20312 29510
rect 20260 29446 20312 29452
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 20272 29102 20300 29446
rect 20456 29170 20484 29446
rect 20444 29164 20496 29170
rect 20444 29106 20496 29112
rect 20168 29096 20220 29102
rect 20168 29038 20220 29044
rect 20260 29096 20312 29102
rect 20260 29038 20312 29044
rect 20076 28688 20128 28694
rect 20076 28630 20128 28636
rect 20180 28490 20208 29038
rect 20272 28626 20300 29038
rect 20260 28620 20312 28626
rect 20260 28562 20312 28568
rect 20168 28484 20220 28490
rect 20168 28426 20220 28432
rect 21008 28150 21036 30058
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 21100 28966 21128 29650
rect 21088 28960 21140 28966
rect 21088 28902 21140 28908
rect 21180 28960 21232 28966
rect 21180 28902 21232 28908
rect 21100 28529 21128 28902
rect 21192 28558 21220 28902
rect 21180 28552 21232 28558
rect 21086 28520 21142 28529
rect 21180 28494 21232 28500
rect 21086 28455 21142 28464
rect 21192 28150 21220 28494
rect 20996 28144 21048 28150
rect 20996 28086 21048 28092
rect 21180 28144 21232 28150
rect 21180 28086 21232 28092
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 20352 27940 20404 27946
rect 20352 27882 20404 27888
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 20364 27674 20392 27882
rect 20352 27668 20404 27674
rect 20352 27610 20404 27616
rect 19892 27532 19944 27538
rect 19892 27474 19944 27480
rect 19904 26858 19932 27474
rect 19892 26852 19944 26858
rect 19892 26794 19944 26800
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19984 26240 20036 26246
rect 19984 26182 20036 26188
rect 19996 25906 20024 26182
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19996 25430 20024 25842
rect 19984 25424 20036 25430
rect 19984 25366 20036 25372
rect 20364 25362 20392 27610
rect 21100 27470 21128 27950
rect 21180 27668 21232 27674
rect 21180 27610 21232 27616
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 20904 26784 20956 26790
rect 20904 26726 20956 26732
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 20352 25356 20404 25362
rect 20352 25298 20404 25304
rect 19444 24954 19472 25298
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19798 24848 19854 24857
rect 20272 24818 20300 25230
rect 19798 24783 19854 24792
rect 20260 24812 20312 24818
rect 19812 24750 19840 24783
rect 20260 24754 20312 24760
rect 20364 24750 20392 25298
rect 19800 24744 19852 24750
rect 20352 24744 20404 24750
rect 19852 24704 19932 24732
rect 19800 24686 19852 24692
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19904 24342 19932 24704
rect 20352 24686 20404 24692
rect 20364 24410 20392 24686
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 19892 24336 19944 24342
rect 19892 24278 19944 24284
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 19076 23798 19104 24210
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 18970 23488 19026 23497
rect 18970 23423 19026 23432
rect 18984 22710 19012 23423
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 20088 22982 20116 24346
rect 20916 24206 20944 26726
rect 21100 26586 21128 27406
rect 21192 26790 21220 27610
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 21192 25770 21220 26726
rect 21284 26450 21312 33106
rect 21364 32768 21416 32774
rect 21468 32756 21496 33272
rect 21416 32728 21496 32756
rect 21364 32710 21416 32716
rect 21376 32280 21404 32710
rect 21456 32292 21508 32298
rect 21376 32252 21456 32280
rect 21376 31686 21404 32252
rect 21456 32234 21508 32240
rect 21560 31890 21588 37216
rect 21732 36644 21784 36650
rect 21732 36586 21784 36592
rect 21640 35760 21692 35766
rect 21640 35702 21692 35708
rect 21652 34066 21680 35702
rect 21640 34060 21692 34066
rect 21640 34002 21692 34008
rect 21652 33114 21680 34002
rect 21640 33108 21692 33114
rect 21640 33050 21692 33056
rect 21744 32434 21772 36586
rect 21836 36582 21864 37334
rect 21928 36786 21956 37810
rect 21916 36780 21968 36786
rect 21916 36722 21968 36728
rect 22008 36780 22060 36786
rect 22008 36722 22060 36728
rect 21916 36644 21968 36650
rect 21916 36586 21968 36592
rect 21824 36576 21876 36582
rect 21824 36518 21876 36524
rect 21928 36378 21956 36586
rect 21916 36372 21968 36378
rect 21916 36314 21968 36320
rect 22020 36106 22048 36722
rect 22008 36100 22060 36106
rect 22008 36042 22060 36048
rect 21824 35080 21876 35086
rect 21824 35022 21876 35028
rect 21836 34474 21864 35022
rect 22020 34678 22048 36042
rect 22192 35692 22244 35698
rect 22192 35634 22244 35640
rect 22204 35290 22232 35634
rect 22192 35284 22244 35290
rect 22192 35226 22244 35232
rect 22008 34672 22060 34678
rect 22008 34614 22060 34620
rect 21824 34468 21876 34474
rect 21824 34410 21876 34416
rect 21916 34468 21968 34474
rect 21916 34410 21968 34416
rect 21836 34202 21864 34410
rect 21824 34196 21876 34202
rect 21824 34138 21876 34144
rect 21928 34134 21956 34410
rect 21916 34128 21968 34134
rect 21916 34070 21968 34076
rect 22388 34066 22416 43386
rect 23204 43376 23256 43382
rect 23204 43318 23256 43324
rect 23020 43104 23072 43110
rect 23020 43046 23072 43052
rect 23032 42226 23060 43046
rect 23112 42764 23164 42770
rect 23112 42706 23164 42712
rect 23020 42220 23072 42226
rect 23020 42162 23072 42168
rect 22744 42084 22796 42090
rect 22744 42026 22796 42032
rect 22652 42016 22704 42022
rect 22652 41958 22704 41964
rect 22468 40996 22520 41002
rect 22468 40938 22520 40944
rect 22480 40526 22508 40938
rect 22468 40520 22520 40526
rect 22468 40462 22520 40468
rect 22480 39642 22508 40462
rect 22560 39908 22612 39914
rect 22560 39850 22612 39856
rect 22468 39636 22520 39642
rect 22468 39578 22520 39584
rect 22468 38752 22520 38758
rect 22468 38694 22520 38700
rect 22480 34649 22508 38694
rect 22572 36854 22600 39850
rect 22664 37330 22692 41958
rect 22756 40526 22784 42026
rect 23124 42022 23152 42706
rect 23216 42090 23244 43318
rect 23480 43308 23532 43314
rect 23480 43250 23532 43256
rect 23204 42084 23256 42090
rect 23204 42026 23256 42032
rect 23112 42016 23164 42022
rect 23112 41958 23164 41964
rect 23124 41177 23152 41958
rect 23492 41818 23520 43250
rect 23584 42838 23612 43590
rect 23860 43178 23888 43590
rect 24044 43314 24072 43590
rect 25056 43450 25084 43794
rect 25412 43648 25464 43654
rect 25412 43590 25464 43596
rect 25596 43648 25648 43654
rect 25596 43590 25648 43596
rect 25044 43444 25096 43450
rect 25044 43386 25096 43392
rect 24032 43308 24084 43314
rect 24032 43250 24084 43256
rect 24216 43308 24268 43314
rect 24216 43250 24268 43256
rect 23848 43172 23900 43178
rect 23848 43114 23900 43120
rect 23572 42832 23624 42838
rect 23572 42774 23624 42780
rect 23664 42832 23716 42838
rect 23664 42774 23716 42780
rect 23584 41818 23612 42774
rect 23676 42294 23704 42774
rect 23756 42560 23808 42566
rect 23756 42502 23808 42508
rect 23664 42288 23716 42294
rect 23664 42230 23716 42236
rect 23676 42004 23704 42230
rect 23768 42226 23796 42502
rect 23756 42220 23808 42226
rect 23756 42162 23808 42168
rect 23756 42016 23808 42022
rect 23676 41976 23756 42004
rect 23756 41958 23808 41964
rect 23480 41812 23532 41818
rect 23480 41754 23532 41760
rect 23572 41812 23624 41818
rect 23572 41754 23624 41760
rect 23296 41744 23348 41750
rect 23296 41686 23348 41692
rect 23664 41744 23716 41750
rect 23664 41686 23716 41692
rect 23110 41168 23166 41177
rect 23110 41103 23166 41112
rect 23112 41064 23164 41070
rect 23112 41006 23164 41012
rect 23204 41064 23256 41070
rect 23204 41006 23256 41012
rect 22928 40656 22980 40662
rect 22928 40598 22980 40604
rect 22744 40520 22796 40526
rect 22744 40462 22796 40468
rect 22940 39846 22968 40598
rect 23020 39976 23072 39982
rect 23020 39918 23072 39924
rect 22928 39840 22980 39846
rect 22928 39782 22980 39788
rect 22940 39574 22968 39782
rect 22928 39568 22980 39574
rect 22928 39510 22980 39516
rect 22940 39302 22968 39510
rect 22928 39296 22980 39302
rect 22928 39238 22980 39244
rect 22940 38758 22968 39238
rect 22928 38752 22980 38758
rect 22928 38694 22980 38700
rect 22940 38486 22968 38694
rect 22836 38480 22888 38486
rect 22836 38422 22888 38428
rect 22928 38480 22980 38486
rect 22928 38422 22980 38428
rect 22848 38010 22876 38422
rect 22836 38004 22888 38010
rect 22836 37946 22888 37952
rect 22940 37398 22968 38422
rect 22928 37392 22980 37398
rect 22928 37334 22980 37340
rect 22652 37324 22704 37330
rect 22652 37266 22704 37272
rect 22560 36848 22612 36854
rect 22560 36790 22612 36796
rect 22664 36786 22692 37266
rect 22652 36780 22704 36786
rect 22652 36722 22704 36728
rect 22664 36689 22692 36722
rect 22650 36680 22706 36689
rect 22650 36615 22706 36624
rect 23032 36242 23060 39918
rect 23020 36236 23072 36242
rect 23020 36178 23072 36184
rect 23032 35834 23060 36178
rect 23020 35828 23072 35834
rect 23020 35770 23072 35776
rect 22836 35148 22888 35154
rect 22836 35090 22888 35096
rect 22848 34746 22876 35090
rect 22836 34740 22888 34746
rect 22836 34682 22888 34688
rect 22466 34640 22522 34649
rect 22466 34575 22522 34584
rect 22376 34060 22428 34066
rect 22376 34002 22428 34008
rect 22388 33658 22416 34002
rect 22376 33652 22428 33658
rect 22376 33594 22428 33600
rect 22388 33114 22416 33594
rect 22848 33134 22876 34682
rect 23032 33998 23060 35770
rect 23124 34066 23152 41006
rect 23216 35766 23244 41006
rect 23308 40730 23336 41686
rect 23676 41274 23704 41686
rect 23480 41268 23532 41274
rect 23480 41210 23532 41216
rect 23664 41268 23716 41274
rect 23664 41210 23716 41216
rect 23296 40724 23348 40730
rect 23296 40666 23348 40672
rect 23296 40452 23348 40458
rect 23296 40394 23348 40400
rect 23308 40186 23336 40394
rect 23296 40180 23348 40186
rect 23296 40122 23348 40128
rect 23492 39098 23520 41210
rect 23572 40112 23624 40118
rect 23572 40054 23624 40060
rect 23480 39092 23532 39098
rect 23480 39034 23532 39040
rect 23388 38820 23440 38826
rect 23388 38762 23440 38768
rect 23400 38554 23428 38762
rect 23492 38758 23520 39034
rect 23584 38826 23612 40054
rect 23664 39840 23716 39846
rect 23664 39782 23716 39788
rect 23676 39438 23704 39782
rect 23664 39432 23716 39438
rect 23664 39374 23716 39380
rect 23676 39098 23704 39374
rect 23664 39092 23716 39098
rect 23664 39034 23716 39040
rect 23572 38820 23624 38826
rect 23572 38762 23624 38768
rect 23480 38752 23532 38758
rect 23480 38694 23532 38700
rect 23388 38548 23440 38554
rect 23388 38490 23440 38496
rect 23492 37466 23520 38694
rect 23768 38010 23796 41958
rect 23860 41274 23888 43114
rect 24228 42838 24256 43250
rect 24216 42832 24268 42838
rect 24216 42774 24268 42780
rect 23848 41268 23900 41274
rect 23848 41210 23900 41216
rect 23848 41132 23900 41138
rect 23848 41074 23900 41080
rect 23860 39001 23888 41074
rect 23940 40996 23992 41002
rect 23940 40938 23992 40944
rect 23846 38992 23902 39001
rect 23846 38927 23902 38936
rect 23756 38004 23808 38010
rect 23756 37946 23808 37952
rect 23860 37670 23888 38927
rect 23848 37664 23900 37670
rect 23848 37606 23900 37612
rect 23480 37460 23532 37466
rect 23480 37402 23532 37408
rect 23860 37398 23888 37606
rect 23848 37392 23900 37398
rect 23848 37334 23900 37340
rect 23860 36786 23888 37334
rect 23848 36780 23900 36786
rect 23848 36722 23900 36728
rect 23572 36576 23624 36582
rect 23572 36518 23624 36524
rect 23584 36378 23612 36518
rect 23572 36372 23624 36378
rect 23572 36314 23624 36320
rect 23204 35760 23256 35766
rect 23204 35702 23256 35708
rect 23216 35154 23244 35702
rect 23204 35148 23256 35154
rect 23204 35090 23256 35096
rect 23756 34944 23808 34950
rect 23756 34886 23808 34892
rect 23296 34672 23348 34678
rect 23296 34614 23348 34620
rect 23112 34060 23164 34066
rect 23112 34002 23164 34008
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 22376 33108 22428 33114
rect 22376 33050 22428 33056
rect 22756 33106 22876 33134
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 22112 32502 22140 32914
rect 22284 32904 22336 32910
rect 22284 32846 22336 32852
rect 22296 32570 22324 32846
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 22100 32496 22152 32502
rect 22100 32438 22152 32444
rect 21732 32428 21784 32434
rect 21732 32370 21784 32376
rect 21548 31884 21600 31890
rect 21548 31826 21600 31832
rect 21364 31680 21416 31686
rect 21364 31622 21416 31628
rect 21376 30394 21404 31622
rect 21560 31482 21588 31826
rect 21548 31476 21600 31482
rect 21548 31418 21600 31424
rect 21744 31414 21772 32370
rect 22112 32026 22140 32438
rect 22296 32212 22324 32506
rect 22376 32224 22428 32230
rect 22296 32184 22376 32212
rect 22376 32166 22428 32172
rect 22100 32020 22152 32026
rect 22100 31962 22152 31968
rect 21732 31408 21784 31414
rect 21732 31350 21784 31356
rect 22112 31278 22140 31962
rect 21916 31272 21968 31278
rect 21916 31214 21968 31220
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 21640 31136 21692 31142
rect 21640 31078 21692 31084
rect 21364 30388 21416 30394
rect 21364 30330 21416 30336
rect 21456 29708 21508 29714
rect 21456 29650 21508 29656
rect 21468 29306 21496 29650
rect 21456 29300 21508 29306
rect 21456 29242 21508 29248
rect 21456 28620 21508 28626
rect 21456 28562 21508 28568
rect 21468 28150 21496 28562
rect 21548 28552 21600 28558
rect 21548 28494 21600 28500
rect 21456 28144 21508 28150
rect 21456 28086 21508 28092
rect 21468 27946 21496 28086
rect 21456 27940 21508 27946
rect 21456 27882 21508 27888
rect 21560 26994 21588 28494
rect 21652 28218 21680 31078
rect 21732 30796 21784 30802
rect 21732 30738 21784 30744
rect 21744 30054 21772 30738
rect 21928 30666 21956 31214
rect 21916 30660 21968 30666
rect 21916 30602 21968 30608
rect 21732 30048 21784 30054
rect 21732 29990 21784 29996
rect 21744 29102 21772 29990
rect 22112 29714 22140 31214
rect 22284 31136 22336 31142
rect 22284 31078 22336 31084
rect 22296 29782 22324 31078
rect 22284 29776 22336 29782
rect 22284 29718 22336 29724
rect 22100 29708 22152 29714
rect 22100 29650 22152 29656
rect 22112 29102 22140 29650
rect 22388 29617 22416 32166
rect 22652 31816 22704 31822
rect 22652 31758 22704 31764
rect 22664 31346 22692 31758
rect 22652 31340 22704 31346
rect 22652 31282 22704 31288
rect 22756 30802 22784 33106
rect 23308 33046 23336 34614
rect 23768 34542 23796 34886
rect 23860 34678 23888 36722
rect 23848 34672 23900 34678
rect 23848 34614 23900 34620
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 23388 33448 23440 33454
rect 23388 33390 23440 33396
rect 23296 33040 23348 33046
rect 23400 33017 23428 33390
rect 23768 33318 23796 34478
rect 23860 34474 23888 34614
rect 23848 34468 23900 34474
rect 23848 34410 23900 34416
rect 23848 33856 23900 33862
rect 23848 33798 23900 33804
rect 23860 33454 23888 33798
rect 23952 33522 23980 40938
rect 24228 39370 24256 42774
rect 24400 42696 24452 42702
rect 24400 42638 24452 42644
rect 24412 42226 24440 42638
rect 24400 42220 24452 42226
rect 24400 42162 24452 42168
rect 24412 41750 24440 42162
rect 24400 41744 24452 41750
rect 24400 41686 24452 41692
rect 24412 40526 24440 41686
rect 24768 41676 24820 41682
rect 24768 41618 24820 41624
rect 24780 41274 24808 41618
rect 24768 41268 24820 41274
rect 24768 41210 24820 41216
rect 24584 40928 24636 40934
rect 24584 40870 24636 40876
rect 24492 40656 24544 40662
rect 24492 40598 24544 40604
rect 24400 40520 24452 40526
rect 24400 40462 24452 40468
rect 24412 40186 24440 40462
rect 24400 40180 24452 40186
rect 24400 40122 24452 40128
rect 24504 39846 24532 40598
rect 24492 39840 24544 39846
rect 24492 39782 24544 39788
rect 24504 39574 24532 39782
rect 24492 39568 24544 39574
rect 24492 39510 24544 39516
rect 24032 39364 24084 39370
rect 24032 39306 24084 39312
rect 24216 39364 24268 39370
rect 24216 39306 24268 39312
rect 24044 38758 24072 39306
rect 24228 38962 24256 39306
rect 24400 39296 24452 39302
rect 24400 39238 24452 39244
rect 24216 38956 24268 38962
rect 24216 38898 24268 38904
rect 24032 38752 24084 38758
rect 24032 38694 24084 38700
rect 24412 38486 24440 39238
rect 24596 38554 24624 40870
rect 24584 38548 24636 38554
rect 24584 38490 24636 38496
rect 24400 38480 24452 38486
rect 24400 38422 24452 38428
rect 24032 37256 24084 37262
rect 24032 37198 24084 37204
rect 24044 36650 24072 37198
rect 24674 36680 24730 36689
rect 24032 36644 24084 36650
rect 24674 36615 24730 36624
rect 24032 36586 24084 36592
rect 24688 36582 24716 36615
rect 24676 36576 24728 36582
rect 24676 36518 24728 36524
rect 25056 36378 25084 43386
rect 25424 42838 25452 43590
rect 25608 43178 25636 43590
rect 26608 43376 26660 43382
rect 26608 43318 26660 43324
rect 25504 43172 25556 43178
rect 25504 43114 25556 43120
rect 25596 43172 25648 43178
rect 25596 43114 25648 43120
rect 25412 42832 25464 42838
rect 25412 42774 25464 42780
rect 25320 42764 25372 42770
rect 25320 42706 25372 42712
rect 25332 42362 25360 42706
rect 25320 42356 25372 42362
rect 25320 42298 25372 42304
rect 25516 41818 25544 43114
rect 25608 42794 25636 43114
rect 26240 42832 26292 42838
rect 25608 42766 25728 42794
rect 26240 42774 26292 42780
rect 25596 42560 25648 42566
rect 25596 42502 25648 42508
rect 25608 42226 25636 42502
rect 25596 42220 25648 42226
rect 25596 42162 25648 42168
rect 25700 42090 25728 42766
rect 25688 42084 25740 42090
rect 25688 42026 25740 42032
rect 25700 41818 25728 42026
rect 26252 41818 26280 42774
rect 26620 42090 26648 43318
rect 27528 43240 27580 43246
rect 27528 43182 27580 43188
rect 27988 43240 28040 43246
rect 27988 43182 28040 43188
rect 26700 42832 26752 42838
rect 26700 42774 26752 42780
rect 26712 42294 26740 42774
rect 27540 42770 27568 43182
rect 27620 43104 27672 43110
rect 27620 43046 27672 43052
rect 27528 42764 27580 42770
rect 27528 42706 27580 42712
rect 26700 42288 26752 42294
rect 26700 42230 26752 42236
rect 26608 42084 26660 42090
rect 26608 42026 26660 42032
rect 25504 41812 25556 41818
rect 25504 41754 25556 41760
rect 25688 41812 25740 41818
rect 25688 41754 25740 41760
rect 26240 41812 26292 41818
rect 26240 41754 26292 41760
rect 26620 41614 26648 42026
rect 26712 42022 26740 42230
rect 27632 42226 27660 43046
rect 28000 42906 28028 43182
rect 27988 42900 28040 42906
rect 27988 42842 28040 42848
rect 27620 42220 27672 42226
rect 27620 42162 27672 42168
rect 26700 42016 26752 42022
rect 26700 41958 26752 41964
rect 27252 42016 27304 42022
rect 27252 41958 27304 41964
rect 26700 41744 26752 41750
rect 26700 41686 26752 41692
rect 26608 41608 26660 41614
rect 26608 41550 26660 41556
rect 26620 41274 26648 41550
rect 26608 41268 26660 41274
rect 26608 41210 26660 41216
rect 26712 41206 26740 41686
rect 26884 41608 26936 41614
rect 26884 41550 26936 41556
rect 26700 41200 26752 41206
rect 26700 41142 26752 41148
rect 25228 41064 25280 41070
rect 25228 41006 25280 41012
rect 25240 40730 25268 41006
rect 25688 40928 25740 40934
rect 25688 40870 25740 40876
rect 25228 40724 25280 40730
rect 25228 40666 25280 40672
rect 25700 39914 25728 40870
rect 26792 40112 26844 40118
rect 26792 40054 26844 40060
rect 25780 40044 25832 40050
rect 25780 39986 25832 39992
rect 25688 39908 25740 39914
rect 25688 39850 25740 39856
rect 25136 39500 25188 39506
rect 25136 39442 25188 39448
rect 25148 38758 25176 39442
rect 25320 39432 25372 39438
rect 25320 39374 25372 39380
rect 25332 38826 25360 39374
rect 25792 39302 25820 39986
rect 26700 39568 26752 39574
rect 26700 39510 26752 39516
rect 26240 39364 26292 39370
rect 26240 39306 26292 39312
rect 25780 39296 25832 39302
rect 25780 39238 25832 39244
rect 25792 38962 25820 39238
rect 25780 38956 25832 38962
rect 25780 38898 25832 38904
rect 25320 38820 25372 38826
rect 25596 38820 25648 38826
rect 25320 38762 25372 38768
rect 25516 38780 25596 38808
rect 25136 38752 25188 38758
rect 25136 38694 25188 38700
rect 25136 38480 25188 38486
rect 25136 38422 25188 38428
rect 25148 38010 25176 38422
rect 25332 38350 25360 38762
rect 25320 38344 25372 38350
rect 25320 38286 25372 38292
rect 25516 38214 25544 38780
rect 25596 38762 25648 38768
rect 25688 38752 25740 38758
rect 25688 38694 25740 38700
rect 25700 38332 25728 38694
rect 25792 38457 25820 38898
rect 26252 38554 26280 39306
rect 26712 39030 26740 39510
rect 26700 39024 26752 39030
rect 26700 38966 26752 38972
rect 26240 38548 26292 38554
rect 26240 38490 26292 38496
rect 26608 38480 26660 38486
rect 25778 38448 25834 38457
rect 26608 38422 26660 38428
rect 26700 38480 26752 38486
rect 26700 38422 26752 38428
rect 25778 38383 25834 38392
rect 25700 38304 25820 38332
rect 25504 38208 25556 38214
rect 25504 38150 25556 38156
rect 25516 38010 25544 38150
rect 25136 38004 25188 38010
rect 25136 37946 25188 37952
rect 25504 38004 25556 38010
rect 25504 37946 25556 37952
rect 25688 37664 25740 37670
rect 25688 37606 25740 37612
rect 25228 37120 25280 37126
rect 25228 37062 25280 37068
rect 25240 36718 25268 37062
rect 25700 36786 25728 37606
rect 25688 36780 25740 36786
rect 25688 36722 25740 36728
rect 25228 36712 25280 36718
rect 25228 36654 25280 36660
rect 25240 36378 25268 36654
rect 25044 36372 25096 36378
rect 25044 36314 25096 36320
rect 25228 36372 25280 36378
rect 25228 36314 25280 36320
rect 24308 36304 24360 36310
rect 24308 36246 24360 36252
rect 24124 36100 24176 36106
rect 24124 36042 24176 36048
rect 24032 36032 24084 36038
rect 24032 35974 24084 35980
rect 24044 35562 24072 35974
rect 24032 35556 24084 35562
rect 24032 35498 24084 35504
rect 24044 34678 24072 35498
rect 24136 35494 24164 36042
rect 24320 35698 24348 36246
rect 24492 36168 24544 36174
rect 24492 36110 24544 36116
rect 24308 35692 24360 35698
rect 24308 35634 24360 35640
rect 24320 35544 24348 35634
rect 24400 35556 24452 35562
rect 24320 35516 24400 35544
rect 24124 35488 24176 35494
rect 24124 35430 24176 35436
rect 24032 34672 24084 34678
rect 24032 34614 24084 34620
rect 24136 34202 24164 35430
rect 24320 35222 24348 35516
rect 24400 35498 24452 35504
rect 24308 35216 24360 35222
rect 24308 35158 24360 35164
rect 24216 35080 24268 35086
rect 24216 35022 24268 35028
rect 24228 34610 24256 35022
rect 24320 34746 24348 35158
rect 24308 34740 24360 34746
rect 24308 34682 24360 34688
rect 24216 34604 24268 34610
rect 24216 34546 24268 34552
rect 24228 34202 24256 34546
rect 24124 34196 24176 34202
rect 24124 34138 24176 34144
rect 24216 34196 24268 34202
rect 24216 34138 24268 34144
rect 24308 33652 24360 33658
rect 24308 33594 24360 33600
rect 23940 33516 23992 33522
rect 23940 33458 23992 33464
rect 23848 33448 23900 33454
rect 23848 33390 23900 33396
rect 23756 33312 23808 33318
rect 23756 33254 23808 33260
rect 23952 33134 23980 33458
rect 24124 33448 24176 33454
rect 24124 33390 24176 33396
rect 23480 33108 23532 33114
rect 23480 33050 23532 33056
rect 23584 33106 23980 33134
rect 23296 32982 23348 32988
rect 23386 33008 23442 33017
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 22848 32570 22876 32846
rect 22836 32564 22888 32570
rect 22836 32506 22888 32512
rect 23308 32230 23336 32982
rect 23386 32943 23442 32952
rect 23492 32910 23520 33050
rect 23480 32904 23532 32910
rect 23480 32846 23532 32852
rect 23020 32224 23072 32230
rect 23020 32166 23072 32172
rect 23296 32224 23348 32230
rect 23296 32166 23348 32172
rect 23032 32026 23060 32166
rect 23020 32020 23072 32026
rect 23020 31962 23072 31968
rect 23032 31142 23060 31962
rect 23020 31136 23072 31142
rect 23020 31078 23072 31084
rect 22744 30796 22796 30802
rect 22744 30738 22796 30744
rect 22756 30394 22784 30738
rect 23020 30592 23072 30598
rect 23020 30534 23072 30540
rect 22744 30388 22796 30394
rect 22744 30330 22796 30336
rect 22374 29608 22430 29617
rect 22374 29543 22430 29552
rect 22468 29572 22520 29578
rect 22468 29514 22520 29520
rect 21732 29096 21784 29102
rect 21732 29038 21784 29044
rect 22008 29096 22060 29102
rect 22008 29038 22060 29044
rect 22100 29096 22152 29102
rect 22100 29038 22152 29044
rect 21640 28212 21692 28218
rect 21640 28154 21692 28160
rect 21744 27849 21772 29038
rect 22020 28801 22048 29038
rect 22006 28792 22062 28801
rect 22112 28762 22140 29038
rect 22006 28727 22062 28736
rect 22100 28756 22152 28762
rect 22100 28698 22152 28704
rect 22480 28626 22508 29514
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22480 28082 22508 28562
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 21824 27940 21876 27946
rect 21824 27882 21876 27888
rect 21916 27940 21968 27946
rect 21916 27882 21968 27888
rect 21730 27840 21786 27849
rect 21730 27775 21786 27784
rect 21836 27316 21864 27882
rect 21928 27674 21956 27882
rect 21916 27668 21968 27674
rect 21916 27610 21968 27616
rect 21916 27328 21968 27334
rect 21836 27288 21916 27316
rect 21916 27270 21968 27276
rect 21548 26988 21600 26994
rect 21548 26930 21600 26936
rect 21560 26586 21588 26930
rect 21548 26580 21600 26586
rect 21548 26522 21600 26528
rect 21272 26444 21324 26450
rect 21272 26386 21324 26392
rect 21284 26042 21312 26386
rect 21824 26240 21876 26246
rect 21824 26182 21876 26188
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 21836 25974 21864 26182
rect 21824 25968 21876 25974
rect 21824 25910 21876 25916
rect 21732 25900 21784 25906
rect 21732 25842 21784 25848
rect 21744 25770 21772 25842
rect 21836 25770 21864 25910
rect 21180 25764 21232 25770
rect 21180 25706 21232 25712
rect 21732 25764 21784 25770
rect 21732 25706 21784 25712
rect 21824 25764 21876 25770
rect 21824 25706 21876 25712
rect 21192 25498 21220 25706
rect 21180 25492 21232 25498
rect 21180 25434 21232 25440
rect 21192 24954 21220 25434
rect 21744 25226 21772 25706
rect 21732 25220 21784 25226
rect 21732 25162 21784 25168
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 21180 24948 21232 24954
rect 21180 24890 21232 24896
rect 21284 24818 21312 25094
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21284 24682 21312 24754
rect 21180 24676 21232 24682
rect 21180 24618 21232 24624
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21088 24336 21140 24342
rect 21088 24278 21140 24284
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 20168 23656 20220 23662
rect 20168 23598 20220 23604
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 18972 22704 19024 22710
rect 18972 22646 19024 22652
rect 19246 22672 19302 22681
rect 19246 22607 19248 22616
rect 19300 22607 19302 22616
rect 19248 22578 19300 22584
rect 19260 22098 19288 22578
rect 19430 22536 19486 22545
rect 19430 22471 19486 22480
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19260 21690 19288 22034
rect 19444 21962 19472 22471
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19432 21956 19484 21962
rect 19432 21898 19484 21904
rect 19444 21690 19472 21898
rect 19248 21684 19300 21690
rect 19248 21626 19300 21632
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 20088 21486 20116 22918
rect 20180 22409 20208 23598
rect 20720 23588 20772 23594
rect 20720 23530 20772 23536
rect 20732 23322 20760 23530
rect 20916 23474 20944 24142
rect 21100 23526 21128 24278
rect 21192 23730 21220 24618
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 20824 23446 20944 23474
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20824 23254 20852 23446
rect 20812 23248 20864 23254
rect 20812 23190 20864 23196
rect 21100 22778 21128 23462
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21284 22778 21312 23122
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21272 22772 21324 22778
rect 21324 22732 21496 22760
rect 21272 22714 21324 22720
rect 20260 22568 20312 22574
rect 20260 22510 20312 22516
rect 20166 22400 20222 22409
rect 20166 22335 20222 22344
rect 20272 21894 20300 22510
rect 21100 22166 21128 22714
rect 21088 22160 21140 22166
rect 21088 22102 21140 22108
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20272 21554 20300 21830
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 20088 21146 20116 21422
rect 20076 21140 20128 21146
rect 20076 21082 20128 21088
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18984 19854 19012 20878
rect 19076 20602 19104 20946
rect 21008 20874 21036 21966
rect 21100 21690 21128 22102
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18984 19446 19012 19790
rect 18972 19440 19024 19446
rect 18972 19382 19024 19388
rect 19444 18902 19472 20198
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 20088 20058 20116 20402
rect 21284 20398 21312 20742
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 20352 20324 20404 20330
rect 20352 20266 20404 20272
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19720 19378 19748 19654
rect 20364 19378 20392 20266
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 21008 19514 21036 19858
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21192 19514 21220 19654
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19352 17882 19380 18838
rect 19444 18426 19472 18838
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 18880 17808 18932 17814
rect 18880 17750 18932 17756
rect 19444 17746 19472 18226
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 18524 16998 18552 17682
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18524 16658 18552 16934
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18524 16114 18552 16594
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18524 16017 18552 16050
rect 18510 16008 18566 16017
rect 18510 15943 18566 15952
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18616 15162 18644 15506
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15948 11218 15976 12378
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15948 10742 15976 11154
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15842 10160 15898 10169
rect 15842 10095 15898 10104
rect 15856 10062 15884 10095
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15856 9722 15884 9998
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15856 8090 15884 9658
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15948 8022 15976 10678
rect 16132 10674 16160 11086
rect 16684 10810 16712 11086
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16132 10266 16160 10610
rect 16672 10532 16724 10538
rect 16776 10520 16804 12582
rect 16960 12442 16988 12718
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17052 12374 17080 13262
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17144 10810 17172 11222
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 16724 10492 16804 10520
rect 16672 10474 16724 10480
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16684 10198 16712 10474
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16500 8838 16528 9998
rect 16684 9722 16712 10134
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8090 16528 8774
rect 16592 8566 16620 9590
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 15120 7313 15148 7958
rect 15948 7546 15976 7958
rect 16592 7954 16620 8502
rect 17236 8090 17264 13670
rect 17512 10810 17540 13806
rect 18432 13786 18552 13814
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17880 11898 17908 12310
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17972 11830 18000 12310
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17696 11150 17724 11630
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17604 9110 17632 9862
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17512 8362 17540 8910
rect 17604 8634 17632 9046
rect 17696 8974 17724 11086
rect 18064 10606 18092 13126
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18248 10674 18276 12650
rect 18340 11898 18368 13466
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18432 12646 18460 12786
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18420 12164 18472 12170
rect 18420 12106 18472 12112
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18432 11694 18460 12106
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18064 10266 18092 10542
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17512 8090 17540 8298
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 16592 7546 16620 7890
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 15106 7304 15162 7313
rect 15106 7239 15162 7248
rect 15120 7002 15148 7239
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14660 6322 14688 6666
rect 15212 6458 15240 6734
rect 15580 6458 15608 7142
rect 17052 6934 17080 7142
rect 17040 6928 17092 6934
rect 17040 6870 17092 6876
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15948 6458 15976 6802
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 17052 6322 17080 6870
rect 17144 6458 17172 7890
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 17420 6866 17448 7210
rect 17696 7206 17724 7822
rect 17788 7342 17816 8366
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 17788 6390 17816 7278
rect 17880 7002 17908 8366
rect 17960 7948 18012 7954
rect 18064 7936 18092 10202
rect 18524 9722 18552 13786
rect 18696 13796 18748 13802
rect 18696 13738 18748 13744
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18616 13190 18644 13330
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18616 12209 18644 13126
rect 18602 12200 18658 12209
rect 18602 12135 18658 12144
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18524 9518 18552 9658
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18012 7908 18092 7936
rect 17960 7890 18012 7896
rect 18524 7886 18552 9318
rect 18708 9042 18736 13738
rect 18800 13462 18828 14418
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18800 11218 18828 13398
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18984 12374 19012 12582
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18892 11558 18920 12242
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 19076 11506 19104 15846
rect 19168 12306 19196 17206
rect 19352 15570 19380 17546
rect 19444 17338 19472 17682
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19444 16794 19472 17274
rect 19628 17066 19656 17682
rect 20364 17678 20392 19314
rect 21008 18970 21036 19450
rect 21192 19174 21220 19450
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19616 17060 19668 17066
rect 19616 17002 19668 17008
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19904 16590 19932 17070
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 20456 16250 20484 18022
rect 20548 17202 20576 18838
rect 21284 18426 21312 20334
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21376 18970 21404 19314
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 20628 18148 20680 18154
rect 20628 18090 20680 18096
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20548 16794 20576 17138
rect 20640 17066 20668 18090
rect 21468 17921 21496 22732
rect 21640 22500 21692 22506
rect 21640 22442 21692 22448
rect 21652 21690 21680 22442
rect 21744 22166 21772 25162
rect 21928 24206 21956 27270
rect 22296 26246 22324 28018
rect 22468 26784 22520 26790
rect 22468 26726 22520 26732
rect 22480 26518 22508 26726
rect 22468 26512 22520 26518
rect 22468 26454 22520 26460
rect 22284 26240 22336 26246
rect 22284 26182 22336 26188
rect 22296 25974 22324 26182
rect 22480 26042 22508 26454
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 22836 26308 22888 26314
rect 22836 26250 22888 26256
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22284 25968 22336 25974
rect 22284 25910 22336 25916
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 22112 24954 22140 25230
rect 22100 24948 22152 24954
rect 22100 24890 22152 24896
rect 22296 24818 22324 25910
rect 22284 24812 22336 24818
rect 22284 24754 22336 24760
rect 22848 24342 22876 26250
rect 22940 26042 22968 26318
rect 22928 26036 22980 26042
rect 22928 25978 22980 25984
rect 22940 25702 22968 25978
rect 22928 25696 22980 25702
rect 22928 25638 22980 25644
rect 23032 24954 23060 30534
rect 23480 30388 23532 30394
rect 23480 30330 23532 30336
rect 23492 29850 23520 30330
rect 23480 29844 23532 29850
rect 23480 29786 23532 29792
rect 23112 29776 23164 29782
rect 23112 29718 23164 29724
rect 23124 29306 23152 29718
rect 23388 29640 23440 29646
rect 23388 29582 23440 29588
rect 23478 29608 23534 29617
rect 23400 29306 23428 29582
rect 23478 29543 23534 29552
rect 23112 29300 23164 29306
rect 23112 29242 23164 29248
rect 23388 29300 23440 29306
rect 23388 29242 23440 29248
rect 23112 28620 23164 28626
rect 23112 28562 23164 28568
rect 23124 28150 23152 28562
rect 23204 28552 23256 28558
rect 23204 28494 23256 28500
rect 23112 28144 23164 28150
rect 23112 28086 23164 28092
rect 23216 27674 23244 28494
rect 23204 27668 23256 27674
rect 23204 27610 23256 27616
rect 23204 25220 23256 25226
rect 23204 25162 23256 25168
rect 23020 24948 23072 24954
rect 23020 24890 23072 24896
rect 22928 24608 22980 24614
rect 22928 24550 22980 24556
rect 22836 24336 22888 24342
rect 22836 24278 22888 24284
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 21928 23050 21956 24142
rect 22848 23866 22876 24278
rect 22940 24206 22968 24550
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 23112 23656 23164 23662
rect 23112 23598 23164 23604
rect 22836 23520 22888 23526
rect 22836 23462 22888 23468
rect 22100 23180 22152 23186
rect 22100 23122 22152 23128
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 21916 22704 21968 22710
rect 21916 22646 21968 22652
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21732 22160 21784 22166
rect 21732 22102 21784 22108
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21652 21418 21680 21626
rect 21744 21622 21772 22102
rect 21836 22001 21864 22374
rect 21822 21992 21878 22001
rect 21822 21927 21878 21936
rect 21732 21616 21784 21622
rect 21732 21558 21784 21564
rect 21732 21480 21784 21486
rect 21732 21422 21784 21428
rect 21640 21412 21692 21418
rect 21640 21354 21692 21360
rect 21744 21146 21772 21422
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21928 21010 21956 22646
rect 22112 22574 22140 23122
rect 22100 22568 22152 22574
rect 22100 22510 22152 22516
rect 22112 21894 22140 22510
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22112 21010 22140 21830
rect 22848 21554 22876 23462
rect 23124 23225 23152 23598
rect 23110 23216 23166 23225
rect 23110 23151 23166 23160
rect 23020 23112 23072 23118
rect 23216 23100 23244 25162
rect 23492 24857 23520 29543
rect 23584 25362 23612 33106
rect 24136 32978 24164 33390
rect 24124 32972 24176 32978
rect 24124 32914 24176 32920
rect 24124 32768 24176 32774
rect 24124 32710 24176 32716
rect 24136 32298 24164 32710
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 24124 32292 24176 32298
rect 24124 32234 24176 32240
rect 24136 32026 24164 32234
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 24228 31754 24256 32370
rect 24216 31748 24268 31754
rect 24216 31690 24268 31696
rect 23756 31136 23808 31142
rect 23756 31078 23808 31084
rect 23768 29753 23796 31078
rect 23848 30864 23900 30870
rect 23848 30806 23900 30812
rect 23860 30394 23888 30806
rect 23940 30728 23992 30734
rect 23940 30670 23992 30676
rect 24124 30728 24176 30734
rect 24228 30716 24256 31690
rect 24176 30688 24256 30716
rect 24124 30670 24176 30676
rect 23952 30394 23980 30670
rect 23848 30388 23900 30394
rect 23848 30330 23900 30336
rect 23940 30388 23992 30394
rect 23940 30330 23992 30336
rect 24136 30258 24164 30670
rect 24124 30252 24176 30258
rect 24124 30194 24176 30200
rect 23848 30116 23900 30122
rect 23848 30058 23900 30064
rect 24124 30116 24176 30122
rect 24124 30058 24176 30064
rect 23754 29744 23810 29753
rect 23754 29679 23810 29688
rect 23768 29578 23796 29679
rect 23860 29578 23888 30058
rect 24136 29714 24164 30058
rect 24124 29708 24176 29714
rect 24124 29650 24176 29656
rect 23940 29640 23992 29646
rect 23940 29582 23992 29588
rect 23756 29572 23808 29578
rect 23756 29514 23808 29520
rect 23848 29572 23900 29578
rect 23848 29514 23900 29520
rect 23952 29306 23980 29582
rect 23940 29300 23992 29306
rect 23940 29242 23992 29248
rect 24320 28994 24348 33594
rect 24504 32026 24532 36110
rect 25792 35018 25820 38304
rect 26620 37942 26648 38422
rect 26608 37936 26660 37942
rect 26608 37878 26660 37884
rect 26516 37800 26568 37806
rect 26516 37742 26568 37748
rect 25964 37664 26016 37670
rect 25964 37606 26016 37612
rect 25976 37466 26004 37606
rect 26528 37466 26556 37742
rect 26712 37738 26740 38422
rect 26700 37732 26752 37738
rect 26700 37674 26752 37680
rect 25964 37460 26016 37466
rect 25964 37402 26016 37408
rect 26516 37460 26568 37466
rect 26516 37402 26568 37408
rect 26608 37324 26660 37330
rect 26608 37266 26660 37272
rect 26620 36854 26648 37266
rect 26608 36848 26660 36854
rect 26608 36790 26660 36796
rect 26804 36718 26832 40054
rect 26896 39438 26924 41550
rect 27264 41002 27292 41958
rect 27344 41132 27396 41138
rect 27344 41074 27396 41080
rect 27252 40996 27304 41002
rect 27252 40938 27304 40944
rect 27356 40390 27384 41074
rect 28000 40594 28028 42842
rect 29184 42764 29236 42770
rect 29184 42706 29236 42712
rect 29552 42764 29604 42770
rect 29552 42706 29604 42712
rect 29196 42090 29224 42706
rect 29460 42152 29512 42158
rect 29460 42094 29512 42100
rect 29184 42084 29236 42090
rect 29184 42026 29236 42032
rect 29472 42022 29500 42094
rect 29460 42016 29512 42022
rect 29460 41958 29512 41964
rect 29276 41676 29328 41682
rect 29276 41618 29328 41624
rect 29288 40934 29316 41618
rect 29472 41274 29500 41958
rect 29564 41682 29592 42706
rect 29644 42696 29696 42702
rect 29644 42638 29696 42644
rect 29656 42226 29684 42638
rect 30300 42226 30328 43823
rect 30380 43648 30432 43654
rect 30380 43590 30432 43596
rect 30392 42838 30420 43590
rect 30472 43444 30524 43450
rect 30472 43386 30524 43392
rect 30484 43081 30512 43386
rect 30564 43376 30616 43382
rect 30564 43318 30616 43324
rect 30470 43072 30526 43081
rect 30470 43007 30526 43016
rect 30380 42832 30432 42838
rect 30380 42774 30432 42780
rect 30392 42294 30420 42774
rect 30380 42288 30432 42294
rect 30380 42230 30432 42236
rect 29644 42220 29696 42226
rect 29644 42162 29696 42168
rect 30288 42220 30340 42226
rect 30288 42162 30340 42168
rect 29656 41818 29684 42162
rect 29644 41812 29696 41818
rect 29644 41754 29696 41760
rect 29552 41676 29604 41682
rect 29552 41618 29604 41624
rect 29460 41268 29512 41274
rect 29460 41210 29512 41216
rect 29564 40934 29592 41618
rect 30576 41614 30604 43318
rect 30760 42158 30788 44270
rect 31024 44192 31076 44198
rect 31024 44134 31076 44140
rect 31036 43994 31064 44134
rect 31024 43988 31076 43994
rect 31024 43930 31076 43936
rect 30840 43852 30892 43858
rect 30840 43794 30892 43800
rect 30852 43450 30880 43794
rect 31208 43716 31260 43722
rect 31208 43658 31260 43664
rect 31024 43648 31076 43654
rect 31024 43590 31076 43596
rect 30840 43444 30892 43450
rect 30840 43386 30892 43392
rect 30748 42152 30800 42158
rect 30748 42094 30800 42100
rect 30656 41744 30708 41750
rect 30656 41686 30708 41692
rect 30104 41608 30156 41614
rect 30104 41550 30156 41556
rect 30564 41608 30616 41614
rect 30564 41550 30616 41556
rect 30116 41138 30144 41550
rect 30576 41206 30604 41550
rect 30668 41274 30696 41686
rect 30656 41268 30708 41274
rect 30656 41210 30708 41216
rect 30564 41200 30616 41206
rect 30564 41142 30616 41148
rect 30104 41132 30156 41138
rect 30104 41074 30156 41080
rect 30472 40996 30524 41002
rect 30472 40938 30524 40944
rect 29276 40928 29328 40934
rect 29276 40870 29328 40876
rect 29552 40928 29604 40934
rect 29552 40870 29604 40876
rect 27620 40588 27672 40594
rect 27620 40530 27672 40536
rect 27988 40588 28040 40594
rect 27988 40530 28040 40536
rect 28724 40588 28776 40594
rect 28724 40530 28776 40536
rect 27344 40384 27396 40390
rect 27344 40326 27396 40332
rect 27356 39846 27384 40326
rect 27632 39914 27660 40530
rect 28000 39982 28028 40530
rect 27988 39976 28040 39982
rect 27988 39918 28040 39924
rect 27620 39908 27672 39914
rect 27620 39850 27672 39856
rect 27344 39840 27396 39846
rect 27344 39782 27396 39788
rect 28000 39642 28028 39918
rect 28736 39846 28764 40530
rect 29288 40458 29316 40870
rect 29276 40452 29328 40458
rect 29276 40394 29328 40400
rect 29288 40050 29316 40394
rect 29564 40390 29592 40870
rect 30484 40662 30512 40938
rect 30576 40730 30604 41142
rect 30564 40724 30616 40730
rect 30564 40666 30616 40672
rect 30472 40656 30524 40662
rect 30472 40598 30524 40604
rect 30012 40520 30064 40526
rect 30012 40462 30064 40468
rect 29552 40384 29604 40390
rect 29552 40326 29604 40332
rect 29276 40044 29328 40050
rect 29276 39986 29328 39992
rect 29564 39982 29592 40326
rect 30024 40050 30052 40462
rect 30012 40044 30064 40050
rect 30012 39986 30064 39992
rect 29552 39976 29604 39982
rect 29552 39918 29604 39924
rect 28724 39840 28776 39846
rect 28724 39782 28776 39788
rect 29460 39840 29512 39846
rect 29460 39782 29512 39788
rect 27988 39636 28040 39642
rect 27988 39578 28040 39584
rect 28172 39636 28224 39642
rect 28172 39578 28224 39584
rect 26884 39432 26936 39438
rect 26884 39374 26936 39380
rect 27252 38752 27304 38758
rect 27252 38694 27304 38700
rect 27264 37670 27292 38694
rect 28000 38554 28028 39578
rect 28184 38962 28212 39578
rect 28356 39500 28408 39506
rect 28356 39442 28408 39448
rect 28172 38956 28224 38962
rect 28172 38898 28224 38904
rect 28368 38758 28396 39442
rect 28356 38752 28408 38758
rect 28356 38694 28408 38700
rect 27988 38548 28040 38554
rect 27988 38490 28040 38496
rect 27252 37664 27304 37670
rect 27252 37606 27304 37612
rect 28000 37330 28028 38490
rect 27988 37324 28040 37330
rect 27988 37266 28040 37272
rect 28356 37324 28408 37330
rect 28356 37266 28408 37272
rect 28000 36922 28028 37266
rect 27988 36916 28040 36922
rect 27988 36858 28040 36864
rect 26792 36712 26844 36718
rect 26792 36654 26844 36660
rect 27620 36712 27672 36718
rect 27620 36654 27672 36660
rect 26424 36304 26476 36310
rect 26424 36246 26476 36252
rect 26332 35556 26384 35562
rect 26332 35498 26384 35504
rect 25780 35012 25832 35018
rect 25780 34954 25832 34960
rect 25596 34400 25648 34406
rect 25596 34342 25648 34348
rect 24676 34060 24728 34066
rect 24676 34002 24728 34008
rect 25412 34060 25464 34066
rect 25412 34002 25464 34008
rect 24688 33658 24716 34002
rect 25424 33658 25452 34002
rect 25608 33833 25636 34342
rect 25594 33824 25650 33833
rect 25594 33759 25650 33768
rect 24676 33652 24728 33658
rect 24676 33594 24728 33600
rect 25412 33652 25464 33658
rect 25412 33594 25464 33600
rect 25424 33134 25452 33594
rect 25502 33144 25558 33153
rect 25424 33106 25502 33134
rect 25502 33079 25558 33088
rect 25608 32978 25636 33759
rect 25792 33425 25820 34954
rect 26344 34950 26372 35498
rect 26436 35494 26464 36246
rect 26424 35488 26476 35494
rect 26424 35430 26476 35436
rect 26436 35222 26464 35430
rect 26424 35216 26476 35222
rect 26424 35158 26476 35164
rect 26332 34944 26384 34950
rect 26332 34886 26384 34892
rect 26146 34640 26202 34649
rect 25872 34604 25924 34610
rect 26146 34575 26202 34584
rect 25872 34546 25924 34552
rect 25884 34202 25912 34546
rect 26160 34542 26188 34575
rect 26148 34536 26200 34542
rect 26148 34478 26200 34484
rect 25872 34196 25924 34202
rect 25872 34138 25924 34144
rect 26056 33448 26108 33454
rect 25778 33416 25834 33425
rect 26056 33390 26108 33396
rect 25778 33351 25834 33360
rect 25964 33380 26016 33386
rect 25596 32972 25648 32978
rect 25596 32914 25648 32920
rect 25228 32768 25280 32774
rect 25228 32710 25280 32716
rect 25240 32366 25268 32710
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 24492 32020 24544 32026
rect 24492 31962 24544 31968
rect 24504 31822 24532 31962
rect 24584 31952 24636 31958
rect 24584 31894 24636 31900
rect 24492 31816 24544 31822
rect 24492 31758 24544 31764
rect 24400 31476 24452 31482
rect 24400 31418 24452 31424
rect 24412 30802 24440 31418
rect 24504 30938 24532 31758
rect 24596 31482 24624 31894
rect 24584 31476 24636 31482
rect 24584 31418 24636 31424
rect 25240 31346 25268 32302
rect 25608 31686 25636 32914
rect 25596 31680 25648 31686
rect 25596 31622 25648 31628
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 24584 31272 24636 31278
rect 24584 31214 24636 31220
rect 24492 30932 24544 30938
rect 24492 30874 24544 30880
rect 24400 30796 24452 30802
rect 24400 30738 24452 30744
rect 24596 30598 24624 31214
rect 24584 30592 24636 30598
rect 24584 30534 24636 30540
rect 24596 29306 24624 30534
rect 24860 29776 24912 29782
rect 24860 29718 24912 29724
rect 24872 29306 24900 29718
rect 25504 29504 25556 29510
rect 25504 29446 25556 29452
rect 24584 29300 24636 29306
rect 24584 29242 24636 29248
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 25516 29170 25544 29446
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 24136 28966 24348 28994
rect 24136 27962 24164 28966
rect 25412 28960 25464 28966
rect 25412 28902 25464 28908
rect 25226 28656 25282 28665
rect 25424 28626 25452 28902
rect 25226 28591 25282 28600
rect 25412 28620 25464 28626
rect 25240 28558 25268 28591
rect 25412 28562 25464 28568
rect 25228 28552 25280 28558
rect 25148 28512 25228 28540
rect 24216 28416 24268 28422
rect 24216 28358 24268 28364
rect 23952 27934 24164 27962
rect 23664 27668 23716 27674
rect 23664 27610 23716 27616
rect 23676 26994 23704 27610
rect 23952 27062 23980 27934
rect 24124 27872 24176 27878
rect 24124 27814 24176 27820
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 23940 27056 23992 27062
rect 23940 26998 23992 27004
rect 23664 26988 23716 26994
rect 23664 26930 23716 26936
rect 23664 26852 23716 26858
rect 23664 26794 23716 26800
rect 23572 25356 23624 25362
rect 23572 25298 23624 25304
rect 23584 24954 23612 25298
rect 23572 24948 23624 24954
rect 23572 24890 23624 24896
rect 23478 24848 23534 24857
rect 23478 24783 23534 24792
rect 23676 23474 23704 26794
rect 23952 26625 23980 26998
rect 23938 26616 23994 26625
rect 24044 26586 24072 27406
rect 23938 26551 23994 26560
rect 24032 26580 24084 26586
rect 24032 26522 24084 26528
rect 24032 25696 24084 25702
rect 24032 25638 24084 25644
rect 24044 25430 24072 25638
rect 24032 25424 24084 25430
rect 24032 25366 24084 25372
rect 23848 24676 23900 24682
rect 23848 24618 23900 24624
rect 23860 24342 23888 24618
rect 24136 24410 24164 27814
rect 24228 25770 24256 28358
rect 25148 28150 25176 28512
rect 25228 28494 25280 28500
rect 25424 28150 25452 28562
rect 25136 28144 25188 28150
rect 25042 28112 25098 28121
rect 25136 28086 25188 28092
rect 25412 28144 25464 28150
rect 25412 28086 25464 28092
rect 25042 28047 25098 28056
rect 25228 28076 25280 28082
rect 25056 28014 25084 28047
rect 25228 28018 25280 28024
rect 25044 28008 25096 28014
rect 25044 27950 25096 27956
rect 25056 27674 25084 27950
rect 25044 27668 25096 27674
rect 25044 27610 25096 27616
rect 24492 27600 24544 27606
rect 24492 27542 24544 27548
rect 24308 27464 24360 27470
rect 24308 27406 24360 27412
rect 24216 25764 24268 25770
rect 24216 25706 24268 25712
rect 24228 25498 24256 25706
rect 24216 25492 24268 25498
rect 24216 25434 24268 25440
rect 24320 25430 24348 27406
rect 24400 27396 24452 27402
rect 24400 27338 24452 27344
rect 24308 25424 24360 25430
rect 24308 25366 24360 25372
rect 24320 24886 24348 25366
rect 24308 24880 24360 24886
rect 24308 24822 24360 24828
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 23848 24336 23900 24342
rect 23848 24278 23900 24284
rect 23860 24070 23888 24278
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23860 23526 23888 24006
rect 23492 23446 23704 23474
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 24412 23474 24440 27338
rect 24504 27130 24532 27542
rect 24492 27124 24544 27130
rect 24492 27066 24544 27072
rect 24504 26586 24532 27066
rect 24860 27056 24912 27062
rect 24860 26998 24912 27004
rect 24492 26580 24544 26586
rect 24492 26522 24544 26528
rect 24504 26042 24532 26522
rect 24492 26036 24544 26042
rect 24492 25978 24544 25984
rect 24504 25770 24532 25978
rect 24676 25968 24728 25974
rect 24676 25910 24728 25916
rect 24492 25764 24544 25770
rect 24492 25706 24544 25712
rect 24504 25430 24532 25706
rect 24492 25424 24544 25430
rect 24492 25366 24544 25372
rect 24504 24954 24532 25366
rect 24492 24948 24544 24954
rect 24492 24890 24544 24896
rect 23296 23248 23348 23254
rect 23296 23190 23348 23196
rect 23072 23072 23244 23100
rect 23020 23054 23072 23060
rect 23032 22778 23060 23054
rect 23020 22772 23072 22778
rect 23020 22714 23072 22720
rect 23308 22710 23336 23190
rect 23296 22704 23348 22710
rect 23296 22646 23348 22652
rect 22928 22500 22980 22506
rect 22928 22442 22980 22448
rect 22940 22030 22968 22442
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 22940 21146 22968 21966
rect 23308 21690 23336 22646
rect 23492 22234 23520 23446
rect 23860 23254 23888 23462
rect 24412 23446 24624 23474
rect 23848 23248 23900 23254
rect 23848 23190 23900 23196
rect 24596 23118 24624 23446
rect 24584 23112 24636 23118
rect 24688 23089 24716 25910
rect 24872 25226 24900 26998
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 24860 25220 24912 25226
rect 24860 25162 24912 25168
rect 24952 25220 25004 25226
rect 24952 25162 25004 25168
rect 24860 24880 24912 24886
rect 24860 24822 24912 24828
rect 24768 24336 24820 24342
rect 24768 24278 24820 24284
rect 24780 23594 24808 24278
rect 24768 23588 24820 23594
rect 24768 23530 24820 23536
rect 24780 23254 24808 23530
rect 24768 23248 24820 23254
rect 24768 23190 24820 23196
rect 24584 23054 24636 23060
rect 24674 23080 24730 23089
rect 24596 22778 24624 23054
rect 24674 23015 24730 23024
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24688 22574 24716 23015
rect 24780 22642 24808 23190
rect 24872 23118 24900 24822
rect 24964 24206 24992 25162
rect 25056 24954 25084 25230
rect 25044 24948 25096 24954
rect 25044 24890 25096 24896
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 25148 23798 25176 26250
rect 25240 25974 25268 28018
rect 25424 27674 25452 28086
rect 25516 28082 25544 29106
rect 25504 28076 25556 28082
rect 25504 28018 25556 28024
rect 25608 27878 25636 31622
rect 25792 30190 25820 33351
rect 25964 33322 26016 33328
rect 25976 32570 26004 33322
rect 25964 32564 26016 32570
rect 25964 32506 26016 32512
rect 25976 31482 26004 32506
rect 26068 32473 26096 33390
rect 26146 33144 26202 33153
rect 26146 33079 26202 33088
rect 26054 32464 26110 32473
rect 26054 32399 26110 32408
rect 25964 31476 26016 31482
rect 25964 31418 26016 31424
rect 25976 31210 26004 31418
rect 25964 31204 26016 31210
rect 25964 31146 26016 31152
rect 25780 30184 25832 30190
rect 25780 30126 25832 30132
rect 25780 30048 25832 30054
rect 25780 29990 25832 29996
rect 26056 30048 26108 30054
rect 26056 29990 26108 29996
rect 25792 29782 25820 29990
rect 25780 29776 25832 29782
rect 25780 29718 25832 29724
rect 25872 29164 25924 29170
rect 25872 29106 25924 29112
rect 25596 27872 25648 27878
rect 25596 27814 25648 27820
rect 25412 27668 25464 27674
rect 25412 27610 25464 27616
rect 25596 27328 25648 27334
rect 25596 27270 25648 27276
rect 25608 26382 25636 27270
rect 25780 26852 25832 26858
rect 25780 26794 25832 26800
rect 25792 26518 25820 26794
rect 25780 26512 25832 26518
rect 25780 26454 25832 26460
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25608 26042 25636 26318
rect 25596 26036 25648 26042
rect 25596 25978 25648 25984
rect 25228 25968 25280 25974
rect 25228 25910 25280 25916
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25148 23474 25176 23734
rect 25148 23446 25268 23474
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 25240 23050 25268 23446
rect 25228 23044 25280 23050
rect 25228 22986 25280 22992
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24676 22568 24728 22574
rect 24676 22510 24728 22516
rect 23848 22432 23900 22438
rect 23848 22374 23900 22380
rect 23860 22273 23888 22374
rect 23846 22264 23902 22273
rect 23480 22228 23532 22234
rect 24780 22234 24808 22578
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 23846 22199 23902 22208
rect 24768 22228 24820 22234
rect 23480 22170 23532 22176
rect 24768 22170 24820 22176
rect 23296 21684 23348 21690
rect 23296 21626 23348 21632
rect 23308 21418 23336 21626
rect 23492 21486 23520 22170
rect 25792 22166 25820 22374
rect 25780 22160 25832 22166
rect 25780 22102 25832 22108
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23296 21412 23348 21418
rect 23296 21354 23348 21360
rect 23756 21412 23808 21418
rect 23756 21354 23808 21360
rect 24216 21412 24268 21418
rect 24216 21354 24268 21360
rect 23768 21146 23796 21354
rect 22928 21140 22980 21146
rect 22928 21082 22980 21088
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 21916 21004 21968 21010
rect 21916 20946 21968 20952
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 23204 21004 23256 21010
rect 23204 20946 23256 20952
rect 21928 20534 21956 20946
rect 22112 20874 22140 20946
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 22112 20602 22140 20810
rect 23216 20602 23244 20946
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 23204 20596 23256 20602
rect 23204 20538 23256 20544
rect 21916 20528 21968 20534
rect 21916 20470 21968 20476
rect 24228 20466 24256 21354
rect 24780 21146 24808 21966
rect 25056 21554 25084 21966
rect 25504 21888 25556 21894
rect 25504 21830 25556 21836
rect 25516 21690 25544 21830
rect 25504 21684 25556 21690
rect 25504 21626 25556 21632
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25148 21350 25176 21422
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 25148 20942 25176 21286
rect 25412 21004 25464 21010
rect 25412 20946 25464 20952
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 24308 20868 24360 20874
rect 24308 20810 24360 20816
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 23020 20392 23072 20398
rect 23020 20334 23072 20340
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22664 19961 22692 20198
rect 22650 19952 22706 19961
rect 22650 19887 22706 19896
rect 22664 19854 22692 19887
rect 22652 19848 22704 19854
rect 22652 19790 22704 19796
rect 22664 19514 22692 19790
rect 22652 19508 22704 19514
rect 22652 19450 22704 19456
rect 21548 19372 21600 19378
rect 21548 19314 21600 19320
rect 21560 18902 21588 19314
rect 23032 18902 23060 20334
rect 23204 19916 23256 19922
rect 23124 19876 23204 19904
rect 23124 19174 23152 19876
rect 23204 19858 23256 19864
rect 24320 19718 24348 20810
rect 25148 20262 25176 20878
rect 25424 20330 25452 20946
rect 25516 20806 25544 21626
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25608 20942 25636 21490
rect 25884 21078 25912 29106
rect 25964 27396 26016 27402
rect 25964 27338 26016 27344
rect 25976 21690 26004 27338
rect 26068 26926 26096 29990
rect 26160 27538 26188 33079
rect 26240 32972 26292 32978
rect 26240 32914 26292 32920
rect 26252 32570 26280 32914
rect 26344 32910 26372 34886
rect 26436 34406 26464 35158
rect 26608 35080 26660 35086
rect 26608 35022 26660 35028
rect 26620 34678 26648 35022
rect 26608 34672 26660 34678
rect 26608 34614 26660 34620
rect 26424 34400 26476 34406
rect 26424 34342 26476 34348
rect 26332 32904 26384 32910
rect 26332 32846 26384 32852
rect 26240 32564 26292 32570
rect 26240 32506 26292 32512
rect 26240 31748 26292 31754
rect 26240 31690 26292 31696
rect 26252 30802 26280 31690
rect 26240 30796 26292 30802
rect 26240 30738 26292 30744
rect 26252 30326 26280 30738
rect 26240 30320 26292 30326
rect 26240 30262 26292 30268
rect 26332 30252 26384 30258
rect 26332 30194 26384 30200
rect 26344 29850 26372 30194
rect 26436 30104 26464 34342
rect 26620 34202 26648 34614
rect 26804 34202 26832 36654
rect 27632 36378 27660 36654
rect 28368 36582 28396 37266
rect 28540 36644 28592 36650
rect 28540 36586 28592 36592
rect 27896 36576 27948 36582
rect 28356 36576 28408 36582
rect 27896 36518 27948 36524
rect 28078 36544 28134 36553
rect 27620 36372 27672 36378
rect 27620 36314 27672 36320
rect 27528 36168 27580 36174
rect 27528 36110 27580 36116
rect 27252 36100 27304 36106
rect 27252 36042 27304 36048
rect 26884 35692 26936 35698
rect 26884 35634 26936 35640
rect 26976 35692 27028 35698
rect 26976 35634 27028 35640
rect 26896 35086 26924 35634
rect 26988 35290 27016 35634
rect 26976 35284 27028 35290
rect 27028 35244 27108 35272
rect 26976 35226 27028 35232
rect 26884 35080 26936 35086
rect 26936 35040 27016 35068
rect 26884 35022 26936 35028
rect 26884 34468 26936 34474
rect 26884 34410 26936 34416
rect 26608 34196 26660 34202
rect 26608 34138 26660 34144
rect 26792 34196 26844 34202
rect 26792 34138 26844 34144
rect 26896 34134 26924 34410
rect 26884 34128 26936 34134
rect 26884 34070 26936 34076
rect 26792 33992 26844 33998
rect 26792 33934 26844 33940
rect 26804 33114 26832 33934
rect 26896 33386 26924 34070
rect 26988 33590 27016 35040
rect 27080 33998 27108 35244
rect 27264 34678 27292 36042
rect 27540 35494 27568 36110
rect 27528 35488 27580 35494
rect 27528 35430 27580 35436
rect 27252 34672 27304 34678
rect 27252 34614 27304 34620
rect 27068 33992 27120 33998
rect 27068 33934 27120 33940
rect 26976 33584 27028 33590
rect 26976 33526 27028 33532
rect 26884 33380 26936 33386
rect 26884 33322 26936 33328
rect 26792 33108 26844 33114
rect 26792 33050 26844 33056
rect 26700 32836 26752 32842
rect 26700 32778 26752 32784
rect 26516 32768 26568 32774
rect 26516 32710 26568 32716
rect 26608 32768 26660 32774
rect 26608 32710 26660 32716
rect 26528 32434 26556 32710
rect 26516 32428 26568 32434
rect 26516 32370 26568 32376
rect 26620 31822 26648 32710
rect 26712 32298 26740 32778
rect 26988 32502 27016 33526
rect 27080 33134 27108 33934
rect 27540 33658 27568 35430
rect 27528 33652 27580 33658
rect 27528 33594 27580 33600
rect 27712 33380 27764 33386
rect 27712 33322 27764 33328
rect 27080 33106 27292 33134
rect 27724 33114 27752 33322
rect 26976 32496 27028 32502
rect 26976 32438 27028 32444
rect 26700 32292 26752 32298
rect 26700 32234 26752 32240
rect 26712 31958 26740 32234
rect 26700 31952 26752 31958
rect 26700 31894 26752 31900
rect 26608 31816 26660 31822
rect 26608 31758 26660 31764
rect 26620 31482 26648 31758
rect 26608 31476 26660 31482
rect 26608 31418 26660 31424
rect 26712 31142 26740 31894
rect 26884 31816 26936 31822
rect 26884 31758 26936 31764
rect 26896 31346 26924 31758
rect 26884 31340 26936 31346
rect 26884 31282 26936 31288
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 26700 31136 26752 31142
rect 26700 31078 26752 31084
rect 26712 30870 26740 31078
rect 26700 30864 26752 30870
rect 26700 30806 26752 30812
rect 26516 30116 26568 30122
rect 26436 30076 26516 30104
rect 26332 29844 26384 29850
rect 26332 29786 26384 29792
rect 26240 29776 26292 29782
rect 26240 29718 26292 29724
rect 26252 28762 26280 29718
rect 26436 29306 26464 30076
rect 26516 30058 26568 30064
rect 26712 29782 26740 30806
rect 27172 30326 27200 31282
rect 27264 30870 27292 33106
rect 27712 33108 27764 33114
rect 27712 33050 27764 33056
rect 27802 33008 27858 33017
rect 27802 32943 27858 32952
rect 27712 32564 27764 32570
rect 27712 32506 27764 32512
rect 27528 32428 27580 32434
rect 27528 32370 27580 32376
rect 27540 32026 27568 32370
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 27252 30864 27304 30870
rect 27252 30806 27304 30812
rect 27264 30394 27292 30806
rect 27252 30388 27304 30394
rect 27252 30330 27304 30336
rect 27160 30320 27212 30326
rect 27160 30262 27212 30268
rect 26700 29776 26752 29782
rect 26700 29718 26752 29724
rect 26712 29306 26740 29718
rect 27172 29578 27200 30262
rect 27160 29572 27212 29578
rect 27160 29514 27212 29520
rect 26424 29300 26476 29306
rect 26424 29242 26476 29248
rect 26700 29300 26752 29306
rect 26700 29242 26752 29248
rect 27160 29096 27212 29102
rect 27160 29038 27212 29044
rect 26606 28792 26662 28801
rect 26240 28756 26292 28762
rect 26606 28727 26662 28736
rect 26240 28698 26292 28704
rect 26514 28656 26570 28665
rect 26514 28591 26570 28600
rect 26148 27532 26200 27538
rect 26148 27474 26200 27480
rect 26056 26920 26108 26926
rect 26056 26862 26108 26868
rect 26240 26920 26292 26926
rect 26240 26862 26292 26868
rect 26068 24750 26096 26862
rect 26056 24744 26108 24750
rect 26056 24686 26108 24692
rect 26252 22778 26280 26862
rect 26528 24274 26556 28591
rect 26620 26926 26648 28727
rect 27172 28694 27200 29038
rect 27160 28688 27212 28694
rect 27160 28630 27212 28636
rect 27528 28620 27580 28626
rect 27528 28562 27580 28568
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27172 28393 27200 28494
rect 27158 28384 27214 28393
rect 27158 28319 27214 28328
rect 27172 28218 27200 28319
rect 27540 28218 27568 28562
rect 27160 28212 27212 28218
rect 27160 28154 27212 28160
rect 27252 28212 27304 28218
rect 27252 28154 27304 28160
rect 27528 28212 27580 28218
rect 27528 28154 27580 28160
rect 26976 27124 27028 27130
rect 26976 27066 27028 27072
rect 26884 26988 26936 26994
rect 26884 26930 26936 26936
rect 26608 26920 26660 26926
rect 26608 26862 26660 26868
rect 26792 26920 26844 26926
rect 26792 26862 26844 26868
rect 26608 25968 26660 25974
rect 26608 25910 26660 25916
rect 26620 25838 26648 25910
rect 26804 25838 26832 26862
rect 26896 26382 26924 26930
rect 26884 26376 26936 26382
rect 26884 26318 26936 26324
rect 26896 26042 26924 26318
rect 26884 26036 26936 26042
rect 26884 25978 26936 25984
rect 26608 25832 26660 25838
rect 26608 25774 26660 25780
rect 26792 25832 26844 25838
rect 26792 25774 26844 25780
rect 26606 24712 26662 24721
rect 26606 24647 26662 24656
rect 26620 24614 26648 24647
rect 26608 24608 26660 24614
rect 26608 24550 26660 24556
rect 26516 24268 26568 24274
rect 26516 24210 26568 24216
rect 26528 23798 26556 24210
rect 26700 24064 26752 24070
rect 26700 24006 26752 24012
rect 26516 23792 26568 23798
rect 26516 23734 26568 23740
rect 26528 23474 26556 23734
rect 26436 23446 26556 23474
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 26252 22574 26280 22714
rect 26436 22710 26464 23446
rect 26608 23180 26660 23186
rect 26608 23122 26660 23128
rect 26620 22778 26648 23122
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 26712 22710 26740 24006
rect 26988 23474 27016 27066
rect 27160 25764 27212 25770
rect 27160 25706 27212 25712
rect 27172 25498 27200 25706
rect 27160 25492 27212 25498
rect 27160 25434 27212 25440
rect 27068 24064 27120 24070
rect 27068 24006 27120 24012
rect 27080 23662 27108 24006
rect 27068 23656 27120 23662
rect 27068 23598 27120 23604
rect 26988 23446 27108 23474
rect 27080 23186 27108 23446
rect 27068 23180 27120 23186
rect 27068 23122 27120 23128
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 26424 22704 26476 22710
rect 26424 22646 26476 22652
rect 26700 22704 26752 22710
rect 26700 22646 26752 22652
rect 27172 22574 27200 22918
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26792 22568 26844 22574
rect 26792 22510 26844 22516
rect 27160 22568 27212 22574
rect 27160 22510 27212 22516
rect 26804 22234 26832 22510
rect 26792 22228 26844 22234
rect 26792 22170 26844 22176
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 26988 21690 27016 22034
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 26976 21684 27028 21690
rect 26976 21626 27028 21632
rect 26516 21412 26568 21418
rect 26516 21354 26568 21360
rect 25872 21072 25924 21078
rect 25872 21014 25924 21020
rect 26528 21010 26556 21354
rect 26516 21004 26568 21010
rect 26516 20946 26568 20952
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25504 20800 25556 20806
rect 25504 20742 25556 20748
rect 25872 20800 25924 20806
rect 25872 20742 25924 20748
rect 25412 20324 25464 20330
rect 25412 20266 25464 20272
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24320 19417 24348 19654
rect 24306 19408 24362 19417
rect 24216 19372 24268 19378
rect 24306 19343 24362 19352
rect 24216 19314 24268 19320
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 21548 18896 21600 18902
rect 21548 18838 21600 18844
rect 23020 18896 23072 18902
rect 23020 18838 23072 18844
rect 21732 18828 21784 18834
rect 21732 18770 21784 18776
rect 21744 18290 21772 18770
rect 23020 18760 23072 18766
rect 23124 18748 23152 19110
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23072 18720 23152 18748
rect 23020 18702 23072 18708
rect 21732 18284 21784 18290
rect 21732 18226 21784 18232
rect 21744 18193 21772 18226
rect 21730 18184 21786 18193
rect 21730 18119 21786 18128
rect 23032 18086 23060 18702
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 23020 18080 23072 18086
rect 23020 18022 23072 18028
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 21454 17912 21510 17921
rect 21454 17847 21510 17856
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17270 21036 17614
rect 21100 17338 21128 17750
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 21100 16794 21128 17274
rect 21192 17202 21220 17614
rect 22020 17542 22048 18022
rect 22008 17536 22060 17542
rect 22006 17504 22008 17513
rect 22060 17504 22062 17513
rect 22006 17439 22062 17448
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 21100 16250 21128 16594
rect 21192 16590 21220 17138
rect 22112 16658 22140 18022
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22756 16794 22784 17274
rect 22834 17232 22890 17241
rect 22834 17167 22890 17176
rect 22848 17134 22876 17167
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19904 15638 19932 15982
rect 22112 15978 22140 16390
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 19892 15632 19944 15638
rect 19892 15574 19944 15580
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19352 15026 19380 15506
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19904 14550 19932 14894
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 13394 19472 13806
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19260 12782 19288 13330
rect 19444 12986 19472 13330
rect 20088 12986 20116 14826
rect 20180 14482 20208 15846
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20824 14550 20852 14758
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20180 14074 20208 14418
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 20088 12714 20116 12922
rect 20180 12850 20208 13262
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20076 12708 20128 12714
rect 20076 12650 20128 12656
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 20088 11898 20116 12650
rect 20272 12374 20300 13738
rect 20364 13734 20392 14350
rect 20824 14074 20852 14486
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20916 14006 20944 15914
rect 22572 15706 22600 16526
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 21744 14822 21772 15506
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 22388 14550 22416 15302
rect 22756 15162 22784 15438
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22926 15056 22982 15065
rect 22926 14991 22982 15000
rect 22940 14958 22968 14991
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 23032 14618 23060 18022
rect 23110 17912 23166 17921
rect 23110 17847 23166 17856
rect 23020 14612 23072 14618
rect 23020 14554 23072 14560
rect 22376 14544 22428 14550
rect 22376 14486 22428 14492
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21086 14240 21142 14249
rect 21086 14175 21142 14184
rect 21100 14006 21128 14175
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20364 12442 20392 13670
rect 21468 13530 21496 13806
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21192 12918 21220 13398
rect 21560 13326 21588 14282
rect 22388 14074 22416 14486
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22848 14006 22876 14486
rect 23124 14074 23152 17847
rect 23216 17814 23244 18022
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23216 17542 23244 17750
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23216 17338 23244 17478
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23492 17105 23520 18226
rect 23676 18154 23704 18770
rect 24228 18766 24256 19314
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24216 18760 24268 18766
rect 24044 18720 24216 18748
rect 23756 18624 23808 18630
rect 23756 18566 23808 18572
rect 23768 18358 23796 18566
rect 23756 18352 23808 18358
rect 23756 18294 23808 18300
rect 23664 18148 23716 18154
rect 23664 18090 23716 18096
rect 24044 17678 24072 18720
rect 24216 18702 24268 18708
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 24032 17672 24084 17678
rect 24032 17614 24084 17620
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23952 17270 23980 17478
rect 24320 17377 24348 18566
rect 24412 18290 24440 19110
rect 24490 18864 24546 18873
rect 24490 18799 24546 18808
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24306 17368 24362 17377
rect 24306 17303 24362 17312
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 24504 17134 24532 18799
rect 25148 18630 25176 20198
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25332 19174 25360 19858
rect 25424 19718 25452 20266
rect 25516 19990 25544 20742
rect 25884 20466 25912 20742
rect 26528 20602 26556 20946
rect 27068 20868 27120 20874
rect 27068 20810 27120 20816
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 26792 20800 26844 20806
rect 26792 20742 26844 20748
rect 26516 20596 26568 20602
rect 26516 20538 26568 20544
rect 25872 20460 25924 20466
rect 25872 20402 25924 20408
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 25504 19984 25556 19990
rect 25504 19926 25556 19932
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 24768 18352 24820 18358
rect 24768 18294 24820 18300
rect 24780 18086 24808 18294
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 25056 18086 25084 18226
rect 25148 18154 25176 18566
rect 25332 18358 25360 19110
rect 25424 18834 25452 19654
rect 26148 19236 26200 19242
rect 26148 19178 26200 19184
rect 25412 18828 25464 18834
rect 25412 18770 25464 18776
rect 25320 18352 25372 18358
rect 25320 18294 25372 18300
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25136 18148 25188 18154
rect 25136 18090 25188 18096
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 24780 17814 24808 18022
rect 24768 17808 24820 17814
rect 24768 17750 24820 17756
rect 24780 17270 24808 17750
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24492 17128 24544 17134
rect 23478 17096 23534 17105
rect 24492 17070 24544 17076
rect 23478 17031 23534 17040
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 24308 17060 24360 17066
rect 24308 17002 24360 17008
rect 23204 16720 23256 16726
rect 23204 16662 23256 16668
rect 23216 16250 23244 16662
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 23216 15638 23244 16186
rect 23584 16182 23612 16458
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 23204 15632 23256 15638
rect 23256 15592 23336 15620
rect 23204 15574 23256 15580
rect 23308 15026 23336 15592
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23204 14952 23256 14958
rect 23204 14894 23256 14900
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 23124 13870 23152 14010
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 23112 13728 23164 13734
rect 23216 13705 23244 14894
rect 23308 14890 23336 14962
rect 23296 14884 23348 14890
rect 23296 14826 23348 14832
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23112 13670 23164 13676
rect 23202 13696 23258 13705
rect 22388 13326 22416 13670
rect 23124 13530 23152 13670
rect 23202 13631 23258 13640
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 21376 12986 21404 13262
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21180 12912 21232 12918
rect 21180 12854 21232 12860
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18800 10810 18828 11154
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18708 8634 18736 8978
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18788 8016 18840 8022
rect 18788 7958 18840 7964
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 7206 18092 7278
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 18064 6458 18092 7142
rect 18524 7002 18552 7822
rect 18800 7274 18828 7958
rect 18892 7410 18920 11494
rect 19076 11478 19196 11506
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19076 10266 19104 11290
rect 19168 11286 19196 11478
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19352 10198 19380 11834
rect 20088 11558 20116 11834
rect 20272 11762 20300 12310
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 21008 11558 21036 12174
rect 21100 11898 21128 12310
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21376 11762 21404 12922
rect 21560 12170 21588 13262
rect 22388 12986 22416 13262
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 23112 12640 23164 12646
rect 23112 12582 23164 12588
rect 22848 12374 22876 12582
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21560 11694 21588 12106
rect 21548 11688 21600 11694
rect 21548 11630 21600 11636
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19444 10606 19472 11154
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19996 10606 20024 10950
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19168 9722 19196 10134
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 19444 9042 19472 10542
rect 20076 10532 20128 10538
rect 20076 10474 20128 10480
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19984 10192 20036 10198
rect 19984 10134 20036 10140
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19904 9110 19932 9454
rect 19996 9382 20024 10134
rect 20088 10062 20116 10474
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19892 9104 19944 9110
rect 19892 9046 19944 9052
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19246 8936 19302 8945
rect 19302 8894 19380 8922
rect 19246 8871 19302 8880
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18800 6934 18828 7210
rect 18892 7002 18920 7346
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18788 6928 18840 6934
rect 18788 6870 18840 6876
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 13818 54 14136 82
rect 19352 82 19380 8894
rect 19444 8634 19472 8978
rect 20456 8634 20484 11494
rect 22848 11354 22876 12310
rect 22940 11558 22968 12378
rect 23124 12345 23152 12582
rect 23110 12336 23166 12345
rect 23110 12271 23166 12280
rect 23216 12102 23244 13631
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 22928 11552 22980 11558
rect 22928 11494 22980 11500
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22940 11218 22968 11494
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 22928 11212 22980 11218
rect 22928 11154 22980 11160
rect 21468 10810 21496 11154
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 22296 10674 22324 11086
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22940 10538 22968 11154
rect 22928 10532 22980 10538
rect 22928 10474 22980 10480
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20640 9110 20668 9318
rect 20628 9104 20680 9110
rect 20628 9046 20680 9052
rect 20640 8634 20668 9046
rect 21008 8634 21036 10406
rect 22928 10192 22980 10198
rect 22928 10134 22980 10140
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21284 9722 21312 9862
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21284 9382 21312 9658
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19628 7274 19656 7890
rect 20364 7546 20392 8366
rect 21192 8294 21220 8910
rect 21376 8362 21404 9862
rect 22480 9722 22508 9998
rect 22940 9722 22968 10134
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23032 9926 23060 9998
rect 23020 9920 23072 9926
rect 23020 9862 23072 9868
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22928 9716 22980 9722
rect 22928 9658 22980 9664
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21560 9178 21588 9522
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21836 9110 21864 9522
rect 23032 9110 23060 9862
rect 23202 9616 23258 9625
rect 23202 9551 23258 9560
rect 23216 9178 23244 9551
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 23020 9104 23072 9110
rect 23020 9046 23072 9052
rect 21836 8566 21864 9046
rect 21824 8560 21876 8566
rect 21824 8502 21876 8508
rect 21364 8356 21416 8362
rect 21364 8298 21416 8304
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21192 8090 21220 8230
rect 21376 8090 21404 8298
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 20916 7546 20944 7890
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 19616 7268 19668 7274
rect 19616 7210 19668 7216
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 23308 4185 23336 14554
rect 23400 14550 23428 15438
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 23400 11286 23428 14486
rect 23480 13456 23532 13462
rect 23480 13398 23532 13404
rect 23492 12986 23520 13398
rect 23584 13326 23612 16118
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 23848 15972 23900 15978
rect 23848 15914 23900 15920
rect 23768 15706 23796 15914
rect 23756 15700 23808 15706
rect 23756 15642 23808 15648
rect 23768 15094 23796 15642
rect 23860 15094 23888 15914
rect 24136 15638 24164 17002
rect 24320 16522 24348 17002
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 24308 16516 24360 16522
rect 24308 16458 24360 16464
rect 24504 16182 24532 16594
rect 24492 16176 24544 16182
rect 24492 16118 24544 16124
rect 24584 15972 24636 15978
rect 24584 15914 24636 15920
rect 24124 15632 24176 15638
rect 24176 15592 24256 15620
rect 24124 15574 24176 15580
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 23848 15088 23900 15094
rect 23848 15030 23900 15036
rect 23860 14074 23888 15030
rect 24032 15020 24084 15026
rect 24084 14980 24164 15008
rect 24032 14962 24084 14968
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23572 13320 23624 13326
rect 23624 13280 23704 13308
rect 23572 13262 23624 13268
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23492 12714 23520 12922
rect 23480 12708 23532 12714
rect 23480 12650 23532 12656
rect 23478 12200 23534 12209
rect 23478 12135 23534 12144
rect 23492 11812 23520 12135
rect 23572 11824 23624 11830
rect 23492 11784 23572 11812
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23400 10742 23428 11222
rect 23492 11150 23520 11784
rect 23572 11766 23624 11772
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23584 10606 23612 11222
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 23480 10532 23532 10538
rect 23480 10474 23532 10480
rect 23388 10464 23440 10470
rect 23388 10406 23440 10412
rect 23400 9586 23428 10406
rect 23492 9674 23520 10474
rect 23584 10266 23612 10542
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23676 10062 23704 13280
rect 23768 13190 23796 13466
rect 24136 13326 24164 14980
rect 24228 14618 24256 15592
rect 24596 15502 24624 15914
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24216 14612 24268 14618
rect 24216 14554 24268 14560
rect 24400 13728 24452 13734
rect 24400 13670 24452 13676
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23768 12850 23796 13126
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 23940 12708 23992 12714
rect 23940 12650 23992 12656
rect 23952 12374 23980 12650
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 23940 12368 23992 12374
rect 23940 12310 23992 12316
rect 24044 11762 24072 12378
rect 24136 11898 24164 13262
rect 24412 12374 24440 13670
rect 24596 12850 24624 15438
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 24964 14074 24992 14418
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 24952 13796 25004 13802
rect 24952 13738 25004 13744
rect 24964 13569 24992 13738
rect 24950 13560 25006 13569
rect 24950 13495 25006 13504
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24872 12850 24900 13330
rect 24584 12844 24636 12850
rect 24584 12786 24636 12792
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24596 12442 24624 12786
rect 24584 12436 24636 12442
rect 24584 12378 24636 12384
rect 24400 12368 24452 12374
rect 24400 12310 24452 12316
rect 24124 11892 24176 11898
rect 24124 11834 24176 11840
rect 24032 11756 24084 11762
rect 24032 11698 24084 11704
rect 24124 11620 24176 11626
rect 24124 11562 24176 11568
rect 24136 11082 24164 11562
rect 24412 11354 24440 12310
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23492 9646 23612 9674
rect 23676 9654 23704 9998
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23400 9178 23428 9522
rect 23584 9518 23612 9646
rect 23664 9648 23716 9654
rect 23768 9625 23796 10542
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24688 10198 24716 10406
rect 24676 10192 24728 10198
rect 24676 10134 24728 10140
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 24688 9722 24716 10134
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 23664 9590 23716 9596
rect 23754 9616 23810 9625
rect 23754 9551 23810 9560
rect 23572 9512 23624 9518
rect 23572 9454 23624 9460
rect 24872 9178 24900 9998
rect 24964 9654 24992 10134
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 23294 4176 23350 4185
rect 23294 4111 23350 4120
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19430 82 19486 480
rect 19352 54 19486 82
rect 2778 0 2834 54
rect 8298 0 8354 54
rect 13818 0 13874 54
rect 19430 0 19486 54
rect 24950 82 25006 480
rect 25056 82 25084 18022
rect 25148 17882 25176 18090
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 25240 17746 25268 18158
rect 25332 17882 25360 18294
rect 25424 17882 25452 18770
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25412 17876 25464 17882
rect 25412 17818 25464 17824
rect 25228 17740 25280 17746
rect 25228 17682 25280 17688
rect 25240 17338 25268 17682
rect 25228 17332 25280 17338
rect 25228 17274 25280 17280
rect 25884 16250 25912 18022
rect 26160 17746 26188 19178
rect 26240 18080 26292 18086
rect 26240 18022 26292 18028
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26252 17134 26280 18022
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26344 16658 26372 20198
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26436 18698 26464 19110
rect 26424 18692 26476 18698
rect 26424 18634 26476 18640
rect 26528 18426 26556 20538
rect 26620 20398 26648 20742
rect 26804 20534 26832 20742
rect 26792 20528 26844 20534
rect 26792 20470 26844 20476
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 26804 20058 26832 20470
rect 27080 20398 27108 20810
rect 27172 20602 27200 22510
rect 27160 20596 27212 20602
rect 27160 20538 27212 20544
rect 27068 20392 27120 20398
rect 27068 20334 27120 20340
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 27264 19922 27292 28154
rect 27528 28008 27580 28014
rect 27528 27950 27580 27956
rect 27344 27532 27396 27538
rect 27344 27474 27396 27480
rect 27356 26994 27384 27474
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27344 26852 27396 26858
rect 27344 26794 27396 26800
rect 27356 26518 27384 26794
rect 27344 26512 27396 26518
rect 27344 26454 27396 26460
rect 27356 25906 27384 26454
rect 27540 26314 27568 27950
rect 27620 27668 27672 27674
rect 27620 27610 27672 27616
rect 27528 26308 27580 26314
rect 27528 26250 27580 26256
rect 27344 25900 27396 25906
rect 27344 25842 27396 25848
rect 27356 25430 27384 25842
rect 27344 25424 27396 25430
rect 27344 25366 27396 25372
rect 27356 24886 27384 25366
rect 27344 24880 27396 24886
rect 27344 24822 27396 24828
rect 27356 24342 27384 24822
rect 27344 24336 27396 24342
rect 27344 24278 27396 24284
rect 27356 23798 27384 24278
rect 27344 23792 27396 23798
rect 27344 23734 27396 23740
rect 27344 23656 27396 23662
rect 27344 23598 27396 23604
rect 27356 23118 27384 23598
rect 27436 23588 27488 23594
rect 27436 23530 27488 23536
rect 27448 23186 27476 23530
rect 27632 23474 27660 27610
rect 27724 26926 27752 32506
rect 27816 28014 27844 32943
rect 27804 28008 27856 28014
rect 27804 27950 27856 27956
rect 27816 27674 27844 27950
rect 27804 27668 27856 27674
rect 27804 27610 27856 27616
rect 27712 26920 27764 26926
rect 27712 26862 27764 26868
rect 27804 26784 27856 26790
rect 27804 26726 27856 26732
rect 27712 24676 27764 24682
rect 27712 24618 27764 24624
rect 27724 24410 27752 24618
rect 27712 24404 27764 24410
rect 27712 24346 27764 24352
rect 27816 23866 27844 26726
rect 27804 23860 27856 23866
rect 27804 23802 27856 23808
rect 27540 23446 27660 23474
rect 27436 23180 27488 23186
rect 27436 23122 27488 23128
rect 27344 23112 27396 23118
rect 27344 23054 27396 23060
rect 27356 22982 27384 23054
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27540 22098 27568 23446
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27356 21049 27384 21830
rect 27540 21554 27568 21830
rect 27908 21690 27936 36518
rect 28356 36518 28408 36524
rect 28078 36479 28134 36488
rect 28092 32978 28120 36479
rect 28264 35488 28316 35494
rect 28264 35430 28316 35436
rect 28276 34105 28304 35430
rect 28262 34096 28318 34105
rect 28552 34066 28580 36586
rect 28262 34031 28318 34040
rect 28540 34060 28592 34066
rect 28080 32972 28132 32978
rect 28080 32914 28132 32920
rect 28092 32502 28120 32914
rect 28080 32496 28132 32502
rect 28080 32438 28132 32444
rect 28172 30592 28224 30598
rect 28172 30534 28224 30540
rect 28184 30122 28212 30534
rect 28276 30394 28304 34031
rect 28540 34002 28592 34008
rect 28552 33658 28580 34002
rect 28540 33652 28592 33658
rect 28540 33594 28592 33600
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28644 31686 28672 32166
rect 28632 31680 28684 31686
rect 28632 31622 28684 31628
rect 28264 30388 28316 30394
rect 28264 30330 28316 30336
rect 28276 30190 28304 30330
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 28540 30184 28592 30190
rect 28540 30126 28592 30132
rect 28172 30116 28224 30122
rect 28172 30058 28224 30064
rect 28080 30048 28132 30054
rect 28080 29990 28132 29996
rect 28092 29782 28120 29990
rect 28080 29776 28132 29782
rect 28080 29718 28132 29724
rect 27986 29608 28042 29617
rect 27986 29543 28042 29552
rect 28000 28626 28028 29543
rect 28092 29306 28120 29718
rect 28184 29714 28212 30058
rect 28172 29708 28224 29714
rect 28172 29650 28224 29656
rect 28080 29300 28132 29306
rect 28080 29242 28132 29248
rect 28080 28960 28132 28966
rect 28184 28948 28212 29650
rect 28264 29028 28316 29034
rect 28264 28970 28316 28976
rect 28132 28920 28212 28948
rect 28080 28902 28132 28908
rect 27988 28620 28040 28626
rect 27988 28562 28040 28568
rect 27986 28520 28042 28529
rect 27986 28455 28042 28464
rect 28000 27538 28028 28455
rect 27988 27532 28040 27538
rect 27988 27474 28040 27480
rect 28000 27130 28028 27474
rect 27988 27124 28040 27130
rect 27988 27066 28040 27072
rect 27988 25696 28040 25702
rect 27988 25638 28040 25644
rect 28000 25430 28028 25638
rect 27988 25424 28040 25430
rect 27988 25366 28040 25372
rect 27988 24200 28040 24206
rect 27988 24142 28040 24148
rect 28000 23866 28028 24142
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 28000 23322 28028 23666
rect 27988 23316 28040 23322
rect 27988 23258 28040 23264
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 27896 21684 27948 21690
rect 27896 21626 27948 21632
rect 27804 21616 27856 21622
rect 27804 21558 27856 21564
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27528 21412 27580 21418
rect 27580 21372 27660 21400
rect 27528 21354 27580 21360
rect 27436 21344 27488 21350
rect 27436 21286 27488 21292
rect 27342 21040 27398 21049
rect 27342 20975 27398 20984
rect 27252 19916 27304 19922
rect 27252 19858 27304 19864
rect 26884 19712 26936 19718
rect 26884 19654 26936 19660
rect 26792 19440 26844 19446
rect 26792 19382 26844 19388
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26516 18420 26568 18426
rect 26516 18362 26568 18368
rect 26620 18136 26648 18770
rect 26700 18148 26752 18154
rect 26620 18108 26700 18136
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26528 17066 26556 17682
rect 26620 17610 26648 18108
rect 26700 18090 26752 18096
rect 26804 17746 26832 19382
rect 26896 18873 26924 19654
rect 27264 19514 27292 19858
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 26882 18864 26938 18873
rect 26882 18799 26938 18808
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 26884 18624 26936 18630
rect 26884 18566 26936 18572
rect 26896 18426 26924 18566
rect 26884 18420 26936 18426
rect 26884 18362 26936 18368
rect 26988 18290 27016 18702
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 26988 18086 27016 18226
rect 26976 18080 27028 18086
rect 26976 18022 27028 18028
rect 26792 17740 26844 17746
rect 26792 17682 26844 17688
rect 26608 17604 26660 17610
rect 26608 17546 26660 17552
rect 26804 17338 26832 17682
rect 26792 17332 26844 17338
rect 26792 17274 26844 17280
rect 26700 17196 26752 17202
rect 26700 17138 26752 17144
rect 26516 17060 26568 17066
rect 26516 17002 26568 17008
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 26332 16652 26384 16658
rect 26332 16594 26384 16600
rect 25872 16244 25924 16250
rect 25872 16186 25924 16192
rect 26436 16114 26464 16934
rect 26608 16788 26660 16794
rect 26608 16730 26660 16736
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 26424 16108 26476 16114
rect 26424 16050 26476 16056
rect 26516 16108 26568 16114
rect 26516 16050 26568 16056
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25332 15638 25360 15846
rect 26068 15706 26096 16050
rect 26332 15972 26384 15978
rect 26332 15914 26384 15920
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 26344 15638 26372 15914
rect 25320 15632 25372 15638
rect 25320 15574 25372 15580
rect 26332 15632 26384 15638
rect 26332 15574 26384 15580
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25240 15026 25268 15302
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 25240 14618 25268 14962
rect 25332 14890 25360 15574
rect 25872 15020 25924 15026
rect 25872 14962 25924 14968
rect 25320 14884 25372 14890
rect 25320 14826 25372 14832
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 25332 13938 25360 14214
rect 25884 13938 25912 14962
rect 26344 14822 26372 15574
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 25228 13796 25280 13802
rect 25228 13738 25280 13744
rect 25240 13462 25268 13738
rect 25332 13530 25360 13874
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25228 13456 25280 13462
rect 25228 13398 25280 13404
rect 25240 13190 25268 13398
rect 25228 13184 25280 13190
rect 25228 13126 25280 13132
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25228 12368 25280 12374
rect 25228 12310 25280 12316
rect 25240 11558 25268 12310
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25136 11008 25188 11014
rect 25136 10950 25188 10956
rect 25148 10606 25176 10950
rect 25240 10810 25268 11494
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 25424 10470 25452 12582
rect 25504 11824 25556 11830
rect 25504 11766 25556 11772
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25424 9722 25452 10406
rect 25516 10198 25544 11766
rect 25700 11626 25728 12582
rect 25792 12238 25820 12718
rect 25884 12374 25912 13874
rect 26344 13462 26372 14758
rect 26424 14476 26476 14482
rect 26528 14464 26556 16050
rect 26620 15570 26648 16730
rect 26712 16726 26740 17138
rect 26700 16720 26752 16726
rect 26700 16662 26752 16668
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26620 15162 26648 15506
rect 26884 15360 26936 15366
rect 26884 15302 26936 15308
rect 26608 15156 26660 15162
rect 26608 15098 26660 15104
rect 26896 15094 26924 15302
rect 26884 15088 26936 15094
rect 26884 15030 26936 15036
rect 26896 14890 26924 15030
rect 26792 14884 26844 14890
rect 26792 14826 26844 14832
rect 26884 14884 26936 14890
rect 26884 14826 26936 14832
rect 26804 14482 26832 14826
rect 26476 14436 26556 14464
rect 26792 14476 26844 14482
rect 26424 14418 26476 14424
rect 26792 14418 26844 14424
rect 26436 14074 26464 14418
rect 26976 14272 27028 14278
rect 26976 14214 27028 14220
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26988 13870 27016 14214
rect 26976 13864 27028 13870
rect 26976 13806 27028 13812
rect 26700 13728 26752 13734
rect 26700 13670 26752 13676
rect 26332 13456 26384 13462
rect 26332 13398 26384 13404
rect 26344 12714 26372 13398
rect 26712 13394 26740 13670
rect 26700 13388 26752 13394
rect 26700 13330 26752 13336
rect 26332 12708 26384 12714
rect 26332 12650 26384 12656
rect 26712 12442 26740 13330
rect 26884 13252 26936 13258
rect 26884 13194 26936 13200
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 25872 12368 25924 12374
rect 25872 12310 25924 12316
rect 25780 12232 25832 12238
rect 25780 12174 25832 12180
rect 25884 11762 25912 12310
rect 26608 12300 26660 12306
rect 26608 12242 26660 12248
rect 26620 11898 26648 12242
rect 26608 11892 26660 11898
rect 26608 11834 26660 11840
rect 25872 11756 25924 11762
rect 25872 11698 25924 11704
rect 25688 11620 25740 11626
rect 25688 11562 25740 11568
rect 25884 11354 25912 11698
rect 26700 11552 26752 11558
rect 26700 11494 26752 11500
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 26712 11286 26740 11494
rect 26700 11280 26752 11286
rect 26700 11222 26752 11228
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26332 11008 26384 11014
rect 26332 10950 26384 10956
rect 26148 10600 26200 10606
rect 26148 10542 26200 10548
rect 25504 10192 25556 10198
rect 25504 10134 25556 10140
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 25332 9178 25360 9454
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 26160 8294 26188 10542
rect 26344 10169 26372 10950
rect 26528 10810 26556 11086
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26712 10470 26740 11222
rect 26896 10606 26924 13194
rect 26988 12306 27016 13806
rect 26976 12300 27028 12306
rect 26976 12242 27028 12248
rect 26988 11354 27016 12242
rect 26976 11348 27028 11354
rect 26976 11290 27028 11296
rect 26988 10606 27016 11290
rect 26884 10600 26936 10606
rect 26804 10560 26884 10588
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26804 10198 26832 10560
rect 26884 10542 26936 10548
rect 26976 10600 27028 10606
rect 26976 10542 27028 10548
rect 26884 10464 26936 10470
rect 26884 10406 26936 10412
rect 26792 10192 26844 10198
rect 26330 10160 26386 10169
rect 26792 10134 26844 10140
rect 26330 10095 26386 10104
rect 26804 9110 26832 10134
rect 26896 9994 26924 10406
rect 27080 10130 27108 18566
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 27172 17814 27200 18158
rect 27160 17808 27212 17814
rect 27160 17750 27212 17756
rect 27160 17128 27212 17134
rect 27160 17070 27212 17076
rect 27172 16658 27200 17070
rect 27252 16720 27304 16726
rect 27252 16662 27304 16668
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 27172 16046 27200 16594
rect 27264 16250 27292 16662
rect 27252 16244 27304 16250
rect 27252 16186 27304 16192
rect 27160 16040 27212 16046
rect 27160 15982 27212 15988
rect 27172 11218 27200 15982
rect 27356 14618 27384 20975
rect 27448 19990 27476 21286
rect 27632 20806 27660 21372
rect 27816 21350 27844 21558
rect 28000 21486 28028 21830
rect 27988 21480 28040 21486
rect 27988 21422 28040 21428
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 27896 21004 27948 21010
rect 27896 20946 27948 20952
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27436 19984 27488 19990
rect 27436 19926 27488 19932
rect 27540 19310 27568 19994
rect 27528 19304 27580 19310
rect 27528 19246 27580 19252
rect 27528 19168 27580 19174
rect 27528 19110 27580 19116
rect 27434 18864 27490 18873
rect 27434 18799 27490 18808
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 27356 14074 27384 14554
rect 27344 14068 27396 14074
rect 27344 14010 27396 14016
rect 27356 13938 27384 14010
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 27448 13814 27476 18799
rect 27540 16096 27568 19110
rect 27632 18970 27660 20742
rect 27908 20262 27936 20946
rect 28000 20806 28028 21422
rect 27988 20800 28040 20806
rect 27988 20742 28040 20748
rect 27896 20256 27948 20262
rect 27896 20198 27948 20204
rect 27712 19304 27764 19310
rect 27712 19246 27764 19252
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 27620 18148 27672 18154
rect 27724 18136 27752 19246
rect 27672 18108 27752 18136
rect 27620 18090 27672 18096
rect 27632 16794 27660 18090
rect 27908 18086 27936 20198
rect 28000 19904 28028 20742
rect 28092 20058 28120 28902
rect 28276 28626 28304 28970
rect 28264 28620 28316 28626
rect 28264 28562 28316 28568
rect 28276 28422 28304 28562
rect 28264 28416 28316 28422
rect 28264 28358 28316 28364
rect 28276 28014 28304 28358
rect 28264 28008 28316 28014
rect 28264 27950 28316 27956
rect 28276 27538 28304 27950
rect 28356 27872 28408 27878
rect 28356 27814 28408 27820
rect 28264 27532 28316 27538
rect 28264 27474 28316 27480
rect 28276 26246 28304 27474
rect 28264 26240 28316 26246
rect 28264 26182 28316 26188
rect 28276 25838 28304 26182
rect 28368 25838 28396 27814
rect 28264 25832 28316 25838
rect 28264 25774 28316 25780
rect 28356 25832 28408 25838
rect 28356 25774 28408 25780
rect 28172 23180 28224 23186
rect 28172 23122 28224 23128
rect 28184 22778 28212 23122
rect 28276 23050 28304 25774
rect 28448 25152 28500 25158
rect 28448 25094 28500 25100
rect 28460 24818 28488 25094
rect 28552 24954 28580 30126
rect 28632 29708 28684 29714
rect 28632 29650 28684 29656
rect 28644 29034 28672 29650
rect 28632 29028 28684 29034
rect 28632 28970 28684 28976
rect 28632 26580 28684 26586
rect 28632 26522 28684 26528
rect 28644 26042 28672 26522
rect 28632 26036 28684 26042
rect 28632 25978 28684 25984
rect 28540 24948 28592 24954
rect 28540 24890 28592 24896
rect 28448 24812 28500 24818
rect 28448 24754 28500 24760
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 28264 23044 28316 23050
rect 28264 22986 28316 22992
rect 28172 22772 28224 22778
rect 28172 22714 28224 22720
rect 28368 22642 28396 23802
rect 28448 23248 28500 23254
rect 28448 23190 28500 23196
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28460 22574 28488 23190
rect 28448 22568 28500 22574
rect 28448 22510 28500 22516
rect 28448 22432 28500 22438
rect 28448 22374 28500 22380
rect 28460 22030 28488 22374
rect 28552 22234 28580 24890
rect 28736 23474 28764 39782
rect 29472 39302 29500 39782
rect 29460 39296 29512 39302
rect 29460 39238 29512 39244
rect 29276 38888 29328 38894
rect 29276 38830 29328 38836
rect 29092 38752 29144 38758
rect 29092 38694 29144 38700
rect 29104 38350 29132 38694
rect 29288 38554 29316 38830
rect 29472 38826 29500 39238
rect 29460 38820 29512 38826
rect 29460 38762 29512 38768
rect 29276 38548 29328 38554
rect 29276 38490 29328 38496
rect 29564 38418 29592 39918
rect 30024 39642 30052 39986
rect 30380 39908 30432 39914
rect 30380 39850 30432 39856
rect 30012 39636 30064 39642
rect 30012 39578 30064 39584
rect 29920 38820 29972 38826
rect 29920 38762 29972 38768
rect 29552 38412 29604 38418
rect 29552 38354 29604 38360
rect 29092 38344 29144 38350
rect 29092 38286 29144 38292
rect 29104 38010 29132 38286
rect 29092 38004 29144 38010
rect 29092 37946 29144 37952
rect 29564 37806 29592 38354
rect 29932 38010 29960 38762
rect 30392 38457 30420 39850
rect 30656 39568 30708 39574
rect 30656 39510 30708 39516
rect 30668 39098 30696 39510
rect 30656 39092 30708 39098
rect 30656 39034 30708 39040
rect 30378 38448 30434 38457
rect 30378 38383 30434 38392
rect 30564 38412 30616 38418
rect 30392 38323 30420 38383
rect 30564 38354 30616 38360
rect 30196 38208 30248 38214
rect 30196 38150 30248 38156
rect 29920 38004 29972 38010
rect 29972 37964 30052 37992
rect 29920 37946 29972 37952
rect 29736 37868 29788 37874
rect 29736 37810 29788 37816
rect 29552 37800 29604 37806
rect 29552 37742 29604 37748
rect 29460 37324 29512 37330
rect 29460 37266 29512 37272
rect 29368 37256 29420 37262
rect 29368 37198 29420 37204
rect 28908 36644 28960 36650
rect 28908 36586 28960 36592
rect 28920 36242 28948 36586
rect 29380 36582 29408 37198
rect 29472 36582 29500 37266
rect 29748 37126 29776 37810
rect 29920 37800 29972 37806
rect 29920 37742 29972 37748
rect 29932 37330 29960 37742
rect 30024 37738 30052 37964
rect 30208 37806 30236 38150
rect 30576 37874 30604 38354
rect 30564 37868 30616 37874
rect 30564 37810 30616 37816
rect 30196 37800 30248 37806
rect 30196 37742 30248 37748
rect 30012 37732 30064 37738
rect 30012 37674 30064 37680
rect 30208 37398 30236 37742
rect 30196 37392 30248 37398
rect 30196 37334 30248 37340
rect 29920 37324 29972 37330
rect 29920 37266 29972 37272
rect 29736 37120 29788 37126
rect 29736 37062 29788 37068
rect 29644 36916 29696 36922
rect 29644 36858 29696 36864
rect 29656 36689 29684 36858
rect 29748 36718 29776 37062
rect 29736 36712 29788 36718
rect 29642 36680 29698 36689
rect 29736 36654 29788 36660
rect 29642 36615 29698 36624
rect 29368 36576 29420 36582
rect 29368 36518 29420 36524
rect 29460 36576 29512 36582
rect 29460 36518 29512 36524
rect 28908 36236 28960 36242
rect 28908 36178 28960 36184
rect 29092 36236 29144 36242
rect 29092 36178 29144 36184
rect 28920 35766 28948 36178
rect 28908 35760 28960 35766
rect 28908 35702 28960 35708
rect 29104 35290 29132 36178
rect 29368 36168 29420 36174
rect 29368 36110 29420 36116
rect 29276 36100 29328 36106
rect 29276 36042 29328 36048
rect 29288 35630 29316 36042
rect 29276 35624 29328 35630
rect 29276 35566 29328 35572
rect 29092 35284 29144 35290
rect 29092 35226 29144 35232
rect 28908 34400 28960 34406
rect 28908 34342 28960 34348
rect 28816 34060 28868 34066
rect 28816 34002 28868 34008
rect 28828 32774 28856 34002
rect 28920 33969 28948 34342
rect 29104 34066 29132 35226
rect 29182 35184 29238 35193
rect 29182 35119 29238 35128
rect 29196 34406 29224 35119
rect 29184 34400 29236 34406
rect 29184 34342 29236 34348
rect 29288 34134 29316 35566
rect 29380 35154 29408 36110
rect 29368 35148 29420 35154
rect 29368 35090 29420 35096
rect 29380 34746 29408 35090
rect 29368 34740 29420 34746
rect 29368 34682 29420 34688
rect 29368 34196 29420 34202
rect 29368 34138 29420 34144
rect 29276 34128 29328 34134
rect 29276 34070 29328 34076
rect 29092 34060 29144 34066
rect 29092 34002 29144 34008
rect 28906 33960 28962 33969
rect 28906 33895 28962 33904
rect 29184 33448 29236 33454
rect 29184 33390 29236 33396
rect 29196 32978 29224 33390
rect 29380 33134 29408 34138
rect 29472 33522 29500 36518
rect 29552 35556 29604 35562
rect 29552 35498 29604 35504
rect 29564 35222 29592 35498
rect 29552 35216 29604 35222
rect 29552 35158 29604 35164
rect 29552 35080 29604 35086
rect 29550 35048 29552 35057
rect 29604 35048 29606 35057
rect 29550 34983 29606 34992
rect 29564 34678 29592 34983
rect 29552 34672 29604 34678
rect 29552 34614 29604 34620
rect 29552 34536 29604 34542
rect 29552 34478 29604 34484
rect 29564 33862 29592 34478
rect 29552 33856 29604 33862
rect 29552 33798 29604 33804
rect 29460 33516 29512 33522
rect 29460 33458 29512 33464
rect 29380 33106 29500 33134
rect 29564 33114 29592 33798
rect 29656 33590 29684 36615
rect 29932 36378 29960 37266
rect 29920 36372 29972 36378
rect 29920 36314 29972 36320
rect 30564 36304 30616 36310
rect 30564 36246 30616 36252
rect 30472 36168 30524 36174
rect 30472 36110 30524 36116
rect 30484 35834 30512 36110
rect 30576 35834 30604 36246
rect 30472 35828 30524 35834
rect 30472 35770 30524 35776
rect 30564 35828 30616 35834
rect 30564 35770 30616 35776
rect 30196 35488 30248 35494
rect 30196 35430 30248 35436
rect 30208 35222 30236 35430
rect 30484 35290 30512 35770
rect 30472 35284 30524 35290
rect 30472 35226 30524 35232
rect 29736 35216 29788 35222
rect 29736 35158 29788 35164
rect 30196 35216 30248 35222
rect 30196 35158 30248 35164
rect 29748 34678 29776 35158
rect 30012 34944 30064 34950
rect 30012 34886 30064 34892
rect 29736 34672 29788 34678
rect 29736 34614 29788 34620
rect 29644 33584 29696 33590
rect 29644 33526 29696 33532
rect 29748 33402 29776 34614
rect 30024 34610 30052 34886
rect 30012 34604 30064 34610
rect 30012 34546 30064 34552
rect 30208 34474 30236 35158
rect 30576 35154 30604 35770
rect 30564 35148 30616 35154
rect 30564 35090 30616 35096
rect 30196 34468 30248 34474
rect 30196 34410 30248 34416
rect 30380 33992 30432 33998
rect 30760 33969 30788 42094
rect 30852 41546 30880 43386
rect 31036 43178 31064 43590
rect 31024 43172 31076 43178
rect 31024 43114 31076 43120
rect 31036 42838 31064 43114
rect 31220 42838 31248 43658
rect 31300 43648 31352 43654
rect 31300 43590 31352 43596
rect 31312 43314 31340 43590
rect 31300 43308 31352 43314
rect 31300 43250 31352 43256
rect 31668 43172 31720 43178
rect 31668 43114 31720 43120
rect 31024 42832 31076 42838
rect 31024 42774 31076 42780
rect 31208 42832 31260 42838
rect 31208 42774 31260 42780
rect 31036 42362 31064 42774
rect 31680 42634 31708 43114
rect 31864 42809 31892 44270
rect 34796 44192 34848 44198
rect 34796 44134 34848 44140
rect 32588 43988 32640 43994
rect 32588 43930 32640 43936
rect 32600 43314 32628 43930
rect 33692 43920 33744 43926
rect 33692 43862 33744 43868
rect 33324 43784 33376 43790
rect 33324 43726 33376 43732
rect 33336 43450 33364 43726
rect 33508 43716 33560 43722
rect 33508 43658 33560 43664
rect 33324 43444 33376 43450
rect 33324 43386 33376 43392
rect 32588 43308 32640 43314
rect 32588 43250 32640 43256
rect 31850 42800 31906 42809
rect 32862 42800 32918 42809
rect 31850 42735 31906 42744
rect 32496 42764 32548 42770
rect 32862 42735 32918 42744
rect 32496 42706 32548 42712
rect 31668 42628 31720 42634
rect 31668 42570 31720 42576
rect 31024 42356 31076 42362
rect 31024 42298 31076 42304
rect 30840 41540 30892 41546
rect 30840 41482 30892 41488
rect 31680 41138 31708 42570
rect 32508 42022 32536 42706
rect 32036 42016 32088 42022
rect 32036 41958 32088 41964
rect 32496 42016 32548 42022
rect 32496 41958 32548 41964
rect 31668 41132 31720 41138
rect 31668 41074 31720 41080
rect 31944 41132 31996 41138
rect 31944 41074 31996 41080
rect 31668 40928 31720 40934
rect 31668 40870 31720 40876
rect 31680 40730 31708 40870
rect 31956 40730 31984 41074
rect 32048 40730 32076 41958
rect 32312 41676 32364 41682
rect 32312 41618 32364 41624
rect 32220 41608 32272 41614
rect 32220 41550 32272 41556
rect 32232 41138 32260 41550
rect 32220 41132 32272 41138
rect 32220 41074 32272 41080
rect 31668 40724 31720 40730
rect 31668 40666 31720 40672
rect 31944 40724 31996 40730
rect 31944 40666 31996 40672
rect 32036 40724 32088 40730
rect 32036 40666 32088 40672
rect 32128 40588 32180 40594
rect 32128 40530 32180 40536
rect 31300 40384 31352 40390
rect 31300 40326 31352 40332
rect 31312 39982 31340 40326
rect 32140 40186 32168 40530
rect 32128 40180 32180 40186
rect 32128 40122 32180 40128
rect 30840 39976 30892 39982
rect 30840 39918 30892 39924
rect 31300 39976 31352 39982
rect 31300 39918 31352 39924
rect 30852 37942 30880 39918
rect 31576 39908 31628 39914
rect 31576 39850 31628 39856
rect 31114 39536 31170 39545
rect 31588 39506 31616 39850
rect 31114 39471 31170 39480
rect 31576 39500 31628 39506
rect 31128 39370 31156 39471
rect 31576 39442 31628 39448
rect 31116 39364 31168 39370
rect 31116 39306 31168 39312
rect 31128 39030 31156 39306
rect 31116 39024 31168 39030
rect 31116 38966 31168 38972
rect 31116 38752 31168 38758
rect 31116 38694 31168 38700
rect 31128 38010 31156 38694
rect 31116 38004 31168 38010
rect 31116 37946 31168 37952
rect 30840 37936 30892 37942
rect 30840 37878 30892 37884
rect 31116 37324 31168 37330
rect 31116 37266 31168 37272
rect 31128 36922 31156 37266
rect 31300 37120 31352 37126
rect 31300 37062 31352 37068
rect 31116 36916 31168 36922
rect 31116 36858 31168 36864
rect 31024 36100 31076 36106
rect 31024 36042 31076 36048
rect 31036 34610 31064 36042
rect 31312 35834 31340 37062
rect 32140 36718 32168 40122
rect 32232 39030 32260 41074
rect 32324 40934 32352 41618
rect 32312 40928 32364 40934
rect 32312 40870 32364 40876
rect 32220 39024 32272 39030
rect 32220 38966 32272 38972
rect 32218 38856 32274 38865
rect 32324 38842 32352 40870
rect 32404 39636 32456 39642
rect 32404 39578 32456 39584
rect 32274 38814 32352 38842
rect 32218 38791 32274 38800
rect 32128 36712 32180 36718
rect 32128 36654 32180 36660
rect 32140 36378 32168 36654
rect 31576 36372 31628 36378
rect 31576 36314 31628 36320
rect 32128 36372 32180 36378
rect 32128 36314 32180 36320
rect 31588 35834 31616 36314
rect 32232 36145 32260 38791
rect 32312 38752 32364 38758
rect 32416 38740 32444 39578
rect 32364 38712 32444 38740
rect 32312 38694 32364 38700
rect 32324 37738 32352 38694
rect 32404 37800 32456 37806
rect 32404 37742 32456 37748
rect 32312 37732 32364 37738
rect 32312 37674 32364 37680
rect 32324 37398 32352 37674
rect 32312 37392 32364 37398
rect 32312 37334 32364 37340
rect 32324 36922 32352 37334
rect 32416 37126 32444 37742
rect 32404 37120 32456 37126
rect 32404 37062 32456 37068
rect 32312 36916 32364 36922
rect 32312 36858 32364 36864
rect 32416 36786 32444 37062
rect 32404 36780 32456 36786
rect 32404 36722 32456 36728
rect 32404 36644 32456 36650
rect 32404 36586 32456 36592
rect 32416 36242 32444 36586
rect 32404 36236 32456 36242
rect 32404 36178 32456 36184
rect 32218 36136 32274 36145
rect 32218 36071 32274 36080
rect 32416 35834 32444 36178
rect 32508 36106 32536 41958
rect 32876 41177 32904 42735
rect 32956 42016 33008 42022
rect 32956 41958 33008 41964
rect 32862 41168 32918 41177
rect 32862 41103 32918 41112
rect 32772 41064 32824 41070
rect 32772 41006 32824 41012
rect 32680 39500 32732 39506
rect 32680 39442 32732 39448
rect 32692 39098 32720 39442
rect 32680 39092 32732 39098
rect 32680 39034 32732 39040
rect 32784 37233 32812 41006
rect 32876 38418 32904 41103
rect 32864 38412 32916 38418
rect 32864 38354 32916 38360
rect 32864 37256 32916 37262
rect 32770 37224 32826 37233
rect 32864 37198 32916 37204
rect 32770 37159 32826 37168
rect 32680 36644 32732 36650
rect 32680 36586 32732 36592
rect 32496 36100 32548 36106
rect 32496 36042 32548 36048
rect 31300 35828 31352 35834
rect 31300 35770 31352 35776
rect 31576 35828 31628 35834
rect 31576 35770 31628 35776
rect 32404 35828 32456 35834
rect 32404 35770 32456 35776
rect 31852 35556 31904 35562
rect 31852 35498 31904 35504
rect 31864 35154 31892 35498
rect 31852 35148 31904 35154
rect 31852 35090 31904 35096
rect 31864 34746 31892 35090
rect 32220 35080 32272 35086
rect 32220 35022 32272 35028
rect 31852 34740 31904 34746
rect 31852 34682 31904 34688
rect 30840 34604 30892 34610
rect 30840 34546 30892 34552
rect 31024 34604 31076 34610
rect 31024 34546 31076 34552
rect 30852 34202 30880 34546
rect 30840 34196 30892 34202
rect 30840 34138 30892 34144
rect 30380 33934 30432 33940
rect 30746 33960 30802 33969
rect 30392 33658 30420 33934
rect 30746 33895 30802 33904
rect 30380 33652 30432 33658
rect 30380 33594 30432 33600
rect 31036 33522 31064 34546
rect 31864 34406 31892 34682
rect 32232 34610 32260 35022
rect 32692 34678 32720 36586
rect 32680 34672 32732 34678
rect 32680 34614 32732 34620
rect 32220 34604 32272 34610
rect 32220 34546 32272 34552
rect 31852 34400 31904 34406
rect 31852 34342 31904 34348
rect 32232 34202 32260 34546
rect 32692 34202 32720 34614
rect 32220 34196 32272 34202
rect 32220 34138 32272 34144
rect 32680 34196 32732 34202
rect 32680 34138 32732 34144
rect 32128 34060 32180 34066
rect 32128 34002 32180 34008
rect 31852 33856 31904 33862
rect 31852 33798 31904 33804
rect 31024 33516 31076 33522
rect 31024 33458 31076 33464
rect 29656 33374 29776 33402
rect 30564 33380 30616 33386
rect 29184 32972 29236 32978
rect 29184 32914 29236 32920
rect 29368 32972 29420 32978
rect 29368 32914 29420 32920
rect 29000 32836 29052 32842
rect 29000 32778 29052 32784
rect 28816 32768 28868 32774
rect 28816 32710 28868 32716
rect 29012 32570 29040 32778
rect 29092 32768 29144 32774
rect 29092 32710 29144 32716
rect 29000 32564 29052 32570
rect 29000 32506 29052 32512
rect 29104 30802 29132 32710
rect 29380 31686 29408 32914
rect 29368 31680 29420 31686
rect 29368 31622 29420 31628
rect 29472 31278 29500 33106
rect 29552 33108 29604 33114
rect 29552 33050 29604 33056
rect 29552 32904 29604 32910
rect 29552 32846 29604 32852
rect 29564 31890 29592 32846
rect 29656 32570 29684 33374
rect 30564 33322 30616 33328
rect 29736 33312 29788 33318
rect 29736 33254 29788 33260
rect 29644 32564 29696 32570
rect 29644 32506 29696 32512
rect 29656 32298 29684 32506
rect 29644 32292 29696 32298
rect 29644 32234 29696 32240
rect 29656 32026 29684 32234
rect 29644 32020 29696 32026
rect 29644 31962 29696 31968
rect 29552 31884 29604 31890
rect 29552 31826 29604 31832
rect 29460 31272 29512 31278
rect 29460 31214 29512 31220
rect 29564 30938 29592 31826
rect 29656 31482 29684 31962
rect 29644 31476 29696 31482
rect 29644 31418 29696 31424
rect 29552 30932 29604 30938
rect 29552 30874 29604 30880
rect 29092 30796 29144 30802
rect 29092 30738 29144 30744
rect 29104 30054 29132 30738
rect 29092 30048 29144 30054
rect 29092 29990 29144 29996
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 28920 28082 28948 29582
rect 28908 28076 28960 28082
rect 28908 28018 28960 28024
rect 29000 27464 29052 27470
rect 29000 27406 29052 27412
rect 29012 27130 29040 27406
rect 29000 27124 29052 27130
rect 29000 27066 29052 27072
rect 29104 27010 29132 29990
rect 29460 28960 29512 28966
rect 29460 28902 29512 28908
rect 29184 28552 29236 28558
rect 29184 28494 29236 28500
rect 29196 27674 29224 28494
rect 29472 28150 29500 28902
rect 29748 28393 29776 33254
rect 30378 33008 30434 33017
rect 30378 32943 30434 32952
rect 29920 32768 29972 32774
rect 29920 32710 29972 32716
rect 29932 32434 29960 32710
rect 29920 32428 29972 32434
rect 29920 32370 29972 32376
rect 29932 31346 29960 32370
rect 30288 31476 30340 31482
rect 30288 31418 30340 31424
rect 29920 31340 29972 31346
rect 29920 31282 29972 31288
rect 30196 30796 30248 30802
rect 30196 30738 30248 30744
rect 30208 30326 30236 30738
rect 30300 30394 30328 31418
rect 30392 31346 30420 32943
rect 30576 32570 30604 33322
rect 31036 33134 31064 33458
rect 30944 33106 31064 33134
rect 30656 33040 30708 33046
rect 30656 32982 30708 32988
rect 30564 32564 30616 32570
rect 30564 32506 30616 32512
rect 30668 32298 30696 32982
rect 30748 32904 30800 32910
rect 30944 32892 30972 33106
rect 30800 32864 30972 32892
rect 30748 32846 30800 32852
rect 30472 32292 30524 32298
rect 30472 32234 30524 32240
rect 30656 32292 30708 32298
rect 30656 32234 30708 32240
rect 30484 32026 30512 32234
rect 30760 32026 30788 32846
rect 31864 32366 31892 33798
rect 32140 33318 32168 34002
rect 32784 33640 32812 37159
rect 32876 36310 32904 37198
rect 32968 36718 32996 41958
rect 33416 41472 33468 41478
rect 33416 41414 33468 41420
rect 33324 40928 33376 40934
rect 33324 40870 33376 40876
rect 33140 40452 33192 40458
rect 33140 40394 33192 40400
rect 33048 39908 33100 39914
rect 33048 39850 33100 39856
rect 33060 39642 33088 39850
rect 33048 39636 33100 39642
rect 33048 39578 33100 39584
rect 33152 39438 33180 40394
rect 33336 40050 33364 40870
rect 33428 40662 33456 41414
rect 33416 40656 33468 40662
rect 33416 40598 33468 40604
rect 33324 40044 33376 40050
rect 33324 39986 33376 39992
rect 33336 39642 33364 39986
rect 33324 39636 33376 39642
rect 33324 39578 33376 39584
rect 33428 39574 33456 40598
rect 33520 40050 33548 43658
rect 33704 43110 33732 43862
rect 33876 43444 33928 43450
rect 33876 43386 33928 43392
rect 33692 43104 33744 43110
rect 33692 43046 33744 43052
rect 33704 42906 33732 43046
rect 33692 42900 33744 42906
rect 33692 42842 33744 42848
rect 33704 42294 33732 42842
rect 33888 42362 33916 43386
rect 34244 43104 34296 43110
rect 34244 43046 34296 43052
rect 34256 42702 34284 43046
rect 34808 42838 34836 44134
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 35440 43104 35492 43110
rect 35440 43046 35492 43052
rect 34796 42832 34848 42838
rect 34796 42774 34848 42780
rect 34244 42696 34296 42702
rect 34244 42638 34296 42644
rect 34060 42628 34112 42634
rect 34060 42570 34112 42576
rect 33876 42356 33928 42362
rect 33876 42298 33928 42304
rect 33692 42288 33744 42294
rect 33744 42248 33824 42276
rect 33692 42230 33744 42236
rect 33692 42084 33744 42090
rect 33692 42026 33744 42032
rect 33704 41750 33732 42026
rect 33692 41744 33744 41750
rect 33692 41686 33744 41692
rect 33704 41274 33732 41686
rect 33692 41268 33744 41274
rect 33692 41210 33744 41216
rect 33692 40996 33744 41002
rect 33692 40938 33744 40944
rect 33704 40662 33732 40938
rect 33692 40656 33744 40662
rect 33612 40616 33692 40644
rect 33508 40044 33560 40050
rect 33508 39986 33560 39992
rect 33416 39568 33468 39574
rect 33416 39510 33468 39516
rect 33140 39432 33192 39438
rect 33140 39374 33192 39380
rect 33048 38752 33100 38758
rect 33048 38694 33100 38700
rect 33060 38554 33088 38694
rect 33048 38548 33100 38554
rect 33048 38490 33100 38496
rect 33048 38412 33100 38418
rect 33048 38354 33100 38360
rect 32956 36712 33008 36718
rect 32956 36654 33008 36660
rect 32864 36304 32916 36310
rect 32864 36246 32916 36252
rect 33060 36242 33088 38354
rect 33048 36236 33100 36242
rect 33048 36178 33100 36184
rect 33048 35488 33100 35494
rect 33048 35430 33100 35436
rect 33060 35290 33088 35430
rect 33048 35284 33100 35290
rect 33048 35226 33100 35232
rect 32864 35012 32916 35018
rect 32864 34954 32916 34960
rect 32692 33612 32812 33640
rect 32128 33312 32180 33318
rect 32128 33254 32180 33260
rect 32140 32502 32168 33254
rect 32586 33144 32642 33153
rect 32692 33134 32720 33612
rect 32772 33516 32824 33522
rect 32772 33458 32824 33464
rect 32642 33106 32720 33134
rect 32784 33114 32812 33458
rect 32772 33108 32824 33114
rect 32586 33079 32642 33088
rect 32404 33040 32456 33046
rect 32404 32982 32456 32988
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 32128 32496 32180 32502
rect 32128 32438 32180 32444
rect 31852 32360 31904 32366
rect 31852 32302 31904 32308
rect 32036 32360 32088 32366
rect 32036 32302 32088 32308
rect 30472 32020 30524 32026
rect 30472 31962 30524 31968
rect 30748 32020 30800 32026
rect 30748 31962 30800 31968
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 30472 31680 30524 31686
rect 30472 31622 30524 31628
rect 30380 31340 30432 31346
rect 30380 31282 30432 31288
rect 30484 31278 30512 31622
rect 30472 31272 30524 31278
rect 30472 31214 30524 31220
rect 30484 30802 30512 31214
rect 31024 31136 31076 31142
rect 31024 31078 31076 31084
rect 31576 31136 31628 31142
rect 31576 31078 31628 31084
rect 30472 30796 30524 30802
rect 30472 30738 30524 30744
rect 30484 30666 30512 30738
rect 30656 30728 30708 30734
rect 30656 30670 30708 30676
rect 30472 30660 30524 30666
rect 30472 30602 30524 30608
rect 30288 30388 30340 30394
rect 30288 30330 30340 30336
rect 30196 30320 30248 30326
rect 30196 30262 30248 30268
rect 30300 30122 30328 30330
rect 30288 30116 30340 30122
rect 30288 30058 30340 30064
rect 30196 29776 30248 29782
rect 30196 29718 30248 29724
rect 30208 29306 30236 29718
rect 30196 29300 30248 29306
rect 30196 29242 30248 29248
rect 30300 29050 30328 30058
rect 30484 29782 30512 30602
rect 30668 30258 30696 30670
rect 30656 30252 30708 30258
rect 30656 30194 30708 30200
rect 30472 29776 30524 29782
rect 30472 29718 30524 29724
rect 31036 29714 31064 31078
rect 31588 30394 31616 31078
rect 31576 30388 31628 30394
rect 31576 30330 31628 30336
rect 30564 29708 30616 29714
rect 30564 29650 30616 29656
rect 31024 29708 31076 29714
rect 31024 29650 31076 29656
rect 30300 29022 30420 29050
rect 30576 29034 30604 29650
rect 31208 29640 31260 29646
rect 31208 29582 31260 29588
rect 31220 29170 31248 29582
rect 31208 29164 31260 29170
rect 31208 29106 31260 29112
rect 30392 28966 30420 29022
rect 30564 29028 30616 29034
rect 30564 28970 30616 28976
rect 30380 28960 30432 28966
rect 30576 28937 30604 28970
rect 31116 28960 31168 28966
rect 30380 28902 30432 28908
rect 30562 28928 30618 28937
rect 30392 28694 30420 28902
rect 31116 28902 31168 28908
rect 30562 28863 30618 28872
rect 30380 28688 30432 28694
rect 30380 28630 30432 28636
rect 31024 28620 31076 28626
rect 31024 28562 31076 28568
rect 30196 28416 30248 28422
rect 29734 28384 29790 28393
rect 30196 28358 30248 28364
rect 30472 28416 30524 28422
rect 30472 28358 30524 28364
rect 29734 28319 29790 28328
rect 29460 28144 29512 28150
rect 29460 28086 29512 28092
rect 29736 27940 29788 27946
rect 29736 27882 29788 27888
rect 29748 27674 29776 27882
rect 29184 27668 29236 27674
rect 29184 27610 29236 27616
rect 29736 27668 29788 27674
rect 29736 27610 29788 27616
rect 29748 27130 29776 27610
rect 29736 27124 29788 27130
rect 29736 27066 29788 27072
rect 29012 26982 29132 27010
rect 28816 26920 28868 26926
rect 28816 26862 28868 26868
rect 28828 23662 28856 26862
rect 28908 24404 28960 24410
rect 28908 24346 28960 24352
rect 28920 23866 28948 24346
rect 28908 23860 28960 23866
rect 28908 23802 28960 23808
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 28736 23446 28856 23474
rect 28540 22228 28592 22234
rect 28540 22170 28592 22176
rect 28724 22160 28776 22166
rect 28724 22102 28776 22108
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 28184 21486 28212 21966
rect 28356 21888 28408 21894
rect 28356 21830 28408 21836
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28368 21350 28396 21830
rect 28460 21554 28488 21966
rect 28736 21690 28764 22102
rect 28724 21684 28776 21690
rect 28724 21626 28776 21632
rect 28448 21548 28500 21554
rect 28448 21490 28500 21496
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 28828 21146 28856 23446
rect 28908 22976 28960 22982
rect 28908 22918 28960 22924
rect 28816 21140 28868 21146
rect 28816 21082 28868 21088
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28724 20392 28776 20398
rect 28724 20334 28776 20340
rect 28736 20262 28764 20334
rect 28264 20256 28316 20262
rect 28264 20198 28316 20204
rect 28724 20256 28776 20262
rect 28724 20198 28776 20204
rect 28080 20052 28132 20058
rect 28080 19994 28132 20000
rect 28276 19990 28304 20198
rect 28264 19984 28316 19990
rect 28264 19926 28316 19932
rect 28080 19916 28132 19922
rect 28000 19876 28080 19904
rect 28080 19858 28132 19864
rect 28092 19825 28120 19858
rect 28078 19816 28134 19825
rect 28078 19751 28134 19760
rect 28276 19514 28304 19926
rect 28540 19916 28592 19922
rect 28540 19858 28592 19864
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28264 19508 28316 19514
rect 28264 19450 28316 19456
rect 28460 19174 28488 19790
rect 27988 19168 28040 19174
rect 27988 19110 28040 19116
rect 28448 19168 28500 19174
rect 28448 19110 28500 19116
rect 28000 18290 28028 19110
rect 28460 18630 28488 19110
rect 28552 18766 28580 19858
rect 28632 18828 28684 18834
rect 28632 18770 28684 18776
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28448 18624 28500 18630
rect 28448 18566 28500 18572
rect 28460 18426 28488 18566
rect 28448 18420 28500 18426
rect 28448 18362 28500 18368
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 27896 18080 27948 18086
rect 27896 18022 27948 18028
rect 28460 17882 28488 18362
rect 28552 18290 28580 18702
rect 28540 18284 28592 18290
rect 28540 18226 28592 18232
rect 28644 18222 28672 18770
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 28448 17876 28500 17882
rect 28448 17818 28500 17824
rect 27896 17740 27948 17746
rect 27896 17682 27948 17688
rect 27908 16998 27936 17682
rect 28170 17504 28226 17513
rect 28170 17439 28226 17448
rect 27896 16992 27948 16998
rect 27896 16934 27948 16940
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27908 16522 27936 16934
rect 27896 16516 27948 16522
rect 27896 16458 27948 16464
rect 27540 16068 27660 16096
rect 27632 15337 27660 16068
rect 27618 15328 27674 15337
rect 27618 15263 27674 15272
rect 27448 13786 27568 13814
rect 27540 11694 27568 13786
rect 27632 12986 27660 15263
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 27632 12782 27660 12922
rect 27620 12776 27672 12782
rect 27620 12718 27672 12724
rect 27632 12374 27660 12718
rect 27620 12368 27672 12374
rect 27620 12310 27672 12316
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 27172 10266 27200 11154
rect 27816 10849 27844 11630
rect 27802 10840 27858 10849
rect 27620 10804 27672 10810
rect 27802 10775 27858 10784
rect 27620 10746 27672 10752
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27264 10266 27292 10542
rect 27160 10260 27212 10266
rect 27160 10202 27212 10208
rect 27252 10260 27304 10266
rect 27252 10202 27304 10208
rect 27068 10124 27120 10130
rect 27068 10066 27120 10072
rect 26884 9988 26936 9994
rect 26884 9930 26936 9936
rect 27080 9722 27108 10066
rect 27068 9716 27120 9722
rect 27068 9658 27120 9664
rect 27264 9518 27292 10202
rect 27632 9586 27660 10746
rect 27620 9580 27672 9586
rect 27620 9522 27672 9528
rect 27252 9512 27304 9518
rect 27252 9454 27304 9460
rect 26792 9104 26844 9110
rect 26792 9046 26844 9052
rect 27264 9042 27292 9454
rect 27816 9450 27844 10775
rect 27804 9444 27856 9450
rect 27804 9386 27856 9392
rect 27252 9036 27304 9042
rect 27252 8978 27304 8984
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 27172 8634 27200 8910
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 27264 8430 27292 8978
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 27252 8424 27304 8430
rect 27252 8366 27304 8372
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 26436 8090 26464 8366
rect 26424 8084 26476 8090
rect 26424 8026 26476 8032
rect 27908 4154 27936 16458
rect 28184 15745 28212 17439
rect 28644 17338 28672 18158
rect 28632 17332 28684 17338
rect 28632 17274 28684 17280
rect 28264 17128 28316 17134
rect 28264 17070 28316 17076
rect 28276 16794 28304 17070
rect 28540 17060 28592 17066
rect 28736 17048 28764 20198
rect 28828 20058 28856 20878
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28828 19854 28856 19994
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28920 18902 28948 22918
rect 29012 22778 29040 26982
rect 29748 26858 29776 27066
rect 30208 27062 30236 28358
rect 30484 28082 30512 28358
rect 30472 28076 30524 28082
rect 30472 28018 30524 28024
rect 31036 27878 31064 28562
rect 31128 27946 31156 28902
rect 31220 28762 31248 29106
rect 31208 28756 31260 28762
rect 31208 28698 31260 28704
rect 31208 28416 31260 28422
rect 31208 28358 31260 28364
rect 31116 27940 31168 27946
rect 31116 27882 31168 27888
rect 30932 27872 30984 27878
rect 30932 27814 30984 27820
rect 31024 27872 31076 27878
rect 31220 27849 31248 28358
rect 31024 27814 31076 27820
rect 31206 27840 31262 27849
rect 30564 27328 30616 27334
rect 30564 27270 30616 27276
rect 30840 27328 30892 27334
rect 30840 27270 30892 27276
rect 30576 27130 30604 27270
rect 30564 27124 30616 27130
rect 30564 27066 30616 27072
rect 30196 27056 30248 27062
rect 30196 26998 30248 27004
rect 29736 26852 29788 26858
rect 29736 26794 29788 26800
rect 30576 26790 30604 27066
rect 30852 26994 30880 27270
rect 30944 27130 30972 27814
rect 31036 27402 31064 27814
rect 31206 27775 31262 27784
rect 31024 27396 31076 27402
rect 31024 27338 31076 27344
rect 31116 27396 31168 27402
rect 31116 27338 31168 27344
rect 30932 27124 30984 27130
rect 30932 27066 30984 27072
rect 31128 26994 31156 27338
rect 30840 26988 30892 26994
rect 30840 26930 30892 26936
rect 31116 26988 31168 26994
rect 31116 26930 31168 26936
rect 30288 26784 30340 26790
rect 30288 26726 30340 26732
rect 30564 26784 30616 26790
rect 30564 26726 30616 26732
rect 29092 26376 29144 26382
rect 29092 26318 29144 26324
rect 29104 25702 29132 26318
rect 29092 25696 29144 25702
rect 29092 25638 29144 25644
rect 29644 25696 29696 25702
rect 29644 25638 29696 25644
rect 29092 25424 29144 25430
rect 29092 25366 29144 25372
rect 29184 25424 29236 25430
rect 29184 25366 29236 25372
rect 29104 24954 29132 25366
rect 29092 24948 29144 24954
rect 29092 24890 29144 24896
rect 29196 24886 29224 25366
rect 29656 25226 29684 25638
rect 29644 25220 29696 25226
rect 29644 25162 29696 25168
rect 29184 24880 29236 24886
rect 29184 24822 29236 24828
rect 29656 24818 29684 25162
rect 29644 24812 29696 24818
rect 29644 24754 29696 24760
rect 29368 24676 29420 24682
rect 29368 24618 29420 24624
rect 29092 24608 29144 24614
rect 29092 24550 29144 24556
rect 29104 24070 29132 24550
rect 29380 24410 29408 24618
rect 29368 24404 29420 24410
rect 29368 24346 29420 24352
rect 29092 24064 29144 24070
rect 29092 24006 29144 24012
rect 29104 23322 29132 24006
rect 29736 23520 29788 23526
rect 29736 23462 29788 23468
rect 29092 23316 29144 23322
rect 29092 23258 29144 23264
rect 29748 23186 29776 23462
rect 30300 23186 30328 26726
rect 30748 26444 30800 26450
rect 30748 26386 30800 26392
rect 30760 25702 30788 26386
rect 30852 25974 30880 26930
rect 31128 26314 31156 26930
rect 31116 26308 31168 26314
rect 31116 26250 31168 26256
rect 31300 26240 31352 26246
rect 31300 26182 31352 26188
rect 30840 25968 30892 25974
rect 30840 25910 30892 25916
rect 31312 25906 31340 26182
rect 31300 25900 31352 25906
rect 31300 25842 31352 25848
rect 31576 25900 31628 25906
rect 31576 25842 31628 25848
rect 31024 25832 31076 25838
rect 31024 25774 31076 25780
rect 30656 25696 30708 25702
rect 30656 25638 30708 25644
rect 30748 25696 30800 25702
rect 30748 25638 30800 25644
rect 30668 25498 30696 25638
rect 30656 25492 30708 25498
rect 30656 25434 30708 25440
rect 30656 25356 30708 25362
rect 30656 25298 30708 25304
rect 30668 24614 30696 25298
rect 30564 24608 30616 24614
rect 30564 24550 30616 24556
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 30576 24342 30604 24550
rect 30564 24336 30616 24342
rect 30564 24278 30616 24284
rect 30760 24206 30788 25638
rect 31036 25226 31064 25774
rect 31208 25696 31260 25702
rect 31208 25638 31260 25644
rect 31024 25220 31076 25226
rect 31024 25162 31076 25168
rect 31220 25158 31248 25638
rect 31208 25152 31260 25158
rect 31208 25094 31260 25100
rect 30564 24200 30616 24206
rect 30564 24142 30616 24148
rect 30748 24200 30800 24206
rect 30748 24142 30800 24148
rect 30576 23798 30604 24142
rect 30564 23792 30616 23798
rect 30564 23734 30616 23740
rect 30760 23225 30788 24142
rect 31220 23866 31248 25094
rect 31588 24750 31616 25842
rect 31772 25362 31800 31758
rect 32048 31686 32076 32302
rect 32036 31680 32088 31686
rect 32036 31622 32088 31628
rect 31944 31340 31996 31346
rect 31944 31282 31996 31288
rect 31956 30938 31984 31282
rect 31944 30932 31996 30938
rect 31944 30874 31996 30880
rect 31944 30728 31996 30734
rect 31944 30670 31996 30676
rect 31956 29850 31984 30670
rect 31944 29844 31996 29850
rect 31944 29786 31996 29792
rect 32034 26616 32090 26625
rect 32034 26551 32090 26560
rect 32048 26518 32076 26551
rect 32036 26512 32088 26518
rect 32036 26454 32088 26460
rect 32048 25974 32076 26454
rect 32140 26450 32168 32438
rect 32324 32298 32352 32846
rect 32416 32434 32444 32982
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 32312 32292 32364 32298
rect 32312 32234 32364 32240
rect 32324 32026 32352 32234
rect 32312 32020 32364 32026
rect 32312 31962 32364 31968
rect 32600 31890 32628 33079
rect 32772 33050 32824 33056
rect 32588 31884 32640 31890
rect 32588 31826 32640 31832
rect 32600 31482 32628 31826
rect 32588 31476 32640 31482
rect 32588 31418 32640 31424
rect 32404 30864 32456 30870
rect 32404 30806 32456 30812
rect 32416 30394 32444 30806
rect 32404 30388 32456 30394
rect 32404 30330 32456 30336
rect 32416 29306 32444 30330
rect 32496 30116 32548 30122
rect 32496 30058 32548 30064
rect 32508 29714 32536 30058
rect 32496 29708 32548 29714
rect 32496 29650 32548 29656
rect 32508 29306 32536 29650
rect 32404 29300 32456 29306
rect 32404 29242 32456 29248
rect 32496 29300 32548 29306
rect 32496 29242 32548 29248
rect 32600 28994 32628 31418
rect 32784 31414 32812 33050
rect 32772 31408 32824 31414
rect 32772 31350 32824 31356
rect 32784 30870 32812 31350
rect 32772 30864 32824 30870
rect 32772 30806 32824 30812
rect 32876 30648 32904 34954
rect 32956 34672 33008 34678
rect 32956 34614 33008 34620
rect 32968 34202 32996 34614
rect 32956 34196 33008 34202
rect 32956 34138 33008 34144
rect 32968 33590 32996 34138
rect 33152 33862 33180 39374
rect 33520 39370 33548 39986
rect 33612 39914 33640 40616
rect 33692 40598 33744 40604
rect 33692 40384 33744 40390
rect 33692 40326 33744 40332
rect 33600 39908 33652 39914
rect 33600 39850 33652 39856
rect 33508 39364 33560 39370
rect 33508 39306 33560 39312
rect 33612 38826 33640 39850
rect 33600 38820 33652 38826
rect 33600 38762 33652 38768
rect 33230 38720 33286 38729
rect 33230 38655 33286 38664
rect 33244 37398 33272 38655
rect 33612 38554 33640 38762
rect 33600 38548 33652 38554
rect 33600 38490 33652 38496
rect 33704 38486 33732 40326
rect 33796 38486 33824 42248
rect 33968 42016 34020 42022
rect 33968 41958 34020 41964
rect 33980 39574 34008 41958
rect 34072 41614 34100 42570
rect 34256 42362 34284 42638
rect 34704 42560 34756 42566
rect 34704 42502 34756 42508
rect 34244 42356 34296 42362
rect 34244 42298 34296 42304
rect 34716 41818 34744 42502
rect 34808 42362 34836 42774
rect 35452 42634 35480 43046
rect 35716 42832 35768 42838
rect 35912 42809 35940 49558
rect 36082 49520 36138 49558
rect 41432 49558 41658 49586
rect 38016 44396 38068 44402
rect 38016 44338 38068 44344
rect 37096 43376 37148 43382
rect 37096 43318 37148 43324
rect 36174 43072 36230 43081
rect 36174 43007 36230 43016
rect 35716 42774 35768 42780
rect 35898 42800 35954 42809
rect 35532 42696 35584 42702
rect 35532 42638 35584 42644
rect 35440 42628 35492 42634
rect 35440 42570 35492 42576
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 34796 42356 34848 42362
rect 34796 42298 34848 42304
rect 35256 42220 35308 42226
rect 35256 42162 35308 42168
rect 34704 41812 34756 41818
rect 34704 41754 34756 41760
rect 34612 41744 34664 41750
rect 34612 41686 34664 41692
rect 34060 41608 34112 41614
rect 34060 41550 34112 41556
rect 34072 40662 34100 41550
rect 34624 40934 34652 41686
rect 34716 41138 34744 41754
rect 35268 41750 35296 42162
rect 35440 42152 35492 42158
rect 35440 42094 35492 42100
rect 35452 42022 35480 42094
rect 35440 42016 35492 42022
rect 35440 41958 35492 41964
rect 35256 41744 35308 41750
rect 35256 41686 35308 41692
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 34704 41132 34756 41138
rect 34704 41074 34756 41080
rect 34612 40928 34664 40934
rect 34612 40870 34664 40876
rect 34060 40656 34112 40662
rect 34060 40598 34112 40604
rect 34520 40180 34572 40186
rect 34520 40122 34572 40128
rect 33968 39568 34020 39574
rect 33968 39510 34020 39516
rect 33980 38554 34008 39510
rect 34336 38820 34388 38826
rect 34336 38762 34388 38768
rect 33968 38548 34020 38554
rect 33968 38490 34020 38496
rect 33692 38480 33744 38486
rect 33692 38422 33744 38428
rect 33784 38480 33836 38486
rect 33784 38422 33836 38428
rect 33704 38010 33732 38422
rect 33692 38004 33744 38010
rect 33692 37946 33744 37952
rect 33796 37942 33824 38422
rect 34348 38350 34376 38762
rect 34336 38344 34388 38350
rect 34336 38286 34388 38292
rect 33784 37936 33836 37942
rect 33784 37878 33836 37884
rect 34348 37874 34376 38286
rect 34336 37868 34388 37874
rect 34336 37810 34388 37816
rect 33232 37392 33284 37398
rect 33232 37334 33284 37340
rect 33784 36916 33836 36922
rect 33784 36858 33836 36864
rect 33796 36825 33824 36858
rect 33782 36816 33838 36825
rect 33782 36751 33838 36760
rect 33796 36718 33824 36751
rect 33784 36712 33836 36718
rect 33704 36672 33784 36700
rect 33232 36236 33284 36242
rect 33232 36178 33284 36184
rect 33244 35766 33272 36178
rect 33506 36136 33562 36145
rect 33506 36071 33562 36080
rect 33232 35760 33284 35766
rect 33232 35702 33284 35708
rect 33140 33856 33192 33862
rect 33244 33833 33272 35702
rect 33324 35556 33376 35562
rect 33324 35498 33376 35504
rect 33416 35556 33468 35562
rect 33416 35498 33468 35504
rect 33336 34950 33364 35498
rect 33428 35290 33456 35498
rect 33416 35284 33468 35290
rect 33416 35226 33468 35232
rect 33324 34944 33376 34950
rect 33324 34886 33376 34892
rect 33520 34066 33548 36071
rect 33704 34649 33732 36672
rect 33784 36654 33836 36660
rect 34060 36100 34112 36106
rect 34060 36042 34112 36048
rect 33784 35080 33836 35086
rect 33784 35022 33836 35028
rect 33796 34746 33824 35022
rect 33968 34944 34020 34950
rect 33968 34886 34020 34892
rect 33980 34746 34008 34886
rect 33784 34740 33836 34746
rect 33784 34682 33836 34688
rect 33968 34740 34020 34746
rect 33968 34682 34020 34688
rect 33690 34640 33746 34649
rect 33690 34575 33746 34584
rect 33600 34468 33652 34474
rect 33600 34410 33652 34416
rect 33508 34060 33560 34066
rect 33508 34002 33560 34008
rect 33322 33960 33378 33969
rect 33322 33895 33378 33904
rect 33140 33798 33192 33804
rect 33230 33824 33286 33833
rect 33230 33759 33286 33768
rect 32956 33584 33008 33590
rect 32956 33526 33008 33532
rect 33232 33584 33284 33590
rect 33232 33526 33284 33532
rect 32968 33402 32996 33526
rect 32968 33374 33180 33402
rect 33048 33312 33100 33318
rect 33048 33254 33100 33260
rect 33060 33114 33088 33254
rect 33048 33108 33100 33114
rect 33048 33050 33100 33056
rect 33152 32842 33180 33374
rect 33140 32836 33192 32842
rect 33140 32778 33192 32784
rect 33140 32224 33192 32230
rect 33140 32166 33192 32172
rect 33152 31414 33180 32166
rect 33140 31408 33192 31414
rect 33140 31350 33192 31356
rect 32956 30660 33008 30666
rect 32876 30620 32956 30648
rect 32956 30602 33008 30608
rect 32864 30184 32916 30190
rect 32864 30126 32916 30132
rect 32876 29782 32904 30126
rect 32864 29776 32916 29782
rect 32864 29718 32916 29724
rect 32772 29708 32824 29714
rect 32772 29650 32824 29656
rect 32784 29306 32812 29650
rect 32772 29300 32824 29306
rect 32772 29242 32824 29248
rect 32956 29164 33008 29170
rect 32956 29106 33008 29112
rect 32416 28966 32628 28994
rect 32312 27600 32364 27606
rect 32312 27542 32364 27548
rect 32220 27464 32272 27470
rect 32220 27406 32272 27412
rect 32128 26444 32180 26450
rect 32128 26386 32180 26392
rect 32232 26314 32260 27406
rect 32324 27062 32352 27542
rect 32312 27056 32364 27062
rect 32312 26998 32364 27004
rect 32220 26308 32272 26314
rect 32220 26250 32272 26256
rect 32036 25968 32088 25974
rect 32036 25910 32088 25916
rect 32312 25968 32364 25974
rect 32312 25910 32364 25916
rect 31760 25356 31812 25362
rect 31760 25298 31812 25304
rect 32128 25356 32180 25362
rect 32128 25298 32180 25304
rect 31668 25152 31720 25158
rect 31668 25094 31720 25100
rect 31680 24818 31708 25094
rect 32140 24818 32168 25298
rect 31668 24812 31720 24818
rect 31668 24754 31720 24760
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 31576 24744 31628 24750
rect 31576 24686 31628 24692
rect 31300 24676 31352 24682
rect 31300 24618 31352 24624
rect 31312 24206 31340 24618
rect 32140 24614 32168 24754
rect 31392 24608 31444 24614
rect 31392 24550 31444 24556
rect 32128 24608 32180 24614
rect 32128 24550 32180 24556
rect 31300 24200 31352 24206
rect 31300 24142 31352 24148
rect 31208 23860 31260 23866
rect 31208 23802 31260 23808
rect 30840 23656 30892 23662
rect 30840 23598 30892 23604
rect 31206 23624 31262 23633
rect 30852 23526 30880 23598
rect 31206 23559 31262 23568
rect 30840 23520 30892 23526
rect 30840 23462 30892 23468
rect 30746 23216 30802 23225
rect 29736 23180 29788 23186
rect 29736 23122 29788 23128
rect 30288 23180 30340 23186
rect 30746 23151 30802 23160
rect 30288 23122 30340 23128
rect 29276 22976 29328 22982
rect 29276 22918 29328 22924
rect 29000 22772 29052 22778
rect 29000 22714 29052 22720
rect 29288 22574 29316 22918
rect 29276 22568 29328 22574
rect 29276 22510 29328 22516
rect 29828 22568 29880 22574
rect 29828 22510 29880 22516
rect 29288 22166 29316 22510
rect 29276 22160 29328 22166
rect 29276 22102 29328 22108
rect 29092 22092 29144 22098
rect 29092 22034 29144 22040
rect 29104 21010 29132 22034
rect 29552 21956 29604 21962
rect 29552 21898 29604 21904
rect 29276 21888 29328 21894
rect 29276 21830 29328 21836
rect 29288 21622 29316 21830
rect 29564 21622 29592 21898
rect 29276 21616 29328 21622
rect 29276 21558 29328 21564
rect 29552 21616 29604 21622
rect 29552 21558 29604 21564
rect 29184 21412 29236 21418
rect 29184 21354 29236 21360
rect 29092 21004 29144 21010
rect 29092 20946 29144 20952
rect 29000 20868 29052 20874
rect 29000 20810 29052 20816
rect 29012 20058 29040 20810
rect 29104 20806 29132 20946
rect 29092 20800 29144 20806
rect 29092 20742 29144 20748
rect 29104 20330 29132 20742
rect 29196 20602 29224 21354
rect 29288 20874 29316 21558
rect 29564 20942 29592 21558
rect 29644 21548 29696 21554
rect 29644 21490 29696 21496
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 29276 20868 29328 20874
rect 29276 20810 29328 20816
rect 29184 20596 29236 20602
rect 29184 20538 29236 20544
rect 29092 20324 29144 20330
rect 29092 20266 29144 20272
rect 29000 20052 29052 20058
rect 29000 19994 29052 20000
rect 29104 19718 29132 20266
rect 29196 19990 29224 20538
rect 29288 20534 29316 20810
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29276 20528 29328 20534
rect 29276 20470 29328 20476
rect 29184 19984 29236 19990
rect 29184 19926 29236 19932
rect 29092 19712 29144 19718
rect 29092 19654 29144 19660
rect 29104 19310 29132 19654
rect 29196 19334 29224 19926
rect 29380 19718 29408 20742
rect 29564 20534 29592 20878
rect 29552 20528 29604 20534
rect 29552 20470 29604 20476
rect 29656 20466 29684 21490
rect 29644 20460 29696 20466
rect 29644 20402 29696 20408
rect 29644 20324 29696 20330
rect 29644 20266 29696 20272
rect 29460 19916 29512 19922
rect 29460 19858 29512 19864
rect 29368 19712 29420 19718
rect 29368 19654 29420 19660
rect 29380 19514 29408 19654
rect 29472 19514 29500 19858
rect 29656 19514 29684 20266
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29368 19508 29420 19514
rect 29368 19450 29420 19456
rect 29460 19508 29512 19514
rect 29460 19450 29512 19456
rect 29644 19508 29696 19514
rect 29644 19450 29696 19456
rect 29092 19304 29144 19310
rect 29196 19306 29316 19334
rect 29092 19246 29144 19252
rect 29288 18970 29316 19306
rect 29656 18970 29684 19450
rect 29748 19378 29776 19790
rect 29736 19372 29788 19378
rect 29736 19314 29788 19320
rect 29276 18964 29328 18970
rect 29276 18906 29328 18912
rect 29644 18964 29696 18970
rect 29644 18906 29696 18912
rect 28908 18896 28960 18902
rect 28908 18838 28960 18844
rect 29288 18222 29316 18906
rect 29368 18624 29420 18630
rect 29368 18566 29420 18572
rect 29276 18216 29328 18222
rect 29276 18158 29328 18164
rect 29184 18148 29236 18154
rect 29184 18090 29236 18096
rect 28908 17808 28960 17814
rect 28908 17750 28960 17756
rect 28592 17020 28764 17048
rect 28540 17002 28592 17008
rect 28356 16992 28408 16998
rect 28356 16934 28408 16940
rect 28264 16788 28316 16794
rect 28264 16730 28316 16736
rect 28368 16658 28396 16934
rect 28356 16652 28408 16658
rect 28356 16594 28408 16600
rect 28170 15736 28226 15745
rect 28170 15671 28226 15680
rect 28264 14952 28316 14958
rect 28264 14894 28316 14900
rect 28276 14550 28304 14894
rect 28264 14544 28316 14550
rect 28264 14486 28316 14492
rect 28080 14476 28132 14482
rect 28080 14418 28132 14424
rect 28092 14074 28120 14418
rect 28080 14068 28132 14074
rect 28080 14010 28132 14016
rect 28092 12782 28120 14010
rect 28080 12776 28132 12782
rect 28080 12718 28132 12724
rect 28092 12442 28120 12718
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 28092 11694 28120 12378
rect 28080 11688 28132 11694
rect 28080 11630 28132 11636
rect 28092 10130 28120 11630
rect 28080 10124 28132 10130
rect 28080 10066 28132 10072
rect 28448 10124 28500 10130
rect 28448 10066 28500 10072
rect 28172 9988 28224 9994
rect 28172 9930 28224 9936
rect 28184 9722 28212 9930
rect 28460 9722 28488 10066
rect 28172 9716 28224 9722
rect 28172 9658 28224 9664
rect 28448 9716 28500 9722
rect 28448 9658 28500 9664
rect 28184 8974 28212 9658
rect 28460 9110 28488 9658
rect 28448 9104 28500 9110
rect 28448 9046 28500 9052
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 28460 8634 28488 9046
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 27908 4126 28212 4154
rect 28184 3913 28212 4126
rect 28170 3904 28226 3913
rect 28170 3839 28226 3848
rect 28552 134 28580 17002
rect 28920 16726 28948 17750
rect 29196 16833 29224 18090
rect 29288 17338 29316 18158
rect 29276 17332 29328 17338
rect 29276 17274 29328 17280
rect 29182 16824 29238 16833
rect 29182 16759 29238 16768
rect 28908 16720 28960 16726
rect 28908 16662 28960 16668
rect 28920 16250 28948 16662
rect 29000 16448 29052 16454
rect 29000 16390 29052 16396
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 28644 16017 28672 16050
rect 28630 16008 28686 16017
rect 28630 15943 28686 15952
rect 29012 14482 29040 16390
rect 29276 15632 29328 15638
rect 29276 15574 29328 15580
rect 29288 15094 29316 15574
rect 29380 15502 29408 18566
rect 29552 18352 29604 18358
rect 29552 18294 29604 18300
rect 29564 17882 29592 18294
rect 29552 17876 29604 17882
rect 29552 17818 29604 17824
rect 29644 17740 29696 17746
rect 29840 17728 29868 22510
rect 29920 22500 29972 22506
rect 29920 22442 29972 22448
rect 29932 18290 29960 22442
rect 30300 22438 30328 23122
rect 30472 22976 30524 22982
rect 30472 22918 30524 22924
rect 30484 22574 30512 22918
rect 30472 22568 30524 22574
rect 30472 22510 30524 22516
rect 30288 22432 30340 22438
rect 30288 22374 30340 22380
rect 30012 20324 30064 20330
rect 30012 20266 30064 20272
rect 30024 20097 30052 20266
rect 30010 20088 30066 20097
rect 30010 20023 30066 20032
rect 30104 19236 30156 19242
rect 30104 19178 30156 19184
rect 30116 19009 30144 19178
rect 30102 19000 30158 19009
rect 30102 18935 30158 18944
rect 30300 18952 30328 22374
rect 30378 22264 30434 22273
rect 30378 22199 30434 22208
rect 30392 22166 30420 22199
rect 30380 22160 30432 22166
rect 30380 22102 30432 22108
rect 30392 21418 30420 22102
rect 30380 21412 30432 21418
rect 30380 21354 30432 21360
rect 30562 21040 30618 21049
rect 30562 20975 30618 20984
rect 30656 21004 30708 21010
rect 30576 20942 30604 20975
rect 30656 20946 30708 20952
rect 30564 20936 30616 20942
rect 30564 20878 30616 20884
rect 30668 20602 30696 20946
rect 30656 20596 30708 20602
rect 30656 20538 30708 20544
rect 30748 20596 30800 20602
rect 30748 20538 30800 20544
rect 30668 19446 30696 20538
rect 30760 20058 30788 20538
rect 30748 20052 30800 20058
rect 30748 19994 30800 20000
rect 30748 19712 30800 19718
rect 30748 19654 30800 19660
rect 30656 19440 30708 19446
rect 30656 19382 30708 19388
rect 30300 18924 30420 18952
rect 30288 18828 30340 18834
rect 30288 18770 30340 18776
rect 30196 18624 30248 18630
rect 30196 18566 30248 18572
rect 30208 18426 30236 18566
rect 30300 18426 30328 18770
rect 30196 18420 30248 18426
rect 30196 18362 30248 18368
rect 30288 18420 30340 18426
rect 30288 18362 30340 18368
rect 29920 18284 29972 18290
rect 29920 18226 29972 18232
rect 30300 18086 30328 18362
rect 29920 18080 29972 18086
rect 29920 18022 29972 18028
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 29696 17700 29868 17728
rect 29644 17682 29696 17688
rect 29656 17202 29684 17682
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29656 16998 29684 17138
rect 29932 17134 29960 18022
rect 30300 17921 30328 18022
rect 30286 17912 30342 17921
rect 30286 17847 30342 17856
rect 30012 17740 30064 17746
rect 30012 17682 30064 17688
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 29644 16992 29696 16998
rect 29644 16934 29696 16940
rect 29656 16182 29684 16934
rect 30024 16794 30052 17682
rect 30104 17672 30156 17678
rect 30104 17614 30156 17620
rect 30116 17202 30144 17614
rect 30104 17196 30156 17202
rect 30104 17138 30156 17144
rect 30288 16992 30340 16998
rect 30288 16934 30340 16940
rect 29736 16788 29788 16794
rect 29736 16730 29788 16736
rect 30012 16788 30064 16794
rect 30012 16730 30064 16736
rect 29644 16176 29696 16182
rect 29644 16118 29696 16124
rect 29748 16046 29776 16730
rect 30300 16726 30328 16934
rect 30288 16720 30340 16726
rect 30288 16662 30340 16668
rect 30196 16584 30248 16590
rect 30196 16526 30248 16532
rect 30208 16114 30236 16526
rect 30196 16108 30248 16114
rect 30196 16050 30248 16056
rect 29736 16040 29788 16046
rect 29736 15982 29788 15988
rect 29748 15706 29776 15982
rect 30300 15910 30328 16662
rect 30392 16017 30420 18924
rect 30760 18193 30788 19654
rect 30746 18184 30802 18193
rect 30746 18119 30802 18128
rect 30378 16008 30434 16017
rect 30378 15943 30434 15952
rect 30288 15904 30340 15910
rect 30288 15846 30340 15852
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 29368 15496 29420 15502
rect 29368 15438 29420 15444
rect 29380 15162 29408 15438
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 29276 15088 29328 15094
rect 29276 15030 29328 15036
rect 29288 14550 29316 15030
rect 30300 14890 30328 15846
rect 30852 15570 30880 23462
rect 30930 23216 30986 23225
rect 30930 23151 30986 23160
rect 30944 19514 30972 23151
rect 31024 22568 31076 22574
rect 31024 22510 31076 22516
rect 31036 22098 31064 22510
rect 31116 22228 31168 22234
rect 31116 22170 31168 22176
rect 31024 22092 31076 22098
rect 31024 22034 31076 22040
rect 31128 21350 31156 22170
rect 31116 21344 31168 21350
rect 31116 21286 31168 21292
rect 31024 20868 31076 20874
rect 31024 20810 31076 20816
rect 31036 20398 31064 20810
rect 31116 20528 31168 20534
rect 31116 20470 31168 20476
rect 31024 20392 31076 20398
rect 31024 20334 31076 20340
rect 31128 19990 31156 20470
rect 31116 19984 31168 19990
rect 31116 19926 31168 19932
rect 31024 19916 31076 19922
rect 31024 19858 31076 19864
rect 30932 19508 30984 19514
rect 30932 19450 30984 19456
rect 30932 19304 30984 19310
rect 30932 19246 30984 19252
rect 30944 17610 30972 19246
rect 31036 17882 31064 19858
rect 31116 18828 31168 18834
rect 31116 18770 31168 18776
rect 31128 18358 31156 18770
rect 31116 18352 31168 18358
rect 31116 18294 31168 18300
rect 31128 18154 31156 18294
rect 31116 18148 31168 18154
rect 31116 18090 31168 18096
rect 31024 17876 31076 17882
rect 31024 17818 31076 17824
rect 30932 17604 30984 17610
rect 30932 17546 30984 17552
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 31128 16250 31156 16390
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 30840 15564 30892 15570
rect 30840 15506 30892 15512
rect 30852 15162 30880 15506
rect 30840 15156 30892 15162
rect 30840 15098 30892 15104
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 30288 14884 30340 14890
rect 30288 14826 30340 14832
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 30208 14550 30236 14758
rect 29276 14544 29328 14550
rect 29276 14486 29328 14492
rect 30196 14544 30248 14550
rect 30196 14486 30248 14492
rect 29000 14476 29052 14482
rect 29000 14418 29052 14424
rect 29184 14408 29236 14414
rect 29184 14350 29236 14356
rect 29196 14074 29224 14350
rect 29184 14068 29236 14074
rect 29184 14010 29236 14016
rect 29092 14000 29144 14006
rect 28814 13968 28870 13977
rect 29092 13942 29144 13948
rect 28814 13903 28870 13912
rect 28828 13870 28856 13903
rect 28816 13864 28868 13870
rect 28816 13806 28868 13812
rect 29104 13802 29132 13942
rect 29092 13796 29144 13802
rect 29092 13738 29144 13744
rect 29196 13530 29224 14010
rect 29288 14006 29316 14486
rect 29276 14000 29328 14006
rect 29276 13942 29328 13948
rect 29828 14000 29880 14006
rect 29828 13942 29880 13948
rect 29460 13796 29512 13802
rect 29460 13738 29512 13744
rect 29472 13530 29500 13738
rect 29184 13524 29236 13530
rect 29184 13466 29236 13472
rect 29460 13524 29512 13530
rect 29460 13466 29512 13472
rect 28816 13388 28868 13394
rect 28816 13330 28868 13336
rect 28828 12850 28856 13330
rect 29736 13184 29788 13190
rect 29736 13126 29788 13132
rect 28816 12844 28868 12850
rect 28816 12786 28868 12792
rect 28828 12753 28856 12786
rect 28814 12744 28870 12753
rect 28632 12708 28684 12714
rect 29748 12714 29776 13126
rect 28814 12679 28870 12688
rect 29736 12708 29788 12714
rect 28632 12650 28684 12656
rect 29736 12650 29788 12656
rect 28644 12238 28672 12650
rect 29748 12442 29776 12650
rect 28908 12436 28960 12442
rect 28908 12378 28960 12384
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 28644 11354 28672 12174
rect 28920 11558 28948 12378
rect 29276 11688 29328 11694
rect 29276 11630 29328 11636
rect 28908 11552 28960 11558
rect 28908 11494 28960 11500
rect 28632 11348 28684 11354
rect 28632 11290 28684 11296
rect 28724 11212 28776 11218
rect 28724 11154 28776 11160
rect 28736 11082 28764 11154
rect 28724 11076 28776 11082
rect 28724 11018 28776 11024
rect 28736 10810 28764 11018
rect 28724 10804 28776 10810
rect 28724 10746 28776 10752
rect 28920 10266 28948 11494
rect 29288 11354 29316 11630
rect 29276 11348 29328 11354
rect 29276 11290 29328 11296
rect 29840 11150 29868 13942
rect 30576 13394 30604 14894
rect 30852 14346 30880 15098
rect 30840 14340 30892 14346
rect 30840 14282 30892 14288
rect 31220 13569 31248 23559
rect 31312 23322 31340 24142
rect 31404 23866 31432 24550
rect 31576 24132 31628 24138
rect 31576 24074 31628 24080
rect 31484 24064 31536 24070
rect 31484 24006 31536 24012
rect 31392 23860 31444 23866
rect 31392 23802 31444 23808
rect 31300 23316 31352 23322
rect 31300 23258 31352 23264
rect 31300 20528 31352 20534
rect 31300 20470 31352 20476
rect 31312 19922 31340 20470
rect 31300 19916 31352 19922
rect 31300 19858 31352 19864
rect 31404 19417 31432 23802
rect 31496 23730 31524 24006
rect 31588 23730 31616 24074
rect 31484 23724 31536 23730
rect 31484 23666 31536 23672
rect 31576 23724 31628 23730
rect 31576 23666 31628 23672
rect 31496 23254 31524 23666
rect 32324 23474 32352 25910
rect 32416 24342 32444 28966
rect 32968 28626 32996 29106
rect 32956 28620 33008 28626
rect 32956 28562 33008 28568
rect 32496 28416 32548 28422
rect 32496 28358 32548 28364
rect 32508 28014 32536 28358
rect 32968 28218 32996 28562
rect 33140 28416 33192 28422
rect 33140 28358 33192 28364
rect 32956 28212 33008 28218
rect 32956 28154 33008 28160
rect 32496 28008 32548 28014
rect 32496 27950 32548 27956
rect 32968 27713 32996 28154
rect 32954 27704 33010 27713
rect 32954 27639 33010 27648
rect 32772 27396 32824 27402
rect 32772 27338 32824 27344
rect 32680 27328 32732 27334
rect 32680 27270 32732 27276
rect 32496 27124 32548 27130
rect 32496 27066 32548 27072
rect 32508 26858 32536 27066
rect 32692 26994 32720 27270
rect 32784 26994 32812 27338
rect 32680 26988 32732 26994
rect 32680 26930 32732 26936
rect 32772 26988 32824 26994
rect 32772 26930 32824 26936
rect 32496 26852 32548 26858
rect 32496 26794 32548 26800
rect 32692 26246 32720 26930
rect 33152 26382 33180 28358
rect 33140 26376 33192 26382
rect 33140 26318 33192 26324
rect 32680 26240 32732 26246
rect 32680 26182 32732 26188
rect 32496 25492 32548 25498
rect 32496 25434 32548 25440
rect 32508 24818 32536 25434
rect 32496 24812 32548 24818
rect 32496 24754 32548 24760
rect 32588 24676 32640 24682
rect 32588 24618 32640 24624
rect 32404 24336 32456 24342
rect 32404 24278 32456 24284
rect 32416 23798 32444 24278
rect 32600 24206 32628 24618
rect 32588 24200 32640 24206
rect 32588 24142 32640 24148
rect 32692 24138 32720 26182
rect 33152 25974 33180 26318
rect 33140 25968 33192 25974
rect 33140 25910 33192 25916
rect 32864 25764 32916 25770
rect 32864 25706 32916 25712
rect 33140 25764 33192 25770
rect 33140 25706 33192 25712
rect 32876 25294 32904 25706
rect 32864 25288 32916 25294
rect 32864 25230 32916 25236
rect 32772 25152 32824 25158
rect 32772 25094 32824 25100
rect 32680 24132 32732 24138
rect 32680 24074 32732 24080
rect 32404 23792 32456 23798
rect 32404 23734 32456 23740
rect 32416 23633 32444 23734
rect 32402 23624 32458 23633
rect 32402 23559 32458 23568
rect 32324 23446 32444 23474
rect 31484 23248 31536 23254
rect 31484 23190 31536 23196
rect 32128 23112 32180 23118
rect 32128 23054 32180 23060
rect 31484 22636 31536 22642
rect 31484 22578 31536 22584
rect 31496 20602 31524 22578
rect 32140 22166 32168 23054
rect 32128 22160 32180 22166
rect 32128 22102 32180 22108
rect 32128 21480 32180 21486
rect 32128 21422 32180 21428
rect 31668 21344 31720 21350
rect 31668 21286 31720 21292
rect 31484 20596 31536 20602
rect 31484 20538 31536 20544
rect 31576 20052 31628 20058
rect 31576 19994 31628 20000
rect 31390 19408 31446 19417
rect 31390 19343 31446 19352
rect 31300 19168 31352 19174
rect 31392 19168 31444 19174
rect 31300 19110 31352 19116
rect 31390 19136 31392 19145
rect 31444 19136 31446 19145
rect 31312 16794 31340 19110
rect 31390 19071 31446 19080
rect 31404 17066 31432 19071
rect 31588 18970 31616 19994
rect 31576 18964 31628 18970
rect 31576 18906 31628 18912
rect 31484 18216 31536 18222
rect 31482 18184 31484 18193
rect 31536 18184 31538 18193
rect 31482 18119 31538 18128
rect 31496 17882 31524 18119
rect 31484 17876 31536 17882
rect 31484 17818 31536 17824
rect 31392 17060 31444 17066
rect 31392 17002 31444 17008
rect 31300 16788 31352 16794
rect 31300 16730 31352 16736
rect 31312 16114 31340 16730
rect 31300 16108 31352 16114
rect 31496 16096 31524 17818
rect 31576 16244 31628 16250
rect 31576 16186 31628 16192
rect 31300 16050 31352 16056
rect 31404 16068 31524 16096
rect 31300 14476 31352 14482
rect 31300 14418 31352 14424
rect 31312 14278 31340 14418
rect 31300 14272 31352 14278
rect 31300 14214 31352 14220
rect 31312 14006 31340 14214
rect 31300 14000 31352 14006
rect 31300 13942 31352 13948
rect 31312 13705 31340 13942
rect 31298 13696 31354 13705
rect 31298 13631 31354 13640
rect 31206 13560 31262 13569
rect 31206 13495 31262 13504
rect 30564 13388 30616 13394
rect 30564 13330 30616 13336
rect 30576 12986 30604 13330
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 30472 12912 30524 12918
rect 30472 12854 30524 12860
rect 29920 12844 29972 12850
rect 29920 12786 29972 12792
rect 29932 12442 29960 12786
rect 29920 12436 29972 12442
rect 29920 12378 29972 12384
rect 30484 12238 30512 12854
rect 30564 12368 30616 12374
rect 30564 12310 30616 12316
rect 30472 12232 30524 12238
rect 30472 12174 30524 12180
rect 30484 11830 30512 12174
rect 30576 11898 30604 12310
rect 30564 11892 30616 11898
rect 30564 11834 30616 11840
rect 30472 11824 30524 11830
rect 30472 11766 30524 11772
rect 31220 11694 31248 13495
rect 31312 13394 31340 13631
rect 31300 13388 31352 13394
rect 31300 13330 31352 13336
rect 31312 12986 31340 13330
rect 31404 13258 31432 16068
rect 31588 15978 31616 16186
rect 31484 15972 31536 15978
rect 31484 15914 31536 15920
rect 31576 15972 31628 15978
rect 31576 15914 31628 15920
rect 31496 14550 31524 15914
rect 31588 15638 31616 15914
rect 31576 15632 31628 15638
rect 31576 15574 31628 15580
rect 31680 15162 31708 21286
rect 32140 20806 32168 21422
rect 32312 21004 32364 21010
rect 32312 20946 32364 20952
rect 31944 20800 31996 20806
rect 31944 20742 31996 20748
rect 32128 20800 32180 20806
rect 32128 20742 32180 20748
rect 31956 20602 31984 20742
rect 31944 20596 31996 20602
rect 31944 20538 31996 20544
rect 31956 20505 31984 20538
rect 31942 20496 31998 20505
rect 31942 20431 31998 20440
rect 31956 20058 31984 20431
rect 31944 20052 31996 20058
rect 31944 19994 31996 20000
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32128 19440 32180 19446
rect 32128 19382 32180 19388
rect 31944 19304 31996 19310
rect 31944 19246 31996 19252
rect 31956 18630 31984 19246
rect 32036 19236 32088 19242
rect 32036 19178 32088 19184
rect 32048 19145 32076 19178
rect 32034 19136 32090 19145
rect 32034 19071 32090 19080
rect 32140 18834 32168 19382
rect 32232 19156 32260 19790
rect 32324 19378 32352 20946
rect 32416 19553 32444 23446
rect 32496 23316 32548 23322
rect 32496 23258 32548 23264
rect 32508 22438 32536 23258
rect 32496 22432 32548 22438
rect 32496 22374 32548 22380
rect 32508 21078 32536 22374
rect 32588 21480 32640 21486
rect 32588 21422 32640 21428
rect 32600 21146 32628 21422
rect 32588 21140 32640 21146
rect 32588 21082 32640 21088
rect 32496 21072 32548 21078
rect 32496 21014 32548 21020
rect 32508 20262 32536 21014
rect 32496 20256 32548 20262
rect 32496 20198 32548 20204
rect 32508 20058 32536 20198
rect 32496 20052 32548 20058
rect 32496 19994 32548 20000
rect 32402 19544 32458 19553
rect 32402 19479 32458 19488
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32508 19242 32536 19994
rect 32496 19236 32548 19242
rect 32496 19178 32548 19184
rect 32404 19168 32456 19174
rect 32232 19128 32404 19156
rect 32232 18970 32260 19128
rect 32404 19110 32456 19116
rect 32220 18964 32272 18970
rect 32220 18906 32272 18912
rect 32600 18834 32628 21082
rect 32784 21010 32812 25094
rect 33152 24818 33180 25706
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 32956 22432 33008 22438
rect 32956 22374 33008 22380
rect 32864 21412 32916 21418
rect 32864 21354 32916 21360
rect 32876 21010 32904 21354
rect 32772 21004 32824 21010
rect 32772 20946 32824 20952
rect 32864 21004 32916 21010
rect 32864 20946 32916 20952
rect 32772 20868 32824 20874
rect 32772 20810 32824 20816
rect 32784 19802 32812 20810
rect 32968 20346 32996 22374
rect 33140 22092 33192 22098
rect 33140 22034 33192 22040
rect 33152 21418 33180 22034
rect 33140 21412 33192 21418
rect 33140 21354 33192 21360
rect 32692 19774 32812 19802
rect 32876 20318 32996 20346
rect 32128 18828 32180 18834
rect 32220 18828 32272 18834
rect 32180 18788 32220 18816
rect 32128 18770 32180 18776
rect 32220 18770 32272 18776
rect 32404 18828 32456 18834
rect 32404 18770 32456 18776
rect 32588 18828 32640 18834
rect 32588 18770 32640 18776
rect 32312 18760 32364 18766
rect 32312 18702 32364 18708
rect 32220 18692 32272 18698
rect 32220 18634 32272 18640
rect 31944 18624 31996 18630
rect 31944 18566 31996 18572
rect 31956 18290 31984 18566
rect 31944 18284 31996 18290
rect 31944 18226 31996 18232
rect 31852 18216 31904 18222
rect 31852 18158 31904 18164
rect 31864 17882 31892 18158
rect 31852 17876 31904 17882
rect 31852 17818 31904 17824
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 31760 17060 31812 17066
rect 31760 17002 31812 17008
rect 31772 15978 31800 17002
rect 31956 16794 31984 17138
rect 31944 16788 31996 16794
rect 31944 16730 31996 16736
rect 32232 16726 32260 18634
rect 32324 17746 32352 18702
rect 32416 18086 32444 18770
rect 32404 18080 32456 18086
rect 32404 18022 32456 18028
rect 32600 17882 32628 18770
rect 32692 18154 32720 19774
rect 32680 18148 32732 18154
rect 32680 18090 32732 18096
rect 32772 18080 32824 18086
rect 32772 18022 32824 18028
rect 32588 17876 32640 17882
rect 32588 17818 32640 17824
rect 32312 17740 32364 17746
rect 32312 17682 32364 17688
rect 32324 17270 32352 17682
rect 32496 17536 32548 17542
rect 32496 17478 32548 17484
rect 32508 17338 32536 17478
rect 32496 17332 32548 17338
rect 32496 17274 32548 17280
rect 32312 17264 32364 17270
rect 32312 17206 32364 17212
rect 32678 17232 32734 17241
rect 32678 17167 32734 17176
rect 32692 17134 32720 17167
rect 32680 17128 32732 17134
rect 32680 17070 32732 17076
rect 32588 17060 32640 17066
rect 32588 17002 32640 17008
rect 32312 16992 32364 16998
rect 32312 16934 32364 16940
rect 32324 16726 32352 16934
rect 32220 16720 32272 16726
rect 32220 16662 32272 16668
rect 32312 16720 32364 16726
rect 32312 16662 32364 16668
rect 31760 15972 31812 15978
rect 31760 15914 31812 15920
rect 32232 15706 32260 16662
rect 32324 16250 32352 16662
rect 32496 16584 32548 16590
rect 32496 16526 32548 16532
rect 32312 16244 32364 16250
rect 32364 16204 32444 16232
rect 32312 16186 32364 16192
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32036 15632 32088 15638
rect 32036 15574 32088 15580
rect 31944 15496 31996 15502
rect 31944 15438 31996 15444
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 31668 15156 31720 15162
rect 31668 15098 31720 15104
rect 31680 14958 31708 15098
rect 31668 14952 31720 14958
rect 31668 14894 31720 14900
rect 31772 14550 31800 15302
rect 31484 14544 31536 14550
rect 31484 14486 31536 14492
rect 31760 14544 31812 14550
rect 31760 14486 31812 14492
rect 31496 14006 31524 14486
rect 31484 14000 31536 14006
rect 31484 13942 31536 13948
rect 31576 13796 31628 13802
rect 31576 13738 31628 13744
rect 31588 13530 31616 13738
rect 31772 13530 31800 14486
rect 31956 14482 31984 15438
rect 32048 15162 32076 15574
rect 32036 15156 32088 15162
rect 32036 15098 32088 15104
rect 31944 14476 31996 14482
rect 31944 14418 31996 14424
rect 31852 14408 31904 14414
rect 31852 14350 31904 14356
rect 31864 13938 31892 14350
rect 31852 13932 31904 13938
rect 31852 13874 31904 13880
rect 32048 13802 32076 15098
rect 32324 14074 32352 16050
rect 32416 14550 32444 16204
rect 32508 16114 32536 16526
rect 32496 16108 32548 16114
rect 32496 16050 32548 16056
rect 32600 15638 32628 17002
rect 32588 15632 32640 15638
rect 32588 15574 32640 15580
rect 32600 15434 32628 15574
rect 32588 15428 32640 15434
rect 32588 15370 32640 15376
rect 32404 14544 32456 14550
rect 32404 14486 32456 14492
rect 32416 14074 32444 14486
rect 32496 14408 32548 14414
rect 32496 14350 32548 14356
rect 32312 14068 32364 14074
rect 32312 14010 32364 14016
rect 32404 14068 32456 14074
rect 32404 14010 32456 14016
rect 32036 13796 32088 13802
rect 32036 13738 32088 13744
rect 31576 13524 31628 13530
rect 31576 13466 31628 13472
rect 31760 13524 31812 13530
rect 31760 13466 31812 13472
rect 31392 13252 31444 13258
rect 31392 13194 31444 13200
rect 31300 12980 31352 12986
rect 31300 12922 31352 12928
rect 31300 12708 31352 12714
rect 31300 12650 31352 12656
rect 31576 12708 31628 12714
rect 31576 12650 31628 12656
rect 31668 12708 31720 12714
rect 31668 12650 31720 12656
rect 31312 12306 31340 12650
rect 31300 12300 31352 12306
rect 31300 12242 31352 12248
rect 31208 11688 31260 11694
rect 31208 11630 31260 11636
rect 30748 11348 30800 11354
rect 30748 11290 30800 11296
rect 29920 11280 29972 11286
rect 29920 11222 29972 11228
rect 29828 11144 29880 11150
rect 29828 11086 29880 11092
rect 29840 10810 29868 11086
rect 29932 10810 29960 11222
rect 29828 10804 29880 10810
rect 29828 10746 29880 10752
rect 29920 10804 29972 10810
rect 29920 10746 29972 10752
rect 28908 10260 28960 10266
rect 28908 10202 28960 10208
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28736 9586 28764 9998
rect 28920 9722 28948 10202
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 28816 9648 28868 9654
rect 28816 9590 28868 9596
rect 28724 9580 28776 9586
rect 28724 9522 28776 9528
rect 28724 9036 28776 9042
rect 28828 9024 28856 9590
rect 28920 9450 28948 9658
rect 29564 9586 29592 9998
rect 29932 9722 29960 10746
rect 30194 10704 30250 10713
rect 30194 10639 30250 10648
rect 30208 10606 30236 10639
rect 30196 10600 30248 10606
rect 30196 10542 30248 10548
rect 30760 10538 30788 11290
rect 31312 11082 31340 12242
rect 31588 12102 31616 12650
rect 31680 12442 31708 12650
rect 31668 12436 31720 12442
rect 31668 12378 31720 12384
rect 32036 12368 32088 12374
rect 32036 12310 32088 12316
rect 31576 12096 31628 12102
rect 31576 12038 31628 12044
rect 32048 11898 32076 12310
rect 32220 12232 32272 12238
rect 32220 12174 32272 12180
rect 32036 11892 32088 11898
rect 32036 11834 32088 11840
rect 31760 11688 31812 11694
rect 31760 11630 31812 11636
rect 31300 11076 31352 11082
rect 31300 11018 31352 11024
rect 31312 10742 31340 11018
rect 31300 10736 31352 10742
rect 31300 10678 31352 10684
rect 30748 10532 30800 10538
rect 30748 10474 30800 10480
rect 30840 10532 30892 10538
rect 30840 10474 30892 10480
rect 30852 10266 30880 10474
rect 30840 10260 30892 10266
rect 30840 10202 30892 10208
rect 31772 10130 31800 11630
rect 32048 11286 32076 11834
rect 32232 11762 32260 12174
rect 32220 11756 32272 11762
rect 32220 11698 32272 11704
rect 32036 11280 32088 11286
rect 32036 11222 32088 11228
rect 31944 11144 31996 11150
rect 31944 11086 31996 11092
rect 31956 10674 31984 11086
rect 32048 10810 32076 11222
rect 32324 11150 32352 14010
rect 32404 13796 32456 13802
rect 32404 13738 32456 13744
rect 32416 13190 32444 13738
rect 32508 13546 32536 14350
rect 32600 13682 32628 15370
rect 32680 14816 32732 14822
rect 32680 14758 32732 14764
rect 32692 14414 32720 14758
rect 32680 14408 32732 14414
rect 32680 14350 32732 14356
rect 32784 13734 32812 18022
rect 32876 14278 32904 20318
rect 32956 20256 33008 20262
rect 32956 20198 33008 20204
rect 32968 19514 32996 20198
rect 33244 19786 33272 33526
rect 33336 33114 33364 33895
rect 33520 33658 33548 34002
rect 33508 33652 33560 33658
rect 33508 33594 33560 33600
rect 33416 33312 33468 33318
rect 33416 33254 33468 33260
rect 33324 33108 33376 33114
rect 33324 33050 33376 33056
rect 33428 32434 33456 33254
rect 33508 33040 33560 33046
rect 33508 32982 33560 32988
rect 33520 32570 33548 32982
rect 33508 32564 33560 32570
rect 33508 32506 33560 32512
rect 33416 32428 33468 32434
rect 33416 32370 33468 32376
rect 33428 31958 33456 32370
rect 33520 32298 33548 32506
rect 33508 32292 33560 32298
rect 33508 32234 33560 32240
rect 33416 31952 33468 31958
rect 33416 31894 33468 31900
rect 33508 31952 33560 31958
rect 33508 31894 33560 31900
rect 33416 31272 33468 31278
rect 33416 31214 33468 31220
rect 33428 29170 33456 31214
rect 33520 31142 33548 31894
rect 33612 31822 33640 34410
rect 34072 33454 34100 36042
rect 34244 35556 34296 35562
rect 34244 35498 34296 35504
rect 34060 33448 34112 33454
rect 34060 33390 34112 33396
rect 33968 32904 34020 32910
rect 33968 32846 34020 32852
rect 33784 32836 33836 32842
rect 33784 32778 33836 32784
rect 33796 32434 33824 32778
rect 33784 32428 33836 32434
rect 33784 32370 33836 32376
rect 33600 31816 33652 31822
rect 33600 31758 33652 31764
rect 33796 31754 33824 32370
rect 33980 32026 34008 32846
rect 34072 32473 34100 33390
rect 34152 33108 34204 33114
rect 34152 33050 34204 33056
rect 34058 32464 34114 32473
rect 34058 32399 34114 32408
rect 33968 32020 34020 32026
rect 33968 31962 34020 31968
rect 33968 31816 34020 31822
rect 33968 31758 34020 31764
rect 33784 31748 33836 31754
rect 33784 31690 33836 31696
rect 33980 31482 34008 31758
rect 33968 31476 34020 31482
rect 33968 31418 34020 31424
rect 33508 31136 33560 31142
rect 33508 31078 33560 31084
rect 33520 30870 33548 31078
rect 33980 30938 34008 31418
rect 33968 30932 34020 30938
rect 33968 30874 34020 30880
rect 33508 30864 33560 30870
rect 33508 30806 33560 30812
rect 33520 30394 33548 30806
rect 33968 30728 34020 30734
rect 33968 30670 34020 30676
rect 33508 30388 33560 30394
rect 33508 30330 33560 30336
rect 33508 30252 33560 30258
rect 33508 30194 33560 30200
rect 33520 30122 33548 30194
rect 33508 30116 33560 30122
rect 33508 30058 33560 30064
rect 33980 29782 34008 30670
rect 33968 29776 34020 29782
rect 33874 29744 33930 29753
rect 33508 29708 33560 29714
rect 33968 29718 34020 29724
rect 33874 29679 33930 29688
rect 33508 29650 33560 29656
rect 33416 29164 33468 29170
rect 33416 29106 33468 29112
rect 33520 29034 33548 29650
rect 33888 29646 33916 29679
rect 33876 29640 33928 29646
rect 33876 29582 33928 29588
rect 33508 29028 33560 29034
rect 33508 28970 33560 28976
rect 33416 28688 33468 28694
rect 33416 28630 33468 28636
rect 33324 28552 33376 28558
rect 33324 28494 33376 28500
rect 33336 28218 33364 28494
rect 33324 28212 33376 28218
rect 33324 28154 33376 28160
rect 33428 27878 33456 28630
rect 33692 28552 33744 28558
rect 33692 28494 33744 28500
rect 33416 27872 33468 27878
rect 33416 27814 33468 27820
rect 33416 27464 33468 27470
rect 33416 27406 33468 27412
rect 33428 27130 33456 27406
rect 33416 27124 33468 27130
rect 33416 27066 33468 27072
rect 33324 26580 33376 26586
rect 33428 26568 33456 27066
rect 33376 26540 33456 26568
rect 33324 26522 33376 26528
rect 33416 26240 33468 26246
rect 33416 26182 33468 26188
rect 33428 25430 33456 26182
rect 33704 25906 33732 28494
rect 33784 27872 33836 27878
rect 33784 27814 33836 27820
rect 33796 27606 33824 27814
rect 33784 27600 33836 27606
rect 33784 27542 33836 27548
rect 33796 26790 33824 27542
rect 33784 26784 33836 26790
rect 33784 26726 33836 26732
rect 33796 26518 33824 26726
rect 33784 26512 33836 26518
rect 33784 26454 33836 26460
rect 33796 26042 33824 26454
rect 33876 26308 33928 26314
rect 33876 26250 33928 26256
rect 33784 26036 33836 26042
rect 33784 25978 33836 25984
rect 33692 25900 33744 25906
rect 33692 25842 33744 25848
rect 33416 25424 33468 25430
rect 33416 25366 33468 25372
rect 33428 24954 33456 25366
rect 33704 25294 33732 25842
rect 33888 25770 33916 26250
rect 34072 25838 34100 32399
rect 34164 31482 34192 33050
rect 34256 32910 34284 35498
rect 34532 35057 34560 40122
rect 34624 39574 34652 40870
rect 35268 40730 35296 41686
rect 35256 40724 35308 40730
rect 35256 40666 35308 40672
rect 34796 40588 34848 40594
rect 34796 40530 34848 40536
rect 34808 40186 34836 40530
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 34796 40180 34848 40186
rect 34796 40122 34848 40128
rect 35256 39976 35308 39982
rect 35256 39918 35308 39924
rect 34612 39568 34664 39574
rect 34612 39510 34664 39516
rect 34624 38962 34652 39510
rect 35268 39438 35296 39918
rect 35256 39432 35308 39438
rect 35256 39374 35308 39380
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 34612 38956 34664 38962
rect 34612 38898 34664 38904
rect 34624 37670 34652 38898
rect 35256 38888 35308 38894
rect 35256 38830 35308 38836
rect 35268 38214 35296 38830
rect 35256 38208 35308 38214
rect 35256 38150 35308 38156
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34796 37732 34848 37738
rect 34796 37674 34848 37680
rect 34612 37664 34664 37670
rect 34612 37606 34664 37612
rect 34624 37466 34652 37606
rect 34612 37460 34664 37466
rect 34612 37402 34664 37408
rect 34808 37126 34836 37674
rect 34796 37120 34848 37126
rect 34796 37062 34848 37068
rect 34612 36236 34664 36242
rect 34612 36178 34664 36184
rect 34624 35494 34652 36178
rect 34704 36032 34756 36038
rect 34704 35974 34756 35980
rect 34612 35488 34664 35494
rect 34612 35430 34664 35436
rect 34518 35048 34574 35057
rect 34518 34983 34574 34992
rect 34426 34096 34482 34105
rect 34426 34031 34428 34040
rect 34480 34031 34482 34040
rect 34428 34002 34480 34008
rect 34440 33658 34468 34002
rect 34428 33652 34480 33658
rect 34428 33594 34480 33600
rect 34244 32904 34296 32910
rect 34244 32846 34296 32852
rect 34152 31476 34204 31482
rect 34152 31418 34204 31424
rect 34164 31278 34192 31418
rect 34256 31346 34284 32846
rect 34440 31754 34468 33594
rect 34624 33590 34652 35430
rect 34716 35222 34744 35974
rect 34704 35216 34756 35222
rect 34704 35158 34756 35164
rect 34808 34202 34836 37062
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34796 34196 34848 34202
rect 34796 34138 34848 34144
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34612 33584 34664 33590
rect 34612 33526 34664 33532
rect 35268 33454 35296 38150
rect 35452 37262 35480 41958
rect 35544 41614 35572 42638
rect 35728 42362 35756 42774
rect 35898 42735 35954 42744
rect 35716 42356 35768 42362
rect 35716 42298 35768 42304
rect 35912 42294 35940 42735
rect 35624 42288 35676 42294
rect 35624 42230 35676 42236
rect 35900 42288 35952 42294
rect 35900 42230 35952 42236
rect 35532 41608 35584 41614
rect 35532 41550 35584 41556
rect 35544 41206 35572 41550
rect 35532 41200 35584 41206
rect 35532 41142 35584 41148
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 35440 36576 35492 36582
rect 35440 36518 35492 36524
rect 35348 35216 35400 35222
rect 35348 35158 35400 35164
rect 35360 34746 35388 35158
rect 35348 34740 35400 34746
rect 35348 34682 35400 34688
rect 35256 33448 35308 33454
rect 35256 33390 35308 33396
rect 35256 33312 35308 33318
rect 35256 33254 35308 33260
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34428 31748 34480 31754
rect 34428 31690 34480 31696
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34244 31340 34296 31346
rect 34244 31282 34296 31288
rect 34152 31272 34204 31278
rect 34152 31214 34204 31220
rect 34256 30734 34284 31282
rect 34244 30728 34296 30734
rect 34244 30670 34296 30676
rect 34612 30728 34664 30734
rect 34612 30670 34664 30676
rect 34152 30388 34204 30394
rect 34152 30330 34204 30336
rect 34164 29850 34192 30330
rect 34624 29850 34652 30670
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 35268 30190 35296 33254
rect 35348 31884 35400 31890
rect 35348 31826 35400 31832
rect 35360 31686 35388 31826
rect 35348 31680 35400 31686
rect 35348 31622 35400 31628
rect 35360 30598 35388 31622
rect 35452 31346 35480 36518
rect 35636 35170 35664 42230
rect 36188 42158 36216 43007
rect 37108 42770 37136 43318
rect 37096 42764 37148 42770
rect 37096 42706 37148 42712
rect 35808 42152 35860 42158
rect 35808 42094 35860 42100
rect 36176 42152 36228 42158
rect 36176 42094 36228 42100
rect 35716 40520 35768 40526
rect 35716 40462 35768 40468
rect 35728 39982 35756 40462
rect 35820 40050 35848 42094
rect 37740 42016 37792 42022
rect 37740 41958 37792 41964
rect 36636 41472 36688 41478
rect 36636 41414 36688 41420
rect 36648 41070 36676 41414
rect 37752 41274 37780 41958
rect 37740 41268 37792 41274
rect 37740 41210 37792 41216
rect 36636 41064 36688 41070
rect 36636 41006 36688 41012
rect 36544 40928 36596 40934
rect 36544 40870 36596 40876
rect 36268 40588 36320 40594
rect 36268 40530 36320 40536
rect 36280 40186 36308 40530
rect 36268 40180 36320 40186
rect 36268 40122 36320 40128
rect 35808 40044 35860 40050
rect 35808 39986 35860 39992
rect 35716 39976 35768 39982
rect 35716 39918 35768 39924
rect 35728 39302 35756 39918
rect 35716 39296 35768 39302
rect 35716 39238 35768 39244
rect 35728 38894 35756 39238
rect 35716 38888 35768 38894
rect 35716 38830 35768 38836
rect 35728 38486 35756 38830
rect 35716 38480 35768 38486
rect 35716 38422 35768 38428
rect 35820 38332 35848 39986
rect 36176 39500 36228 39506
rect 36176 39442 36228 39448
rect 35900 38820 35952 38826
rect 35900 38762 35952 38768
rect 35912 38350 35940 38762
rect 36188 38758 36216 39442
rect 36176 38752 36228 38758
rect 36176 38694 36228 38700
rect 36084 38412 36136 38418
rect 36084 38354 36136 38360
rect 35728 38304 35848 38332
rect 35900 38344 35952 38350
rect 35728 36553 35756 38304
rect 35900 38286 35952 38292
rect 36096 37942 36124 38354
rect 36084 37936 36136 37942
rect 36084 37878 36136 37884
rect 36096 37670 36124 37878
rect 36084 37664 36136 37670
rect 36084 37606 36136 37612
rect 35898 37360 35954 37369
rect 35808 37324 35860 37330
rect 35898 37295 35954 37304
rect 35992 37324 36044 37330
rect 35808 37266 35860 37272
rect 35820 36922 35848 37266
rect 35912 37262 35940 37295
rect 35992 37266 36044 37272
rect 35900 37256 35952 37262
rect 35900 37198 35952 37204
rect 35808 36916 35860 36922
rect 35808 36858 35860 36864
rect 35714 36544 35770 36553
rect 35714 36479 35770 36488
rect 35820 35834 35848 36858
rect 36004 36718 36032 37266
rect 35992 36712 36044 36718
rect 35992 36654 36044 36660
rect 35900 36372 35952 36378
rect 35900 36314 35952 36320
rect 35808 35828 35860 35834
rect 35808 35770 35860 35776
rect 35544 35142 35664 35170
rect 35716 35216 35768 35222
rect 35716 35158 35768 35164
rect 35544 34542 35572 35142
rect 35624 35080 35676 35086
rect 35624 35022 35676 35028
rect 35636 34678 35664 35022
rect 35728 34678 35756 35158
rect 35624 34672 35676 34678
rect 35624 34614 35676 34620
rect 35716 34672 35768 34678
rect 35716 34614 35768 34620
rect 35532 34536 35584 34542
rect 35532 34478 35584 34484
rect 35532 33856 35584 33862
rect 35532 33798 35584 33804
rect 35544 32910 35572 33798
rect 35820 33134 35848 35770
rect 35912 35630 35940 36314
rect 36096 36242 36124 37606
rect 36176 37256 36228 37262
rect 36176 37198 36228 37204
rect 36188 36922 36216 37198
rect 36176 36916 36228 36922
rect 36176 36858 36228 36864
rect 36280 36378 36308 40122
rect 36556 39846 36584 40870
rect 36648 40662 36676 41006
rect 36636 40656 36688 40662
rect 36636 40598 36688 40604
rect 38028 40594 38056 44338
rect 41142 44296 41198 44305
rect 41142 44231 41198 44240
rect 38200 42764 38252 42770
rect 38200 42706 38252 42712
rect 39856 42764 39908 42770
rect 39856 42706 39908 42712
rect 38212 42022 38240 42706
rect 39764 42628 39816 42634
rect 39764 42570 39816 42576
rect 38476 42560 38528 42566
rect 38476 42502 38528 42508
rect 38568 42560 38620 42566
rect 38568 42502 38620 42508
rect 38488 42226 38516 42502
rect 38476 42220 38528 42226
rect 38476 42162 38528 42168
rect 38580 42090 38608 42502
rect 38292 42084 38344 42090
rect 38292 42026 38344 42032
rect 38568 42084 38620 42090
rect 38568 42026 38620 42032
rect 38200 42016 38252 42022
rect 38200 41958 38252 41964
rect 38016 40588 38068 40594
rect 38016 40530 38068 40536
rect 38028 40186 38056 40530
rect 38016 40180 38068 40186
rect 38016 40122 38068 40128
rect 36912 39976 36964 39982
rect 36912 39918 36964 39924
rect 36544 39840 36596 39846
rect 36544 39782 36596 39788
rect 36924 39642 36952 39918
rect 37004 39840 37056 39846
rect 37004 39782 37056 39788
rect 37740 39840 37792 39846
rect 37740 39782 37792 39788
rect 36912 39636 36964 39642
rect 36912 39578 36964 39584
rect 36636 39432 36688 39438
rect 36636 39374 36688 39380
rect 36648 38962 36676 39374
rect 36636 38956 36688 38962
rect 36636 38898 36688 38904
rect 36360 38752 36412 38758
rect 36360 38694 36412 38700
rect 36372 38457 36400 38694
rect 36648 38554 36676 38898
rect 36912 38752 36964 38758
rect 37016 38740 37044 39782
rect 37752 39574 37780 39782
rect 37740 39568 37792 39574
rect 37740 39510 37792 39516
rect 37096 38752 37148 38758
rect 36964 38720 37096 38740
rect 36964 38712 37002 38720
rect 36912 38694 36964 38700
rect 37058 38712 37096 38720
rect 37096 38694 37148 38700
rect 37002 38655 37058 38664
rect 36636 38548 36688 38554
rect 36636 38490 36688 38496
rect 37016 38486 37044 38655
rect 37004 38480 37056 38486
rect 36358 38448 36414 38457
rect 37004 38422 37056 38428
rect 36358 38383 36414 38392
rect 36544 38412 36596 38418
rect 36268 36372 36320 36378
rect 36268 36314 36320 36320
rect 36084 36236 36136 36242
rect 36084 36178 36136 36184
rect 35900 35624 35952 35630
rect 35900 35566 35952 35572
rect 35912 33386 35940 35566
rect 36096 34950 36124 36178
rect 36084 34944 36136 34950
rect 36084 34886 36136 34892
rect 35900 33380 35952 33386
rect 35900 33322 35952 33328
rect 35728 33106 35848 33134
rect 35532 32904 35584 32910
rect 35532 32846 35584 32852
rect 35544 32570 35572 32846
rect 35624 32768 35676 32774
rect 35624 32710 35676 32716
rect 35532 32564 35584 32570
rect 35532 32506 35584 32512
rect 35636 32502 35664 32710
rect 35624 32496 35676 32502
rect 35624 32438 35676 32444
rect 35440 31340 35492 31346
rect 35440 31282 35492 31288
rect 35452 30938 35480 31282
rect 35440 30932 35492 30938
rect 35440 30874 35492 30880
rect 35348 30592 35400 30598
rect 35348 30534 35400 30540
rect 35256 30184 35308 30190
rect 35256 30126 35308 30132
rect 34152 29844 34204 29850
rect 34152 29786 34204 29792
rect 34612 29844 34664 29850
rect 34612 29786 34664 29792
rect 35256 29844 35308 29850
rect 35256 29786 35308 29792
rect 34624 29306 34652 29786
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34612 29300 34664 29306
rect 34612 29242 34664 29248
rect 35268 29102 35296 29786
rect 34152 29096 34204 29102
rect 34152 29038 34204 29044
rect 35256 29096 35308 29102
rect 35256 29038 35308 29044
rect 34164 28966 34192 29038
rect 34152 28960 34204 28966
rect 34152 28902 34204 28908
rect 34164 28014 34192 28902
rect 35268 28694 35296 29038
rect 35256 28688 35308 28694
rect 34610 28656 34666 28665
rect 35256 28630 35308 28636
rect 34610 28591 34612 28600
rect 34664 28591 34666 28600
rect 34612 28562 34664 28568
rect 34624 28150 34652 28562
rect 34794 28384 34850 28393
rect 34794 28319 34850 28328
rect 34612 28144 34664 28150
rect 34612 28086 34664 28092
rect 34152 28008 34204 28014
rect 34152 27950 34204 27956
rect 34428 27464 34480 27470
rect 34428 27406 34480 27412
rect 34440 27334 34468 27406
rect 34428 27328 34480 27334
rect 34428 27270 34480 27276
rect 34060 25832 34112 25838
rect 34060 25774 34112 25780
rect 33876 25764 33928 25770
rect 33876 25706 33928 25712
rect 33692 25288 33744 25294
rect 33692 25230 33744 25236
rect 33416 24948 33468 24954
rect 33416 24890 33468 24896
rect 34336 24880 34388 24886
rect 34336 24822 34388 24828
rect 33598 24712 33654 24721
rect 33598 24647 33654 24656
rect 34152 24676 34204 24682
rect 33416 24336 33468 24342
rect 33416 24278 33468 24284
rect 33428 23594 33456 24278
rect 33324 23588 33376 23594
rect 33324 23530 33376 23536
rect 33416 23588 33468 23594
rect 33416 23530 33468 23536
rect 33336 23118 33364 23530
rect 33428 23322 33456 23530
rect 33416 23316 33468 23322
rect 33416 23258 33468 23264
rect 33508 23248 33560 23254
rect 33508 23190 33560 23196
rect 33324 23112 33376 23118
rect 33324 23054 33376 23060
rect 33336 22234 33364 23054
rect 33520 22778 33548 23190
rect 33508 22772 33560 22778
rect 33508 22714 33560 22720
rect 33612 22574 33640 24647
rect 34152 24618 34204 24624
rect 34164 23746 34192 24618
rect 34244 24268 34296 24274
rect 34244 24210 34296 24216
rect 34256 23866 34284 24210
rect 34244 23860 34296 23866
rect 34244 23802 34296 23808
rect 34164 23718 34284 23746
rect 34152 23588 34204 23594
rect 34152 23530 34204 23536
rect 34164 23118 34192 23530
rect 33968 23112 34020 23118
rect 33968 23054 34020 23060
rect 34152 23112 34204 23118
rect 34152 23054 34204 23060
rect 33980 22778 34008 23054
rect 33968 22772 34020 22778
rect 33968 22714 34020 22720
rect 33600 22568 33652 22574
rect 33600 22510 33652 22516
rect 33324 22228 33376 22234
rect 33324 22170 33376 22176
rect 34164 22030 34192 23054
rect 34256 22438 34284 23718
rect 34348 23526 34376 24822
rect 34440 24818 34468 27270
rect 34808 26450 34836 28319
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 35360 27538 35388 30534
rect 35452 28762 35480 30874
rect 35440 28756 35492 28762
rect 35440 28698 35492 28704
rect 35348 27532 35400 27538
rect 35348 27474 35400 27480
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 35360 26586 35388 27474
rect 35452 26926 35480 28698
rect 35636 28626 35664 32438
rect 35728 31890 35756 33106
rect 35808 32904 35860 32910
rect 35808 32846 35860 32852
rect 35716 31884 35768 31890
rect 35716 31826 35768 31832
rect 35820 30734 35848 32846
rect 35992 31884 36044 31890
rect 35992 31826 36044 31832
rect 36004 31482 36032 31826
rect 35992 31476 36044 31482
rect 35992 31418 36044 31424
rect 36004 31278 36032 31418
rect 35992 31272 36044 31278
rect 35992 31214 36044 31220
rect 35808 30728 35860 30734
rect 35808 30670 35860 30676
rect 35992 30048 36044 30054
rect 35992 29990 36044 29996
rect 36004 29782 36032 29990
rect 36096 29850 36124 34886
rect 36372 34066 36400 38383
rect 36544 38354 36596 38360
rect 36556 37738 36584 38354
rect 37016 38010 37044 38422
rect 37924 38344 37976 38350
rect 37924 38286 37976 38292
rect 37004 38004 37056 38010
rect 37004 37946 37056 37952
rect 37016 37806 37044 37946
rect 37556 37868 37608 37874
rect 37556 37810 37608 37816
rect 37832 37868 37884 37874
rect 37832 37810 37884 37816
rect 37004 37800 37056 37806
rect 37004 37742 37056 37748
rect 36544 37732 36596 37738
rect 36544 37674 36596 37680
rect 36636 36576 36688 36582
rect 36636 36518 36688 36524
rect 36728 36576 36780 36582
rect 36728 36518 36780 36524
rect 36648 36242 36676 36518
rect 36544 36236 36596 36242
rect 36544 36178 36596 36184
rect 36636 36236 36688 36242
rect 36636 36178 36688 36184
rect 36556 35494 36584 36178
rect 36544 35488 36596 35494
rect 36544 35430 36596 35436
rect 36556 34066 36584 35430
rect 36360 34060 36412 34066
rect 36360 34002 36412 34008
rect 36544 34060 36596 34066
rect 36544 34002 36596 34008
rect 36372 33658 36400 34002
rect 36360 33652 36412 33658
rect 36360 33594 36412 33600
rect 36372 33134 36400 33594
rect 36556 33454 36584 34002
rect 36544 33448 36596 33454
rect 36544 33390 36596 33396
rect 36188 33106 36400 33134
rect 36188 31686 36216 33106
rect 36556 32842 36584 33390
rect 36544 32836 36596 32842
rect 36544 32778 36596 32784
rect 36452 32360 36504 32366
rect 36556 32348 36584 32778
rect 36740 32774 36768 36518
rect 36820 36168 36872 36174
rect 36820 36110 36872 36116
rect 36832 35698 36860 36110
rect 37016 35834 37044 37742
rect 37096 37732 37148 37738
rect 37096 37674 37148 37680
rect 37108 37126 37136 37674
rect 37568 37126 37596 37810
rect 37844 37777 37872 37810
rect 37830 37768 37886 37777
rect 37830 37703 37886 37712
rect 37936 37466 37964 38286
rect 37924 37460 37976 37466
rect 37924 37402 37976 37408
rect 37096 37120 37148 37126
rect 37096 37062 37148 37068
rect 37556 37120 37608 37126
rect 37556 37062 37608 37068
rect 37108 36718 37136 37062
rect 37568 36786 37596 37062
rect 37556 36780 37608 36786
rect 37556 36722 37608 36728
rect 37096 36712 37148 36718
rect 37096 36654 37148 36660
rect 37924 36712 37976 36718
rect 37924 36654 37976 36660
rect 37936 36378 37964 36654
rect 37924 36372 37976 36378
rect 37924 36314 37976 36320
rect 37004 35828 37056 35834
rect 37004 35770 37056 35776
rect 36820 35692 36872 35698
rect 36820 35634 36872 35640
rect 37016 35562 37044 35770
rect 38028 35630 38056 40122
rect 38108 38752 38160 38758
rect 38108 38694 38160 38700
rect 38120 38010 38148 38694
rect 38108 38004 38160 38010
rect 38108 37946 38160 37952
rect 37280 35624 37332 35630
rect 37280 35566 37332 35572
rect 38016 35624 38068 35630
rect 38016 35566 38068 35572
rect 37004 35556 37056 35562
rect 37004 35498 37056 35504
rect 37016 34746 37044 35498
rect 37292 35290 37320 35566
rect 37280 35284 37332 35290
rect 37280 35226 37332 35232
rect 38212 35222 38240 41958
rect 38304 36718 38332 42026
rect 38580 41750 38608 42026
rect 38568 41744 38620 41750
rect 38488 41704 38568 41732
rect 38488 41002 38516 41704
rect 38568 41686 38620 41692
rect 38568 41608 38620 41614
rect 38568 41550 38620 41556
rect 38580 41138 38608 41550
rect 38660 41540 38712 41546
rect 38660 41482 38712 41488
rect 38568 41132 38620 41138
rect 38568 41074 38620 41080
rect 38476 40996 38528 41002
rect 38476 40938 38528 40944
rect 38488 40594 38516 40938
rect 38580 40730 38608 41074
rect 38568 40724 38620 40730
rect 38568 40666 38620 40672
rect 38476 40588 38528 40594
rect 38476 40530 38528 40536
rect 38568 39568 38620 39574
rect 38568 39510 38620 39516
rect 38580 39098 38608 39510
rect 38672 39438 38700 41482
rect 39120 40996 39172 41002
rect 39120 40938 39172 40944
rect 38752 40384 38804 40390
rect 38752 40326 38804 40332
rect 38764 39914 38792 40326
rect 39132 40186 39160 40938
rect 39776 40594 39804 42570
rect 39868 42362 39896 42706
rect 40316 42560 40368 42566
rect 40316 42502 40368 42508
rect 39856 42356 39908 42362
rect 39856 42298 39908 42304
rect 40132 42084 40184 42090
rect 40132 42026 40184 42032
rect 40144 41614 40172 42026
rect 40328 41750 40356 42502
rect 40776 42016 40828 42022
rect 40776 41958 40828 41964
rect 40316 41744 40368 41750
rect 40316 41686 40368 41692
rect 40408 41744 40460 41750
rect 40408 41686 40460 41692
rect 40132 41608 40184 41614
rect 40184 41568 40264 41596
rect 40132 41550 40184 41556
rect 39948 40928 40000 40934
rect 39948 40870 40000 40876
rect 39764 40588 39816 40594
rect 39764 40530 39816 40536
rect 39120 40180 39172 40186
rect 39120 40122 39172 40128
rect 39776 40118 39804 40530
rect 39764 40112 39816 40118
rect 39764 40054 39816 40060
rect 38752 39908 38804 39914
rect 38752 39850 38804 39856
rect 39304 39908 39356 39914
rect 39304 39850 39356 39856
rect 38660 39432 38712 39438
rect 38660 39374 38712 39380
rect 38568 39092 38620 39098
rect 38568 39034 38620 39040
rect 38672 38350 38700 39374
rect 38764 39030 38792 39850
rect 39316 39370 39344 39850
rect 39304 39364 39356 39370
rect 39304 39306 39356 39312
rect 39316 39030 39344 39306
rect 38752 39024 38804 39030
rect 38752 38966 38804 38972
rect 39304 39024 39356 39030
rect 39304 38966 39356 38972
rect 38752 38820 38804 38826
rect 38752 38762 38804 38768
rect 38764 38486 38792 38762
rect 38752 38480 38804 38486
rect 38752 38422 38804 38428
rect 39120 38480 39172 38486
rect 39120 38422 39172 38428
rect 38660 38344 38712 38350
rect 38660 38286 38712 38292
rect 38660 37256 38712 37262
rect 38660 37198 38712 37204
rect 38672 36854 38700 37198
rect 38764 36854 38792 38422
rect 39132 37738 39160 38422
rect 39316 38010 39344 38966
rect 39488 38412 39540 38418
rect 39488 38354 39540 38360
rect 39500 38010 39528 38354
rect 39304 38004 39356 38010
rect 39304 37946 39356 37952
rect 39488 38004 39540 38010
rect 39488 37946 39540 37952
rect 39120 37732 39172 37738
rect 39120 37674 39172 37680
rect 39132 37398 39160 37674
rect 39960 37466 39988 40870
rect 40132 39568 40184 39574
rect 40052 39528 40132 39556
rect 40052 38758 40080 39528
rect 40132 39510 40184 39516
rect 40236 39438 40264 41568
rect 40328 40730 40356 41686
rect 40420 40934 40448 41686
rect 40788 41138 40816 41958
rect 40868 41540 40920 41546
rect 40868 41482 40920 41488
rect 40880 41138 40908 41482
rect 40776 41132 40828 41138
rect 40776 41074 40828 41080
rect 40868 41132 40920 41138
rect 40868 41074 40920 41080
rect 40408 40928 40460 40934
rect 40408 40870 40460 40876
rect 40788 40730 40816 41074
rect 40316 40724 40368 40730
rect 40316 40666 40368 40672
rect 40776 40724 40828 40730
rect 40776 40666 40828 40672
rect 40880 40050 40908 41074
rect 40868 40044 40920 40050
rect 40868 39986 40920 39992
rect 41156 39982 41184 44231
rect 41432 42634 41460 49558
rect 41602 49520 41658 49558
rect 46952 49558 47178 49586
rect 41420 42628 41472 42634
rect 41420 42570 41472 42576
rect 42248 41744 42300 41750
rect 42248 41686 42300 41692
rect 42064 41676 42116 41682
rect 42064 41618 42116 41624
rect 41696 40996 41748 41002
rect 41696 40938 41748 40944
rect 41708 40662 41736 40938
rect 42076 40934 42104 41618
rect 42156 41472 42208 41478
rect 42156 41414 42208 41420
rect 42064 40928 42116 40934
rect 42064 40870 42116 40876
rect 41696 40656 41748 40662
rect 41696 40598 41748 40604
rect 41788 40656 41840 40662
rect 41788 40598 41840 40604
rect 41604 40452 41656 40458
rect 41604 40394 41656 40400
rect 41328 40112 41380 40118
rect 41328 40054 41380 40060
rect 41144 39976 41196 39982
rect 41064 39936 41144 39964
rect 40960 39840 41012 39846
rect 40960 39782 41012 39788
rect 40972 39574 41000 39782
rect 40960 39568 41012 39574
rect 40960 39510 41012 39516
rect 40224 39432 40276 39438
rect 40224 39374 40276 39380
rect 40236 39098 40264 39374
rect 40224 39092 40276 39098
rect 40224 39034 40276 39040
rect 40040 38752 40092 38758
rect 40040 38694 40092 38700
rect 40052 38554 40080 38694
rect 40040 38548 40092 38554
rect 40040 38490 40092 38496
rect 40408 37800 40460 37806
rect 40408 37742 40460 37748
rect 39948 37460 40000 37466
rect 39948 37402 40000 37408
rect 39120 37392 39172 37398
rect 39120 37334 39172 37340
rect 38660 36848 38712 36854
rect 38660 36790 38712 36796
rect 38752 36848 38804 36854
rect 38752 36790 38804 36796
rect 39132 36786 39160 37334
rect 40420 37233 40448 37742
rect 40684 37460 40736 37466
rect 40684 37402 40736 37408
rect 40406 37224 40462 37233
rect 40406 37159 40462 37168
rect 40592 37188 40644 37194
rect 40592 37130 40644 37136
rect 40604 36786 40632 37130
rect 39120 36780 39172 36786
rect 39120 36722 39172 36728
rect 40592 36780 40644 36786
rect 40592 36722 40644 36728
rect 38292 36712 38344 36718
rect 38292 36654 38344 36660
rect 38936 36576 38988 36582
rect 38936 36518 38988 36524
rect 38948 36310 38976 36518
rect 38936 36304 38988 36310
rect 38936 36246 38988 36252
rect 38476 36236 38528 36242
rect 38476 36178 38528 36184
rect 38488 35834 38516 36178
rect 38948 35834 38976 36246
rect 38476 35828 38528 35834
rect 38476 35770 38528 35776
rect 38936 35828 38988 35834
rect 38936 35770 38988 35776
rect 39132 35494 39160 36722
rect 40696 36650 40724 37402
rect 40776 37256 40828 37262
rect 40776 37198 40828 37204
rect 40788 36922 40816 37198
rect 40776 36916 40828 36922
rect 40776 36858 40828 36864
rect 40684 36644 40736 36650
rect 40684 36586 40736 36592
rect 39580 36576 39632 36582
rect 39580 36518 39632 36524
rect 39212 36304 39264 36310
rect 39212 36246 39264 36252
rect 39224 35562 39252 36246
rect 39396 36168 39448 36174
rect 39396 36110 39448 36116
rect 39212 35556 39264 35562
rect 39212 35498 39264 35504
rect 39120 35488 39172 35494
rect 39120 35430 39172 35436
rect 39224 35222 39252 35498
rect 38200 35216 38252 35222
rect 38200 35158 38252 35164
rect 39212 35216 39264 35222
rect 39212 35158 39264 35164
rect 37004 34740 37056 34746
rect 37004 34682 37056 34688
rect 36820 34536 36872 34542
rect 36820 34478 36872 34484
rect 36832 34134 36860 34478
rect 37016 34406 37044 34682
rect 38212 34406 38240 35158
rect 39120 35080 39172 35086
rect 38382 35048 38438 35057
rect 39120 35022 39172 35028
rect 38382 34983 38438 34992
rect 38844 35012 38896 35018
rect 37004 34400 37056 34406
rect 37004 34342 37056 34348
rect 37924 34400 37976 34406
rect 37924 34342 37976 34348
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 37016 34134 37044 34342
rect 36820 34128 36872 34134
rect 36820 34070 36872 34076
rect 37004 34128 37056 34134
rect 37004 34070 37056 34076
rect 37832 34128 37884 34134
rect 37832 34070 37884 34076
rect 37740 33992 37792 33998
rect 37740 33934 37792 33940
rect 37752 33522 37780 33934
rect 37844 33658 37872 34070
rect 37936 33658 37964 34342
rect 37832 33652 37884 33658
rect 37832 33594 37884 33600
rect 37924 33652 37976 33658
rect 37924 33594 37976 33600
rect 37740 33516 37792 33522
rect 37740 33458 37792 33464
rect 36912 33380 36964 33386
rect 36912 33322 36964 33328
rect 36924 33046 36952 33322
rect 36912 33040 36964 33046
rect 36912 32982 36964 32988
rect 36728 32768 36780 32774
rect 36728 32710 36780 32716
rect 36504 32320 36584 32348
rect 36452 32302 36504 32308
rect 36176 31680 36228 31686
rect 36176 31622 36228 31628
rect 36084 29844 36136 29850
rect 36084 29786 36136 29792
rect 35992 29776 36044 29782
rect 35992 29718 36044 29724
rect 36004 29102 36032 29718
rect 36084 29708 36136 29714
rect 36188 29696 36216 31622
rect 36464 31482 36492 32302
rect 36452 31476 36504 31482
rect 36452 31418 36504 31424
rect 36452 31272 36504 31278
rect 36452 31214 36504 31220
rect 36464 30938 36492 31214
rect 36452 30932 36504 30938
rect 36452 30874 36504 30880
rect 36464 30666 36492 30874
rect 36452 30660 36504 30666
rect 36452 30602 36504 30608
rect 36464 30394 36492 30602
rect 36452 30388 36504 30394
rect 36452 30330 36504 30336
rect 36464 30190 36492 30330
rect 36924 30326 36952 32982
rect 37740 32972 37792 32978
rect 37740 32914 37792 32920
rect 37372 32360 37424 32366
rect 37372 32302 37424 32308
rect 37384 32026 37412 32302
rect 37372 32020 37424 32026
rect 37372 31962 37424 31968
rect 37752 31958 37780 32914
rect 37844 32230 37872 33594
rect 38108 33312 38160 33318
rect 38108 33254 38160 33260
rect 38120 33153 38148 33254
rect 38106 33144 38162 33153
rect 38028 33102 38106 33130
rect 37832 32224 37884 32230
rect 37832 32166 37884 32172
rect 37844 31958 37872 32166
rect 37740 31952 37792 31958
rect 37740 31894 37792 31900
rect 37832 31952 37884 31958
rect 37832 31894 37884 31900
rect 37740 31816 37792 31822
rect 37740 31758 37792 31764
rect 37752 31482 37780 31758
rect 37740 31476 37792 31482
rect 37740 31418 37792 31424
rect 37832 31136 37884 31142
rect 37832 31078 37884 31084
rect 37740 30796 37792 30802
rect 37740 30738 37792 30744
rect 36912 30320 36964 30326
rect 36912 30262 36964 30268
rect 36452 30184 36504 30190
rect 36452 30126 36504 30132
rect 36136 29668 36216 29696
rect 36084 29650 36136 29656
rect 35992 29096 36044 29102
rect 35992 29038 36044 29044
rect 35716 29028 35768 29034
rect 35716 28970 35768 28976
rect 35624 28620 35676 28626
rect 35624 28562 35676 28568
rect 35636 28218 35664 28562
rect 35624 28212 35676 28218
rect 35624 28154 35676 28160
rect 35728 28082 35756 28970
rect 36004 28626 36032 29038
rect 36096 29034 36124 29650
rect 36820 29640 36872 29646
rect 36820 29582 36872 29588
rect 36084 29028 36136 29034
rect 36084 28970 36136 28976
rect 36096 28937 36124 28970
rect 36082 28928 36138 28937
rect 36082 28863 36138 28872
rect 36832 28626 36860 29582
rect 36924 29102 36952 30262
rect 37280 30116 37332 30122
rect 37280 30058 37332 30064
rect 37556 30116 37608 30122
rect 37556 30058 37608 30064
rect 37188 29640 37240 29646
rect 37188 29582 37240 29588
rect 37200 29170 37228 29582
rect 37292 29170 37320 30058
rect 37568 29714 37596 30058
rect 37752 30054 37780 30738
rect 37740 30048 37792 30054
rect 37740 29990 37792 29996
rect 37648 29844 37700 29850
rect 37648 29786 37700 29792
rect 37556 29708 37608 29714
rect 37556 29650 37608 29656
rect 37568 29306 37596 29650
rect 37556 29300 37608 29306
rect 37556 29242 37608 29248
rect 37188 29164 37240 29170
rect 37188 29106 37240 29112
rect 37280 29164 37332 29170
rect 37280 29106 37332 29112
rect 37568 29102 37596 29242
rect 36912 29096 36964 29102
rect 36912 29038 36964 29044
rect 37556 29096 37608 29102
rect 37556 29038 37608 29044
rect 36924 28762 36952 29038
rect 37660 28966 37688 29786
rect 37648 28960 37700 28966
rect 37648 28902 37700 28908
rect 36912 28756 36964 28762
rect 36912 28698 36964 28704
rect 35992 28620 36044 28626
rect 35992 28562 36044 28568
rect 36820 28620 36872 28626
rect 36820 28562 36872 28568
rect 35808 28144 35860 28150
rect 35808 28086 35860 28092
rect 35716 28076 35768 28082
rect 35716 28018 35768 28024
rect 35716 27532 35768 27538
rect 35716 27474 35768 27480
rect 35728 26926 35756 27474
rect 35440 26920 35492 26926
rect 35440 26862 35492 26868
rect 35716 26920 35768 26926
rect 35716 26862 35768 26868
rect 35728 26586 35756 26862
rect 35348 26580 35400 26586
rect 35348 26522 35400 26528
rect 35716 26580 35768 26586
rect 35716 26522 35768 26528
rect 34796 26444 34848 26450
rect 34796 26386 34848 26392
rect 34808 26042 34836 26386
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34796 26036 34848 26042
rect 34796 25978 34848 25984
rect 35348 26036 35400 26042
rect 35348 25978 35400 25984
rect 35164 25764 35216 25770
rect 35164 25706 35216 25712
rect 34704 25696 34756 25702
rect 34704 25638 34756 25644
rect 34716 25294 34744 25638
rect 35176 25294 35204 25706
rect 35256 25424 35308 25430
rect 35256 25366 35308 25372
rect 34704 25288 34756 25294
rect 34704 25230 34756 25236
rect 35164 25288 35216 25294
rect 35164 25230 35216 25236
rect 34520 25152 34572 25158
rect 34520 25094 34572 25100
rect 34428 24812 34480 24818
rect 34428 24754 34480 24760
rect 34532 24682 34560 25094
rect 34520 24676 34572 24682
rect 34520 24618 34572 24624
rect 34532 24410 34560 24618
rect 34716 24410 34744 25230
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 35268 24682 35296 25366
rect 35256 24676 35308 24682
rect 35256 24618 35308 24624
rect 34520 24404 34572 24410
rect 34520 24346 34572 24352
rect 34704 24404 34756 24410
rect 34704 24346 34756 24352
rect 34612 24336 34664 24342
rect 34612 24278 34664 24284
rect 34624 23866 34652 24278
rect 35256 24132 35308 24138
rect 35256 24074 35308 24080
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34612 23860 34664 23866
rect 34612 23802 34664 23808
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34336 23520 34388 23526
rect 34336 23462 34388 23468
rect 34624 22506 34652 23666
rect 34796 23588 34848 23594
rect 34796 23530 34848 23536
rect 34704 23520 34756 23526
rect 34704 23462 34756 23468
rect 34716 23254 34744 23462
rect 34704 23248 34756 23254
rect 34704 23190 34756 23196
rect 34716 22778 34744 23190
rect 34808 23050 34836 23530
rect 35268 23322 35296 24074
rect 35256 23316 35308 23322
rect 35256 23258 35308 23264
rect 34796 23044 34848 23050
rect 34796 22986 34848 22992
rect 34808 22778 34836 22986
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 34704 22772 34756 22778
rect 34704 22714 34756 22720
rect 34796 22772 34848 22778
rect 34796 22714 34848 22720
rect 35360 22624 35388 25978
rect 35820 25344 35848 28086
rect 36004 27674 36032 28562
rect 36452 28552 36504 28558
rect 36452 28494 36504 28500
rect 36176 27872 36228 27878
rect 36176 27814 36228 27820
rect 35992 27668 36044 27674
rect 35992 27610 36044 27616
rect 35900 27464 35952 27470
rect 35900 27406 35952 27412
rect 35912 26450 35940 27406
rect 35992 27328 36044 27334
rect 35992 27270 36044 27276
rect 35900 26444 35952 26450
rect 35900 26386 35952 26392
rect 35728 25316 35848 25344
rect 35440 24132 35492 24138
rect 35440 24074 35492 24080
rect 35452 23730 35480 24074
rect 35440 23724 35492 23730
rect 35440 23666 35492 23672
rect 35452 23474 35480 23666
rect 35728 23474 35756 25316
rect 35808 25220 35860 25226
rect 35808 25162 35860 25168
rect 35820 24274 35848 25162
rect 35912 24954 35940 26386
rect 35900 24948 35952 24954
rect 35900 24890 35952 24896
rect 35808 24268 35860 24274
rect 35808 24210 35860 24216
rect 35452 23446 35664 23474
rect 35728 23446 35940 23474
rect 35268 22596 35388 22624
rect 34612 22500 34664 22506
rect 34612 22442 34664 22448
rect 34244 22432 34296 22438
rect 34244 22374 34296 22380
rect 33876 22024 33928 22030
rect 33876 21966 33928 21972
rect 34152 22024 34204 22030
rect 34152 21966 34204 21972
rect 33888 21690 33916 21966
rect 33876 21684 33928 21690
rect 33876 21626 33928 21632
rect 33600 21548 33652 21554
rect 33600 21490 33652 21496
rect 33612 21457 33640 21490
rect 33598 21448 33654 21457
rect 33598 21383 33654 21392
rect 33416 21004 33468 21010
rect 33416 20946 33468 20952
rect 33428 20058 33456 20946
rect 33784 20528 33836 20534
rect 33784 20470 33836 20476
rect 33796 20330 33824 20470
rect 34164 20466 34192 21966
rect 34152 20460 34204 20466
rect 34152 20402 34204 20408
rect 33784 20324 33836 20330
rect 33784 20266 33836 20272
rect 33416 20052 33468 20058
rect 33416 19994 33468 20000
rect 33600 19984 33652 19990
rect 33600 19926 33652 19932
rect 33232 19780 33284 19786
rect 33232 19722 33284 19728
rect 33046 19544 33102 19553
rect 32956 19508 33008 19514
rect 33612 19514 33640 19926
rect 33796 19786 33824 20266
rect 34060 20052 34112 20058
rect 34164 20040 34192 20402
rect 34112 20012 34192 20040
rect 34060 19994 34112 20000
rect 34256 19938 34284 22374
rect 34520 22160 34572 22166
rect 34520 22102 34572 22108
rect 34532 21350 34560 22102
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 35164 21412 35216 21418
rect 35164 21354 35216 21360
rect 34520 21344 34572 21350
rect 35176 21321 35204 21354
rect 34520 21286 34572 21292
rect 35162 21312 35218 21321
rect 34532 21146 34560 21286
rect 35162 21247 35218 21256
rect 34520 21140 34572 21146
rect 34520 21082 34572 21088
rect 35268 21010 35296 22596
rect 35348 21888 35400 21894
rect 35348 21830 35400 21836
rect 35360 21554 35388 21830
rect 35636 21554 35664 23446
rect 35808 23112 35860 23118
rect 35808 23054 35860 23060
rect 35820 22778 35848 23054
rect 35808 22772 35860 22778
rect 35808 22714 35860 22720
rect 35348 21548 35400 21554
rect 35348 21490 35400 21496
rect 35624 21548 35676 21554
rect 35624 21490 35676 21496
rect 35360 21146 35388 21490
rect 35348 21140 35400 21146
rect 35348 21082 35400 21088
rect 35256 21004 35308 21010
rect 35256 20946 35308 20952
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 35162 20360 35218 20369
rect 35268 20346 35296 20946
rect 35218 20318 35296 20346
rect 35162 20295 35218 20304
rect 35176 20262 35204 20295
rect 35164 20256 35216 20262
rect 35164 20198 35216 20204
rect 34072 19910 34284 19938
rect 33784 19780 33836 19786
rect 33784 19722 33836 19728
rect 33046 19479 33102 19488
rect 33600 19508 33652 19514
rect 32956 19450 33008 19456
rect 32956 19304 33008 19310
rect 32956 19246 33008 19252
rect 32968 17270 32996 19246
rect 33060 18290 33088 19479
rect 33600 19450 33652 19456
rect 33230 19408 33286 19417
rect 33230 19343 33286 19352
rect 33048 18284 33100 18290
rect 33048 18226 33100 18232
rect 33048 18148 33100 18154
rect 33048 18090 33100 18096
rect 32956 17264 33008 17270
rect 32956 17206 33008 17212
rect 32956 16992 33008 16998
rect 32956 16934 33008 16940
rect 32968 15502 32996 16934
rect 32956 15496 33008 15502
rect 32956 15438 33008 15444
rect 32956 14952 33008 14958
rect 32956 14894 33008 14900
rect 32968 14793 32996 14894
rect 32954 14784 33010 14793
rect 32954 14719 33010 14728
rect 32864 14272 32916 14278
rect 32864 14214 32916 14220
rect 32956 13932 33008 13938
rect 32956 13874 33008 13880
rect 32968 13814 32996 13874
rect 33060 13841 33088 18090
rect 33140 17332 33192 17338
rect 33140 17274 33192 17280
rect 33152 16250 33180 17274
rect 33244 17134 33272 19343
rect 33324 19168 33376 19174
rect 33324 19110 33376 19116
rect 33336 17202 33364 19110
rect 33600 18964 33652 18970
rect 33600 18906 33652 18912
rect 33612 18873 33640 18906
rect 33598 18864 33654 18873
rect 33598 18799 33654 18808
rect 33612 18426 33640 18799
rect 33508 18420 33560 18426
rect 33508 18362 33560 18368
rect 33600 18420 33652 18426
rect 33600 18362 33652 18368
rect 33520 18329 33548 18362
rect 34072 18358 34100 19910
rect 35636 19854 35664 21490
rect 35912 20398 35940 23446
rect 36004 22681 36032 27270
rect 36084 26852 36136 26858
rect 36084 26794 36136 26800
rect 36096 25838 36124 26794
rect 36188 26790 36216 27814
rect 36464 27130 36492 28494
rect 37752 28121 37780 29990
rect 37738 28112 37794 28121
rect 36636 28076 36688 28082
rect 37738 28047 37794 28056
rect 36636 28018 36688 28024
rect 36648 27674 36676 28018
rect 36636 27668 36688 27674
rect 36636 27610 36688 27616
rect 37844 27334 37872 31078
rect 38028 28150 38056 33102
rect 38106 33079 38162 33088
rect 38212 29850 38240 34342
rect 38396 33114 38424 34983
rect 38844 34954 38896 34960
rect 38856 34610 38884 34954
rect 38844 34604 38896 34610
rect 38844 34546 38896 34552
rect 38936 34604 38988 34610
rect 38936 34546 38988 34552
rect 38844 34468 38896 34474
rect 38948 34456 38976 34546
rect 38896 34428 38976 34456
rect 38844 34410 38896 34416
rect 38660 34400 38712 34406
rect 38660 34342 38712 34348
rect 38672 34202 38700 34342
rect 39132 34202 39160 35022
rect 39224 34746 39252 35158
rect 39212 34740 39264 34746
rect 39212 34682 39264 34688
rect 39408 34202 39436 36110
rect 39488 34468 39540 34474
rect 39488 34410 39540 34416
rect 38660 34196 38712 34202
rect 38660 34138 38712 34144
rect 39120 34196 39172 34202
rect 39120 34138 39172 34144
rect 39396 34196 39448 34202
rect 39396 34138 39448 34144
rect 38936 33652 38988 33658
rect 38936 33594 38988 33600
rect 38948 33386 38976 33594
rect 39408 33590 39436 34138
rect 39396 33584 39448 33590
rect 39396 33526 39448 33532
rect 39500 33522 39528 34410
rect 39212 33516 39264 33522
rect 39212 33458 39264 33464
rect 39488 33516 39540 33522
rect 39488 33458 39540 33464
rect 38936 33380 38988 33386
rect 38936 33322 38988 33328
rect 38384 33108 38436 33114
rect 38384 33050 38436 33056
rect 39028 33040 39080 33046
rect 39028 32982 39080 32988
rect 38752 32972 38804 32978
rect 38752 32914 38804 32920
rect 38764 32230 38792 32914
rect 38936 32904 38988 32910
rect 38936 32846 38988 32852
rect 38844 32768 38896 32774
rect 38844 32710 38896 32716
rect 38752 32224 38804 32230
rect 38752 32166 38804 32172
rect 38476 31952 38528 31958
rect 38476 31894 38528 31900
rect 38488 31346 38516 31894
rect 38568 31748 38620 31754
rect 38568 31690 38620 31696
rect 38580 31346 38608 31690
rect 38476 31340 38528 31346
rect 38476 31282 38528 31288
rect 38568 31340 38620 31346
rect 38568 31282 38620 31288
rect 38292 31272 38344 31278
rect 38292 31214 38344 31220
rect 38304 30938 38332 31214
rect 38292 30932 38344 30938
rect 38292 30874 38344 30880
rect 38384 30048 38436 30054
rect 38384 29990 38436 29996
rect 38200 29844 38252 29850
rect 38200 29786 38252 29792
rect 38108 29164 38160 29170
rect 38108 29106 38160 29112
rect 38120 28762 38148 29106
rect 38200 28960 38252 28966
rect 38200 28902 38252 28908
rect 38108 28756 38160 28762
rect 38108 28698 38160 28704
rect 38212 28694 38240 28902
rect 38200 28688 38252 28694
rect 38200 28630 38252 28636
rect 38016 28144 38068 28150
rect 38016 28086 38068 28092
rect 38292 28008 38344 28014
rect 38292 27950 38344 27956
rect 38016 27872 38068 27878
rect 38016 27814 38068 27820
rect 38028 27606 38056 27814
rect 38304 27606 38332 27950
rect 38016 27600 38068 27606
rect 38016 27542 38068 27548
rect 38292 27600 38344 27606
rect 38292 27542 38344 27548
rect 37832 27328 37884 27334
rect 37832 27270 37884 27276
rect 38028 27130 38056 27542
rect 36452 27124 36504 27130
rect 36452 27066 36504 27072
rect 38016 27124 38068 27130
rect 38016 27066 38068 27072
rect 38304 27062 38332 27542
rect 38292 27056 38344 27062
rect 38292 26998 38344 27004
rect 36176 26784 36228 26790
rect 36176 26726 36228 26732
rect 36188 26586 36216 26726
rect 36176 26580 36228 26586
rect 36176 26522 36228 26528
rect 36084 25832 36136 25838
rect 36084 25774 36136 25780
rect 36096 25498 36124 25774
rect 36188 25770 36216 26522
rect 38304 26518 38332 26998
rect 38292 26512 38344 26518
rect 38292 26454 38344 26460
rect 37740 26240 37792 26246
rect 37740 26182 37792 26188
rect 37752 26042 37780 26182
rect 37740 26036 37792 26042
rect 37740 25978 37792 25984
rect 37752 25770 37780 25978
rect 38396 25906 38424 29990
rect 38488 29782 38516 31282
rect 38580 30190 38608 31282
rect 38568 30184 38620 30190
rect 38568 30126 38620 30132
rect 38476 29776 38528 29782
rect 38476 29718 38528 29724
rect 38488 28948 38516 29718
rect 38568 28960 38620 28966
rect 38488 28920 38568 28948
rect 38488 28694 38516 28920
rect 38568 28902 38620 28908
rect 38476 28688 38528 28694
rect 38476 28630 38528 28636
rect 38488 27946 38516 28630
rect 38476 27940 38528 27946
rect 38476 27882 38528 27888
rect 38568 27464 38620 27470
rect 38568 27406 38620 27412
rect 38580 26994 38608 27406
rect 38660 27328 38712 27334
rect 38660 27270 38712 27276
rect 38568 26988 38620 26994
rect 38568 26930 38620 26936
rect 38476 26376 38528 26382
rect 38476 26318 38528 26324
rect 38488 25906 38516 26318
rect 38580 26314 38608 26930
rect 38672 26858 38700 27270
rect 38660 26852 38712 26858
rect 38660 26794 38712 26800
rect 38568 26308 38620 26314
rect 38568 26250 38620 26256
rect 38580 25974 38608 26250
rect 38568 25968 38620 25974
rect 38568 25910 38620 25916
rect 37832 25900 37884 25906
rect 37832 25842 37884 25848
rect 38384 25900 38436 25906
rect 38384 25842 38436 25848
rect 38476 25900 38528 25906
rect 38476 25842 38528 25848
rect 36176 25764 36228 25770
rect 36176 25706 36228 25712
rect 37740 25764 37792 25770
rect 37740 25706 37792 25712
rect 36084 25492 36136 25498
rect 36084 25434 36136 25440
rect 36188 25430 36216 25706
rect 37004 25696 37056 25702
rect 37004 25638 37056 25644
rect 37372 25696 37424 25702
rect 37372 25638 37424 25644
rect 37016 25430 37044 25638
rect 36176 25424 36228 25430
rect 36176 25366 36228 25372
rect 37004 25424 37056 25430
rect 37004 25366 37056 25372
rect 36360 25220 36412 25226
rect 36360 25162 36412 25168
rect 36176 25152 36228 25158
rect 36176 25094 36228 25100
rect 36188 23118 36216 25094
rect 36372 24886 36400 25162
rect 36360 24880 36412 24886
rect 36360 24822 36412 24828
rect 36820 24812 36872 24818
rect 36820 24754 36872 24760
rect 36360 24268 36412 24274
rect 36360 24210 36412 24216
rect 36372 23866 36400 24210
rect 36636 24064 36688 24070
rect 36636 24006 36688 24012
rect 36360 23860 36412 23866
rect 36360 23802 36412 23808
rect 36648 23730 36676 24006
rect 36636 23724 36688 23730
rect 36636 23666 36688 23672
rect 36268 23520 36320 23526
rect 36268 23462 36320 23468
rect 36280 23254 36308 23462
rect 36648 23322 36676 23666
rect 36636 23316 36688 23322
rect 36636 23258 36688 23264
rect 36268 23248 36320 23254
rect 36268 23190 36320 23196
rect 36176 23112 36228 23118
rect 36176 23054 36228 23060
rect 36832 23050 36860 24754
rect 36912 24676 36964 24682
rect 36912 24618 36964 24624
rect 36924 24342 36952 24618
rect 37384 24342 37412 25638
rect 37648 24676 37700 24682
rect 37648 24618 37700 24624
rect 37556 24608 37608 24614
rect 37556 24550 37608 24556
rect 36912 24336 36964 24342
rect 36912 24278 36964 24284
rect 37372 24336 37424 24342
rect 37372 24278 37424 24284
rect 36924 24070 36952 24278
rect 36912 24064 36964 24070
rect 36912 24006 36964 24012
rect 37464 23792 37516 23798
rect 37464 23734 37516 23740
rect 37476 23594 37504 23734
rect 37464 23588 37516 23594
rect 37464 23530 37516 23536
rect 36820 23044 36872 23050
rect 36820 22986 36872 22992
rect 35990 22672 36046 22681
rect 35990 22607 36046 22616
rect 36728 22568 36780 22574
rect 36728 22510 36780 22516
rect 36176 22432 36228 22438
rect 36176 22374 36228 22380
rect 36188 22166 36216 22374
rect 36176 22160 36228 22166
rect 36176 22102 36228 22108
rect 36268 22160 36320 22166
rect 36268 22102 36320 22108
rect 36280 21350 36308 22102
rect 36740 21593 36768 22510
rect 36832 22030 36860 22986
rect 37188 22976 37240 22982
rect 37188 22918 37240 22924
rect 37200 22574 37228 22918
rect 37188 22568 37240 22574
rect 37188 22510 37240 22516
rect 36820 22024 36872 22030
rect 36820 21966 36872 21972
rect 36726 21584 36782 21593
rect 36360 21548 36412 21554
rect 36726 21519 36782 21528
rect 36360 21490 36412 21496
rect 36268 21344 36320 21350
rect 36268 21286 36320 21292
rect 36176 21072 36228 21078
rect 36176 21014 36228 21020
rect 36084 20936 36136 20942
rect 36084 20878 36136 20884
rect 36096 20602 36124 20878
rect 36188 20602 36216 21014
rect 36372 20942 36400 21490
rect 36360 20936 36412 20942
rect 36360 20878 36412 20884
rect 36832 20856 36860 21966
rect 36912 21888 36964 21894
rect 36912 21830 36964 21836
rect 36924 21554 36952 21830
rect 37476 21622 37504 23530
rect 37568 22778 37596 24550
rect 37660 24274 37688 24618
rect 37844 24449 37872 25842
rect 38396 25498 38424 25842
rect 38384 25492 38436 25498
rect 38384 25434 38436 25440
rect 38764 24886 38792 32166
rect 38856 30598 38884 32710
rect 38948 32337 38976 32846
rect 39040 32570 39068 32982
rect 39224 32842 39252 33458
rect 39592 33318 39620 36518
rect 40776 36304 40828 36310
rect 40776 36246 40828 36252
rect 40316 36168 40368 36174
rect 40316 36110 40368 36116
rect 40328 35834 40356 36110
rect 40788 35834 40816 36246
rect 40316 35828 40368 35834
rect 40316 35770 40368 35776
rect 40776 35828 40828 35834
rect 40776 35770 40828 35776
rect 40592 35148 40644 35154
rect 41064 35136 41092 39936
rect 41144 39918 41196 39924
rect 41144 38752 41196 38758
rect 41144 38694 41196 38700
rect 41156 36106 41184 38694
rect 41340 37448 41368 40054
rect 41616 39642 41644 40394
rect 41696 40384 41748 40390
rect 41696 40326 41748 40332
rect 41708 39914 41736 40326
rect 41800 39914 41828 40598
rect 41696 39908 41748 39914
rect 41696 39850 41748 39856
rect 41788 39908 41840 39914
rect 41788 39850 41840 39856
rect 41604 39636 41656 39642
rect 41604 39578 41656 39584
rect 41512 39568 41564 39574
rect 41512 39510 41564 39516
rect 41420 38820 41472 38826
rect 41420 38762 41472 38768
rect 41432 38282 41460 38762
rect 41524 38554 41552 39510
rect 41708 39098 41736 39850
rect 41696 39092 41748 39098
rect 41696 39034 41748 39040
rect 41800 38808 41828 39850
rect 41880 38820 41932 38826
rect 41800 38780 41880 38808
rect 41880 38762 41932 38768
rect 41604 38752 41656 38758
rect 41604 38694 41656 38700
rect 41512 38548 41564 38554
rect 41512 38490 41564 38496
rect 41420 38276 41472 38282
rect 41420 38218 41472 38224
rect 41432 38010 41460 38218
rect 41420 38004 41472 38010
rect 41420 37946 41472 37952
rect 41616 37466 41644 38694
rect 41892 38554 41920 38762
rect 41880 38548 41932 38554
rect 41880 38490 41932 38496
rect 41892 38418 41920 38490
rect 41880 38412 41932 38418
rect 41880 38354 41932 38360
rect 41696 38344 41748 38350
rect 41696 38286 41748 38292
rect 41708 38010 41736 38286
rect 41696 38004 41748 38010
rect 41696 37946 41748 37952
rect 41788 37936 41840 37942
rect 41788 37878 41840 37884
rect 41604 37460 41656 37466
rect 41340 37420 41460 37448
rect 41328 36168 41380 36174
rect 41328 36110 41380 36116
rect 41144 36100 41196 36106
rect 41144 36042 41196 36048
rect 41236 35692 41288 35698
rect 41236 35634 41288 35640
rect 41248 35290 41276 35634
rect 41236 35284 41288 35290
rect 41236 35226 41288 35232
rect 41064 35108 41276 35136
rect 40592 35090 40644 35096
rect 39854 34776 39910 34785
rect 39854 34711 39910 34720
rect 39580 33312 39632 33318
rect 39580 33254 39632 33260
rect 39868 33114 39896 34711
rect 40604 34678 40632 35090
rect 40868 35080 40920 35086
rect 40868 35022 40920 35028
rect 40592 34672 40644 34678
rect 40592 34614 40644 34620
rect 40776 34400 40828 34406
rect 40776 34342 40828 34348
rect 40592 34128 40644 34134
rect 40592 34070 40644 34076
rect 40604 33658 40632 34070
rect 40592 33652 40644 33658
rect 40592 33594 40644 33600
rect 40604 33368 40632 33594
rect 40788 33522 40816 34342
rect 40880 33998 40908 35022
rect 41144 35012 41196 35018
rect 41144 34954 41196 34960
rect 41156 34134 41184 34954
rect 41144 34128 41196 34134
rect 41144 34070 41196 34076
rect 41248 34066 41276 35108
rect 41236 34060 41288 34066
rect 41236 34002 41288 34008
rect 40868 33992 40920 33998
rect 40868 33934 40920 33940
rect 40776 33516 40828 33522
rect 40776 33458 40828 33464
rect 40684 33380 40736 33386
rect 40420 33340 40684 33368
rect 39856 33108 39908 33114
rect 39856 33050 39908 33056
rect 39212 32836 39264 32842
rect 39212 32778 39264 32784
rect 39028 32564 39080 32570
rect 39028 32506 39080 32512
rect 38934 32328 38990 32337
rect 38934 32263 38990 32272
rect 38948 31958 38976 32263
rect 38936 31952 38988 31958
rect 38936 31894 38988 31900
rect 39120 31272 39172 31278
rect 39120 31214 39172 31220
rect 38936 30796 38988 30802
rect 38936 30738 38988 30744
rect 38844 30592 38896 30598
rect 38844 30534 38896 30540
rect 38948 30054 38976 30738
rect 38936 30048 38988 30054
rect 38936 29990 38988 29996
rect 38948 28801 38976 29990
rect 38934 28792 38990 28801
rect 38934 28727 38990 28736
rect 38844 28620 38896 28626
rect 38844 28562 38896 28568
rect 38856 28218 38884 28562
rect 39132 28529 39160 31214
rect 39224 30938 39252 32778
rect 39868 32570 39896 33050
rect 40420 32570 40448 33340
rect 40684 33322 40736 33328
rect 41340 33134 41368 36110
rect 41432 34746 41460 37420
rect 41604 37402 41656 37408
rect 41512 37392 41564 37398
rect 41512 37334 41564 37340
rect 41524 36922 41552 37334
rect 41616 36922 41644 37402
rect 41512 36916 41564 36922
rect 41512 36858 41564 36864
rect 41604 36916 41656 36922
rect 41604 36858 41656 36864
rect 41800 36854 41828 37878
rect 41892 37738 41920 38354
rect 41880 37732 41932 37738
rect 41880 37674 41932 37680
rect 41892 37466 41920 37674
rect 41880 37460 41932 37466
rect 41880 37402 41932 37408
rect 41788 36848 41840 36854
rect 41972 36848 42024 36854
rect 41840 36808 41972 36836
rect 41788 36790 41840 36796
rect 42076 36825 42104 40870
rect 42168 40730 42196 41414
rect 42260 41002 42288 41686
rect 46952 41682 46980 49558
rect 47122 49520 47178 49558
rect 46940 41676 46992 41682
rect 46940 41618 46992 41624
rect 42432 41132 42484 41138
rect 42432 41074 42484 41080
rect 42248 40996 42300 41002
rect 42248 40938 42300 40944
rect 42156 40724 42208 40730
rect 42156 40666 42208 40672
rect 42444 40662 42472 41074
rect 43260 40724 43312 40730
rect 43260 40666 43312 40672
rect 42432 40656 42484 40662
rect 42432 40598 42484 40604
rect 42444 40186 42472 40598
rect 42432 40180 42484 40186
rect 42432 40122 42484 40128
rect 42444 39506 42472 40122
rect 43272 40050 43300 40666
rect 43260 40044 43312 40050
rect 43260 39986 43312 39992
rect 43076 39908 43128 39914
rect 43076 39850 43128 39856
rect 43088 39574 43116 39850
rect 43076 39568 43128 39574
rect 43076 39510 43128 39516
rect 42432 39500 42484 39506
rect 42432 39442 42484 39448
rect 42708 39092 42760 39098
rect 42708 39034 42760 39040
rect 42432 37664 42484 37670
rect 42432 37606 42484 37612
rect 42444 37466 42472 37606
rect 42432 37460 42484 37466
rect 42432 37402 42484 37408
rect 41972 36790 42024 36796
rect 42062 36816 42118 36825
rect 42062 36751 42118 36760
rect 42340 36780 42392 36786
rect 41696 36236 41748 36242
rect 41696 36178 41748 36184
rect 41708 36106 41736 36178
rect 41696 36100 41748 36106
rect 41696 36042 41748 36048
rect 41788 36100 41840 36106
rect 41788 36042 41840 36048
rect 41708 35834 41736 36042
rect 41696 35828 41748 35834
rect 41696 35770 41748 35776
rect 41800 35086 41828 36042
rect 41880 35488 41932 35494
rect 41880 35430 41932 35436
rect 41892 35222 41920 35430
rect 41880 35216 41932 35222
rect 41880 35158 41932 35164
rect 41788 35080 41840 35086
rect 41788 35022 41840 35028
rect 41420 34740 41472 34746
rect 41420 34682 41472 34688
rect 41432 34542 41460 34682
rect 41420 34536 41472 34542
rect 41420 34478 41472 34484
rect 41800 34202 41828 35022
rect 41892 34746 41920 35158
rect 41880 34740 41932 34746
rect 41880 34682 41932 34688
rect 41788 34196 41840 34202
rect 41788 34138 41840 34144
rect 41512 33992 41564 33998
rect 41512 33934 41564 33940
rect 41524 33658 41552 33934
rect 41512 33652 41564 33658
rect 41512 33594 41564 33600
rect 41248 33106 41368 33134
rect 41970 33144 42026 33153
rect 40592 33040 40644 33046
rect 40592 32982 40644 32988
rect 39856 32564 39908 32570
rect 39856 32506 39908 32512
rect 40408 32564 40460 32570
rect 40408 32506 40460 32512
rect 39868 32366 39896 32506
rect 39856 32360 39908 32366
rect 39856 32302 39908 32308
rect 40420 32298 40448 32506
rect 40408 32292 40460 32298
rect 40408 32234 40460 32240
rect 39672 31952 39724 31958
rect 39672 31894 39724 31900
rect 39488 31816 39540 31822
rect 39488 31758 39540 31764
rect 39396 31680 39448 31686
rect 39396 31622 39448 31628
rect 39408 31482 39436 31622
rect 39396 31476 39448 31482
rect 39396 31418 39448 31424
rect 39500 31210 39528 31758
rect 39684 31414 39712 31894
rect 40420 31890 40448 32234
rect 40604 32026 40632 32982
rect 41248 32910 41276 33106
rect 42076 33134 42104 36751
rect 42444 36768 42472 37402
rect 42614 37224 42670 37233
rect 42614 37159 42670 37168
rect 42392 36740 42472 36768
rect 42340 36722 42392 36728
rect 42524 34944 42576 34950
rect 42524 34886 42576 34892
rect 42536 34610 42564 34886
rect 42628 34746 42656 37159
rect 42720 36242 42748 39034
rect 43088 39030 43116 39510
rect 43168 39500 43220 39506
rect 43168 39442 43220 39448
rect 43180 39098 43208 39442
rect 43168 39092 43220 39098
rect 43168 39034 43220 39040
rect 43076 39024 43128 39030
rect 43076 38966 43128 38972
rect 43444 39024 43496 39030
rect 43444 38966 43496 38972
rect 43456 38826 43484 38966
rect 43444 38820 43496 38826
rect 43444 38762 43496 38768
rect 43536 38752 43588 38758
rect 43536 38694 43588 38700
rect 43548 38554 43576 38694
rect 43536 38548 43588 38554
rect 43536 38490 43588 38496
rect 43812 38412 43864 38418
rect 43812 38354 43864 38360
rect 43628 37800 43680 37806
rect 43628 37742 43680 37748
rect 43352 37324 43404 37330
rect 43352 37266 43404 37272
rect 43364 36582 43392 37266
rect 43352 36576 43404 36582
rect 43352 36518 43404 36524
rect 42708 36236 42760 36242
rect 42708 36178 42760 36184
rect 42720 36145 42748 36178
rect 43260 36168 43312 36174
rect 42706 36136 42762 36145
rect 43260 36110 43312 36116
rect 42706 36071 42762 36080
rect 43076 36032 43128 36038
rect 43076 35974 43128 35980
rect 43088 35698 43116 35974
rect 43272 35698 43300 36110
rect 43076 35692 43128 35698
rect 43076 35634 43128 35640
rect 43260 35692 43312 35698
rect 43260 35634 43312 35640
rect 43260 35148 43312 35154
rect 43260 35090 43312 35096
rect 42892 35080 42944 35086
rect 42892 35022 42944 35028
rect 42616 34740 42668 34746
rect 42616 34682 42668 34688
rect 42524 34604 42576 34610
rect 42524 34546 42576 34552
rect 42800 34604 42852 34610
rect 42800 34546 42852 34552
rect 42812 34134 42840 34546
rect 42800 34128 42852 34134
rect 42800 34070 42852 34076
rect 42248 34060 42300 34066
rect 42248 34002 42300 34008
rect 42260 33658 42288 34002
rect 42708 33856 42760 33862
rect 42708 33798 42760 33804
rect 42248 33652 42300 33658
rect 42248 33594 42300 33600
rect 42720 33522 42748 33798
rect 42812 33522 42840 34070
rect 42904 33930 42932 35022
rect 43272 34746 43300 35090
rect 43364 34785 43392 36518
rect 43350 34776 43406 34785
rect 43260 34740 43312 34746
rect 43350 34711 43406 34720
rect 43260 34682 43312 34688
rect 43536 34128 43588 34134
rect 43536 34070 43588 34076
rect 43076 33992 43128 33998
rect 43076 33934 43128 33940
rect 42892 33924 42944 33930
rect 42892 33866 42944 33872
rect 42904 33590 42932 33866
rect 42892 33584 42944 33590
rect 42892 33526 42944 33532
rect 42708 33516 42760 33522
rect 42708 33458 42760 33464
rect 42800 33516 42852 33522
rect 42800 33458 42852 33464
rect 42076 33106 42196 33134
rect 42720 33114 42748 33458
rect 42800 33380 42852 33386
rect 42800 33322 42852 33328
rect 41970 33079 42026 33088
rect 41236 32904 41288 32910
rect 41236 32846 41288 32852
rect 40776 32428 40828 32434
rect 40776 32370 40828 32376
rect 40592 32020 40644 32026
rect 40592 31962 40644 31968
rect 40408 31884 40460 31890
rect 40408 31826 40460 31832
rect 40788 31482 40816 32370
rect 41248 32298 41276 32846
rect 41236 32292 41288 32298
rect 41236 32234 41288 32240
rect 41248 31754 41276 32234
rect 41512 31952 41564 31958
rect 41512 31894 41564 31900
rect 41236 31748 41288 31754
rect 41236 31690 41288 31696
rect 40776 31476 40828 31482
rect 40776 31418 40828 31424
rect 41524 31414 41552 31894
rect 41880 31816 41932 31822
rect 41880 31758 41932 31764
rect 41892 31482 41920 31758
rect 41880 31476 41932 31482
rect 41880 31418 41932 31424
rect 39672 31408 39724 31414
rect 39672 31350 39724 31356
rect 41512 31408 41564 31414
rect 41512 31350 41564 31356
rect 39488 31204 39540 31210
rect 39488 31146 39540 31152
rect 39212 30932 39264 30938
rect 39212 30874 39264 30880
rect 39212 30592 39264 30598
rect 39212 30534 39264 30540
rect 39224 30190 39252 30534
rect 39684 30394 39712 31350
rect 41052 31136 41104 31142
rect 41052 31078 41104 31084
rect 39764 30796 39816 30802
rect 39764 30738 39816 30744
rect 39672 30388 39724 30394
rect 39672 30330 39724 30336
rect 39212 30184 39264 30190
rect 39212 30126 39264 30132
rect 39118 28520 39174 28529
rect 39118 28455 39174 28464
rect 38844 28212 38896 28218
rect 38844 28154 38896 28160
rect 39026 27704 39082 27713
rect 39224 27674 39252 30126
rect 39776 30054 39804 30738
rect 40960 30592 41012 30598
rect 40960 30534 41012 30540
rect 40972 30258 41000 30534
rect 40960 30252 41012 30258
rect 40960 30194 41012 30200
rect 39764 30048 39816 30054
rect 39764 29990 39816 29996
rect 39672 29640 39724 29646
rect 39776 29617 39804 29990
rect 40592 29776 40644 29782
rect 40592 29718 40644 29724
rect 39672 29582 39724 29588
rect 39762 29608 39818 29617
rect 39580 29504 39632 29510
rect 39580 29446 39632 29452
rect 39592 29306 39620 29446
rect 39580 29300 39632 29306
rect 39580 29242 39632 29248
rect 39684 29238 39712 29582
rect 39762 29543 39818 29552
rect 40316 29504 40368 29510
rect 40316 29446 40368 29452
rect 39672 29232 39724 29238
rect 39672 29174 39724 29180
rect 40040 29164 40092 29170
rect 40040 29106 40092 29112
rect 40052 28694 40080 29106
rect 40132 28756 40184 28762
rect 40132 28698 40184 28704
rect 40040 28688 40092 28694
rect 40040 28630 40092 28636
rect 39948 28484 40000 28490
rect 39948 28426 40000 28432
rect 39764 27940 39816 27946
rect 39764 27882 39816 27888
rect 39580 27872 39632 27878
rect 39580 27814 39632 27820
rect 39672 27872 39724 27878
rect 39672 27814 39724 27820
rect 39026 27639 39082 27648
rect 39212 27668 39264 27674
rect 38844 25356 38896 25362
rect 38844 25298 38896 25304
rect 38752 24880 38804 24886
rect 38752 24822 38804 24828
rect 38016 24744 38068 24750
rect 38016 24686 38068 24692
rect 37830 24440 37886 24449
rect 37830 24375 37886 24384
rect 37648 24268 37700 24274
rect 37648 24210 37700 24216
rect 37648 24132 37700 24138
rect 37648 24074 37700 24080
rect 37660 23866 37688 24074
rect 37648 23860 37700 23866
rect 37648 23802 37700 23808
rect 37556 22772 37608 22778
rect 37556 22714 37608 22720
rect 37844 22098 37872 24375
rect 38028 22642 38056 24686
rect 38856 24614 38884 25298
rect 38844 24608 38896 24614
rect 38844 24550 38896 24556
rect 38108 24132 38160 24138
rect 38108 24074 38160 24080
rect 38120 23730 38148 24074
rect 38200 24064 38252 24070
rect 38200 24006 38252 24012
rect 38108 23724 38160 23730
rect 38108 23666 38160 23672
rect 38212 23594 38240 24006
rect 38568 23724 38620 23730
rect 38568 23666 38620 23672
rect 38200 23588 38252 23594
rect 38200 23530 38252 23536
rect 38580 23254 38608 23666
rect 38568 23248 38620 23254
rect 38568 23190 38620 23196
rect 38856 23186 38884 24550
rect 38292 23180 38344 23186
rect 38292 23122 38344 23128
rect 38844 23180 38896 23186
rect 38844 23122 38896 23128
rect 38108 23112 38160 23118
rect 38108 23054 38160 23060
rect 38120 22778 38148 23054
rect 38108 22772 38160 22778
rect 38108 22714 38160 22720
rect 38304 22710 38332 23122
rect 39040 22710 39068 27639
rect 39212 27610 39264 27616
rect 39224 27577 39252 27610
rect 39210 27568 39266 27577
rect 39210 27503 39266 27512
rect 39592 26518 39620 27814
rect 39580 26512 39632 26518
rect 39580 26454 39632 26460
rect 39592 26042 39620 26454
rect 39580 26036 39632 26042
rect 39580 25978 39632 25984
rect 39304 25288 39356 25294
rect 39304 25230 39356 25236
rect 39212 25152 39264 25158
rect 39212 25094 39264 25100
rect 39120 24200 39172 24206
rect 39120 24142 39172 24148
rect 39132 23730 39160 24142
rect 39120 23724 39172 23730
rect 39120 23666 39172 23672
rect 38292 22704 38344 22710
rect 38292 22646 38344 22652
rect 39028 22704 39080 22710
rect 39028 22646 39080 22652
rect 38016 22636 38068 22642
rect 38016 22578 38068 22584
rect 38384 22568 38436 22574
rect 38384 22510 38436 22516
rect 38396 22234 38424 22510
rect 38384 22228 38436 22234
rect 38384 22170 38436 22176
rect 37832 22092 37884 22098
rect 37832 22034 37884 22040
rect 38292 22092 38344 22098
rect 38292 22034 38344 22040
rect 38200 22024 38252 22030
rect 38200 21966 38252 21972
rect 37464 21616 37516 21622
rect 37464 21558 37516 21564
rect 36912 21548 36964 21554
rect 36912 21490 36964 21496
rect 36924 21146 36952 21490
rect 36912 21140 36964 21146
rect 36912 21082 36964 21088
rect 36832 20828 36952 20856
rect 36084 20596 36136 20602
rect 36084 20538 36136 20544
rect 36176 20596 36228 20602
rect 36176 20538 36228 20544
rect 35900 20392 35952 20398
rect 35900 20334 35952 20340
rect 36084 20392 36136 20398
rect 36084 20334 36136 20340
rect 35898 20224 35954 20233
rect 35898 20159 35954 20168
rect 34796 19848 34848 19854
rect 34796 19790 34848 19796
rect 35624 19848 35676 19854
rect 35624 19790 35676 19796
rect 34428 19712 34480 19718
rect 34428 19654 34480 19660
rect 34440 19310 34468 19654
rect 34428 19304 34480 19310
rect 34428 19246 34480 19252
rect 34440 18902 34468 19246
rect 34808 18970 34836 19790
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35348 19236 35400 19242
rect 35348 19178 35400 19184
rect 34796 18964 34848 18970
rect 34796 18906 34848 18912
rect 35360 18902 35388 19178
rect 34428 18896 34480 18902
rect 34428 18838 34480 18844
rect 35348 18896 35400 18902
rect 35348 18838 35400 18844
rect 34704 18828 34756 18834
rect 34704 18770 34756 18776
rect 34060 18352 34112 18358
rect 33506 18320 33562 18329
rect 34060 18294 34112 18300
rect 33506 18255 33562 18264
rect 33416 17740 33468 17746
rect 33416 17682 33468 17688
rect 33784 17740 33836 17746
rect 33784 17682 33836 17688
rect 33324 17196 33376 17202
rect 33324 17138 33376 17144
rect 33232 17128 33284 17134
rect 33232 17070 33284 17076
rect 33428 16794 33456 17682
rect 33796 17338 33824 17682
rect 33784 17332 33836 17338
rect 33784 17274 33836 17280
rect 33416 16788 33468 16794
rect 33416 16730 33468 16736
rect 33968 16584 34020 16590
rect 33968 16526 34020 16532
rect 33140 16244 33192 16250
rect 33140 16186 33192 16192
rect 33152 15162 33180 16186
rect 33980 16114 34008 16526
rect 33968 16108 34020 16114
rect 33968 16050 34020 16056
rect 34072 16046 34100 18294
rect 34152 18284 34204 18290
rect 34152 18226 34204 18232
rect 33508 16040 33560 16046
rect 33508 15982 33560 15988
rect 34060 16040 34112 16046
rect 34060 15982 34112 15988
rect 33520 15502 33548 15982
rect 34164 15570 34192 18226
rect 34716 18086 34744 18770
rect 35256 18624 35308 18630
rect 35256 18566 35308 18572
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34704 18080 34756 18086
rect 34704 18022 34756 18028
rect 34716 17814 34744 18022
rect 35268 17882 35296 18566
rect 35360 18426 35388 18838
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 35360 18154 35388 18362
rect 35348 18148 35400 18154
rect 35348 18090 35400 18096
rect 35808 18148 35860 18154
rect 35808 18090 35860 18096
rect 35820 17882 35848 18090
rect 35256 17876 35308 17882
rect 35256 17818 35308 17824
rect 35808 17876 35860 17882
rect 35808 17818 35860 17824
rect 34704 17808 34756 17814
rect 34704 17750 34756 17756
rect 34336 17536 34388 17542
rect 34336 17478 34388 17484
rect 34348 17066 34376 17478
rect 34716 17338 34744 17750
rect 35256 17672 35308 17678
rect 35256 17614 35308 17620
rect 35348 17672 35400 17678
rect 35348 17614 35400 17620
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 34704 17332 34756 17338
rect 34704 17274 34756 17280
rect 34796 17332 34848 17338
rect 34796 17274 34848 17280
rect 34336 17060 34388 17066
rect 34336 17002 34388 17008
rect 34612 16992 34664 16998
rect 34612 16934 34664 16940
rect 34336 16788 34388 16794
rect 34336 16730 34388 16736
rect 34348 15978 34376 16730
rect 34336 15972 34388 15978
rect 34336 15914 34388 15920
rect 34520 15904 34572 15910
rect 34520 15846 34572 15852
rect 34152 15564 34204 15570
rect 34152 15506 34204 15512
rect 33508 15496 33560 15502
rect 33508 15438 33560 15444
rect 33140 15156 33192 15162
rect 33140 15098 33192 15104
rect 33876 15156 33928 15162
rect 33876 15098 33928 15104
rect 33324 14068 33376 14074
rect 33324 14010 33376 14016
rect 32876 13786 32996 13814
rect 33046 13832 33102 13841
rect 32772 13728 32824 13734
rect 32600 13654 32720 13682
rect 32772 13670 32824 13676
rect 32508 13518 32628 13546
rect 32496 13456 32548 13462
rect 32496 13398 32548 13404
rect 32404 13184 32456 13190
rect 32404 13126 32456 13132
rect 32508 12986 32536 13398
rect 32496 12980 32548 12986
rect 32496 12922 32548 12928
rect 32600 12850 32628 13518
rect 32692 12918 32720 13654
rect 32876 13462 32904 13786
rect 33336 13802 33364 14010
rect 33888 13841 33916 15098
rect 34164 14822 34192 15506
rect 33968 14816 34020 14822
rect 33968 14758 34020 14764
rect 34152 14816 34204 14822
rect 34152 14758 34204 14764
rect 33874 13832 33930 13841
rect 33046 13767 33102 13776
rect 33324 13796 33376 13802
rect 33874 13767 33930 13776
rect 33324 13738 33376 13744
rect 32956 13728 33008 13734
rect 32956 13670 33008 13676
rect 32864 13456 32916 13462
rect 32784 13416 32864 13444
rect 32680 12912 32732 12918
rect 32680 12854 32732 12860
rect 32588 12844 32640 12850
rect 32588 12786 32640 12792
rect 32600 12238 32628 12786
rect 32588 12232 32640 12238
rect 32588 12174 32640 12180
rect 32784 11354 32812 13416
rect 32864 13398 32916 13404
rect 32864 13320 32916 13326
rect 32864 13262 32916 13268
rect 32876 12986 32904 13262
rect 32864 12980 32916 12986
rect 32864 12922 32916 12928
rect 32772 11348 32824 11354
rect 32772 11290 32824 11296
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32036 10804 32088 10810
rect 32036 10746 32088 10752
rect 31944 10668 31996 10674
rect 31944 10610 31996 10616
rect 31956 10198 31984 10610
rect 32048 10470 32076 10746
rect 32784 10674 32812 11290
rect 32772 10668 32824 10674
rect 32772 10610 32824 10616
rect 32128 10532 32180 10538
rect 32128 10474 32180 10480
rect 32036 10464 32088 10470
rect 32036 10406 32088 10412
rect 31944 10192 31996 10198
rect 31944 10134 31996 10140
rect 31760 10124 31812 10130
rect 31760 10066 31812 10072
rect 32048 9722 32076 10406
rect 32140 10266 32168 10474
rect 32588 10464 32640 10470
rect 32588 10406 32640 10412
rect 32600 10266 32628 10406
rect 32128 10260 32180 10266
rect 32128 10202 32180 10208
rect 32588 10260 32640 10266
rect 32588 10202 32640 10208
rect 32968 9994 32996 13670
rect 33888 13394 33916 13767
rect 33980 13394 34008 14758
rect 34164 13938 34192 14758
rect 34428 14544 34480 14550
rect 34428 14486 34480 14492
rect 34440 14074 34468 14486
rect 34428 14068 34480 14074
rect 34428 14010 34480 14016
rect 34532 14006 34560 15846
rect 34624 15570 34652 16934
rect 34808 16572 34836 17274
rect 35268 16658 35296 17614
rect 35360 17338 35388 17614
rect 35348 17332 35400 17338
rect 35348 17274 35400 17280
rect 35256 16652 35308 16658
rect 35256 16594 35308 16600
rect 34716 16544 34836 16572
rect 34612 15564 34664 15570
rect 34612 15506 34664 15512
rect 34624 15094 34652 15506
rect 34716 15337 34744 16544
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35268 16250 35296 16594
rect 35256 16244 35308 16250
rect 35256 16186 35308 16192
rect 35072 15564 35124 15570
rect 35072 15506 35124 15512
rect 35084 15473 35112 15506
rect 35070 15464 35126 15473
rect 35070 15399 35126 15408
rect 34796 15360 34848 15366
rect 34702 15328 34758 15337
rect 34796 15302 34848 15308
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 34702 15263 34758 15272
rect 34612 15088 34664 15094
rect 34610 15056 34612 15065
rect 34664 15056 34666 15065
rect 34610 14991 34666 15000
rect 34520 14000 34572 14006
rect 34520 13942 34572 13948
rect 34152 13932 34204 13938
rect 34152 13874 34204 13880
rect 33876 13388 33928 13394
rect 33876 13330 33928 13336
rect 33968 13388 34020 13394
rect 33968 13330 34020 13336
rect 33888 12986 33916 13330
rect 33876 12980 33928 12986
rect 33876 12922 33928 12928
rect 33784 12776 33836 12782
rect 33784 12718 33836 12724
rect 33796 12345 33824 12718
rect 33782 12336 33838 12345
rect 33782 12271 33838 12280
rect 33784 12096 33836 12102
rect 33784 12038 33836 12044
rect 33232 11688 33284 11694
rect 33232 11630 33284 11636
rect 33244 11121 33272 11630
rect 33508 11552 33560 11558
rect 33508 11494 33560 11500
rect 33520 11218 33548 11494
rect 33600 11280 33652 11286
rect 33600 11222 33652 11228
rect 33508 11212 33560 11218
rect 33508 11154 33560 11160
rect 33230 11112 33286 11121
rect 33230 11047 33286 11056
rect 33244 11014 33272 11047
rect 33232 11008 33284 11014
rect 33232 10950 33284 10956
rect 33140 10464 33192 10470
rect 33140 10406 33192 10412
rect 33152 10198 33180 10406
rect 33140 10192 33192 10198
rect 33140 10134 33192 10140
rect 32956 9988 33008 9994
rect 32956 9930 33008 9936
rect 29920 9716 29972 9722
rect 29920 9658 29972 9664
rect 32036 9716 32088 9722
rect 32036 9658 32088 9664
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 28908 9444 28960 9450
rect 28908 9386 28960 9392
rect 29288 9178 29316 9522
rect 29276 9172 29328 9178
rect 29276 9114 29328 9120
rect 29564 9110 29592 9522
rect 31024 9512 31076 9518
rect 31024 9454 31076 9460
rect 29552 9104 29604 9110
rect 29552 9046 29604 9052
rect 28776 8996 28856 9024
rect 29736 9036 29788 9042
rect 28724 8978 28776 8984
rect 29736 8978 29788 8984
rect 28736 8634 28764 8978
rect 28724 8628 28776 8634
rect 28724 8570 28776 8576
rect 29748 8430 29776 8978
rect 31036 8838 31064 9454
rect 33152 9450 33180 10134
rect 33140 9444 33192 9450
rect 33140 9386 33192 9392
rect 30012 8832 30064 8838
rect 30012 8774 30064 8780
rect 31024 8832 31076 8838
rect 31024 8774 31076 8780
rect 30024 8498 30052 8774
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 29736 8424 29788 8430
rect 29736 8366 29788 8372
rect 29368 8356 29420 8362
rect 29368 8298 29420 8304
rect 29380 8090 29408 8298
rect 29748 8090 29776 8366
rect 33244 8362 33272 10950
rect 33520 10810 33548 11154
rect 33508 10804 33560 10810
rect 33508 10746 33560 10752
rect 33612 10470 33640 11222
rect 33796 10810 33824 12038
rect 33980 11694 34008 13330
rect 34164 12753 34192 13874
rect 34532 13802 34560 13942
rect 34520 13796 34572 13802
rect 34520 13738 34572 13744
rect 34520 13388 34572 13394
rect 34520 13330 34572 13336
rect 34336 13252 34388 13258
rect 34336 13194 34388 13200
rect 34348 12986 34376 13194
rect 34532 12986 34560 13330
rect 34336 12980 34388 12986
rect 34336 12922 34388 12928
rect 34520 12980 34572 12986
rect 34520 12922 34572 12928
rect 34348 12782 34376 12922
rect 34716 12918 34744 15263
rect 34808 13326 34836 15302
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35256 15020 35308 15026
rect 35256 14962 35308 14968
rect 34980 14884 35032 14890
rect 34980 14826 35032 14832
rect 34992 14414 35020 14826
rect 35268 14550 35296 14962
rect 35360 14890 35388 15302
rect 35348 14884 35400 14890
rect 35348 14826 35400 14832
rect 35256 14544 35308 14550
rect 35256 14486 35308 14492
rect 34980 14408 35032 14414
rect 34980 14350 35032 14356
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34888 13864 34940 13870
rect 34888 13806 34940 13812
rect 34900 13462 34928 13806
rect 34888 13456 34940 13462
rect 34888 13398 34940 13404
rect 34796 13320 34848 13326
rect 34796 13262 34848 13268
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34704 12912 34756 12918
rect 34704 12854 34756 12860
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 34336 12776 34388 12782
rect 34150 12744 34206 12753
rect 34336 12718 34388 12724
rect 34150 12679 34206 12688
rect 34244 12164 34296 12170
rect 34244 12106 34296 12112
rect 33968 11688 34020 11694
rect 33968 11630 34020 11636
rect 33784 10804 33836 10810
rect 33784 10746 33836 10752
rect 33692 10736 33744 10742
rect 33692 10678 33744 10684
rect 33600 10464 33652 10470
rect 33600 10406 33652 10412
rect 33600 9036 33652 9042
rect 33704 9024 33732 10678
rect 33784 10056 33836 10062
rect 33784 9998 33836 10004
rect 33796 9586 33824 9998
rect 33784 9580 33836 9586
rect 33784 9522 33836 9528
rect 33980 9518 34008 11630
rect 34256 11558 34284 12106
rect 34244 11552 34296 11558
rect 34244 11494 34296 11500
rect 33968 9512 34020 9518
rect 33968 9454 34020 9460
rect 33980 9178 34008 9454
rect 33968 9172 34020 9178
rect 33968 9114 34020 9120
rect 33652 8996 33732 9024
rect 33600 8978 33652 8984
rect 33416 8832 33468 8838
rect 33416 8774 33468 8780
rect 33232 8356 33284 8362
rect 33232 8298 33284 8304
rect 29368 8084 29420 8090
rect 29368 8026 29420 8032
rect 29736 8084 29788 8090
rect 29736 8026 29788 8032
rect 33428 7313 33456 8774
rect 33612 8634 33640 8978
rect 33980 8634 34008 9114
rect 33600 8628 33652 8634
rect 33600 8570 33652 8576
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 34256 8498 34284 11494
rect 34348 10810 34376 12718
rect 34440 12374 34468 12786
rect 34716 12782 34744 12854
rect 34704 12776 34756 12782
rect 35268 12730 35296 14486
rect 35912 14056 35940 20159
rect 35992 17060 36044 17066
rect 35992 17002 36044 17008
rect 36004 16969 36032 17002
rect 35990 16960 36046 16969
rect 35990 16895 36046 16904
rect 35912 14028 36032 14056
rect 35900 13932 35952 13938
rect 35900 13874 35952 13880
rect 35912 13841 35940 13874
rect 35898 13832 35954 13841
rect 36004 13814 36032 14028
rect 36096 13977 36124 20334
rect 36268 19984 36320 19990
rect 36268 19926 36320 19932
rect 36176 19848 36228 19854
rect 36176 19790 36228 19796
rect 36188 19718 36216 19790
rect 36176 19712 36228 19718
rect 36176 19654 36228 19660
rect 36188 18834 36216 19654
rect 36280 19514 36308 19926
rect 36820 19848 36872 19854
rect 36820 19790 36872 19796
rect 36268 19508 36320 19514
rect 36268 19450 36320 19456
rect 36832 19446 36860 19790
rect 36820 19440 36872 19446
rect 36820 19382 36872 19388
rect 36924 19242 36952 20828
rect 37004 20392 37056 20398
rect 37004 20334 37056 20340
rect 36912 19236 36964 19242
rect 36912 19178 36964 19184
rect 36636 19168 36688 19174
rect 36636 19110 36688 19116
rect 36648 18970 36676 19110
rect 36636 18964 36688 18970
rect 36636 18906 36688 18912
rect 36176 18828 36228 18834
rect 36176 18770 36228 18776
rect 36924 18698 36952 19178
rect 36912 18692 36964 18698
rect 36912 18634 36964 18640
rect 37016 18329 37044 20334
rect 37280 20256 37332 20262
rect 37280 20198 37332 20204
rect 37292 19990 37320 20198
rect 37280 19984 37332 19990
rect 37280 19926 37332 19932
rect 37476 19854 37504 21558
rect 37648 21412 37700 21418
rect 37648 21354 37700 21360
rect 37464 19848 37516 19854
rect 37464 19790 37516 19796
rect 37660 19514 37688 21354
rect 38212 21350 38240 21966
rect 38304 21486 38332 22034
rect 38292 21480 38344 21486
rect 38292 21422 38344 21428
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 20942 38240 21286
rect 38200 20936 38252 20942
rect 38200 20878 38252 20884
rect 37924 20596 37976 20602
rect 37924 20538 37976 20544
rect 38108 20596 38160 20602
rect 38108 20538 38160 20544
rect 37740 20256 37792 20262
rect 37740 20198 37792 20204
rect 37752 19825 37780 20198
rect 37936 19990 37964 20538
rect 38120 20505 38148 20538
rect 38106 20496 38162 20505
rect 38106 20431 38162 20440
rect 37832 19984 37884 19990
rect 37832 19926 37884 19932
rect 37924 19984 37976 19990
rect 37924 19926 37976 19932
rect 37738 19816 37794 19825
rect 37738 19751 37794 19760
rect 37844 19514 37872 19926
rect 37648 19508 37700 19514
rect 37648 19450 37700 19456
rect 37832 19508 37884 19514
rect 37832 19450 37884 19456
rect 37936 19446 37964 19926
rect 37924 19440 37976 19446
rect 37924 19382 37976 19388
rect 37556 19304 37608 19310
rect 37556 19246 37608 19252
rect 37002 18320 37058 18329
rect 37002 18255 37058 18264
rect 36268 17740 36320 17746
rect 36268 17682 36320 17688
rect 36280 17270 36308 17682
rect 36728 17536 36780 17542
rect 36728 17478 36780 17484
rect 36912 17536 36964 17542
rect 36912 17478 36964 17484
rect 36268 17264 36320 17270
rect 36268 17206 36320 17212
rect 36636 17264 36688 17270
rect 36636 17206 36688 17212
rect 36648 17066 36676 17206
rect 36636 17060 36688 17066
rect 36636 17002 36688 17008
rect 36452 16992 36504 16998
rect 36452 16934 36504 16940
rect 36176 16720 36228 16726
rect 36176 16662 36228 16668
rect 36188 16250 36216 16662
rect 36360 16448 36412 16454
rect 36360 16390 36412 16396
rect 36176 16244 36228 16250
rect 36176 16186 36228 16192
rect 36188 15910 36216 16186
rect 36266 16008 36322 16017
rect 36266 15943 36322 15952
rect 36176 15904 36228 15910
rect 36176 15846 36228 15852
rect 36280 15570 36308 15943
rect 36372 15910 36400 16390
rect 36360 15904 36412 15910
rect 36360 15846 36412 15852
rect 36268 15564 36320 15570
rect 36268 15506 36320 15512
rect 36280 15201 36308 15506
rect 36266 15192 36322 15201
rect 36266 15127 36322 15136
rect 36280 15094 36308 15127
rect 36268 15088 36320 15094
rect 36268 15030 36320 15036
rect 36268 14544 36320 14550
rect 36372 14532 36400 15846
rect 36464 15706 36492 16934
rect 36648 16454 36676 17002
rect 36740 16726 36768 17478
rect 36924 17202 36952 17478
rect 36912 17196 36964 17202
rect 36912 17138 36964 17144
rect 36728 16720 36780 16726
rect 36728 16662 36780 16668
rect 36636 16448 36688 16454
rect 36636 16390 36688 16396
rect 36544 15972 36596 15978
rect 36544 15914 36596 15920
rect 36556 15706 36584 15914
rect 36452 15700 36504 15706
rect 36452 15642 36504 15648
rect 36544 15700 36596 15706
rect 36544 15642 36596 15648
rect 36648 15366 36676 16390
rect 36544 15360 36596 15366
rect 36544 15302 36596 15308
rect 36636 15360 36688 15366
rect 36636 15302 36688 15308
rect 36556 15026 36584 15302
rect 36544 15020 36596 15026
rect 36544 14962 36596 14968
rect 36648 14890 36676 15302
rect 36820 15020 36872 15026
rect 36820 14962 36872 14968
rect 36636 14884 36688 14890
rect 36636 14826 36688 14832
rect 36832 14550 36860 14962
rect 36820 14544 36872 14550
rect 36320 14504 36400 14532
rect 36648 14504 36820 14532
rect 36268 14486 36320 14492
rect 36280 14074 36308 14486
rect 36268 14068 36320 14074
rect 36268 14010 36320 14016
rect 36082 13968 36138 13977
rect 36082 13903 36138 13912
rect 36004 13786 36124 13814
rect 35898 13767 35954 13776
rect 35348 12980 35400 12986
rect 35348 12922 35400 12928
rect 35360 12782 35388 12922
rect 34704 12718 34756 12724
rect 34716 12442 34744 12718
rect 35176 12702 35296 12730
rect 35348 12776 35400 12782
rect 35348 12718 35400 12724
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 35176 12374 35204 12702
rect 35256 12640 35308 12646
rect 35256 12582 35308 12588
rect 34428 12368 34480 12374
rect 34428 12310 34480 12316
rect 34796 12368 34848 12374
rect 34796 12310 34848 12316
rect 35164 12368 35216 12374
rect 35164 12310 35216 12316
rect 34440 11898 34468 12310
rect 34428 11892 34480 11898
rect 34428 11834 34480 11840
rect 34440 11354 34468 11834
rect 34428 11348 34480 11354
rect 34428 11290 34480 11296
rect 34518 10840 34574 10849
rect 34336 10804 34388 10810
rect 34518 10775 34574 10784
rect 34336 10746 34388 10752
rect 34348 10606 34376 10746
rect 34336 10600 34388 10606
rect 34336 10542 34388 10548
rect 34532 9654 34560 10775
rect 34808 10674 34836 12310
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 35268 11762 35296 12582
rect 36096 12306 36124 13786
rect 36268 13728 36320 13734
rect 36268 13670 36320 13676
rect 36280 13462 36308 13670
rect 36268 13456 36320 13462
rect 36268 13398 36320 13404
rect 36176 13320 36228 13326
rect 36176 13262 36228 13268
rect 36188 12442 36216 13262
rect 36280 12986 36308 13398
rect 36648 13326 36676 14504
rect 36820 14486 36872 14492
rect 36820 13932 36872 13938
rect 36820 13874 36872 13880
rect 36728 13796 36780 13802
rect 36728 13738 36780 13744
rect 36740 13530 36768 13738
rect 36728 13524 36780 13530
rect 36728 13466 36780 13472
rect 36636 13320 36688 13326
rect 36636 13262 36688 13268
rect 36268 12980 36320 12986
rect 36268 12922 36320 12928
rect 36544 12708 36596 12714
rect 36544 12650 36596 12656
rect 36176 12436 36228 12442
rect 36176 12378 36228 12384
rect 36084 12300 36136 12306
rect 36084 12242 36136 12248
rect 35256 11756 35308 11762
rect 35256 11698 35308 11704
rect 35072 11552 35124 11558
rect 35072 11494 35124 11500
rect 35084 11286 35112 11494
rect 35268 11354 35296 11698
rect 35256 11348 35308 11354
rect 35256 11290 35308 11296
rect 35072 11280 35124 11286
rect 35072 11222 35124 11228
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 36096 10713 36124 12242
rect 36556 11762 36584 12650
rect 36728 12300 36780 12306
rect 36728 12242 36780 12248
rect 36740 11830 36768 12242
rect 36728 11824 36780 11830
rect 36728 11766 36780 11772
rect 36544 11756 36596 11762
rect 36544 11698 36596 11704
rect 36176 11552 36228 11558
rect 36176 11494 36228 11500
rect 36188 11286 36216 11494
rect 36176 11280 36228 11286
rect 36176 11222 36228 11228
rect 36188 10810 36216 11222
rect 36832 11082 36860 13874
rect 37016 13705 37044 18255
rect 37568 17678 37596 19246
rect 37936 18902 37964 19382
rect 37924 18896 37976 18902
rect 37844 18856 37924 18884
rect 37844 18426 37872 18856
rect 37924 18838 37976 18844
rect 37924 18760 37976 18766
rect 37924 18702 37976 18708
rect 37832 18420 37884 18426
rect 37832 18362 37884 18368
rect 37936 18154 37964 18702
rect 38108 18420 38160 18426
rect 38108 18362 38160 18368
rect 37924 18148 37976 18154
rect 37924 18090 37976 18096
rect 37648 18080 37700 18086
rect 37648 18022 37700 18028
rect 37556 17672 37608 17678
rect 37556 17614 37608 17620
rect 37372 17536 37424 17542
rect 37660 17490 37688 18022
rect 37936 17882 37964 18090
rect 37924 17876 37976 17882
rect 37924 17818 37976 17824
rect 37372 17478 37424 17484
rect 37188 17060 37240 17066
rect 37188 17002 37240 17008
rect 37200 16114 37228 17002
rect 37188 16108 37240 16114
rect 37188 16050 37240 16056
rect 37200 13938 37228 16050
rect 37384 15745 37412 17478
rect 37568 17462 37688 17490
rect 37464 16720 37516 16726
rect 37464 16662 37516 16668
rect 37370 15736 37426 15745
rect 37476 15706 37504 16662
rect 37370 15671 37426 15680
rect 37464 15700 37516 15706
rect 37464 15642 37516 15648
rect 37188 13932 37240 13938
rect 37188 13874 37240 13880
rect 37568 13841 37596 17462
rect 38016 16720 38068 16726
rect 38016 16662 38068 16668
rect 38028 15910 38056 16662
rect 37832 15904 37884 15910
rect 37832 15846 37884 15852
rect 38016 15904 38068 15910
rect 38016 15846 38068 15852
rect 37844 15706 37872 15846
rect 37832 15700 37884 15706
rect 37832 15642 37884 15648
rect 37648 14340 37700 14346
rect 37648 14282 37700 14288
rect 37660 14074 37688 14282
rect 37648 14068 37700 14074
rect 37648 14010 37700 14016
rect 37554 13832 37610 13841
rect 37554 13767 37610 13776
rect 37002 13696 37058 13705
rect 37002 13631 37058 13640
rect 38014 13696 38070 13705
rect 38014 13631 38070 13640
rect 37830 13424 37886 13433
rect 37830 13359 37832 13368
rect 37884 13359 37886 13368
rect 37832 13330 37884 13336
rect 37188 13320 37240 13326
rect 37188 13262 37240 13268
rect 37200 12850 37228 13262
rect 37844 12986 37872 13330
rect 37832 12980 37884 12986
rect 37832 12922 37884 12928
rect 37096 12844 37148 12850
rect 37096 12786 37148 12792
rect 37188 12844 37240 12850
rect 37188 12786 37240 12792
rect 37004 12708 37056 12714
rect 37004 12650 37056 12656
rect 36912 12096 36964 12102
rect 36912 12038 36964 12044
rect 36924 11286 36952 12038
rect 37016 11558 37044 12650
rect 37108 12102 37136 12786
rect 37096 12096 37148 12102
rect 37096 12038 37148 12044
rect 37004 11552 37056 11558
rect 37004 11494 37056 11500
rect 37016 11354 37044 11494
rect 37004 11348 37056 11354
rect 37004 11290 37056 11296
rect 36912 11280 36964 11286
rect 36912 11222 36964 11228
rect 36912 11144 36964 11150
rect 36912 11086 36964 11092
rect 36728 11076 36780 11082
rect 36728 11018 36780 11024
rect 36820 11076 36872 11082
rect 36820 11018 36872 11024
rect 36176 10804 36228 10810
rect 36176 10746 36228 10752
rect 36740 10742 36768 11018
rect 36728 10736 36780 10742
rect 36082 10704 36138 10713
rect 34796 10668 34848 10674
rect 36728 10678 36780 10684
rect 36832 10674 36860 11018
rect 36082 10639 36138 10648
rect 36820 10668 36872 10674
rect 34796 10610 34848 10616
rect 36820 10610 36872 10616
rect 34612 10464 34664 10470
rect 34612 10406 34664 10412
rect 34624 10266 34652 10406
rect 34808 10266 34836 10610
rect 36728 10464 36780 10470
rect 36728 10406 36780 10412
rect 34612 10260 34664 10266
rect 34612 10202 34664 10208
rect 34796 10260 34848 10266
rect 34796 10202 34848 10208
rect 36084 10260 36136 10266
rect 36084 10202 36136 10208
rect 35716 10056 35768 10062
rect 35716 9998 35768 10004
rect 34704 9988 34756 9994
rect 34704 9930 34756 9936
rect 34520 9648 34572 9654
rect 34520 9590 34572 9596
rect 34244 8492 34296 8498
rect 34244 8434 34296 8440
rect 34532 8430 34560 9590
rect 34716 9586 34744 9930
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34704 9580 34756 9586
rect 34704 9522 34756 9528
rect 34716 9042 34744 9522
rect 35728 9178 35756 9998
rect 35808 9512 35860 9518
rect 35808 9454 35860 9460
rect 35716 9172 35768 9178
rect 35716 9114 35768 9120
rect 34704 9036 34756 9042
rect 34704 8978 34756 8984
rect 34520 8424 34572 8430
rect 34520 8366 34572 8372
rect 34716 8090 34744 8978
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 35728 8498 35756 9114
rect 35820 9110 35848 9454
rect 36096 9450 36124 10202
rect 36544 10124 36596 10130
rect 36544 10066 36596 10072
rect 36084 9444 36136 9450
rect 36084 9386 36136 9392
rect 35808 9104 35860 9110
rect 35808 9046 35860 9052
rect 36556 9042 36584 10066
rect 36740 9722 36768 10406
rect 36832 10130 36860 10610
rect 36924 10198 36952 11086
rect 36912 10192 36964 10198
rect 36912 10134 36964 10140
rect 36820 10124 36872 10130
rect 36820 10066 36872 10072
rect 36728 9716 36780 9722
rect 36728 9658 36780 9664
rect 37108 9178 37136 12038
rect 37200 11150 37228 12786
rect 38028 12306 38056 13631
rect 38016 12300 38068 12306
rect 38016 12242 38068 12248
rect 38028 11898 38056 12242
rect 38016 11892 38068 11898
rect 38016 11834 38068 11840
rect 37464 11756 37516 11762
rect 37464 11698 37516 11704
rect 37924 11756 37976 11762
rect 37924 11698 37976 11704
rect 37476 11354 37504 11698
rect 37740 11552 37792 11558
rect 37740 11494 37792 11500
rect 37752 11354 37780 11494
rect 37464 11348 37516 11354
rect 37464 11290 37516 11296
rect 37740 11348 37792 11354
rect 37740 11290 37792 11296
rect 37188 11144 37240 11150
rect 37188 11086 37240 11092
rect 37752 10810 37780 11290
rect 37832 11280 37884 11286
rect 37832 11222 37884 11228
rect 37844 10810 37872 11222
rect 37740 10804 37792 10810
rect 37740 10746 37792 10752
rect 37832 10804 37884 10810
rect 37832 10746 37884 10752
rect 37740 10260 37792 10266
rect 37740 10202 37792 10208
rect 37752 9722 37780 10202
rect 37936 10062 37964 11698
rect 38120 11121 38148 18362
rect 38200 17264 38252 17270
rect 38200 17206 38252 17212
rect 38212 17066 38240 17206
rect 38200 17060 38252 17066
rect 38200 17002 38252 17008
rect 38200 15564 38252 15570
rect 38200 15506 38252 15512
rect 38212 15094 38240 15506
rect 38200 15088 38252 15094
rect 38200 15030 38252 15036
rect 38200 14000 38252 14006
rect 38200 13942 38252 13948
rect 38212 13190 38240 13942
rect 38304 13569 38332 21422
rect 38396 17746 38424 22170
rect 38476 20868 38528 20874
rect 38476 20810 38528 20816
rect 38488 20466 38516 20810
rect 39040 20534 39068 22646
rect 39224 22098 39252 25094
rect 39316 24954 39344 25230
rect 39304 24948 39356 24954
rect 39304 24890 39356 24896
rect 39304 24336 39356 24342
rect 39304 24278 39356 24284
rect 39316 23526 39344 24278
rect 39684 23594 39712 27814
rect 39776 27606 39804 27882
rect 39764 27600 39816 27606
rect 39764 27542 39816 27548
rect 39856 27600 39908 27606
rect 39856 27542 39908 27548
rect 39776 27130 39804 27542
rect 39764 27124 39816 27130
rect 39764 27066 39816 27072
rect 39764 26784 39816 26790
rect 39868 26772 39896 27542
rect 39960 26858 39988 28426
rect 40052 27470 40080 28630
rect 40144 28218 40172 28698
rect 40132 28212 40184 28218
rect 40132 28154 40184 28160
rect 40040 27464 40092 27470
rect 40040 27406 40092 27412
rect 39948 26852 40000 26858
rect 39948 26794 40000 26800
rect 39816 26744 39896 26772
rect 39764 26726 39816 26732
rect 39776 26518 39804 26726
rect 39764 26512 39816 26518
rect 39764 26454 39816 26460
rect 39776 25702 39804 26454
rect 39764 25696 39816 25702
rect 39764 25638 39816 25644
rect 39776 25430 39804 25638
rect 39764 25424 39816 25430
rect 39764 25366 39816 25372
rect 39776 24954 39804 25366
rect 39764 24948 39816 24954
rect 39764 24890 39816 24896
rect 39960 24818 39988 26794
rect 40328 26314 40356 29446
rect 40604 29306 40632 29718
rect 40592 29300 40644 29306
rect 40592 29242 40644 29248
rect 40684 28552 40736 28558
rect 40736 28512 40816 28540
rect 40684 28494 40736 28500
rect 40408 28008 40460 28014
rect 40408 27950 40460 27956
rect 40316 26308 40368 26314
rect 40316 26250 40368 26256
rect 40328 25430 40356 26250
rect 40316 25424 40368 25430
rect 40316 25366 40368 25372
rect 39948 24812 40000 24818
rect 39948 24754 40000 24760
rect 40420 24750 40448 27950
rect 40788 27402 40816 28512
rect 41064 28014 41092 31078
rect 41144 30796 41196 30802
rect 41144 30738 41196 30744
rect 41156 29850 41184 30738
rect 41788 30592 41840 30598
rect 41788 30534 41840 30540
rect 41328 30252 41380 30258
rect 41328 30194 41380 30200
rect 41144 29844 41196 29850
rect 41144 29786 41196 29792
rect 41144 29640 41196 29646
rect 41144 29582 41196 29588
rect 41156 29050 41184 29582
rect 41236 29572 41288 29578
rect 41236 29514 41288 29520
rect 41248 29170 41276 29514
rect 41236 29164 41288 29170
rect 41236 29106 41288 29112
rect 41156 29034 41276 29050
rect 41156 29028 41288 29034
rect 41156 29022 41236 29028
rect 41236 28970 41288 28976
rect 41144 28960 41196 28966
rect 41144 28902 41196 28908
rect 41156 28762 41184 28902
rect 41144 28756 41196 28762
rect 41144 28698 41196 28704
rect 41248 28490 41276 28970
rect 41236 28484 41288 28490
rect 41236 28426 41288 28432
rect 41052 28008 41104 28014
rect 41052 27950 41104 27956
rect 40776 27396 40828 27402
rect 40776 27338 40828 27344
rect 40788 26518 40816 27338
rect 41340 26926 41368 30194
rect 41696 29708 41748 29714
rect 41696 29650 41748 29656
rect 41708 28966 41736 29650
rect 41696 28960 41748 28966
rect 41696 28902 41748 28908
rect 41512 27872 41564 27878
rect 41512 27814 41564 27820
rect 41524 27606 41552 27814
rect 41708 27713 41736 28902
rect 41800 28694 41828 30534
rect 41984 30190 42012 33079
rect 42064 32768 42116 32774
rect 42064 32710 42116 32716
rect 42076 32502 42104 32710
rect 42064 32496 42116 32502
rect 42064 32438 42116 32444
rect 42168 31278 42196 33106
rect 42708 33108 42760 33114
rect 42708 33050 42760 33056
rect 42812 33046 42840 33322
rect 43088 33114 43116 33934
rect 43548 33386 43576 34070
rect 43536 33380 43588 33386
rect 43536 33322 43588 33328
rect 43076 33108 43128 33114
rect 43076 33050 43128 33056
rect 42800 33040 42852 33046
rect 42800 32982 42852 32988
rect 43352 32972 43404 32978
rect 43352 32914 43404 32920
rect 42432 32428 42484 32434
rect 42432 32370 42484 32376
rect 42444 32337 42472 32370
rect 42430 32328 42486 32337
rect 42430 32263 42486 32272
rect 43364 32230 43392 32914
rect 43536 32428 43588 32434
rect 43536 32370 43588 32376
rect 43352 32224 43404 32230
rect 43352 32166 43404 32172
rect 42156 31272 42208 31278
rect 42156 31214 42208 31220
rect 42708 31136 42760 31142
rect 42708 31078 42760 31084
rect 41972 30184 42024 30190
rect 41972 30126 42024 30132
rect 41880 30048 41932 30054
rect 41880 29990 41932 29996
rect 42524 30048 42576 30054
rect 42524 29990 42576 29996
rect 41892 29306 41920 29990
rect 42536 29850 42564 29990
rect 42524 29844 42576 29850
rect 42524 29786 42576 29792
rect 42340 29572 42392 29578
rect 42340 29514 42392 29520
rect 41880 29300 41932 29306
rect 41880 29242 41932 29248
rect 41892 29016 41920 29242
rect 41972 29028 42024 29034
rect 41892 28988 41972 29016
rect 41892 28694 41920 28988
rect 41972 28970 42024 28976
rect 41788 28688 41840 28694
rect 41788 28630 41840 28636
rect 41880 28688 41932 28694
rect 41880 28630 41932 28636
rect 41694 27704 41750 27713
rect 41800 27674 41828 28630
rect 41694 27639 41750 27648
rect 41788 27668 41840 27674
rect 41788 27610 41840 27616
rect 41512 27600 41564 27606
rect 41512 27542 41564 27548
rect 41524 27062 41552 27542
rect 42352 27062 42380 29514
rect 42536 29238 42564 29786
rect 42524 29232 42576 29238
rect 42524 29174 42576 29180
rect 42432 29164 42484 29170
rect 42432 29106 42484 29112
rect 42444 27606 42472 29106
rect 42524 28552 42576 28558
rect 42524 28494 42576 28500
rect 42536 27946 42564 28494
rect 42524 27940 42576 27946
rect 42524 27882 42576 27888
rect 42432 27600 42484 27606
rect 42432 27542 42484 27548
rect 42444 27402 42472 27542
rect 42432 27396 42484 27402
rect 42432 27338 42484 27344
rect 41512 27056 41564 27062
rect 42340 27056 42392 27062
rect 41512 26998 41564 27004
rect 42260 27016 42340 27044
rect 40868 26920 40920 26926
rect 40868 26862 40920 26868
rect 41328 26920 41380 26926
rect 41328 26862 41380 26868
rect 40776 26512 40828 26518
rect 40776 26454 40828 26460
rect 40776 25696 40828 25702
rect 40776 25638 40828 25644
rect 40408 24744 40460 24750
rect 40408 24686 40460 24692
rect 39764 24608 39816 24614
rect 39764 24550 39816 24556
rect 39776 24206 39804 24550
rect 39764 24200 39816 24206
rect 39764 24142 39816 24148
rect 39672 23588 39724 23594
rect 39672 23530 39724 23536
rect 40408 23588 40460 23594
rect 40408 23530 40460 23536
rect 39304 23520 39356 23526
rect 39304 23462 39356 23468
rect 39316 23254 39344 23462
rect 39304 23248 39356 23254
rect 39304 23190 39356 23196
rect 39316 22438 39344 23190
rect 39396 23112 39448 23118
rect 39396 23054 39448 23060
rect 39408 22642 39436 23054
rect 39396 22636 39448 22642
rect 39396 22578 39448 22584
rect 40420 22574 40448 23530
rect 40788 23118 40816 25638
rect 40880 24585 40908 26862
rect 41524 26858 41552 26998
rect 41604 26988 41656 26994
rect 41604 26930 41656 26936
rect 41512 26852 41564 26858
rect 41512 26794 41564 26800
rect 41052 26784 41104 26790
rect 41052 26726 41104 26732
rect 41064 26586 41092 26726
rect 41052 26580 41104 26586
rect 41052 26522 41104 26528
rect 41616 26518 41644 26930
rect 41604 26512 41656 26518
rect 41604 26454 41656 26460
rect 41880 26512 41932 26518
rect 41880 26454 41932 26460
rect 41788 26376 41840 26382
rect 41788 26318 41840 26324
rect 41800 26042 41828 26318
rect 41788 26036 41840 26042
rect 41788 25978 41840 25984
rect 40960 25832 41012 25838
rect 40960 25774 41012 25780
rect 40972 25673 41000 25774
rect 41892 25770 41920 26454
rect 42260 25974 42288 27016
rect 42340 26998 42392 27004
rect 42444 26518 42472 27338
rect 42432 26512 42484 26518
rect 42432 26454 42484 26460
rect 42536 26314 42564 27882
rect 42524 26308 42576 26314
rect 42524 26250 42576 26256
rect 42340 26036 42392 26042
rect 42340 25978 42392 25984
rect 42248 25968 42300 25974
rect 42248 25910 42300 25916
rect 41696 25764 41748 25770
rect 41696 25706 41748 25712
rect 41880 25764 41932 25770
rect 41880 25706 41932 25712
rect 41604 25696 41656 25702
rect 40958 25664 41014 25673
rect 41604 25638 41656 25644
rect 40958 25599 41014 25608
rect 40972 24721 41000 25599
rect 41616 25498 41644 25638
rect 41708 25498 41736 25706
rect 41604 25492 41656 25498
rect 41604 25434 41656 25440
rect 41696 25492 41748 25498
rect 41696 25434 41748 25440
rect 41972 25356 42024 25362
rect 41972 25298 42024 25304
rect 42064 25356 42116 25362
rect 42064 25298 42116 25304
rect 41052 25152 41104 25158
rect 41052 25094 41104 25100
rect 41144 25152 41196 25158
rect 41144 25094 41196 25100
rect 40958 24712 41014 24721
rect 41064 24682 41092 25094
rect 40958 24647 41014 24656
rect 41052 24676 41104 24682
rect 41052 24618 41104 24624
rect 40866 24576 40922 24585
rect 40866 24511 40922 24520
rect 40500 23112 40552 23118
rect 40500 23054 40552 23060
rect 40776 23112 40828 23118
rect 40776 23054 40828 23060
rect 40512 22778 40540 23054
rect 40500 22772 40552 22778
rect 40500 22714 40552 22720
rect 40408 22568 40460 22574
rect 40408 22510 40460 22516
rect 40880 22506 40908 24511
rect 41064 22778 41092 24618
rect 41156 23730 41184 25094
rect 41984 24954 42012 25298
rect 41972 24948 42024 24954
rect 41972 24890 42024 24896
rect 41788 24676 41840 24682
rect 41788 24618 41840 24624
rect 41328 24608 41380 24614
rect 41328 24550 41380 24556
rect 41420 24608 41472 24614
rect 41420 24550 41472 24556
rect 41340 24342 41368 24550
rect 41328 24336 41380 24342
rect 41328 24278 41380 24284
rect 41144 23724 41196 23730
rect 41144 23666 41196 23672
rect 41340 23594 41368 24278
rect 41432 23866 41460 24550
rect 41512 24200 41564 24206
rect 41512 24142 41564 24148
rect 41524 23866 41552 24142
rect 41420 23860 41472 23866
rect 41420 23802 41472 23808
rect 41512 23860 41564 23866
rect 41512 23802 41564 23808
rect 41328 23588 41380 23594
rect 41328 23530 41380 23536
rect 41696 23588 41748 23594
rect 41696 23530 41748 23536
rect 41340 23254 41368 23530
rect 41328 23248 41380 23254
rect 41328 23190 41380 23196
rect 41340 22778 41368 23190
rect 41708 23118 41736 23530
rect 41696 23112 41748 23118
rect 41696 23054 41748 23060
rect 41052 22772 41104 22778
rect 41052 22714 41104 22720
rect 41328 22772 41380 22778
rect 41328 22714 41380 22720
rect 40868 22500 40920 22506
rect 40868 22442 40920 22448
rect 39304 22432 39356 22438
rect 39304 22374 39356 22380
rect 40316 22432 40368 22438
rect 40316 22374 40368 22380
rect 41144 22432 41196 22438
rect 41144 22374 41196 22380
rect 39212 22092 39264 22098
rect 39212 22034 39264 22040
rect 39224 21486 39252 22034
rect 39488 22024 39540 22030
rect 39488 21966 39540 21972
rect 39212 21480 39264 21486
rect 39212 21422 39264 21428
rect 39224 21078 39252 21422
rect 39212 21072 39264 21078
rect 39212 21014 39264 21020
rect 39028 20528 39080 20534
rect 39028 20470 39080 20476
rect 38476 20460 38528 20466
rect 38476 20402 38528 20408
rect 38476 20324 38528 20330
rect 38476 20266 38528 20272
rect 38488 18086 38516 20266
rect 39224 19990 39252 21014
rect 39500 21010 39528 21966
rect 40328 21350 40356 22374
rect 40592 21956 40644 21962
rect 40592 21898 40644 21904
rect 40960 21956 41012 21962
rect 40960 21898 41012 21904
rect 40500 21888 40552 21894
rect 40500 21830 40552 21836
rect 40512 21554 40540 21830
rect 40500 21548 40552 21554
rect 40500 21490 40552 21496
rect 40316 21344 40368 21350
rect 40316 21286 40368 21292
rect 40328 21078 40356 21286
rect 40316 21072 40368 21078
rect 40316 21014 40368 21020
rect 39488 21004 39540 21010
rect 39488 20946 39540 20952
rect 39304 20800 39356 20806
rect 39304 20742 39356 20748
rect 39212 19984 39264 19990
rect 39212 19926 39264 19932
rect 39224 19310 39252 19926
rect 39316 19922 39344 20742
rect 39500 20602 39528 20946
rect 39488 20596 39540 20602
rect 39488 20538 39540 20544
rect 40328 20262 40356 21014
rect 40316 20256 40368 20262
rect 40316 20198 40368 20204
rect 39304 19916 39356 19922
rect 39304 19858 39356 19864
rect 39316 19514 39344 19858
rect 39304 19508 39356 19514
rect 39304 19450 39356 19456
rect 39212 19304 39264 19310
rect 39212 19246 39264 19252
rect 39224 18970 39252 19246
rect 39212 18964 39264 18970
rect 39212 18906 39264 18912
rect 39224 18222 39252 18906
rect 39316 18426 39344 19450
rect 40328 19174 40356 20198
rect 40604 19718 40632 21898
rect 40776 20936 40828 20942
rect 40776 20878 40828 20884
rect 40788 20602 40816 20878
rect 40776 20596 40828 20602
rect 40776 20538 40828 20544
rect 40972 20330 41000 21898
rect 41052 21072 41104 21078
rect 41052 21014 41104 21020
rect 41064 20806 41092 21014
rect 41052 20800 41104 20806
rect 41052 20742 41104 20748
rect 41064 20602 41092 20742
rect 41052 20596 41104 20602
rect 41052 20538 41104 20544
rect 40960 20324 41012 20330
rect 40960 20266 41012 20272
rect 40972 20058 41000 20266
rect 40960 20052 41012 20058
rect 40960 19994 41012 20000
rect 40500 19712 40552 19718
rect 40500 19654 40552 19660
rect 40592 19712 40644 19718
rect 40592 19654 40644 19660
rect 40512 19378 40540 19654
rect 40500 19372 40552 19378
rect 40500 19314 40552 19320
rect 40316 19168 40368 19174
rect 40316 19110 40368 19116
rect 40328 18902 40356 19110
rect 40316 18896 40368 18902
rect 40316 18838 40368 18844
rect 39580 18624 39632 18630
rect 39580 18566 39632 18572
rect 40132 18624 40184 18630
rect 40132 18566 40184 18572
rect 39304 18420 39356 18426
rect 39304 18362 39356 18368
rect 39592 18290 39620 18566
rect 40040 18352 40092 18358
rect 40040 18294 40092 18300
rect 39580 18284 39632 18290
rect 39580 18226 39632 18232
rect 38660 18216 38712 18222
rect 38658 18184 38660 18193
rect 39028 18216 39080 18222
rect 38712 18184 38714 18193
rect 39028 18158 39080 18164
rect 39212 18216 39264 18222
rect 39212 18158 39264 18164
rect 38658 18119 38714 18128
rect 38672 18086 38700 18119
rect 38476 18080 38528 18086
rect 38476 18022 38528 18028
rect 38660 18080 38712 18086
rect 38660 18022 38712 18028
rect 38384 17740 38436 17746
rect 38384 17682 38436 17688
rect 38844 17740 38896 17746
rect 38844 17682 38896 17688
rect 38396 17610 38424 17682
rect 38384 17604 38436 17610
rect 38384 17546 38436 17552
rect 38856 17270 38884 17682
rect 38844 17264 38896 17270
rect 38844 17206 38896 17212
rect 38476 17196 38528 17202
rect 38476 17138 38528 17144
rect 38488 16726 38516 17138
rect 38568 17060 38620 17066
rect 38568 17002 38620 17008
rect 38476 16720 38528 16726
rect 38476 16662 38528 16668
rect 38384 14068 38436 14074
rect 38384 14010 38436 14016
rect 38396 13802 38424 14010
rect 38488 13938 38516 16662
rect 38580 16182 38608 17002
rect 38568 16176 38620 16182
rect 38568 16118 38620 16124
rect 38568 16040 38620 16046
rect 38568 15982 38620 15988
rect 38580 15706 38608 15982
rect 38568 15700 38620 15706
rect 38568 15642 38620 15648
rect 38752 15564 38804 15570
rect 38752 15506 38804 15512
rect 38764 15162 38792 15506
rect 38752 15156 38804 15162
rect 38752 15098 38804 15104
rect 38476 13932 38528 13938
rect 38476 13874 38528 13880
rect 38384 13796 38436 13802
rect 38384 13738 38436 13744
rect 38290 13560 38346 13569
rect 38290 13495 38346 13504
rect 38304 13258 38332 13495
rect 38292 13252 38344 13258
rect 38292 13194 38344 13200
rect 38200 13184 38252 13190
rect 38200 13126 38252 13132
rect 38212 12442 38240 13126
rect 38200 12436 38252 12442
rect 38200 12378 38252 12384
rect 38488 11762 38516 13874
rect 38660 11892 38712 11898
rect 38660 11834 38712 11840
rect 38476 11756 38528 11762
rect 38476 11698 38528 11704
rect 38672 11694 38700 11834
rect 38660 11688 38712 11694
rect 38580 11648 38660 11676
rect 38106 11112 38162 11121
rect 38106 11047 38162 11056
rect 38108 10668 38160 10674
rect 38108 10610 38160 10616
rect 38120 10062 38148 10610
rect 37924 10056 37976 10062
rect 37924 9998 37976 10004
rect 38108 10056 38160 10062
rect 38108 9998 38160 10004
rect 37936 9722 37964 9998
rect 37740 9716 37792 9722
rect 37740 9658 37792 9664
rect 37924 9716 37976 9722
rect 37924 9658 37976 9664
rect 38580 9654 38608 11648
rect 38660 11630 38712 11636
rect 39040 11014 39068 18158
rect 39224 17814 39252 18158
rect 39672 18080 39724 18086
rect 39672 18022 39724 18028
rect 39212 17808 39264 17814
rect 39212 17750 39264 17756
rect 39224 17270 39252 17750
rect 39488 17740 39540 17746
rect 39488 17682 39540 17688
rect 39212 17264 39264 17270
rect 39212 17206 39264 17212
rect 39500 16998 39528 17682
rect 39488 16992 39540 16998
rect 39488 16934 39540 16940
rect 39302 16824 39358 16833
rect 39302 16759 39358 16768
rect 39316 16658 39344 16759
rect 39304 16652 39356 16658
rect 39304 16594 39356 16600
rect 39316 16250 39344 16594
rect 39500 16454 39528 16934
rect 39488 16448 39540 16454
rect 39488 16390 39540 16396
rect 39304 16244 39356 16250
rect 39304 16186 39356 16192
rect 39500 15570 39528 16390
rect 39684 15978 39712 18022
rect 40052 17746 40080 18294
rect 40144 17882 40172 18566
rect 40328 18086 40356 18838
rect 40500 18216 40552 18222
rect 40500 18158 40552 18164
rect 40316 18080 40368 18086
rect 40316 18022 40368 18028
rect 40512 17882 40540 18158
rect 40132 17876 40184 17882
rect 40132 17818 40184 17824
rect 40500 17876 40552 17882
rect 40500 17818 40552 17824
rect 40040 17740 40092 17746
rect 40040 17682 40092 17688
rect 40052 17270 40080 17682
rect 40040 17264 40092 17270
rect 40040 17206 40092 17212
rect 40868 17060 40920 17066
rect 40868 17002 40920 17008
rect 40316 16992 40368 16998
rect 40316 16934 40368 16940
rect 40328 16794 40356 16934
rect 40316 16788 40368 16794
rect 40316 16730 40368 16736
rect 40328 16114 40356 16730
rect 40880 16726 40908 17002
rect 41156 16998 41184 22374
rect 41696 22160 41748 22166
rect 41696 22102 41748 22108
rect 41328 22024 41380 22030
rect 41328 21966 41380 21972
rect 41340 21146 41368 21966
rect 41708 21350 41736 22102
rect 41800 22030 41828 24618
rect 42076 24410 42104 25298
rect 42352 25294 42380 25978
rect 42720 25838 42748 31078
rect 43364 30258 43392 32166
rect 43444 31816 43496 31822
rect 43444 31758 43496 31764
rect 43456 31482 43484 31758
rect 43444 31476 43496 31482
rect 43444 31418 43496 31424
rect 43548 31346 43576 32370
rect 43640 31482 43668 37742
rect 43824 37670 43852 38354
rect 43812 37664 43864 37670
rect 43812 37606 43864 37612
rect 43824 37369 43852 37606
rect 43810 37360 43866 37369
rect 43810 37295 43866 37304
rect 43824 34785 43852 37295
rect 43904 36236 43956 36242
rect 43904 36178 43956 36184
rect 43916 35494 43944 36178
rect 43904 35488 43956 35494
rect 43904 35430 43956 35436
rect 43810 34776 43866 34785
rect 43810 34711 43866 34720
rect 43824 32978 43852 34711
rect 43812 32972 43864 32978
rect 43812 32914 43864 32920
rect 43628 31476 43680 31482
rect 43628 31418 43680 31424
rect 43536 31340 43588 31346
rect 43536 31282 43588 31288
rect 43640 31278 43668 31418
rect 43628 31272 43680 31278
rect 43628 31214 43680 31220
rect 43352 30252 43404 30258
rect 43352 30194 43404 30200
rect 43536 29776 43588 29782
rect 43536 29718 43588 29724
rect 43444 29640 43496 29646
rect 43444 29582 43496 29588
rect 43456 29170 43484 29582
rect 43548 29306 43576 29718
rect 43536 29300 43588 29306
rect 43536 29242 43588 29248
rect 43444 29164 43496 29170
rect 43444 29106 43496 29112
rect 42800 28688 42852 28694
rect 42800 28630 42852 28636
rect 42812 28218 42840 28630
rect 42800 28212 42852 28218
rect 42800 28154 42852 28160
rect 43916 27538 43944 35430
rect 44364 34468 44416 34474
rect 44364 34410 44416 34416
rect 44376 33386 44404 34410
rect 44548 33516 44600 33522
rect 44548 33458 44600 33464
rect 44088 33380 44140 33386
rect 44088 33322 44140 33328
rect 44364 33380 44416 33386
rect 44364 33322 44416 33328
rect 43996 33312 44048 33318
rect 43996 33254 44048 33260
rect 44008 32910 44036 33254
rect 43996 32904 44048 32910
rect 43996 32846 44048 32852
rect 44100 32774 44128 33322
rect 44376 33114 44404 33322
rect 44364 33108 44416 33114
rect 44364 33050 44416 33056
rect 44088 32768 44140 32774
rect 44088 32710 44140 32716
rect 44100 32298 44128 32710
rect 44560 32502 44588 33458
rect 44548 32496 44600 32502
rect 44548 32438 44600 32444
rect 44088 32292 44140 32298
rect 44088 32234 44140 32240
rect 44100 31958 44128 32234
rect 44088 31952 44140 31958
rect 44088 31894 44140 31900
rect 44100 31482 44128 31894
rect 44088 31476 44140 31482
rect 44088 31418 44140 31424
rect 44824 27872 44876 27878
rect 44824 27814 44876 27820
rect 44546 27568 44602 27577
rect 43904 27532 43956 27538
rect 44546 27503 44602 27512
rect 43904 27474 43956 27480
rect 43168 27328 43220 27334
rect 43168 27270 43220 27276
rect 43180 27130 43208 27270
rect 43916 27130 43944 27474
rect 43168 27124 43220 27130
rect 43168 27066 43220 27072
rect 43904 27124 43956 27130
rect 43904 27066 43956 27072
rect 42984 26920 43036 26926
rect 42984 26862 43036 26868
rect 42708 25832 42760 25838
rect 42708 25774 42760 25780
rect 42340 25288 42392 25294
rect 42340 25230 42392 25236
rect 42720 24750 42748 25774
rect 42708 24744 42760 24750
rect 42708 24686 42760 24692
rect 42996 24449 43024 26862
rect 43076 26580 43128 26586
rect 43076 26522 43128 26528
rect 43088 26042 43116 26522
rect 43536 26512 43588 26518
rect 43536 26454 43588 26460
rect 43076 26036 43128 26042
rect 43076 25978 43128 25984
rect 43548 25770 43576 26454
rect 43536 25764 43588 25770
rect 43536 25706 43588 25712
rect 43076 25696 43128 25702
rect 43076 25638 43128 25644
rect 43088 25498 43116 25638
rect 44560 25498 44588 27503
rect 44640 25832 44692 25838
rect 44640 25774 44692 25780
rect 44652 25673 44680 25774
rect 44638 25664 44694 25673
rect 44638 25599 44694 25608
rect 43076 25492 43128 25498
rect 43076 25434 43128 25440
rect 44548 25492 44600 25498
rect 44548 25434 44600 25440
rect 43260 25356 43312 25362
rect 43260 25298 43312 25304
rect 44640 25356 44692 25362
rect 44640 25298 44692 25304
rect 43272 24954 43300 25298
rect 43260 24948 43312 24954
rect 43260 24890 43312 24896
rect 43996 24880 44048 24886
rect 43996 24822 44048 24828
rect 43168 24608 43220 24614
rect 43168 24550 43220 24556
rect 43536 24608 43588 24614
rect 43536 24550 43588 24556
rect 42982 24440 43038 24449
rect 42064 24404 42116 24410
rect 42982 24375 43038 24384
rect 42064 24346 42116 24352
rect 41880 24132 41932 24138
rect 41880 24074 41932 24080
rect 41892 23254 41920 24074
rect 42076 23866 42104 24346
rect 42064 23860 42116 23866
rect 42064 23802 42116 23808
rect 42524 23860 42576 23866
rect 42524 23802 42576 23808
rect 41880 23248 41932 23254
rect 41880 23190 41932 23196
rect 42064 23112 42116 23118
rect 42064 23054 42116 23060
rect 41880 22432 41932 22438
rect 41880 22374 41932 22380
rect 41892 22234 41920 22374
rect 41880 22228 41932 22234
rect 41880 22170 41932 22176
rect 41788 22024 41840 22030
rect 41788 21966 41840 21972
rect 41420 21344 41472 21350
rect 41420 21286 41472 21292
rect 41696 21344 41748 21350
rect 41696 21286 41748 21292
rect 41328 21140 41380 21146
rect 41328 21082 41380 21088
rect 41432 20330 41460 21286
rect 41708 21078 41736 21286
rect 42076 21078 42104 23054
rect 42340 22228 42392 22234
rect 42340 22170 42392 22176
rect 42352 21554 42380 22170
rect 42340 21548 42392 21554
rect 42340 21490 42392 21496
rect 41696 21072 41748 21078
rect 41696 21014 41748 21020
rect 42064 21072 42116 21078
rect 42064 21014 42116 21020
rect 42076 20534 42104 21014
rect 42064 20528 42116 20534
rect 42064 20470 42116 20476
rect 41420 20324 41472 20330
rect 41420 20266 41472 20272
rect 41972 20324 42024 20330
rect 41972 20266 42024 20272
rect 41432 20058 41460 20266
rect 41420 20052 41472 20058
rect 41420 19994 41472 20000
rect 41788 19984 41840 19990
rect 41788 19926 41840 19932
rect 41512 19848 41564 19854
rect 41512 19790 41564 19796
rect 41524 19378 41552 19790
rect 41800 19514 41828 19926
rect 41984 19854 42012 20266
rect 41972 19848 42024 19854
rect 41972 19790 42024 19796
rect 41880 19712 41932 19718
rect 41880 19654 41932 19660
rect 41788 19508 41840 19514
rect 41788 19450 41840 19456
rect 41512 19372 41564 19378
rect 41512 19314 41564 19320
rect 41892 18834 41920 19654
rect 41880 18828 41932 18834
rect 41880 18770 41932 18776
rect 41892 18426 41920 18770
rect 41880 18420 41932 18426
rect 41880 18362 41932 18368
rect 41984 18068 42012 19790
rect 42076 19786 42104 20470
rect 42064 19780 42116 19786
rect 42064 19722 42116 19728
rect 42432 19372 42484 19378
rect 42432 19314 42484 19320
rect 42444 18902 42472 19314
rect 42432 18896 42484 18902
rect 42432 18838 42484 18844
rect 42340 18692 42392 18698
rect 42392 18652 42472 18680
rect 42340 18634 42392 18640
rect 42340 18284 42392 18290
rect 42340 18226 42392 18232
rect 42352 18154 42380 18226
rect 42444 18154 42472 18652
rect 42340 18148 42392 18154
rect 42340 18090 42392 18096
rect 42432 18148 42484 18154
rect 42432 18090 42484 18096
rect 42064 18080 42116 18086
rect 41984 18040 42064 18068
rect 41984 17746 42012 18040
rect 42064 18022 42116 18028
rect 42352 17882 42380 18090
rect 42340 17876 42392 17882
rect 42340 17818 42392 17824
rect 42444 17746 42472 18090
rect 41972 17740 42024 17746
rect 41972 17682 42024 17688
rect 42432 17740 42484 17746
rect 42432 17682 42484 17688
rect 41984 17338 42012 17682
rect 42064 17672 42116 17678
rect 42064 17614 42116 17620
rect 41972 17332 42024 17338
rect 41972 17274 42024 17280
rect 41144 16992 41196 16998
rect 41144 16934 41196 16940
rect 40868 16720 40920 16726
rect 40868 16662 40920 16668
rect 41052 16720 41104 16726
rect 41052 16662 41104 16668
rect 40316 16108 40368 16114
rect 40316 16050 40368 16056
rect 41064 15978 41092 16662
rect 42076 16114 42104 17614
rect 42536 16969 42564 23802
rect 42892 23520 42944 23526
rect 42892 23462 42944 23468
rect 42904 22982 42932 23462
rect 42892 22976 42944 22982
rect 42892 22918 42944 22924
rect 42904 22438 42932 22918
rect 42892 22432 42944 22438
rect 42892 22374 42944 22380
rect 42996 22098 43024 24375
rect 43180 23730 43208 24550
rect 43260 24200 43312 24206
rect 43260 24142 43312 24148
rect 43444 24200 43496 24206
rect 43444 24142 43496 24148
rect 43272 23730 43300 24142
rect 43456 23798 43484 24142
rect 43444 23792 43496 23798
rect 43444 23734 43496 23740
rect 43168 23724 43220 23730
rect 43168 23666 43220 23672
rect 43260 23724 43312 23730
rect 43260 23666 43312 23672
rect 43180 23322 43208 23666
rect 43168 23316 43220 23322
rect 43168 23258 43220 23264
rect 43168 22636 43220 22642
rect 43168 22578 43220 22584
rect 43180 22234 43208 22578
rect 43168 22228 43220 22234
rect 43168 22170 43220 22176
rect 42984 22092 43036 22098
rect 42984 22034 43036 22040
rect 43272 21554 43300 23666
rect 43456 23474 43484 23734
rect 43364 23446 43484 23474
rect 43364 23322 43392 23446
rect 43352 23316 43404 23322
rect 43352 23258 43404 23264
rect 43444 23112 43496 23118
rect 43548 23100 43576 24550
rect 44008 24410 44036 24822
rect 44272 24676 44324 24682
rect 44272 24618 44324 24624
rect 44284 24585 44312 24618
rect 44652 24614 44680 25298
rect 44836 24857 44864 27814
rect 44822 24848 44878 24857
rect 44822 24783 44878 24792
rect 44640 24608 44692 24614
rect 44270 24576 44326 24585
rect 44640 24550 44692 24556
rect 44732 24608 44784 24614
rect 44732 24550 44784 24556
rect 44270 24511 44326 24520
rect 43996 24404 44048 24410
rect 43996 24346 44048 24352
rect 43628 24336 43680 24342
rect 43628 24278 43680 24284
rect 43640 23594 43668 24278
rect 43812 24200 43864 24206
rect 43812 24142 43864 24148
rect 43628 23588 43680 23594
rect 43628 23530 43680 23536
rect 43628 23248 43680 23254
rect 43628 23190 43680 23196
rect 43496 23072 43576 23100
rect 43444 23054 43496 23060
rect 43456 22778 43484 23054
rect 43444 22772 43496 22778
rect 43444 22714 43496 22720
rect 43640 22438 43668 23190
rect 43824 22624 43852 24142
rect 44180 23520 44232 23526
rect 44652 23497 44680 24550
rect 44180 23462 44232 23468
rect 44638 23488 44694 23497
rect 44192 22642 44220 23462
rect 44638 23423 44694 23432
rect 43732 22596 43852 22624
rect 44180 22636 44232 22642
rect 43628 22432 43680 22438
rect 43628 22374 43680 22380
rect 43352 22092 43404 22098
rect 43352 22034 43404 22040
rect 43364 21690 43392 22034
rect 43352 21684 43404 21690
rect 43352 21626 43404 21632
rect 43442 21584 43498 21593
rect 43260 21548 43312 21554
rect 43442 21519 43498 21528
rect 43260 21490 43312 21496
rect 42616 20936 42668 20942
rect 42616 20878 42668 20884
rect 42628 20602 42656 20878
rect 42616 20596 42668 20602
rect 42616 20538 42668 20544
rect 42800 20528 42852 20534
rect 42800 20470 42852 20476
rect 42812 18970 42840 20470
rect 42892 19848 42944 19854
rect 42892 19790 42944 19796
rect 42800 18964 42852 18970
rect 42800 18906 42852 18912
rect 42800 18284 42852 18290
rect 42904 18272 42932 19790
rect 43272 18766 43300 21490
rect 43456 19174 43484 21519
rect 43536 21072 43588 21078
rect 43536 21014 43588 21020
rect 43548 20602 43576 21014
rect 43536 20596 43588 20602
rect 43536 20538 43588 20544
rect 43548 20330 43576 20538
rect 43732 20516 43760 22596
rect 44180 22578 44232 22584
rect 43812 22500 43864 22506
rect 43812 22442 43864 22448
rect 43824 22030 43852 22442
rect 44744 22409 44772 24550
rect 44730 22400 44786 22409
rect 44730 22335 44786 22344
rect 44836 22216 44864 24783
rect 44916 24268 44968 24274
rect 44916 24210 44968 24216
rect 44928 23866 44956 24210
rect 44916 23860 44968 23866
rect 44916 23802 44968 23808
rect 45468 23860 45520 23866
rect 45468 23802 45520 23808
rect 44916 23180 44968 23186
rect 44916 23122 44968 23128
rect 44928 22438 44956 23122
rect 44916 22432 44968 22438
rect 44916 22374 44968 22380
rect 44744 22188 44864 22216
rect 43812 22024 43864 22030
rect 43812 21966 43864 21972
rect 43996 22024 44048 22030
rect 43996 21966 44048 21972
rect 43824 21078 43852 21966
rect 43904 21888 43956 21894
rect 43904 21830 43956 21836
rect 43916 21554 43944 21830
rect 43904 21548 43956 21554
rect 43904 21490 43956 21496
rect 44008 21418 44036 21966
rect 44548 21888 44600 21894
rect 44548 21830 44600 21836
rect 43996 21412 44048 21418
rect 43996 21354 44048 21360
rect 44008 21146 44036 21354
rect 43996 21140 44048 21146
rect 43996 21082 44048 21088
rect 43812 21072 43864 21078
rect 43812 21014 43864 21020
rect 43732 20488 43852 20516
rect 43536 20324 43588 20330
rect 43536 20266 43588 20272
rect 43548 19972 43576 20266
rect 43720 20052 43772 20058
rect 43720 19994 43772 20000
rect 43628 19984 43680 19990
rect 43548 19944 43628 19972
rect 43548 19514 43576 19944
rect 43628 19926 43680 19932
rect 43732 19514 43760 19994
rect 43824 19854 43852 20488
rect 44456 20460 44508 20466
rect 44456 20402 44508 20408
rect 44468 19990 44496 20402
rect 44456 19984 44508 19990
rect 44456 19926 44508 19932
rect 43812 19848 43864 19854
rect 43812 19790 43864 19796
rect 44560 19718 44588 21830
rect 44744 21593 44772 22188
rect 44824 22092 44876 22098
rect 44824 22034 44876 22040
rect 44730 21584 44786 21593
rect 44730 21519 44786 21528
rect 44836 21350 44864 22034
rect 44824 21344 44876 21350
rect 44928 21321 44956 22374
rect 45480 21457 45508 23802
rect 45466 21448 45522 21457
rect 45466 21383 45522 21392
rect 44824 21286 44876 21292
rect 44914 21312 44970 21321
rect 44548 19712 44600 19718
rect 44548 19654 44600 19660
rect 43536 19508 43588 19514
rect 43536 19450 43588 19456
rect 43720 19508 43772 19514
rect 43720 19450 43772 19456
rect 43444 19168 43496 19174
rect 43444 19110 43496 19116
rect 43996 19168 44048 19174
rect 43996 19110 44048 19116
rect 43536 18896 43588 18902
rect 43536 18838 43588 18844
rect 43260 18760 43312 18766
rect 43260 18702 43312 18708
rect 43272 18358 43300 18702
rect 43548 18426 43576 18838
rect 43720 18760 43772 18766
rect 43720 18702 43772 18708
rect 43536 18420 43588 18426
rect 43536 18362 43588 18368
rect 43260 18352 43312 18358
rect 43260 18294 43312 18300
rect 43732 18290 43760 18702
rect 42852 18244 42932 18272
rect 43720 18284 43772 18290
rect 42800 18226 42852 18232
rect 43720 18226 43772 18232
rect 43536 17128 43588 17134
rect 43536 17070 43588 17076
rect 43548 16969 43576 17070
rect 42522 16960 42578 16969
rect 42522 16895 42578 16904
rect 43534 16960 43590 16969
rect 43534 16895 43590 16904
rect 43168 16720 43220 16726
rect 43168 16662 43220 16668
rect 43628 16720 43680 16726
rect 43628 16662 43680 16668
rect 42248 16516 42300 16522
rect 42248 16458 42300 16464
rect 42156 16176 42208 16182
rect 42156 16118 42208 16124
rect 42064 16108 42116 16114
rect 42064 16050 42116 16056
rect 39672 15972 39724 15978
rect 39672 15914 39724 15920
rect 40316 15972 40368 15978
rect 40316 15914 40368 15920
rect 41052 15972 41104 15978
rect 41052 15914 41104 15920
rect 39488 15564 39540 15570
rect 39488 15506 39540 15512
rect 39120 14952 39172 14958
rect 39120 14894 39172 14900
rect 39132 14618 39160 14894
rect 39580 14884 39632 14890
rect 39580 14826 39632 14832
rect 39120 14612 39172 14618
rect 39120 14554 39172 14560
rect 39132 12782 39160 14554
rect 39592 14414 39620 14826
rect 39684 14550 39712 15914
rect 40040 15360 40092 15366
rect 40040 15302 40092 15308
rect 40052 14958 40080 15302
rect 40328 15162 40356 15914
rect 41064 15638 41092 15914
rect 42076 15706 42104 16050
rect 42064 15700 42116 15706
rect 42064 15642 42116 15648
rect 41052 15632 41104 15638
rect 41052 15574 41104 15580
rect 40960 15496 41012 15502
rect 40960 15438 41012 15444
rect 40592 15360 40644 15366
rect 40592 15302 40644 15308
rect 40316 15156 40368 15162
rect 40316 15098 40368 15104
rect 40040 14952 40092 14958
rect 40040 14894 40092 14900
rect 40328 14890 40356 15098
rect 40604 15026 40632 15302
rect 40592 15020 40644 15026
rect 40592 14962 40644 14968
rect 40316 14884 40368 14890
rect 40316 14826 40368 14832
rect 39672 14544 39724 14550
rect 39672 14486 39724 14492
rect 39580 14408 39632 14414
rect 39580 14350 39632 14356
rect 39212 14272 39264 14278
rect 39212 14214 39264 14220
rect 39224 14074 39252 14214
rect 39592 14074 39620 14350
rect 39212 14068 39264 14074
rect 39212 14010 39264 14016
rect 39580 14068 39632 14074
rect 39580 14010 39632 14016
rect 39684 14006 39712 14486
rect 40972 14482 41000 15438
rect 41696 14884 41748 14890
rect 41696 14826 41748 14832
rect 41420 14544 41472 14550
rect 41420 14486 41472 14492
rect 40960 14476 41012 14482
rect 40960 14418 41012 14424
rect 40500 14272 40552 14278
rect 40500 14214 40552 14220
rect 41328 14272 41380 14278
rect 41328 14214 41380 14220
rect 40512 14006 40540 14214
rect 41340 14074 41368 14214
rect 41328 14068 41380 14074
rect 41328 14010 41380 14016
rect 41432 14006 41460 14486
rect 39672 14000 39724 14006
rect 39672 13942 39724 13948
rect 40500 14000 40552 14006
rect 40500 13942 40552 13948
rect 41420 14000 41472 14006
rect 41420 13942 41472 13948
rect 39684 13462 39712 13942
rect 40960 13932 41012 13938
rect 40960 13874 41012 13880
rect 40972 13705 41000 13874
rect 41604 13796 41656 13802
rect 41604 13738 41656 13744
rect 40958 13696 41014 13705
rect 40958 13631 41014 13640
rect 41616 13462 41644 13738
rect 39672 13456 39724 13462
rect 39672 13398 39724 13404
rect 41604 13456 41656 13462
rect 41604 13398 41656 13404
rect 39580 13320 39632 13326
rect 39580 13262 39632 13268
rect 39592 12850 39620 13262
rect 39684 12986 39712 13398
rect 40868 13252 40920 13258
rect 40868 13194 40920 13200
rect 39672 12980 39724 12986
rect 39672 12922 39724 12928
rect 39580 12844 39632 12850
rect 39580 12786 39632 12792
rect 39120 12776 39172 12782
rect 39120 12718 39172 12724
rect 39132 12442 39160 12718
rect 39120 12436 39172 12442
rect 39120 12378 39172 12384
rect 39132 11694 39160 12378
rect 39684 12374 39712 12922
rect 40880 12714 40908 13194
rect 40960 13184 41012 13190
rect 40960 13126 41012 13132
rect 40972 12714 41000 13126
rect 41616 12986 41644 13398
rect 41708 13258 41736 14826
rect 42168 14006 42196 16118
rect 42260 14550 42288 16458
rect 42616 15904 42668 15910
rect 42616 15846 42668 15852
rect 42524 14952 42576 14958
rect 42524 14894 42576 14900
rect 42536 14793 42564 14894
rect 42522 14784 42578 14793
rect 42522 14719 42578 14728
rect 42628 14618 42656 15846
rect 43180 15706 43208 16662
rect 43640 15910 43668 16662
rect 43628 15904 43680 15910
rect 43628 15846 43680 15852
rect 43168 15700 43220 15706
rect 43168 15642 43220 15648
rect 43640 15638 43668 15846
rect 43628 15632 43680 15638
rect 43628 15574 43680 15580
rect 43640 15162 43668 15574
rect 43720 15428 43772 15434
rect 43720 15370 43772 15376
rect 43628 15156 43680 15162
rect 43628 15098 43680 15104
rect 43640 14890 43668 15098
rect 43536 14884 43588 14890
rect 43536 14826 43588 14832
rect 43628 14884 43680 14890
rect 43628 14826 43680 14832
rect 43548 14618 43576 14826
rect 42616 14612 42668 14618
rect 42616 14554 42668 14560
rect 43536 14612 43588 14618
rect 43536 14554 43588 14560
rect 42248 14544 42300 14550
rect 42248 14486 42300 14492
rect 42156 14000 42208 14006
rect 42156 13942 42208 13948
rect 41696 13252 41748 13258
rect 41696 13194 41748 13200
rect 41604 12980 41656 12986
rect 41604 12922 41656 12928
rect 41512 12912 41564 12918
rect 41512 12854 41564 12860
rect 40868 12708 40920 12714
rect 40868 12650 40920 12656
rect 40960 12708 41012 12714
rect 40960 12650 41012 12656
rect 40880 12374 40908 12650
rect 39672 12368 39724 12374
rect 39672 12310 39724 12316
rect 39948 12368 40000 12374
rect 39948 12310 40000 12316
rect 40868 12368 40920 12374
rect 40868 12310 40920 12316
rect 39672 12232 39724 12238
rect 39672 12174 39724 12180
rect 39684 11762 39712 12174
rect 39960 11898 39988 12310
rect 41524 12238 41552 12854
rect 41880 12708 41932 12714
rect 41880 12650 41932 12656
rect 41892 12238 41920 12650
rect 40776 12232 40828 12238
rect 40776 12174 40828 12180
rect 41512 12232 41564 12238
rect 41512 12174 41564 12180
rect 41880 12232 41932 12238
rect 41880 12174 41932 12180
rect 40788 11898 40816 12174
rect 41328 12164 41380 12170
rect 41328 12106 41380 12112
rect 39948 11892 40000 11898
rect 39948 11834 40000 11840
rect 40776 11892 40828 11898
rect 40776 11834 40828 11840
rect 39672 11756 39724 11762
rect 39672 11698 39724 11704
rect 39120 11688 39172 11694
rect 39120 11630 39172 11636
rect 39132 11354 39160 11630
rect 39120 11348 39172 11354
rect 39120 11290 39172 11296
rect 38660 11008 38712 11014
rect 38660 10950 38712 10956
rect 39028 11008 39080 11014
rect 39028 10950 39080 10956
rect 38672 10810 38700 10950
rect 38660 10804 38712 10810
rect 38660 10746 38712 10752
rect 38672 10606 38700 10746
rect 39132 10606 39160 11290
rect 39304 11212 39356 11218
rect 39304 11154 39356 11160
rect 39316 11121 39344 11154
rect 39302 11112 39358 11121
rect 39302 11047 39358 11056
rect 39316 10810 39344 11047
rect 39304 10804 39356 10810
rect 39304 10746 39356 10752
rect 39960 10742 39988 11834
rect 41340 11762 41368 12106
rect 41892 11830 41920 12174
rect 42168 12170 42196 13942
rect 42260 12850 42288 14486
rect 42628 13977 42656 14554
rect 43536 14476 43588 14482
rect 43536 14418 43588 14424
rect 42984 14272 43036 14278
rect 42984 14214 43036 14220
rect 42996 14074 43024 14214
rect 42984 14068 43036 14074
rect 42984 14010 43036 14016
rect 42614 13968 42670 13977
rect 42614 13903 42670 13912
rect 43548 13734 43576 14418
rect 42616 13728 42668 13734
rect 42616 13670 42668 13676
rect 43536 13728 43588 13734
rect 43536 13670 43588 13676
rect 42628 13326 42656 13670
rect 43258 13560 43314 13569
rect 43258 13495 43314 13504
rect 43272 13394 43300 13495
rect 43548 13433 43576 13670
rect 43534 13424 43590 13433
rect 43260 13388 43312 13394
rect 43534 13359 43590 13368
rect 43260 13330 43312 13336
rect 42616 13320 42668 13326
rect 42616 13262 42668 13268
rect 42628 12986 42656 13262
rect 43168 13184 43220 13190
rect 43168 13126 43220 13132
rect 42616 12980 42668 12986
rect 42616 12922 42668 12928
rect 43180 12850 43208 13126
rect 43272 12986 43300 13330
rect 43260 12980 43312 12986
rect 43260 12922 43312 12928
rect 42248 12844 42300 12850
rect 42248 12786 42300 12792
rect 43168 12844 43220 12850
rect 43168 12786 43220 12792
rect 43180 12442 43208 12786
rect 43536 12640 43588 12646
rect 43536 12582 43588 12588
rect 43168 12436 43220 12442
rect 43168 12378 43220 12384
rect 43548 12374 43576 12582
rect 42248 12368 42300 12374
rect 42248 12310 42300 12316
rect 43536 12368 43588 12374
rect 43536 12310 43588 12316
rect 42156 12164 42208 12170
rect 42156 12106 42208 12112
rect 42260 11898 42288 12310
rect 43352 12164 43404 12170
rect 43352 12106 43404 12112
rect 42248 11892 42300 11898
rect 42248 11834 42300 11840
rect 43076 11892 43128 11898
rect 43076 11834 43128 11840
rect 41880 11824 41932 11830
rect 41880 11766 41932 11772
rect 41328 11756 41380 11762
rect 41328 11698 41380 11704
rect 41696 11756 41748 11762
rect 41696 11698 41748 11704
rect 41512 11620 41564 11626
rect 41512 11562 41564 11568
rect 41420 11280 41472 11286
rect 41420 11222 41472 11228
rect 40040 11144 40092 11150
rect 40040 11086 40092 11092
rect 41328 11144 41380 11150
rect 41328 11086 41380 11092
rect 39948 10736 40000 10742
rect 39948 10678 40000 10684
rect 38660 10600 38712 10606
rect 38660 10542 38712 10548
rect 39120 10600 39172 10606
rect 39120 10542 39172 10548
rect 39132 10266 39160 10542
rect 39580 10532 39632 10538
rect 39580 10474 39632 10480
rect 39120 10260 39172 10266
rect 39120 10202 39172 10208
rect 38568 9648 38620 9654
rect 38568 9590 38620 9596
rect 39132 9518 39160 10202
rect 39592 10130 39620 10474
rect 39960 10198 39988 10678
rect 40052 10674 40080 11086
rect 40040 10668 40092 10674
rect 40040 10610 40092 10616
rect 40498 10568 40554 10577
rect 40498 10503 40554 10512
rect 40512 10470 40540 10503
rect 40500 10464 40552 10470
rect 40500 10406 40552 10412
rect 41340 10198 41368 11086
rect 41432 10810 41460 11222
rect 41420 10804 41472 10810
rect 41420 10746 41472 10752
rect 41432 10266 41460 10746
rect 41420 10260 41472 10266
rect 41420 10202 41472 10208
rect 39948 10192 40000 10198
rect 39948 10134 40000 10140
rect 41328 10192 41380 10198
rect 41328 10134 41380 10140
rect 39580 10124 39632 10130
rect 39580 10066 39632 10072
rect 39960 9722 39988 10134
rect 40132 10124 40184 10130
rect 40132 10066 40184 10072
rect 39948 9716 40000 9722
rect 39948 9658 40000 9664
rect 39120 9512 39172 9518
rect 39120 9454 39172 9460
rect 39132 9178 39160 9454
rect 39960 9450 39988 9658
rect 39948 9444 40000 9450
rect 39948 9386 40000 9392
rect 37096 9172 37148 9178
rect 37096 9114 37148 9120
rect 39120 9172 39172 9178
rect 39120 9114 39172 9120
rect 39960 9042 39988 9386
rect 40144 9178 40172 10066
rect 41524 9722 41552 11562
rect 41512 9716 41564 9722
rect 41512 9658 41564 9664
rect 40500 9512 40552 9518
rect 40500 9454 40552 9460
rect 40512 9178 40540 9454
rect 40132 9172 40184 9178
rect 40132 9114 40184 9120
rect 40500 9172 40552 9178
rect 40500 9114 40552 9120
rect 36544 9036 36596 9042
rect 36544 8978 36596 8984
rect 39948 9036 40000 9042
rect 39948 8978 40000 8984
rect 36556 8634 36584 8978
rect 36544 8628 36596 8634
rect 36544 8570 36596 8576
rect 35716 8492 35768 8498
rect 35716 8434 35768 8440
rect 35072 8424 35124 8430
rect 35072 8366 35124 8372
rect 35084 8090 35112 8366
rect 34704 8084 34756 8090
rect 34704 8026 34756 8032
rect 35072 8084 35124 8090
rect 35072 8026 35124 8032
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 33414 7304 33470 7313
rect 33414 7239 33470 7248
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 36174 3904 36230 3913
rect 36174 3839 36230 3848
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 24950 54 25084 82
rect 28540 128 28592 134
rect 28540 70 28592 76
rect 30470 128 30526 480
rect 30470 76 30472 128
rect 30524 76 30526 128
rect 24950 0 25006 54
rect 30470 0 30526 76
rect 36082 82 36138 480
rect 36188 82 36216 3839
rect 36082 54 36216 82
rect 41602 82 41658 480
rect 41708 82 41736 11698
rect 41892 11082 41920 11766
rect 43088 11762 43116 11834
rect 43364 11762 43392 12106
rect 43076 11756 43128 11762
rect 43076 11698 43128 11704
rect 43352 11756 43404 11762
rect 43352 11698 43404 11704
rect 42892 11552 42944 11558
rect 42892 11494 42944 11500
rect 41880 11076 41932 11082
rect 41880 11018 41932 11024
rect 41892 10606 41920 11018
rect 42904 10810 42932 11494
rect 43088 11354 43116 11698
rect 43548 11558 43576 12310
rect 43536 11552 43588 11558
rect 43536 11494 43588 11500
rect 43076 11348 43128 11354
rect 43076 11290 43128 11296
rect 43732 11150 43760 15370
rect 43904 13932 43956 13938
rect 43904 13874 43956 13880
rect 43916 13841 43944 13874
rect 43902 13832 43958 13841
rect 43902 13767 43958 13776
rect 44008 12782 44036 19110
rect 44836 19009 44864 21286
rect 44914 21247 44970 21256
rect 44822 19000 44878 19009
rect 44822 18935 44878 18944
rect 44088 16992 44140 16998
rect 44088 16934 44140 16940
rect 44100 16114 44128 16934
rect 44088 16108 44140 16114
rect 44088 16050 44140 16056
rect 44100 15706 44128 16050
rect 44088 15700 44140 15706
rect 44088 15642 44140 15648
rect 44824 15564 44876 15570
rect 44928 15552 44956 21247
rect 45468 21004 45520 21010
rect 45468 20946 45520 20952
rect 45480 20466 45508 20946
rect 45468 20460 45520 20466
rect 45468 20402 45520 20408
rect 45480 20369 45508 20402
rect 45466 20360 45522 20369
rect 45466 20295 45522 20304
rect 45008 20256 45060 20262
rect 45008 20198 45060 20204
rect 45020 20058 45048 20198
rect 45008 20052 45060 20058
rect 45008 19994 45060 20000
rect 45008 19916 45060 19922
rect 45008 19858 45060 19864
rect 45020 19174 45048 19858
rect 45008 19168 45060 19174
rect 45008 19110 45060 19116
rect 45008 16652 45060 16658
rect 45008 16594 45060 16600
rect 45020 15910 45048 16594
rect 45008 15904 45060 15910
rect 45008 15846 45060 15852
rect 44876 15524 44956 15552
rect 44824 15506 44876 15512
rect 44456 15496 44508 15502
rect 44456 15438 44508 15444
rect 44468 15162 44496 15438
rect 44730 15192 44786 15201
rect 44456 15156 44508 15162
rect 44730 15127 44786 15136
rect 44456 15098 44508 15104
rect 44744 15026 44772 15127
rect 44732 15020 44784 15026
rect 44732 14962 44784 14968
rect 44836 14890 44864 15506
rect 45020 15473 45048 15846
rect 45006 15464 45062 15473
rect 45006 15399 45062 15408
rect 49514 14920 49570 14929
rect 44180 14884 44232 14890
rect 44180 14826 44232 14832
rect 44824 14884 44876 14890
rect 44824 14826 44876 14832
rect 46940 14884 46992 14890
rect 49514 14855 49570 14864
rect 46940 14826 46992 14832
rect 44192 13258 44220 14826
rect 44916 14816 44968 14822
rect 44916 14758 44968 14764
rect 44928 14618 44956 14758
rect 44916 14612 44968 14618
rect 44916 14554 44968 14560
rect 44180 13252 44232 13258
rect 44180 13194 44232 13200
rect 43996 12776 44048 12782
rect 43996 12718 44048 12724
rect 44192 12374 44220 13194
rect 44456 12640 44508 12646
rect 44456 12582 44508 12588
rect 44180 12368 44232 12374
rect 44180 12310 44232 12316
rect 44468 12238 44496 12582
rect 44456 12232 44508 12238
rect 44456 12174 44508 12180
rect 44468 11898 44496 12174
rect 44456 11892 44508 11898
rect 44456 11834 44508 11840
rect 44180 11552 44232 11558
rect 44180 11494 44232 11500
rect 44192 11286 44220 11494
rect 44180 11280 44232 11286
rect 44180 11222 44232 11228
rect 43444 11144 43496 11150
rect 43444 11086 43496 11092
rect 43720 11144 43772 11150
rect 43720 11086 43772 11092
rect 43456 10810 43484 11086
rect 44192 10810 44220 11222
rect 42892 10804 42944 10810
rect 42892 10746 42944 10752
rect 43444 10804 43496 10810
rect 43444 10746 43496 10752
rect 44180 10804 44232 10810
rect 44180 10746 44232 10752
rect 41972 10668 42024 10674
rect 41972 10610 42024 10616
rect 41880 10600 41932 10606
rect 41880 10542 41932 10548
rect 41984 10266 42012 10610
rect 41972 10260 42024 10266
rect 41972 10202 42024 10208
rect 41602 54 41736 82
rect 46952 82 46980 14826
rect 49528 13977 49556 14855
rect 49514 13968 49570 13977
rect 49514 13903 49570 13912
rect 47122 82 47178 480
rect 46952 54 47178 82
rect 36082 0 36138 54
rect 41602 0 41658 54
rect 47122 0 47178 54
<< via2 >>
rect 110 46416 166 46472
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 110 39752 166 39808
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 2778 39344 2834 39400
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 2594 38664 2650 38720
rect 110 24928 166 24984
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 12990 39480 13046 39536
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 3330 31592 3386 31648
rect 2594 18808 2650 18864
rect 1950 18400 2006 18456
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 3974 28908 3976 28928
rect 3976 28908 4028 28928
rect 4028 28908 4030 28928
rect 3974 28872 4030 28908
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4526 28872 4582 28928
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 23110 43852 23166 43888
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 23110 43832 23112 43852
rect 23112 43832 23164 43852
rect 23164 43832 23166 43852
rect 30286 43832 30342 43888
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 17314 39752 17370 39808
rect 4986 30096 5042 30152
rect 5354 29552 5410 29608
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 3422 19896 3478 19952
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4894 23568 4950 23624
rect 5998 23568 6054 23624
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 8390 30232 8446 30288
rect 9862 29028 9918 29064
rect 9862 29008 9864 29028
rect 9864 29008 9916 29028
rect 9916 29008 9918 29028
rect 9678 28872 9734 28928
rect 8942 23568 8998 23624
rect 8758 22480 8814 22536
rect 7562 20440 7618 20496
rect 7562 18944 7618 19000
rect 8850 18400 8906 18456
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 9954 23024 10010 23080
rect 12070 31728 12126 31784
rect 14462 30232 14518 30288
rect 14554 30096 14610 30152
rect 1490 11192 1546 11248
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 13358 21936 13414 21992
rect 14370 19352 14426 19408
rect 14370 17040 14426 17096
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 15842 37712 15898 37768
rect 17774 38412 17830 38448
rect 17774 38392 17776 38412
rect 17776 38392 17828 38412
rect 17828 38392 17830 38412
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 19062 39344 19118 39400
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 21178 38800 21234 38856
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 17222 35148 17278 35184
rect 17222 35128 17224 35148
rect 17224 35128 17276 35148
rect 17276 35128 17278 35148
rect 17222 32952 17278 33008
rect 15474 31728 15530 31784
rect 15474 29008 15530 29064
rect 16946 29552 17002 29608
rect 16578 28872 16634 28928
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 22190 38936 22246 38992
rect 21178 34584 21234 34640
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 18970 28056 19026 28112
rect 17498 23432 17554 23488
rect 16946 20440 17002 20496
rect 17222 18944 17278 19000
rect 16946 18400 17002 18456
rect 18050 17312 18106 17368
rect 14830 10512 14886 10568
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 1398 4120 1454 4176
rect 3054 4120 3110 4176
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 13174 4120 13230 4176
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 20902 33396 20904 33416
rect 20904 33396 20956 33416
rect 20956 33396 20958 33416
rect 20902 33360 20958 33396
rect 21086 28464 21142 28520
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19798 24792 19854 24848
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 18970 23432 19026 23488
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 23110 41112 23166 41168
rect 22650 36624 22706 36680
rect 22466 34584 22522 34640
rect 23846 38936 23902 38992
rect 24674 36624 24730 36680
rect 25778 38392 25834 38448
rect 23386 32952 23442 33008
rect 22374 29552 22430 29608
rect 22006 28736 22062 28792
rect 21730 27784 21786 27840
rect 19246 22636 19302 22672
rect 19246 22616 19248 22636
rect 19248 22616 19300 22636
rect 19300 22616 19302 22636
rect 19430 22480 19486 22536
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 20166 22344 20222 22400
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 18510 15952 18566 16008
rect 15842 10104 15898 10160
rect 15106 7248 15162 7304
rect 18602 12144 18658 12200
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 23478 29552 23534 29608
rect 21822 21936 21878 21992
rect 23110 23160 23166 23216
rect 23754 29688 23810 29744
rect 30470 43016 30526 43072
rect 25594 33768 25650 33824
rect 25502 33088 25558 33144
rect 26146 34584 26202 34640
rect 25778 33360 25834 33416
rect 25226 28600 25282 28656
rect 23478 24792 23534 24848
rect 23938 26560 23994 26616
rect 25042 28056 25098 28112
rect 24674 23024 24730 23080
rect 26146 33088 26202 33144
rect 26054 32408 26110 32464
rect 23846 22208 23902 22264
rect 22650 19896 22706 19952
rect 27802 32952 27858 33008
rect 26606 28736 26662 28792
rect 26514 28600 26570 28656
rect 27158 28328 27214 28384
rect 26606 24656 26662 24712
rect 24306 19352 24362 19408
rect 21730 18128 21786 18184
rect 21454 17856 21510 17912
rect 22006 17484 22008 17504
rect 22008 17484 22060 17504
rect 22060 17484 22062 17504
rect 22006 17448 22062 17484
rect 22834 17176 22890 17232
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 22926 15000 22982 15056
rect 23110 17856 23166 17912
rect 21086 14184 21142 14240
rect 24490 18808 24546 18864
rect 24306 17312 24362 17368
rect 23478 17040 23534 17096
rect 23202 13640 23258 13696
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19246 8880 19302 8936
rect 23110 12280 23166 12336
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 23202 9560 23258 9616
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 23478 12144 23534 12200
rect 24950 13504 25006 13560
rect 23754 9560 23810 9616
rect 23294 4120 23350 4176
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 28078 36488 28134 36544
rect 28262 34040 28318 34096
rect 27986 29552 28042 29608
rect 27986 28464 28042 28520
rect 27342 20984 27398 21040
rect 26882 18808 26938 18864
rect 26330 10104 26386 10160
rect 27434 18808 27490 18864
rect 30378 38392 30434 38448
rect 29642 36624 29698 36680
rect 29182 35128 29238 35184
rect 28906 33904 28962 33960
rect 29550 35028 29552 35048
rect 29552 35028 29604 35048
rect 29604 35028 29606 35048
rect 29550 34992 29606 35028
rect 31850 42744 31906 42800
rect 32862 42744 32918 42800
rect 31114 39480 31170 39536
rect 32218 38800 32274 38856
rect 32218 36080 32274 36136
rect 32862 41112 32918 41168
rect 32770 37168 32826 37224
rect 30746 33904 30802 33960
rect 30378 32952 30434 33008
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 32586 33088 32642 33144
rect 30562 28872 30618 28928
rect 29734 28328 29790 28384
rect 28078 19760 28134 19816
rect 28170 17448 28226 17504
rect 27618 15272 27674 15328
rect 27802 10784 27858 10840
rect 31206 27784 31262 27840
rect 32034 26560 32090 26616
rect 33230 38664 33286 38720
rect 36174 43016 36230 43072
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 33782 36760 33838 36816
rect 33506 36080 33562 36136
rect 33690 34584 33746 34640
rect 33322 33904 33378 33960
rect 33230 33768 33286 33824
rect 31206 23568 31262 23624
rect 30746 23160 30802 23216
rect 28170 15680 28226 15736
rect 28170 3848 28226 3904
rect 29182 16768 29238 16824
rect 28630 15952 28686 16008
rect 30010 20032 30066 20088
rect 30102 18944 30158 19000
rect 30378 22208 30434 22264
rect 30562 20984 30618 21040
rect 30286 17856 30342 17912
rect 30746 18128 30802 18184
rect 30378 15952 30434 16008
rect 30930 23160 30986 23216
rect 28814 13912 28870 13968
rect 28814 12688 28870 12744
rect 32954 27648 33010 27704
rect 32402 23568 32458 23624
rect 31390 19352 31446 19408
rect 31390 19116 31392 19136
rect 31392 19116 31444 19136
rect 31444 19116 31446 19136
rect 31390 19080 31446 19116
rect 31482 18164 31484 18184
rect 31484 18164 31536 18184
rect 31536 18164 31538 18184
rect 31482 18128 31538 18164
rect 31298 13640 31354 13696
rect 31206 13504 31262 13560
rect 31942 20440 31998 20496
rect 32034 19080 32090 19136
rect 32402 19488 32458 19544
rect 32678 17176 32734 17232
rect 30194 10648 30250 10704
rect 34058 32408 34114 32464
rect 33874 29688 33930 29744
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 34518 34992 34574 35048
rect 34426 34060 34482 34096
rect 34426 34040 34428 34060
rect 34428 34040 34480 34060
rect 34480 34040 34482 34060
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 35898 42744 35954 42800
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 35898 37304 35954 37360
rect 35714 36488 35770 36544
rect 41142 44240 41198 44296
rect 37002 38664 37058 38720
rect 36358 38392 36414 38448
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34610 28620 34666 28656
rect 34610 28600 34612 28620
rect 34612 28600 34664 28620
rect 34664 28600 34666 28620
rect 34794 28328 34850 28384
rect 33598 24656 33654 24712
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 37830 37712 37886 37768
rect 40406 37168 40462 37224
rect 38382 34992 38438 35048
rect 36082 28872 36138 28928
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 33598 21392 33654 21448
rect 33046 19488 33102 19544
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 35162 21256 35218 21312
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 35162 20304 35218 20360
rect 33230 19352 33286 19408
rect 32954 14728 33010 14784
rect 33598 18808 33654 18864
rect 37738 28056 37794 28112
rect 38106 33088 38162 33144
rect 35990 22616 36046 22672
rect 36726 21528 36782 21584
rect 39854 34720 39910 34776
rect 38934 32272 38990 32328
rect 38934 28736 38990 28792
rect 42062 36760 42118 36816
rect 41970 33088 42026 33144
rect 42614 37168 42670 37224
rect 42706 36080 42762 36136
rect 43350 34720 43406 34776
rect 39118 28464 39174 28520
rect 39026 27648 39082 27704
rect 39762 29552 39818 29608
rect 37830 24384 37886 24440
rect 39210 27512 39266 27568
rect 35898 20168 35954 20224
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 33506 18264 33562 18320
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 33046 13776 33102 13832
rect 33874 13776 33930 13832
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 35070 15408 35126 15464
rect 34702 15272 34758 15328
rect 34610 15036 34612 15056
rect 34612 15036 34664 15056
rect 34664 15036 34666 15056
rect 34610 15000 34666 15036
rect 33782 12280 33838 12336
rect 33230 11056 33286 11112
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34150 12688 34206 12744
rect 35990 16904 36046 16960
rect 35898 13776 35954 13832
rect 38106 20440 38162 20496
rect 37738 19760 37794 19816
rect 37002 18264 37058 18320
rect 36266 15952 36322 16008
rect 36266 15136 36322 15192
rect 36082 13912 36138 13968
rect 34518 10784 34574 10840
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 37370 15680 37426 15736
rect 37554 13776 37610 13832
rect 37002 13640 37058 13696
rect 38014 13640 38070 13696
rect 37830 13388 37886 13424
rect 37830 13368 37832 13388
rect 37832 13368 37884 13388
rect 37884 13368 37886 13388
rect 36082 10648 36138 10704
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 42430 32272 42486 32328
rect 41694 27648 41750 27704
rect 40958 25608 41014 25664
rect 40958 24656 41014 24712
rect 40866 24520 40922 24576
rect 38658 18164 38660 18184
rect 38660 18164 38712 18184
rect 38712 18164 38714 18184
rect 38658 18128 38714 18164
rect 38290 13504 38346 13560
rect 38106 11056 38162 11112
rect 39302 16768 39358 16824
rect 43810 37304 43866 37360
rect 43810 34720 43866 34776
rect 44546 27512 44602 27568
rect 44638 25608 44694 25664
rect 42982 24384 43038 24440
rect 44822 24792 44878 24848
rect 44270 24520 44326 24576
rect 44638 23432 44694 23488
rect 43442 21528 43498 21584
rect 44730 22344 44786 22400
rect 44730 21528 44786 21584
rect 45466 21392 45522 21448
rect 42522 16904 42578 16960
rect 43534 16904 43590 16960
rect 40958 13640 41014 13696
rect 42522 14728 42578 14784
rect 39302 11056 39358 11112
rect 42614 13912 42670 13968
rect 43258 13504 43314 13560
rect 43534 13368 43590 13424
rect 40498 10512 40554 10568
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 33414 7248 33470 7304
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 36174 3848 36230 3904
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 43902 13776 43958 13832
rect 44914 21256 44970 21312
rect 44822 18944 44878 19000
rect 45466 20304 45522 20360
rect 44730 15136 44786 15192
rect 45006 15408 45062 15464
rect 49514 14864 49570 14920
rect 49514 13912 49570 13968
<< metal3 >>
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 0 46472 480 46504
rect 0 46416 110 46472
rect 166 46416 480 46472
rect 0 46384 480 46416
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 19568 45184 19888 45185
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 49520 44888 50000 45008
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 41137 44298 41203 44301
rect 49558 44298 49618 44888
rect 41137 44296 49618 44298
rect 41137 44240 41142 44296
rect 41198 44240 49618 44296
rect 41137 44238 49618 44240
rect 41137 44235 41203 44238
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 23105 43890 23171 43893
rect 30281 43890 30347 43893
rect 23105 43888 30347 43890
rect 23105 43832 23110 43888
rect 23166 43832 30286 43888
rect 30342 43832 30347 43888
rect 23105 43830 30347 43832
rect 23105 43827 23171 43830
rect 30281 43827 30347 43830
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 30465 43074 30531 43077
rect 36169 43074 36235 43077
rect 30465 43072 36235 43074
rect 30465 43016 30470 43072
rect 30526 43016 36174 43072
rect 36230 43016 36235 43072
rect 30465 43014 36235 43016
rect 30465 43011 30531 43014
rect 36169 43011 36235 43014
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 31845 42802 31911 42805
rect 32857 42802 32923 42805
rect 35893 42802 35959 42805
rect 31845 42800 35959 42802
rect 31845 42744 31850 42800
rect 31906 42744 32862 42800
rect 32918 42744 35898 42800
rect 35954 42744 35959 42800
rect 31845 42742 35959 42744
rect 31845 42739 31911 42742
rect 32857 42739 32923 42742
rect 35893 42739 35959 42742
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 19568 41920 19888 41921
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 23105 41170 23171 41173
rect 32857 41170 32923 41173
rect 23105 41168 32923 41170
rect 23105 41112 23110 41168
rect 23166 41112 32862 41168
rect 32918 41112 32923 41168
rect 23105 41110 32923 41112
rect 23105 41107 23171 41110
rect 32857 41107 32923 41110
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 105 39810 171 39813
rect 17309 39810 17375 39813
rect 105 39808 17375 39810
rect 105 39752 110 39808
rect 166 39752 17314 39808
rect 17370 39752 17375 39808
rect 105 39750 17375 39752
rect 105 39747 171 39750
rect 17309 39747 17375 39750
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 12985 39538 13051 39541
rect 31109 39538 31175 39541
rect 12985 39536 31175 39538
rect 12985 39480 12990 39536
rect 13046 39480 31114 39536
rect 31170 39480 31175 39536
rect 12985 39478 31175 39480
rect 12985 39475 13051 39478
rect 31109 39475 31175 39478
rect 2773 39402 2839 39405
rect 19057 39402 19123 39405
rect 2773 39400 19123 39402
rect 2773 39344 2778 39400
rect 2834 39344 19062 39400
rect 19118 39344 19123 39400
rect 2773 39342 19123 39344
rect 2773 39339 2839 39342
rect 19057 39339 19123 39342
rect 0 39176 480 39296
rect 4208 39200 4528 39201
rect 62 38722 122 39176
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 22185 38994 22251 38997
rect 23841 38994 23907 38997
rect 22185 38992 23907 38994
rect 22185 38936 22190 38992
rect 22246 38936 23846 38992
rect 23902 38936 23907 38992
rect 22185 38934 23907 38936
rect 22185 38931 22251 38934
rect 23841 38931 23907 38934
rect 21173 38858 21239 38861
rect 32213 38858 32279 38861
rect 21173 38856 32279 38858
rect 21173 38800 21178 38856
rect 21234 38800 32218 38856
rect 32274 38800 32279 38856
rect 21173 38798 32279 38800
rect 21173 38795 21239 38798
rect 32213 38795 32279 38798
rect 2589 38722 2655 38725
rect 62 38720 2655 38722
rect 62 38664 2594 38720
rect 2650 38664 2655 38720
rect 62 38662 2655 38664
rect 2589 38659 2655 38662
rect 33225 38722 33291 38725
rect 36997 38722 37063 38725
rect 33225 38720 37063 38722
rect 33225 38664 33230 38720
rect 33286 38664 37002 38720
rect 37058 38664 37063 38720
rect 33225 38662 37063 38664
rect 33225 38659 33291 38662
rect 36997 38659 37063 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 17769 38450 17835 38453
rect 25773 38450 25839 38453
rect 17769 38448 25839 38450
rect 17769 38392 17774 38448
rect 17830 38392 25778 38448
rect 25834 38392 25839 38448
rect 17769 38390 25839 38392
rect 17769 38387 17835 38390
rect 25773 38387 25839 38390
rect 30373 38450 30439 38453
rect 36353 38450 36419 38453
rect 30373 38448 36419 38450
rect 30373 38392 30378 38448
rect 30434 38392 36358 38448
rect 36414 38392 36419 38448
rect 30373 38390 36419 38392
rect 30373 38387 30439 38390
rect 36353 38387 36419 38390
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 15837 37770 15903 37773
rect 37825 37770 37891 37773
rect 15837 37768 37891 37770
rect 15837 37712 15842 37768
rect 15898 37712 37830 37768
rect 37886 37712 37891 37768
rect 15837 37710 37891 37712
rect 15837 37707 15903 37710
rect 37825 37707 37891 37710
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 35893 37362 35959 37365
rect 43805 37362 43871 37365
rect 35893 37360 43871 37362
rect 35893 37304 35898 37360
rect 35954 37304 43810 37360
rect 43866 37304 43871 37360
rect 35893 37302 43871 37304
rect 35893 37299 35959 37302
rect 43805 37299 43871 37302
rect 32765 37226 32831 37229
rect 40401 37226 40467 37229
rect 42609 37226 42675 37229
rect 32765 37224 42675 37226
rect 32765 37168 32770 37224
rect 32826 37168 40406 37224
rect 40462 37168 42614 37224
rect 42670 37168 42675 37224
rect 32765 37166 42675 37168
rect 32765 37163 32831 37166
rect 40401 37163 40467 37166
rect 42609 37163 42675 37166
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 33777 36818 33843 36821
rect 42057 36818 42123 36821
rect 33777 36816 42123 36818
rect 33777 36760 33782 36816
rect 33838 36760 42062 36816
rect 42118 36760 42123 36816
rect 33777 36758 42123 36760
rect 33777 36755 33843 36758
rect 42057 36755 42123 36758
rect 22645 36682 22711 36685
rect 24669 36682 24735 36685
rect 29637 36682 29703 36685
rect 22645 36680 23490 36682
rect 22645 36624 22650 36680
rect 22706 36624 23490 36680
rect 22645 36622 23490 36624
rect 22645 36619 22711 36622
rect 23430 36546 23490 36622
rect 24669 36680 29703 36682
rect 24669 36624 24674 36680
rect 24730 36624 29642 36680
rect 29698 36624 29703 36680
rect 24669 36622 29703 36624
rect 24669 36619 24735 36622
rect 29637 36619 29703 36622
rect 28073 36546 28139 36549
rect 35709 36546 35775 36549
rect 23430 36544 35775 36546
rect 23430 36488 28078 36544
rect 28134 36488 35714 36544
rect 35770 36488 35775 36544
rect 23430 36486 35775 36488
rect 28073 36483 28139 36486
rect 35709 36483 35775 36486
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 32213 36138 32279 36141
rect 33501 36138 33567 36141
rect 42701 36138 42767 36141
rect 32213 36136 42767 36138
rect 32213 36080 32218 36136
rect 32274 36080 33506 36136
rect 33562 36080 42706 36136
rect 42762 36080 42767 36136
rect 32213 36078 42767 36080
rect 32213 36075 32279 36078
rect 33501 36075 33567 36078
rect 42701 36075 42767 36078
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 17217 35186 17283 35189
rect 29177 35186 29243 35189
rect 17217 35184 29243 35186
rect 17217 35128 17222 35184
rect 17278 35128 29182 35184
rect 29238 35128 29243 35184
rect 17217 35126 29243 35128
rect 17217 35123 17283 35126
rect 29177 35123 29243 35126
rect 29545 35050 29611 35053
rect 34513 35050 34579 35053
rect 38377 35050 38443 35053
rect 29545 35048 38443 35050
rect 29545 34992 29550 35048
rect 29606 34992 34518 35048
rect 34574 34992 38382 35048
rect 38438 34992 38443 35048
rect 29545 34990 38443 34992
rect 29545 34987 29611 34990
rect 34513 34987 34579 34990
rect 38377 34987 38443 34990
rect 49520 34916 50000 34944
rect 49520 34914 49556 34916
rect 49428 34854 49556 34914
rect 49520 34852 49556 34854
rect 49620 34852 50000 34916
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 49520 34824 50000 34852
rect 34928 34783 35248 34784
rect 39849 34778 39915 34781
rect 43345 34778 43411 34781
rect 39849 34776 43411 34778
rect 39849 34720 39854 34776
rect 39910 34720 43350 34776
rect 43406 34720 43411 34776
rect 39849 34718 43411 34720
rect 39849 34715 39915 34718
rect 43345 34715 43411 34718
rect 43805 34778 43871 34781
rect 43805 34776 48330 34778
rect 43805 34720 43810 34776
rect 43866 34720 48330 34776
rect 43805 34718 48330 34720
rect 43805 34715 43871 34718
rect 21173 34642 21239 34645
rect 22461 34642 22527 34645
rect 26141 34642 26207 34645
rect 33685 34642 33751 34645
rect 21173 34640 33751 34642
rect 21173 34584 21178 34640
rect 21234 34584 22466 34640
rect 22522 34584 26146 34640
rect 26202 34584 33690 34640
rect 33746 34584 33751 34640
rect 21173 34582 33751 34584
rect 48270 34642 48330 34718
rect 49550 34642 49556 34644
rect 48270 34582 49556 34642
rect 21173 34579 21239 34582
rect 22461 34579 22527 34582
rect 26141 34579 26207 34582
rect 33685 34579 33751 34582
rect 49550 34580 49556 34582
rect 49620 34580 49626 34644
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 28257 34098 28323 34101
rect 34421 34098 34487 34101
rect 28257 34096 34487 34098
rect 28257 34040 28262 34096
rect 28318 34040 34426 34096
rect 34482 34040 34487 34096
rect 28257 34038 34487 34040
rect 28257 34035 28323 34038
rect 34421 34035 34487 34038
rect 28901 33962 28967 33965
rect 30741 33962 30807 33965
rect 33317 33962 33383 33965
rect 28901 33960 33383 33962
rect 28901 33904 28906 33960
rect 28962 33904 30746 33960
rect 30802 33904 33322 33960
rect 33378 33904 33383 33960
rect 28901 33902 33383 33904
rect 28901 33899 28967 33902
rect 30741 33899 30807 33902
rect 33317 33899 33383 33902
rect 25589 33826 25655 33829
rect 33225 33826 33291 33829
rect 25589 33824 33291 33826
rect 25589 33768 25594 33824
rect 25650 33768 33230 33824
rect 33286 33768 33291 33824
rect 25589 33766 33291 33768
rect 25589 33763 25655 33766
rect 33225 33763 33291 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 20897 33418 20963 33421
rect 25773 33418 25839 33421
rect 20897 33416 25839 33418
rect 20897 33360 20902 33416
rect 20958 33360 25778 33416
rect 25834 33360 25839 33416
rect 20897 33358 25839 33360
rect 20897 33355 20963 33358
rect 25773 33355 25839 33358
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 25497 33146 25563 33149
rect 26141 33146 26207 33149
rect 32581 33146 32647 33149
rect 25497 33144 32647 33146
rect 25497 33088 25502 33144
rect 25558 33088 26146 33144
rect 26202 33088 32586 33144
rect 32642 33088 32647 33144
rect 25497 33086 32647 33088
rect 25497 33083 25563 33086
rect 26141 33083 26207 33086
rect 32581 33083 32647 33086
rect 38101 33146 38167 33149
rect 41965 33146 42031 33149
rect 38101 33144 42031 33146
rect 38101 33088 38106 33144
rect 38162 33088 41970 33144
rect 42026 33088 42031 33144
rect 38101 33086 42031 33088
rect 38101 33083 38167 33086
rect 41965 33083 42031 33086
rect 17217 33010 17283 33013
rect 23381 33010 23447 33013
rect 27797 33010 27863 33013
rect 30373 33010 30439 33013
rect 17217 33008 30439 33010
rect 17217 32952 17222 33008
rect 17278 32952 23386 33008
rect 23442 32952 27802 33008
rect 27858 32952 30378 33008
rect 30434 32952 30439 33008
rect 17217 32950 30439 32952
rect 17217 32947 17283 32950
rect 23381 32947 23447 32950
rect 27797 32947 27863 32950
rect 30373 32947 30439 32950
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 26049 32466 26115 32469
rect 34053 32466 34119 32469
rect 26049 32464 34119 32466
rect 26049 32408 26054 32464
rect 26110 32408 34058 32464
rect 34114 32408 34119 32464
rect 26049 32406 34119 32408
rect 26049 32403 26115 32406
rect 34053 32403 34119 32406
rect 38929 32330 38995 32333
rect 42425 32330 42491 32333
rect 38929 32328 42491 32330
rect 38929 32272 38934 32328
rect 38990 32272 42430 32328
rect 42486 32272 42491 32328
rect 38929 32270 42491 32272
rect 38929 32267 38995 32270
rect 42425 32267 42491 32270
rect 0 32104 480 32224
rect 19568 32128 19888 32129
rect 62 31650 122 32104
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 12065 31786 12131 31789
rect 15469 31786 15535 31789
rect 12065 31784 15535 31786
rect 12065 31728 12070 31784
rect 12126 31728 15474 31784
rect 15530 31728 15535 31784
rect 12065 31726 15535 31728
rect 12065 31723 12131 31726
rect 15469 31723 15535 31726
rect 3325 31650 3391 31653
rect 62 31648 3391 31650
rect 62 31592 3330 31648
rect 3386 31592 3391 31648
rect 62 31590 3391 31592
rect 3325 31587 3391 31590
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 8385 30290 8451 30293
rect 14457 30290 14523 30293
rect 8385 30288 14523 30290
rect 8385 30232 8390 30288
rect 8446 30232 14462 30288
rect 14518 30232 14523 30288
rect 8385 30230 14523 30232
rect 8385 30227 8451 30230
rect 14457 30227 14523 30230
rect 4981 30154 5047 30157
rect 14549 30154 14615 30157
rect 4981 30152 14615 30154
rect 4981 30096 4986 30152
rect 5042 30096 14554 30152
rect 14610 30096 14615 30152
rect 4981 30094 14615 30096
rect 4981 30091 5047 30094
rect 14549 30091 14615 30094
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 23749 29746 23815 29749
rect 33869 29746 33935 29749
rect 23749 29744 33935 29746
rect 23749 29688 23754 29744
rect 23810 29688 33874 29744
rect 33930 29688 33935 29744
rect 23749 29686 33935 29688
rect 23749 29683 23815 29686
rect 33869 29683 33935 29686
rect 5349 29610 5415 29613
rect 16941 29610 17007 29613
rect 5349 29608 17007 29610
rect 5349 29552 5354 29608
rect 5410 29552 16946 29608
rect 17002 29552 17007 29608
rect 5349 29550 17007 29552
rect 5349 29547 5415 29550
rect 16941 29547 17007 29550
rect 22369 29610 22435 29613
rect 23473 29610 23539 29613
rect 27981 29610 28047 29613
rect 39757 29610 39823 29613
rect 22369 29608 39823 29610
rect 22369 29552 22374 29608
rect 22430 29552 23478 29608
rect 23534 29552 27986 29608
rect 28042 29552 39762 29608
rect 39818 29552 39823 29608
rect 22369 29550 39823 29552
rect 22369 29547 22435 29550
rect 23473 29547 23539 29550
rect 27981 29547 28047 29550
rect 39757 29547 39823 29550
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 9857 29066 9923 29069
rect 15469 29066 15535 29069
rect 9857 29064 15535 29066
rect 9857 29008 9862 29064
rect 9918 29008 15474 29064
rect 15530 29008 15535 29064
rect 9857 29006 15535 29008
rect 9857 29003 9923 29006
rect 15469 29003 15535 29006
rect 3969 28930 4035 28933
rect 4521 28930 4587 28933
rect 3969 28928 4587 28930
rect 3969 28872 3974 28928
rect 4030 28872 4526 28928
rect 4582 28872 4587 28928
rect 3969 28870 4587 28872
rect 3969 28867 4035 28870
rect 4521 28867 4587 28870
rect 9673 28930 9739 28933
rect 16573 28930 16639 28933
rect 9673 28928 16639 28930
rect 9673 28872 9678 28928
rect 9734 28872 16578 28928
rect 16634 28872 16639 28928
rect 9673 28870 16639 28872
rect 9673 28867 9739 28870
rect 16573 28867 16639 28870
rect 30557 28930 30623 28933
rect 36077 28930 36143 28933
rect 30557 28928 36143 28930
rect 30557 28872 30562 28928
rect 30618 28872 36082 28928
rect 36138 28872 36143 28928
rect 30557 28870 36143 28872
rect 30557 28867 30623 28870
rect 36077 28867 36143 28870
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 22001 28794 22067 28797
rect 26601 28794 26667 28797
rect 38929 28794 38995 28797
rect 22001 28792 38995 28794
rect 22001 28736 22006 28792
rect 22062 28736 26606 28792
rect 26662 28736 38934 28792
rect 38990 28736 38995 28792
rect 22001 28734 38995 28736
rect 22001 28731 22067 28734
rect 26601 28731 26667 28734
rect 38929 28731 38995 28734
rect 25221 28658 25287 28661
rect 26509 28658 26575 28661
rect 34605 28658 34671 28661
rect 25221 28656 34671 28658
rect 25221 28600 25226 28656
rect 25282 28600 26514 28656
rect 26570 28600 34610 28656
rect 34666 28600 34671 28656
rect 25221 28598 34671 28600
rect 25221 28595 25287 28598
rect 26509 28595 26575 28598
rect 34605 28595 34671 28598
rect 21081 28522 21147 28525
rect 27981 28522 28047 28525
rect 39113 28522 39179 28525
rect 21081 28520 39179 28522
rect 21081 28464 21086 28520
rect 21142 28464 27986 28520
rect 28042 28464 39118 28520
rect 39174 28464 39179 28520
rect 21081 28462 39179 28464
rect 21081 28459 21147 28462
rect 27981 28459 28047 28462
rect 39113 28459 39179 28462
rect 27153 28386 27219 28389
rect 29729 28386 29795 28389
rect 34789 28386 34855 28389
rect 27153 28384 34855 28386
rect 27153 28328 27158 28384
rect 27214 28328 29734 28384
rect 29790 28328 34794 28384
rect 34850 28328 34855 28384
rect 27153 28326 34855 28328
rect 27153 28323 27219 28326
rect 29729 28323 29795 28326
rect 34789 28323 34855 28326
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 18965 28114 19031 28117
rect 25037 28114 25103 28117
rect 37733 28114 37799 28117
rect 18965 28112 37799 28114
rect 18965 28056 18970 28112
rect 19026 28056 25042 28112
rect 25098 28056 37738 28112
rect 37794 28056 37799 28112
rect 18965 28054 37799 28056
rect 18965 28051 19031 28054
rect 25037 28051 25103 28054
rect 37733 28051 37799 28054
rect 21725 27842 21791 27845
rect 31201 27842 31267 27845
rect 21725 27840 31267 27842
rect 21725 27784 21730 27840
rect 21786 27784 31206 27840
rect 31262 27784 31267 27840
rect 21725 27782 31267 27784
rect 21725 27779 21791 27782
rect 31201 27779 31267 27782
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 32949 27706 33015 27709
rect 39021 27706 39087 27709
rect 41689 27706 41755 27709
rect 32949 27704 41755 27706
rect 32949 27648 32954 27704
rect 33010 27648 39026 27704
rect 39082 27648 41694 27704
rect 41750 27648 41755 27704
rect 32949 27646 41755 27648
rect 32949 27643 33015 27646
rect 39021 27643 39087 27646
rect 41689 27643 41755 27646
rect 39205 27570 39271 27573
rect 44541 27570 44607 27573
rect 39205 27568 44607 27570
rect 39205 27512 39210 27568
rect 39266 27512 44546 27568
rect 44602 27512 44607 27568
rect 39205 27510 44607 27512
rect 39205 27507 39271 27510
rect 44541 27507 44607 27510
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 23933 26618 23999 26621
rect 32029 26618 32095 26621
rect 23933 26616 32095 26618
rect 23933 26560 23938 26616
rect 23994 26560 32034 26616
rect 32090 26560 32095 26616
rect 23933 26558 32095 26560
rect 23933 26555 23999 26558
rect 32029 26555 32095 26558
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 40953 25666 41019 25669
rect 44633 25666 44699 25669
rect 40953 25664 44699 25666
rect 40953 25608 40958 25664
rect 41014 25608 44638 25664
rect 44694 25608 44699 25664
rect 40953 25606 44699 25608
rect 40953 25603 41019 25606
rect 44633 25603 44699 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 4208 25056 4528 25057
rect 0 24984 480 25016
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 49520 24988 50000 25016
rect 49520 24986 49556 24988
rect 0 24928 110 24984
rect 166 24928 480 24984
rect 0 24896 480 24928
rect 49428 24926 49556 24986
rect 49520 24924 49556 24926
rect 49620 24924 50000 24988
rect 49520 24896 50000 24924
rect 19793 24850 19859 24853
rect 23473 24850 23539 24853
rect 19793 24848 23539 24850
rect 19793 24792 19798 24848
rect 19854 24792 23478 24848
rect 23534 24792 23539 24848
rect 19793 24790 23539 24792
rect 19793 24787 19859 24790
rect 23473 24787 23539 24790
rect 44817 24850 44883 24853
rect 49366 24850 49372 24852
rect 44817 24848 49372 24850
rect 44817 24792 44822 24848
rect 44878 24792 49372 24848
rect 44817 24790 49372 24792
rect 44817 24787 44883 24790
rect 49366 24788 49372 24790
rect 49436 24788 49442 24852
rect 26601 24714 26667 24717
rect 33593 24714 33659 24717
rect 40953 24714 41019 24717
rect 26601 24712 41019 24714
rect 26601 24656 26606 24712
rect 26662 24656 33598 24712
rect 33654 24656 40958 24712
rect 41014 24656 41019 24712
rect 26601 24654 41019 24656
rect 26601 24651 26667 24654
rect 33593 24651 33659 24654
rect 40953 24651 41019 24654
rect 40861 24578 40927 24581
rect 44265 24578 44331 24581
rect 40861 24576 44331 24578
rect 40861 24520 40866 24576
rect 40922 24520 44270 24576
rect 44326 24520 44331 24576
rect 40861 24518 44331 24520
rect 40861 24515 40927 24518
rect 44265 24515 44331 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 37825 24442 37891 24445
rect 42977 24442 43043 24445
rect 37825 24440 43043 24442
rect 37825 24384 37830 24440
rect 37886 24384 42982 24440
rect 43038 24384 43043 24440
rect 37825 24382 43043 24384
rect 37825 24379 37891 24382
rect 42977 24379 43043 24382
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 4889 23626 4955 23629
rect 5993 23626 6059 23629
rect 8937 23626 9003 23629
rect 4889 23624 9003 23626
rect 4889 23568 4894 23624
rect 4950 23568 5998 23624
rect 6054 23568 8942 23624
rect 8998 23568 9003 23624
rect 4889 23566 9003 23568
rect 4889 23563 4955 23566
rect 5993 23563 6059 23566
rect 8937 23563 9003 23566
rect 31201 23626 31267 23629
rect 32397 23626 32463 23629
rect 31201 23624 32463 23626
rect 31201 23568 31206 23624
rect 31262 23568 32402 23624
rect 32458 23568 32463 23624
rect 31201 23566 32463 23568
rect 31201 23563 31267 23566
rect 32397 23563 32463 23566
rect 17493 23490 17559 23493
rect 18965 23490 19031 23493
rect 17493 23488 19031 23490
rect 17493 23432 17498 23488
rect 17554 23432 18970 23488
rect 19026 23432 19031 23488
rect 17493 23430 19031 23432
rect 17493 23427 17559 23430
rect 18965 23427 19031 23430
rect 43846 23428 43852 23492
rect 43916 23490 43922 23492
rect 44633 23490 44699 23493
rect 43916 23488 44699 23490
rect 43916 23432 44638 23488
rect 44694 23432 44699 23488
rect 43916 23430 44699 23432
rect 43916 23428 43922 23430
rect 44633 23427 44699 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 23105 23218 23171 23221
rect 23422 23218 23428 23220
rect 23105 23216 23428 23218
rect 23105 23160 23110 23216
rect 23166 23160 23428 23216
rect 23105 23158 23428 23160
rect 23105 23155 23171 23158
rect 23422 23156 23428 23158
rect 23492 23218 23498 23220
rect 30741 23218 30807 23221
rect 30925 23218 30991 23221
rect 23492 23216 30991 23218
rect 23492 23160 30746 23216
rect 30802 23160 30930 23216
rect 30986 23160 30991 23216
rect 23492 23158 30991 23160
rect 23492 23156 23498 23158
rect 30741 23155 30807 23158
rect 30925 23155 30991 23158
rect 9949 23082 10015 23085
rect 24669 23082 24735 23085
rect 9949 23080 24735 23082
rect 9949 23024 9954 23080
rect 10010 23024 24674 23080
rect 24730 23024 24735 23080
rect 9949 23022 24735 23024
rect 9949 23019 10015 23022
rect 24669 23019 24735 23022
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 19241 22674 19307 22677
rect 35985 22674 36051 22677
rect 19241 22672 36051 22674
rect 19241 22616 19246 22672
rect 19302 22616 35990 22672
rect 36046 22616 36051 22672
rect 19241 22614 36051 22616
rect 19241 22611 19307 22614
rect 35985 22611 36051 22614
rect 8753 22538 8819 22541
rect 19425 22538 19491 22541
rect 8753 22536 19491 22538
rect 8753 22480 8758 22536
rect 8814 22480 19430 22536
rect 19486 22480 19491 22536
rect 8753 22478 19491 22480
rect 8753 22475 8819 22478
rect 19425 22475 19491 22478
rect 20161 22402 20227 22405
rect 44725 22402 44791 22405
rect 20161 22400 44791 22402
rect 20161 22344 20166 22400
rect 20222 22344 44730 22400
rect 44786 22344 44791 22400
rect 20161 22342 44791 22344
rect 20161 22339 20227 22342
rect 44725 22339 44791 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 23841 22266 23907 22269
rect 30373 22266 30439 22269
rect 23841 22264 30439 22266
rect 23841 22208 23846 22264
rect 23902 22208 30378 22264
rect 30434 22208 30439 22264
rect 23841 22206 30439 22208
rect 23841 22203 23907 22206
rect 30373 22203 30439 22206
rect 13353 21994 13419 21997
rect 21817 21994 21883 21997
rect 13353 21992 21883 21994
rect 13353 21936 13358 21992
rect 13414 21936 21822 21992
rect 21878 21936 21883 21992
rect 13353 21934 21883 21936
rect 13353 21931 13419 21934
rect 21817 21931 21883 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 36721 21586 36787 21589
rect 43437 21586 43503 21589
rect 44725 21586 44791 21589
rect 36721 21584 44791 21586
rect 36721 21528 36726 21584
rect 36782 21528 43442 21584
rect 43498 21528 44730 21584
rect 44786 21528 44791 21584
rect 36721 21526 44791 21528
rect 36721 21523 36787 21526
rect 43437 21523 43503 21526
rect 44725 21523 44791 21526
rect 33593 21450 33659 21453
rect 45461 21450 45527 21453
rect 33593 21448 45527 21450
rect 33593 21392 33598 21448
rect 33654 21392 45466 21448
rect 45522 21392 45527 21448
rect 33593 21390 45527 21392
rect 33593 21387 33659 21390
rect 45461 21387 45527 21390
rect 35157 21314 35223 21317
rect 44909 21314 44975 21317
rect 35157 21312 44975 21314
rect 35157 21256 35162 21312
rect 35218 21256 44914 21312
rect 44970 21256 44975 21312
rect 35157 21254 44975 21256
rect 35157 21251 35223 21254
rect 44909 21251 44975 21254
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 27337 21042 27403 21045
rect 30557 21042 30623 21045
rect 27337 21040 30623 21042
rect 27337 20984 27342 21040
rect 27398 20984 30562 21040
rect 30618 20984 30623 21040
rect 27337 20982 30623 20984
rect 27337 20979 27403 20982
rect 30557 20979 30623 20982
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 7557 20498 7623 20501
rect 16941 20498 17007 20501
rect 7557 20496 17007 20498
rect 7557 20440 7562 20496
rect 7618 20440 16946 20496
rect 17002 20440 17007 20496
rect 7557 20438 17007 20440
rect 7557 20435 7623 20438
rect 16941 20435 17007 20438
rect 31937 20498 32003 20501
rect 38101 20498 38167 20501
rect 31937 20496 38167 20498
rect 31937 20440 31942 20496
rect 31998 20440 38106 20496
rect 38162 20440 38167 20496
rect 31937 20438 38167 20440
rect 31937 20435 32003 20438
rect 38101 20435 38167 20438
rect 35157 20362 35223 20365
rect 45461 20362 45527 20365
rect 35157 20360 45527 20362
rect 35157 20304 35162 20360
rect 35218 20304 45466 20360
rect 45522 20304 45527 20360
rect 35157 20302 45527 20304
rect 35157 20299 35223 20302
rect 35896 20229 35956 20302
rect 45461 20299 45527 20302
rect 35893 20224 35959 20229
rect 35893 20168 35898 20224
rect 35954 20168 35959 20224
rect 35893 20163 35959 20168
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 30005 20090 30071 20093
rect 43846 20090 43852 20092
rect 30005 20088 43852 20090
rect 30005 20032 30010 20088
rect 30066 20032 43852 20088
rect 30005 20030 43852 20032
rect 30005 20027 30071 20030
rect 43846 20028 43852 20030
rect 43916 20028 43922 20092
rect 3417 19954 3483 19957
rect 22645 19954 22711 19957
rect 3417 19952 22711 19954
rect 3417 19896 3422 19952
rect 3478 19896 22650 19952
rect 22706 19896 22711 19952
rect 3417 19894 22711 19896
rect 3417 19891 3483 19894
rect 22645 19891 22711 19894
rect 28073 19818 28139 19821
rect 37733 19818 37799 19821
rect 28073 19816 37799 19818
rect 28073 19760 28078 19816
rect 28134 19760 37738 19816
rect 37794 19760 37799 19816
rect 28073 19758 37799 19760
rect 28073 19755 28139 19758
rect 37733 19755 37799 19758
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 32397 19546 32463 19549
rect 33041 19546 33107 19549
rect 32397 19544 33107 19546
rect 32397 19488 32402 19544
rect 32458 19488 33046 19544
rect 33102 19488 33107 19544
rect 32397 19486 33107 19488
rect 32397 19483 32463 19486
rect 33041 19483 33107 19486
rect 14365 19410 14431 19413
rect 24301 19410 24367 19413
rect 14365 19408 24367 19410
rect 14365 19352 14370 19408
rect 14426 19352 24306 19408
rect 24362 19352 24367 19408
rect 14365 19350 24367 19352
rect 14365 19347 14431 19350
rect 24301 19347 24367 19350
rect 31385 19410 31451 19413
rect 33225 19410 33291 19413
rect 31385 19408 33291 19410
rect 31385 19352 31390 19408
rect 31446 19352 33230 19408
rect 33286 19352 33291 19408
rect 31385 19350 33291 19352
rect 31385 19347 31451 19350
rect 33225 19347 33291 19350
rect 31385 19138 31451 19141
rect 32029 19138 32095 19141
rect 31385 19136 32095 19138
rect 31385 19080 31390 19136
rect 31446 19080 32034 19136
rect 32090 19080 32095 19136
rect 31385 19078 32095 19080
rect 31385 19075 31451 19078
rect 32029 19075 32095 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 7557 19002 7623 19005
rect 17217 19002 17283 19005
rect 7557 19000 17283 19002
rect 7557 18944 7562 19000
rect 7618 18944 17222 19000
rect 17278 18944 17283 19000
rect 7557 18942 17283 18944
rect 7557 18939 7623 18942
rect 17217 18939 17283 18942
rect 30097 19002 30163 19005
rect 44817 19002 44883 19005
rect 30097 19000 44883 19002
rect 30097 18944 30102 19000
rect 30158 18944 44822 19000
rect 44878 18944 44883 19000
rect 30097 18942 44883 18944
rect 30097 18939 30163 18942
rect 44817 18939 44883 18942
rect 2589 18866 2655 18869
rect 24485 18866 24551 18869
rect 2589 18864 24551 18866
rect 2589 18808 2594 18864
rect 2650 18808 24490 18864
rect 24546 18808 24551 18864
rect 2589 18806 24551 18808
rect 2589 18803 2655 18806
rect 24485 18803 24551 18806
rect 26877 18866 26943 18869
rect 27429 18866 27495 18869
rect 33593 18866 33659 18869
rect 26877 18864 33659 18866
rect 26877 18808 26882 18864
rect 26938 18808 27434 18864
rect 27490 18808 33598 18864
rect 33654 18808 33659 18864
rect 26877 18806 33659 18808
rect 26877 18803 26943 18806
rect 27429 18803 27495 18806
rect 33593 18803 33659 18806
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 1945 18458 2011 18461
rect 62 18456 2011 18458
rect 62 18400 1950 18456
rect 2006 18400 2011 18456
rect 62 18398 2011 18400
rect 62 17944 122 18398
rect 1945 18395 2011 18398
rect 8845 18458 8911 18461
rect 16941 18458 17007 18461
rect 8845 18456 17007 18458
rect 8845 18400 8850 18456
rect 8906 18400 16946 18456
rect 17002 18400 17007 18456
rect 8845 18398 17007 18400
rect 8845 18395 8911 18398
rect 16941 18395 17007 18398
rect 33501 18322 33567 18325
rect 36997 18322 37063 18325
rect 33501 18320 37063 18322
rect 33501 18264 33506 18320
rect 33562 18264 37002 18320
rect 37058 18264 37063 18320
rect 33501 18262 37063 18264
rect 33501 18259 33567 18262
rect 36997 18259 37063 18262
rect 21725 18186 21791 18189
rect 30741 18186 30807 18189
rect 21725 18184 30807 18186
rect 21725 18128 21730 18184
rect 21786 18128 30746 18184
rect 30802 18128 30807 18184
rect 21725 18126 30807 18128
rect 21725 18123 21791 18126
rect 30741 18123 30807 18126
rect 31477 18186 31543 18189
rect 38653 18186 38719 18189
rect 31477 18184 38719 18186
rect 31477 18128 31482 18184
rect 31538 18128 38658 18184
rect 38714 18128 38719 18184
rect 31477 18126 38719 18128
rect 31477 18123 31543 18126
rect 38653 18123 38719 18126
rect 19568 17984 19888 17985
rect 0 17824 480 17944
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 21449 17914 21515 17917
rect 23105 17914 23171 17917
rect 30281 17914 30347 17917
rect 21449 17912 30347 17914
rect 21449 17856 21454 17912
rect 21510 17856 23110 17912
rect 23166 17856 30286 17912
rect 30342 17856 30347 17912
rect 21449 17854 30347 17856
rect 21449 17851 21515 17854
rect 23105 17851 23171 17854
rect 30281 17851 30347 17854
rect 22001 17506 22067 17509
rect 28165 17506 28231 17509
rect 22001 17504 28231 17506
rect 22001 17448 22006 17504
rect 22062 17448 28170 17504
rect 28226 17448 28231 17504
rect 22001 17446 28231 17448
rect 22001 17443 22067 17446
rect 28165 17443 28231 17446
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 18045 17370 18111 17373
rect 24301 17370 24367 17373
rect 18045 17368 24367 17370
rect 18045 17312 18050 17368
rect 18106 17312 24306 17368
rect 24362 17312 24367 17368
rect 18045 17310 24367 17312
rect 18045 17307 18111 17310
rect 24301 17307 24367 17310
rect 22829 17234 22895 17237
rect 32673 17234 32739 17237
rect 22829 17232 32739 17234
rect 22829 17176 22834 17232
rect 22890 17176 32678 17232
rect 32734 17176 32739 17232
rect 22829 17174 32739 17176
rect 22829 17171 22895 17174
rect 32673 17171 32739 17174
rect 14365 17098 14431 17101
rect 23473 17098 23539 17101
rect 14365 17096 23539 17098
rect 14365 17040 14370 17096
rect 14426 17040 23478 17096
rect 23534 17040 23539 17096
rect 14365 17038 23539 17040
rect 14365 17035 14431 17038
rect 23473 17035 23539 17038
rect 35985 16962 36051 16965
rect 42517 16962 42583 16965
rect 43529 16962 43595 16965
rect 35985 16960 43595 16962
rect 35985 16904 35990 16960
rect 36046 16904 42522 16960
rect 42578 16904 43534 16960
rect 43590 16904 43595 16960
rect 35985 16902 43595 16904
rect 35985 16899 36051 16902
rect 42517 16899 42583 16902
rect 43529 16899 43595 16902
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 29177 16826 29243 16829
rect 39297 16826 39363 16829
rect 29177 16824 39363 16826
rect 29177 16768 29182 16824
rect 29238 16768 39302 16824
rect 39358 16768 39363 16824
rect 29177 16766 39363 16768
rect 29177 16763 29243 16766
rect 39297 16763 39363 16766
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 18505 16010 18571 16013
rect 19374 16010 19380 16012
rect 18505 16008 19380 16010
rect 18505 15952 18510 16008
rect 18566 15952 19380 16008
rect 18505 15950 19380 15952
rect 18505 15947 18571 15950
rect 19374 15948 19380 15950
rect 19444 15948 19450 16012
rect 28625 16010 28691 16013
rect 30373 16010 30439 16013
rect 36261 16010 36327 16013
rect 28625 16008 36327 16010
rect 28625 15952 28630 16008
rect 28686 15952 30378 16008
rect 30434 15952 36266 16008
rect 36322 15952 36327 16008
rect 28625 15950 36327 15952
rect 28625 15947 28691 15950
rect 30373 15947 30439 15950
rect 36261 15947 36327 15950
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 28165 15738 28231 15741
rect 37365 15738 37431 15741
rect 28165 15736 37431 15738
rect 28165 15680 28170 15736
rect 28226 15680 37370 15736
rect 37426 15680 37431 15736
rect 28165 15678 37431 15680
rect 28165 15675 28231 15678
rect 37365 15675 37431 15678
rect 35065 15466 35131 15469
rect 45001 15466 45067 15469
rect 35065 15464 45067 15466
rect 35065 15408 35070 15464
rect 35126 15408 45006 15464
rect 45062 15408 45067 15464
rect 35065 15406 45067 15408
rect 35065 15403 35131 15406
rect 45001 15403 45067 15406
rect 27613 15330 27679 15333
rect 34697 15330 34763 15333
rect 27613 15328 34763 15330
rect 27613 15272 27618 15328
rect 27674 15272 34702 15328
rect 34758 15272 34763 15328
rect 27613 15270 34763 15272
rect 27613 15267 27679 15270
rect 34697 15267 34763 15270
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 36261 15194 36327 15197
rect 44725 15194 44791 15197
rect 36261 15192 44791 15194
rect 36261 15136 36266 15192
rect 36322 15136 44730 15192
rect 44786 15136 44791 15192
rect 36261 15134 44791 15136
rect 36261 15131 36327 15134
rect 44725 15131 44791 15134
rect 22921 15058 22987 15061
rect 34605 15058 34671 15061
rect 22921 15056 34671 15058
rect 22921 15000 22926 15056
rect 22982 15000 34610 15056
rect 34666 15000 34671 15056
rect 22921 14998 34671 15000
rect 22921 14995 22987 14998
rect 34605 14995 34671 14998
rect 49520 14925 50000 14952
rect 49509 14922 50000 14925
rect 49428 14920 50000 14922
rect 49428 14864 49514 14920
rect 49570 14864 50000 14920
rect 49428 14862 50000 14864
rect 49509 14859 50000 14862
rect 49520 14832 50000 14859
rect 32949 14786 33015 14789
rect 42517 14786 42583 14789
rect 32949 14784 42583 14786
rect 32949 14728 32954 14784
rect 33010 14728 42522 14784
rect 42578 14728 42583 14784
rect 32949 14726 42583 14728
rect 32949 14723 33015 14726
rect 42517 14723 42583 14726
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 21081 14242 21147 14245
rect 23422 14242 23428 14244
rect 21081 14240 23428 14242
rect 21081 14184 21086 14240
rect 21142 14184 23428 14240
rect 21081 14182 23428 14184
rect 21081 14179 21147 14182
rect 23422 14180 23428 14182
rect 23492 14180 23498 14244
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 28809 13970 28875 13973
rect 36077 13970 36143 13973
rect 28809 13968 36143 13970
rect 28809 13912 28814 13968
rect 28870 13912 36082 13968
rect 36138 13912 36143 13968
rect 28809 13910 36143 13912
rect 28809 13907 28875 13910
rect 33041 13834 33107 13837
rect 33869 13834 33935 13837
rect 33041 13832 33935 13834
rect 33041 13776 33046 13832
rect 33102 13776 33874 13832
rect 33930 13776 33935 13832
rect 33041 13774 33935 13776
rect 33041 13771 33107 13774
rect 33869 13771 33935 13774
rect 23197 13698 23263 13701
rect 31293 13698 31359 13701
rect 23197 13696 31359 13698
rect 23197 13640 23202 13696
rect 23258 13640 31298 13696
rect 31354 13640 31359 13696
rect 23197 13638 31359 13640
rect 23197 13635 23263 13638
rect 31293 13635 31359 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 24945 13562 25011 13565
rect 31201 13562 31267 13565
rect 24945 13560 31267 13562
rect 24945 13504 24950 13560
rect 25006 13504 31206 13560
rect 31262 13504 31267 13560
rect 24945 13502 31267 13504
rect 24945 13499 25011 13502
rect 31201 13499 31267 13502
rect 35758 13426 35818 13910
rect 36077 13907 36143 13910
rect 42609 13970 42675 13973
rect 49509 13970 49575 13973
rect 42609 13968 49575 13970
rect 42609 13912 42614 13968
rect 42670 13912 49514 13968
rect 49570 13912 49575 13968
rect 42609 13910 49575 13912
rect 42609 13907 42675 13910
rect 49509 13907 49575 13910
rect 35893 13834 35959 13837
rect 37549 13834 37615 13837
rect 43897 13834 43963 13837
rect 35893 13832 43963 13834
rect 35893 13776 35898 13832
rect 35954 13776 37554 13832
rect 37610 13776 43902 13832
rect 43958 13776 43963 13832
rect 35893 13774 43963 13776
rect 35893 13771 35959 13774
rect 37549 13771 37615 13774
rect 43897 13771 43963 13774
rect 36997 13698 37063 13701
rect 38009 13698 38075 13701
rect 40953 13698 41019 13701
rect 36997 13696 41019 13698
rect 36997 13640 37002 13696
rect 37058 13640 38014 13696
rect 38070 13640 40958 13696
rect 41014 13640 41019 13696
rect 36997 13638 41019 13640
rect 36997 13635 37063 13638
rect 38009 13635 38075 13638
rect 40953 13635 41019 13638
rect 38285 13562 38351 13565
rect 43253 13562 43319 13565
rect 38285 13560 43319 13562
rect 38285 13504 38290 13560
rect 38346 13504 43258 13560
rect 43314 13504 43319 13560
rect 38285 13502 43319 13504
rect 38285 13499 38351 13502
rect 43253 13499 43319 13502
rect 37825 13426 37891 13429
rect 43529 13426 43595 13429
rect 35758 13424 43595 13426
rect 35758 13368 37830 13424
rect 37886 13368 43534 13424
rect 43590 13368 43595 13424
rect 35758 13366 43595 13368
rect 37825 13363 37891 13366
rect 43529 13363 43595 13366
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 28809 12746 28875 12749
rect 34145 12746 34211 12749
rect 28809 12744 34211 12746
rect 28809 12688 28814 12744
rect 28870 12688 34150 12744
rect 34206 12688 34211 12744
rect 28809 12686 34211 12688
rect 28809 12683 28875 12686
rect 34145 12683 34211 12686
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 23105 12338 23171 12341
rect 33777 12338 33843 12341
rect 23105 12336 33843 12338
rect 23105 12280 23110 12336
rect 23166 12280 33782 12336
rect 33838 12280 33843 12336
rect 23105 12278 33843 12280
rect 23105 12275 23171 12278
rect 33777 12275 33843 12278
rect 18597 12202 18663 12205
rect 23473 12202 23539 12205
rect 18597 12200 23539 12202
rect 18597 12144 18602 12200
rect 18658 12144 23478 12200
rect 23534 12144 23539 12200
rect 18597 12142 23539 12144
rect 18597 12139 18663 12142
rect 23473 12139 23539 12142
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 1485 11250 1551 11253
rect 62 11248 1551 11250
rect 62 11192 1490 11248
rect 1546 11192 1551 11248
rect 62 11190 1551 11192
rect 62 10736 122 11190
rect 1485 11187 1551 11190
rect 33225 11114 33291 11117
rect 38101 11114 38167 11117
rect 39297 11114 39363 11117
rect 33225 11112 39363 11114
rect 33225 11056 33230 11112
rect 33286 11056 38106 11112
rect 38162 11056 39302 11112
rect 39358 11056 39363 11112
rect 33225 11054 39363 11056
rect 33225 11051 33291 11054
rect 38101 11051 38167 11054
rect 39297 11051 39363 11054
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 27797 10842 27863 10845
rect 34513 10842 34579 10845
rect 27797 10840 34579 10842
rect 27797 10784 27802 10840
rect 27858 10784 34518 10840
rect 34574 10784 34579 10840
rect 27797 10782 34579 10784
rect 27797 10779 27863 10782
rect 34513 10779 34579 10782
rect 0 10616 480 10736
rect 30189 10706 30255 10709
rect 36077 10706 36143 10709
rect 30189 10704 36143 10706
rect 30189 10648 30194 10704
rect 30250 10648 36082 10704
rect 36138 10648 36143 10704
rect 30189 10646 36143 10648
rect 30189 10643 30255 10646
rect 36077 10643 36143 10646
rect 14825 10570 14891 10573
rect 40493 10570 40559 10573
rect 14825 10568 40559 10570
rect 14825 10512 14830 10568
rect 14886 10512 40498 10568
rect 40554 10512 40559 10568
rect 14825 10510 40559 10512
rect 14825 10507 14891 10510
rect 40493 10507 40559 10510
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 15837 10162 15903 10165
rect 26325 10162 26391 10165
rect 15837 10160 26391 10162
rect 15837 10104 15842 10160
rect 15898 10104 26330 10160
rect 26386 10104 26391 10160
rect 15837 10102 26391 10104
rect 15837 10099 15903 10102
rect 26325 10099 26391 10102
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 23197 9618 23263 9621
rect 23749 9618 23815 9621
rect 23197 9616 23815 9618
rect 23197 9560 23202 9616
rect 23258 9560 23754 9616
rect 23810 9560 23815 9616
rect 23197 9558 23815 9560
rect 23197 9555 23263 9558
rect 23749 9555 23815 9558
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 19241 8938 19307 8941
rect 19374 8938 19380 8940
rect 19241 8936 19380 8938
rect 19241 8880 19246 8936
rect 19302 8880 19380 8936
rect 19241 8878 19380 8880
rect 19241 8875 19307 8878
rect 19374 8876 19380 8878
rect 19444 8876 19450 8940
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 15101 7306 15167 7309
rect 33409 7306 33475 7309
rect 15101 7304 33475 7306
rect 15101 7248 15106 7304
rect 15162 7248 33414 7304
rect 33470 7248 33475 7304
rect 15101 7246 33475 7248
rect 15101 7243 15167 7246
rect 33409 7243 33475 7246
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 49520 4904 50000 5024
rect 19568 4863 19888 4864
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 1393 4178 1459 4181
rect 62 4176 1459 4178
rect 62 4120 1398 4176
rect 1454 4120 1459 4176
rect 62 4118 1459 4120
rect 62 3664 122 4118
rect 1393 4115 1459 4118
rect 3049 4178 3115 4181
rect 13169 4178 13235 4181
rect 3049 4176 13235 4178
rect 3049 4120 3054 4176
rect 3110 4120 13174 4176
rect 13230 4120 13235 4176
rect 3049 4118 13235 4120
rect 3049 4115 3115 4118
rect 13169 4115 13235 4118
rect 23289 4178 23355 4181
rect 49558 4178 49618 4904
rect 23289 4176 49618 4178
rect 23289 4120 23294 4176
rect 23350 4120 49618 4176
rect 23289 4118 49618 4120
rect 23289 4115 23355 4118
rect 28165 3906 28231 3909
rect 36169 3906 36235 3909
rect 28165 3904 36235 3906
rect 28165 3848 28170 3904
rect 28226 3848 36174 3904
rect 36230 3848 36235 3904
rect 28165 3846 36235 3848
rect 28165 3843 28231 3846
rect 36169 3843 36235 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 0 3544 480 3664
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
<< via3 >>
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 49556 34852 49620 34916
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 49556 34580 49620 34644
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 49556 24924 49620 24988
rect 49372 24788 49436 24852
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 43852 23428 43916 23492
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 23428 23156 23492 23220
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 43852 20028 43916 20092
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19380 15948 19444 16012
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 23428 14180 23492 14244
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 19380 8876 19444 8940
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 46816 4528 47376
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 19568 47360 19888 47376
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 34928 46816 35248 47376
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 49555 34916 49621 34917
rect 49555 34852 49556 34916
rect 49620 34852 49621 34916
rect 49555 34851 49621 34852
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 49558 34645 49618 34851
rect 49555 34644 49621 34645
rect 49555 34580 49556 34644
rect 49620 34580 49621 34644
rect 49555 34579 49621 34580
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 49555 24988 49621 24989
rect 49555 24924 49556 24988
rect 49620 24924 49621 24988
rect 49555 24923 49621 24924
rect 49371 24852 49437 24853
rect 49371 24788 49372 24852
rect 49436 24850 49437 24852
rect 49558 24850 49618 24923
rect 49436 24790 49618 24850
rect 49436 24788 49437 24790
rect 49371 24787 49437 24788
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 23427 23220 23493 23221
rect 23427 23156 23428 23220
rect 23492 23156 23493 23220
rect 23427 23155 23493 23156
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19379 16012 19445 16013
rect 19379 15948 19380 16012
rect 19444 15948 19445 16012
rect 19379 15947 19445 15948
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 19382 8941 19442 15947
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 23430 14245 23490 23155
rect 34928 22880 35248 23904
rect 43851 23492 43917 23493
rect 43851 23428 43852 23492
rect 43916 23428 43917 23492
rect 43851 23427 43917 23428
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 43854 20093 43914 23427
rect 43851 20092 43917 20093
rect 43851 20028 43852 20092
rect 43916 20028 43917 20092
rect 43851 20027 43917 20028
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 23427 14244 23493 14245
rect 23427 14180 23428 14244
rect 23492 14180 23493 14244
rect 23427 14179 23493 14180
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19379 8940 19445 8941
rect 19379 8876 19380 8940
rect 19444 8876 19445 8940
rect 19379 8875 19445 8876
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_281
timestamp 1586364061
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_293
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_304
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_330
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_342
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_416
timestamp 1586364061
transform 1 0 39376 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_428
timestamp 1586364061
transform 1 0 40480 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_415
timestamp 1586364061
transform 1 0 39284 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_428
timestamp 1586364061
transform 1 0 40480 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_435
timestamp 1586364061
transform 1 0 41124 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_447
timestamp 1586364061
transform 1 0 42228 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_440
timestamp 1586364061
transform 1 0 41584 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_452
timestamp 1586364061
transform 1 0 42688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_459
timestamp 1586364061
transform 1 0 43332 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_466
timestamp 1586364061
transform 1 0 43976 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_478
timestamp 1586364061
transform 1 0 45080 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_464
timestamp 1586364061
transform 1 0 43792 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_476
timestamp 1586364061
transform 1 0 44896 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_490
timestamp 1586364061
transform 1 0 46184 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_497
timestamp 1586364061
transform 1 0 46828 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_509
timestamp 1586364061
transform 1 0 47932 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_489
timestamp 1586364061
transform 1 0 46092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_501
timestamp 1586364061
transform 1 0 47196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 48852 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 48852 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_515 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 48484 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_513
timestamp 1586364061
transform 1 0 48300 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_324
timestamp 1586364061
transform 1 0 30912 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_410
timestamp 1586364061
transform 1 0 38824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_422
timestamp 1586364061
transform 1 0 39928 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_434
timestamp 1586364061
transform 1 0 41032 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_446
timestamp 1586364061
transform 1 0 42136 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_459
timestamp 1586364061
transform 1 0 43332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_471
timestamp 1586364061
transform 1 0 44436 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_483
timestamp 1586364061
transform 1 0 45540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_495
timestamp 1586364061
transform 1 0 46644 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_507
timestamp 1586364061
transform 1 0 47748 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 48852 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_515
timestamp 1586364061
transform 1 0 48484 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_318
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_415
timestamp 1586364061
transform 1 0 39284 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_428
timestamp 1586364061
transform 1 0 40480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_440
timestamp 1586364061
transform 1 0 41584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_452
timestamp 1586364061
transform 1 0 42688 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_464
timestamp 1586364061
transform 1 0 43792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_476
timestamp 1586364061
transform 1 0 44896 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_489
timestamp 1586364061
transform 1 0 46092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_501
timestamp 1586364061
transform 1 0 47196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 48852 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_513
timestamp 1586364061
transform 1 0 48300 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_288
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_300
timestamp 1586364061
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_312
timestamp 1586364061
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_410
timestamp 1586364061
transform 1 0 38824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_422
timestamp 1586364061
transform 1 0 39928 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_434
timestamp 1586364061
transform 1 0 41032 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_446
timestamp 1586364061
transform 1 0 42136 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_459
timestamp 1586364061
transform 1 0 43332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_471
timestamp 1586364061
transform 1 0 44436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_483
timestamp 1586364061
transform 1 0 45540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_495
timestamp 1586364061
transform 1 0 46644 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_507
timestamp 1586364061
transform 1 0 47748 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 48852 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_515
timestamp 1586364061
transform 1 0 48484 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_281
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_293
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_342
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_415
timestamp 1586364061
transform 1 0 39284 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_428
timestamp 1586364061
transform 1 0 40480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_440
timestamp 1586364061
transform 1 0 41584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_452
timestamp 1586364061
transform 1 0 42688 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_464
timestamp 1586364061
transform 1 0 43792 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_476
timestamp 1586364061
transform 1 0 44896 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_489
timestamp 1586364061
transform 1 0 46092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_501
timestamp 1586364061
transform 1 0 47196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 48852 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_513
timestamp 1586364061
transform 1 0 48300 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_137
timestamp 1586364061
transform 1 0 13708 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_clkbuf_1_0_0_clk_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_155
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_167
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_188
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_192
timestamp 1586364061
transform 1 0 18768 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_216
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_228
timestamp 1586364061
transform 1 0 22080 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_288
timestamp 1586364061
transform 1 0 27600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_281
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_293
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_300
timestamp 1586364061
transform 1 0 28704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_330
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_379
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_410
timestamp 1586364061
transform 1 0 38824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_422
timestamp 1586364061
transform 1 0 39928 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_415
timestamp 1586364061
transform 1 0 39284 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_428
timestamp 1586364061
transform 1 0 40480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_434
timestamp 1586364061
transform 1 0 41032 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_446
timestamp 1586364061
transform 1 0 42136 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_440
timestamp 1586364061
transform 1 0 41584 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_452
timestamp 1586364061
transform 1 0 42688 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_459
timestamp 1586364061
transform 1 0 43332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_471
timestamp 1586364061
transform 1 0 44436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_483
timestamp 1586364061
transform 1 0 45540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_464
timestamp 1586364061
transform 1 0 43792 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_476
timestamp 1586364061
transform 1 0 44896 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_495
timestamp 1586364061
transform 1 0 46644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_507
timestamp 1586364061
transform 1 0 47748 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_489
timestamp 1586364061
transform 1 0 46092 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_501
timestamp 1586364061
transform 1 0 47196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 48852 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 48852 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_515
timestamp 1586364061
transform 1 0 48484 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_513
timestamp 1586364061
transform 1 0 48300 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 2430 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_clkbuf_1  clkbuf_1_0_0_clk tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 18124 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_183
timestamp 1586364061
transform 1 0 17940 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_187
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_191
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_195
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_207
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_300
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_373
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_410
timestamp 1586364061
transform 1 0 38824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_422
timestamp 1586364061
transform 1 0 39928 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_434
timestamp 1586364061
transform 1 0 41032 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_446
timestamp 1586364061
transform 1 0 42136 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_459
timestamp 1586364061
transform 1 0 43332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_471
timestamp 1586364061
transform 1 0 44436 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_483
timestamp 1586364061
transform 1 0 45540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_495
timestamp 1586364061
transform 1 0 46644 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_507
timestamp 1586364061
transform 1 0 47748 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 48852 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_515
timestamp 1586364061
transform 1 0 48484 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 2430 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__603__B
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_166
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__603__A
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_176
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_clkbuf_1  clkbuf_1_1_0_clk
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 2430 592
use scs8hd_decap_4  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_214
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_229
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_281
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_293
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_330
timestamp 1586364061
transform 1 0 31464 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_342
timestamp 1586364061
transform 1 0 32568 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_354
timestamp 1586364061
transform 1 0 33672 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_379
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_391
timestamp 1586364061
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 40388 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_403
timestamp 1586364061
transform 1 0 38180 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_415
timestamp 1586364061
transform 1 0 39284 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_428
timestamp 1586364061
transform 1 0 40480 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_440
timestamp 1586364061
transform 1 0 41584 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_452
timestamp 1586364061
transform 1 0 42688 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_464
timestamp 1586364061
transform 1 0 43792 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_476
timestamp 1586364061
transform 1 0 44896 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 46000 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_489
timestamp 1586364061
transform 1 0 46092 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_501
timestamp 1586364061
transform 1 0 47196 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 48852 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_513
timestamp 1586364061
transform 1 0 48300 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_160
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _603_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16192 0 -1 8160
box -38 -48 866 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 2430 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_176
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_218
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_222
timestamp 1586364061
transform 1 0 21528 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_234
timestamp 1586364061
transform 1 0 22632 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_246
timestamp 1586364061
transform 1 0 23736 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__377__B
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__373__B
timestamp 1586364061
transform 1 0 26680 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_273
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_280
timestamp 1586364061
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_292
timestamp 1586364061
transform 1 0 27968 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__366__A
timestamp 1586364061
transform 1 0 29256 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__366__B
timestamp 1586364061
transform 1 0 29624 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_304
timestamp 1586364061
transform 1 0 29072 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_308
timestamp 1586364061
transform 1 0 29440 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_312
timestamp 1586364061
transform 1 0 29808 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__326__A
timestamp 1586364061
transform 1 0 34684 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__329__A
timestamp 1586364061
transform 1 0 35052 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_349
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_361
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_367
timestamp 1586364061
transform 1 0 34868 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_371
timestamp 1586364061
transform 1 0 35236 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_383
timestamp 1586364061
transform 1 0 36340 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_10_395
timestamp 1586364061
transform 1 0 37444 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_410
timestamp 1586364061
transform 1 0 38824 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_422
timestamp 1586364061
transform 1 0 39928 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_434
timestamp 1586364061
transform 1 0 41032 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_446
timestamp 1586364061
transform 1 0 42136 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 43240 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_459
timestamp 1586364061
transform 1 0 43332 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_471
timestamp 1586364061
transform 1 0 44436 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_483
timestamp 1586364061
transform 1 0 45540 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_495
timestamp 1586364061
transform 1 0 46644 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_507
timestamp 1586364061
transform 1 0 47748 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 48852 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_515
timestamp 1586364061
transform 1 0 48484 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _610_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 866 592
use scs8hd_clkbuf_16  clkbuf_0_clk tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 1878 592
use scs8hd_diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__610__A
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_153
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_187
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_191
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__312__A
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_200
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__312__B
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_207
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_211
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_235
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_nor2_4  _377_
timestamp 1586364061
transform 1 0 26036 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__373__A
timestamp 1586364061
transform 1 0 27048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__377__A
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_280
timestamp 1586364061
transform 1 0 26864 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_284
timestamp 1586364061
transform 1 0 27232 0 1 8160
box -38 -48 1142 592
use scs8hd_nor2_4  _366_
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__361__A
timestamp 1586364061
transform 1 0 28704 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__361__B
timestamp 1586364061
transform 1 0 28336 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_298
timestamp 1586364061
transform 1 0 28520 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_302
timestamp 1586364061
transform 1 0 28888 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_315
timestamp 1586364061
transform 1 0 30084 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_327
timestamp 1586364061
transform 1 0 31188 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_339
timestamp 1586364061
transform 1 0 32292 0 1 8160
box -38 -48 1142 592
use scs8hd_nor2_4  _329_
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use scs8hd_conb_1  _655_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 33764 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__329__B
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__326__B
timestamp 1586364061
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_351
timestamp 1586364061
transform 1 0 33396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_358
timestamp 1586364061
transform 1 0 34040 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_362
timestamp 1586364061
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36524 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_11_384
timestamp 1586364061
transform 1 0 36432 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_387
timestamp 1586364061
transform 1 0 36708 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_399
timestamp 1586364061
transform 1 0 37812 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 40388 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_411
timestamp 1586364061
transform 1 0 38916 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_423
timestamp 1586364061
transform 1 0 40020 0 1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_11_428
timestamp 1586364061
transform 1 0 40480 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_440
timestamp 1586364061
transform 1 0 41584 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_452
timestamp 1586364061
transform 1 0 42688 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_464
timestamp 1586364061
transform 1 0 43792 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_476
timestamp 1586364061
transform 1 0 44896 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 46000 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_489
timestamp 1586364061
transform 1 0 46092 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_501
timestamp 1586364061
transform 1 0 47196 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 48852 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_513
timestamp 1586364061
transform 1 0 48300 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_101
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_4  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 406 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15732 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_157
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_161
timestamp 1586364061
transform 1 0 15916 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_171
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_183
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 774 592
use scs8hd_nor2_4  _312_
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_191
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_207
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_12_235
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_240
timestamp 1586364061
transform 1 0 23184 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24748 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_244
timestamp 1586364061
transform 1 0 23552 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_255
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_259
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_265
timestamp 1586364061
transform 1 0 25484 0 -1 9248
box -38 -48 774 592
use scs8hd_nor2_4  _373_
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_273
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_285
timestamp 1586364061
transform 1 0 27324 0 -1 9248
box -38 -48 1142 592
use scs8hd_nor2_4  _361_
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29716 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_297
timestamp 1586364061
transform 1 0 28428 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_309
timestamp 1586364061
transform 1 0 29532 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_313
timestamp 1586364061
transform 1 0 29900 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__323__B
timestamp 1586364061
transform 1 0 33028 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31004 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_327
timestamp 1586364061
transform 1 0 31188 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_335
timestamp 1586364061
transform 1 0 31924 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_345
timestamp 1586364061
transform 1 0 32844 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _326_
timestamp 1586364061
transform 1 0 34684 0 -1 9248
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33580 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_349
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_356
timestamp 1586364061
transform 1 0 33856 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_364
timestamp 1586364061
transform 1 0 34592 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_374
timestamp 1586364061
transform 1 0 35512 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36524 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35696 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36064 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_378
timestamp 1586364061
transform 1 0 35880 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_382
timestamp 1586364061
transform 1 0 36248 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_388
timestamp 1586364061
transform 1 0 36800 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_396
timestamp 1586364061
transform 1 0 37536 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 40480 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__350__B
timestamp 1586364061
transform 1 0 38824 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40112 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_412
timestamp 1586364061
transform 1 0 39008 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_426
timestamp 1586364061
transform 1 0 40296 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40848 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_430
timestamp 1586364061
transform 1 0 40664 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_434
timestamp 1586364061
transform 1 0 41032 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_446
timestamp 1586364061
transform 1 0 42136 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 43240 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_459
timestamp 1586364061
transform 1 0 43332 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_471
timestamp 1586364061
transform 1 0 44436 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_483
timestamp 1586364061
transform 1 0 45540 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_495
timestamp 1586364061
transform 1 0 46644 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_507
timestamp 1586364061
transform 1 0 47748 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 48852 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_515
timestamp 1586364061
transform 1 0 48484 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_286
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_287
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__550__B
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__550__A
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _550_
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_112
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__551__A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _551_
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_124
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_126
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__551__B
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_134
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_130
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__609__A
timestamp 1586364061
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_151
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__611__A
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_288
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_161
timestamp 1586364061
transform 1 0 15916 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_8  _611_
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_168
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_164
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_180
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_187
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_192
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_191
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_13_213
timestamp 1586364061
transform 1 0 20700 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_289
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_226
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_234
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_230
timestamp 1586364061
transform 1 0 22264 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 23000 0 -1 10336
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_14_249
timestamp 1586364061
transform 1 0 24012 0 -1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24748 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_266
timestamp 1586364061
transform 1 0 25576 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__371__A
timestamp 1586364061
transform 1 0 25760 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_270
timestamp 1586364061
transform 1 0 25944 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_278
timestamp 1586364061
transform 1 0 26680 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_274
timestamp 1586364061
transform 1 0 26312 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__370__A
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_290
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_288
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_284
timestamp 1586364061
transform 1 0 27232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__374__B
timestamp 1586364061
transform 1 0 27416 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__374__A
timestamp 1586364061
transform 1 0 26864 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__372__A
timestamp 1586364061
transform 1 0 26772 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _374_
timestamp 1586364061
transform 1 0 27048 0 1 9248
box -38 -48 866 592
use scs8hd_buf_1  _370_
timestamp 1586364061
transform 1 0 26956 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_295
timestamp 1586364061
transform 1 0 28244 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_291
timestamp 1586364061
transform 1 0 27876 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__362__A
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _362_
timestamp 1586364061
transform 1 0 27968 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_305
timestamp 1586364061
transform 1 0 29164 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_301
timestamp 1586364061
transform 1 0 28796 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_299
timestamp 1586364061
transform 1 0 28612 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__362__B
timestamp 1586364061
transform 1 0 28428 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 29256 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_14_308
timestamp 1586364061
transform 1 0 29440 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_317
timestamp 1586364061
transform 1 0 30268 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 29532 0 -1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_320
timestamp 1586364061
transform 1 0 30544 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_321
timestamp 1586364061
transform 1 0 30636 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30452 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30728 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_324
timestamp 1586364061
transform 1 0 30912 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 30820 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 31004 0 1 9248
box -38 -48 1050 592
use scs8hd_conb_1  _653_
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_291
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_340
timestamp 1586364061
transform 1 0 32384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__323__A
timestamp 1586364061
transform 1 0 32844 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32568 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32936 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_344
timestamp 1586364061
transform 1 0 32752 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_344
timestamp 1586364061
transform 1 0 32752 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _323_
timestamp 1586364061
transform 1 0 33028 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_13_336
timestamp 1586364061
transform 1 0 32016 0 1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_348
timestamp 1586364061
transform 1 0 33120 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_360
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_356
timestamp 1586364061
transform 1 0 33856 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 33488 0 -1 10336
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_14_369
timestamp 1586364061
transform 1 0 35052 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_4  FILLER_14_363
timestamp 1586364061
transform 1 0 34500 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_364
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 35236 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_375
timestamp 1586364061
transform 1 0 35604 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_373
timestamp 1586364061
transform 1 0 35420 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 35604 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_387
timestamp 1586364061
transform 1 0 36708 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 35788 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 35696 0 -1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_395
timestamp 1586364061
transform 1 0 37444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_391
timestamp 1586364061
transform 1 0 37076 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_396
timestamp 1586364061
transform 1 0 37536 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_388
timestamp 1586364061
transform 1 0 36800 0 1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37260 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36892 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37720 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_292
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_400
timestamp 1586364061
transform 1 0 37904 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38088 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_412
timestamp 1586364061
transform 1 0 39008 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_407
timestamp 1586364061
transform 1 0 38548 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_404
timestamp 1586364061
transform 1 0 38272 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__349__B
timestamp 1586364061
transform 1 0 38824 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__350__A
timestamp 1586364061
transform 1 0 38640 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _350_
timestamp 1586364061
transform 1 0 38824 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_423
timestamp 1586364061
transform 1 0 40020 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_417
timestamp 1586364061
transform 1 0 39468 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_426
timestamp 1586364061
transform 1 0 40296 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_423
timestamp 1586364061
transform 1 0 40020 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_419
timestamp 1586364061
transform 1 0 39652 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__354__B
timestamp 1586364061
transform 1 0 39284 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 40112 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 40112 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 40388 0 1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 40480 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41952 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41308 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_439
timestamp 1586364061
transform 1 0 41492 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_451
timestamp 1586364061
transform 1 0 42596 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_435
timestamp 1586364061
transform 1 0 41124 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_439
timestamp 1586364061
transform 1 0 41492 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_443
timestamp 1586364061
transform 1 0 41860 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_446
timestamp 1586364061
transform 1 0 42136 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_293
timestamp 1586364061
transform 1 0 43240 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_463
timestamp 1586364061
transform 1 0 43700 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_475
timestamp 1586364061
transform 1 0 44804 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_459
timestamp 1586364061
transform 1 0 43332 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_471
timestamp 1586364061
transform 1 0 44436 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_483
timestamp 1586364061
transform 1 0 45540 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 46000 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_487
timestamp 1586364061
transform 1 0 45908 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_489
timestamp 1586364061
transform 1 0 46092 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_501
timestamp 1586364061
transform 1 0 47196 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_495
timestamp 1586364061
transform 1 0 46644 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_507
timestamp 1586364061
transform 1 0 47748 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 48852 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 48852 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_513
timestamp 1586364061
transform 1 0 48300 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_515
timestamp 1586364061
transform 1 0 48484 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_294
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_conb_1  _639_
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__549__A
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__549__B
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_295
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_130
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _609_
timestamp 1586364061
transform 1 0 13156 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__602__A
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__602__B
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_140
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_146
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_296
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_187
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _310_
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__311__A
timestamp 1586364061
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__310__A
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__311__B
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_192
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_207
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_211
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_223
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_219
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_215
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__309__A
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _636_
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 866 592
use scs8hd_fill_1  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_252
timestamp 1586364061
transform 1 0 24288 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_248
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_243
timestamp 1586364061
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_297
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_256
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 1050 592
use scs8hd_nor2_4  _372_
timestamp 1586364061
transform 1 0 26772 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__372__B
timestamp 1586364061
transform 1 0 27784 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28152 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_271
timestamp 1586364061
transform 1 0 26036 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_278
timestamp 1586364061
transform 1 0 26680 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_288
timestamp 1586364061
transform 1 0 27600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_292
timestamp 1586364061
transform 1 0 27968 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_302
timestamp 1586364061
transform 1 0 28888 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_296
timestamp 1586364061
transform 1 0 28336 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28704 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_298
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_313
timestamp 1586364061
transform 1 0 29900 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29440 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29624 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_317
timestamp 1586364061
transform 1 0 30268 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30084 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30636 0 1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32200 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32016 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31648 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_334
timestamp 1586364061
transform 1 0 31832 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_347
timestamp 1586364061
transform 1 0 33028 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_358
timestamp 1586364061
transform 1 0 34040 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_351
timestamp 1586364061
transform 1 0 33396 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33212 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 33580 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_362
timestamp 1586364061
transform 1 0 34408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_299
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36708 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37720 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36064 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36524 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38088 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_376
timestamp 1586364061
transform 1 0 35696 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_15_382
timestamp 1586364061
transform 1 0 36248 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_396
timestamp 1586364061
transform 1 0 37536 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_400
timestamp 1586364061
transform 1 0 37904 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _349_
timestamp 1586364061
transform 1 0 38824 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_300
timestamp 1586364061
transform 1 0 40388 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__349__A
timestamp 1586364061
transform 1 0 38640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__354__A
timestamp 1586364061
transform 1 0 39836 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40204 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_404
timestamp 1586364061
transform 1 0 38272 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_419
timestamp 1586364061
transform 1 0 39652 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_423
timestamp 1586364061
transform 1 0 40020 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 41952 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 41768 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41216 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_431
timestamp 1586364061
transform 1 0 40756 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_435
timestamp 1586364061
transform 1 0 41124 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_438
timestamp 1586364061
transform 1 0 41400 0 1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_15_455
timestamp 1586364061
transform 1 0 42964 0 1 10336
box -38 -48 406 592
use scs8hd_conb_1  _654_
timestamp 1586364061
transform 1 0 43700 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43332 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44160 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_461
timestamp 1586364061
transform 1 0 43516 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_466
timestamp 1586364061
transform 1 0 43976 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_470
timestamp 1586364061
transform 1 0 44344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_15_482
timestamp 1586364061
transform 1 0 45448 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_301
timestamp 1586364061
transform 1 0 46000 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_489
timestamp 1586364061
transform 1 0 46092 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_501
timestamp 1586364061
transform 1 0 47196 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 48852 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_513
timestamp 1586364061
transform 1 0 48300 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_302
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_nor2_4  _549_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_303
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_119
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_127
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _602_
timestamp 1586364061
transform 1 0 15364 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_304
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_164
timestamp 1586364061
transform 1 0 16192 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_181
timestamp 1586364061
transform 1 0 17756 0 -1 11424
box -38 -48 1142 592
use scs8hd_nor2_4  _311_
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_305
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__310__B
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_203
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_207
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_218
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_1  _309_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_233
timestamp 1586364061
transform 1 0 22540 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_229
timestamp 1586364061
transform 1 0 22172 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_226
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use scs8hd_conb_1  _652_
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 866 592
use scs8hd_buf_1  _371_
timestamp 1586364061
transform 1 0 25392 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25024 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_250
timestamp 1586364061
transform 1 0 24104 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_254
timestamp 1586364061
transform 1 0 24472 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_258
timestamp 1586364061
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_262
timestamp 1586364061
transform 1 0 25208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_267
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_306
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__375__B
timestamp 1586364061
transform 1 0 26220 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_287
timestamp 1586364061
transform 1 0 27508 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28704 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29164 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29532 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30728 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_299
timestamp 1586364061
transform 1 0 28612 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_303
timestamp 1586364061
transform 1 0 28980 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_307
timestamp 1586364061
transform 1 0 29348 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_320
timestamp 1586364061
transform 1 0 30544 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_307
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_324
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_346
timestamp 1586364061
transform 1 0 32936 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 33672 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__338__A
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35236 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_351
timestamp 1586364061
transform 1 0 33396 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_16_365
timestamp 1586364061
transform 1 0 34684 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_6  FILLER_16_373
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_308
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37076 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_379
timestamp 1586364061
transform 1 0 35972 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_393
timestamp 1586364061
transform 1 0 37260 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _354_
timestamp 1586364061
transform 1 0 39284 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__351__B
timestamp 1586364061
transform 1 0 38824 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_407
timestamp 1586364061
transform 1 0 38548 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_412
timestamp 1586364061
transform 1 0 39008 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_424
timestamp 1586364061
transform 1 0 40112 0 -1 11424
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41216 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_445
timestamp 1586364061
transform 1 0 42044 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_453
timestamp 1586364061
transform 1 0 42780 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_309
timestamp 1586364061
transform 1 0 43240 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_457
timestamp 1586364061
transform 1 0 43148 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_468
timestamp 1586364061
transform 1 0 44160 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_480
timestamp 1586364061
transform 1 0 45264 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_492
timestamp 1586364061
transform 1 0 46368 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_504
timestamp 1586364061
transform 1 0 47472 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 48852 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_310
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_70
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_78
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 314 592
use scs8hd_buf_1  _548_
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_83
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_109
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__548__A
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_311
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _608_
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__607__A
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__608__A
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_148
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_312
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_165
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_190
timestamp 1586364061
transform 1 0 18584 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_194
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_198
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_213
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _638_
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_224
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_239
timestamp 1586364061
transform 1 0 23092 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_235
timestamp 1586364061
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23276 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_313
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_243
timestamp 1586364061
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_261
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _363_
timestamp 1586364061
transform 1 0 27600 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__363__A
timestamp 1586364061
transform 1 0 27416 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__375__A
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__363__B
timestamp 1586364061
transform 1 0 27048 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_274
timestamp 1586364061
transform 1 0 26312 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_278
timestamp 1586364061
transform 1 0 26680 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_284
timestamp 1586364061
transform 1 0 27232 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_314
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_297
timestamp 1586364061
transform 1 0 28428 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_301
timestamp 1586364061
transform 1 0 28796 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_317
timestamp 1586364061
transform 1 0 30268 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_321
timestamp 1586364061
transform 1 0 30636 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_325
timestamp 1586364061
transform 1 0 31004 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30820 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_331
timestamp 1586364061
transform 1 0 31556 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_335
timestamp 1586364061
transform 1 0 31924 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_339
timestamp 1586364061
transform 1 0 32292 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32476 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32108 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_343
timestamp 1586364061
transform 1 0 32660 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__338__B
timestamp 1586364061
transform 1 0 33028 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _338_
timestamp 1586364061
transform 1 0 33212 0 1 11424
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 35236 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_315
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 35052 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34224 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_358
timestamp 1586364061
transform 1 0 34040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_362
timestamp 1586364061
transform 1 0 34408 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36984 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36616 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37996 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_382
timestamp 1586364061
transform 1 0 36248 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_388
timestamp 1586364061
transform 1 0 36800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_399
timestamp 1586364061
transform 1 0 37812 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_407
timestamp 1586364061
transform 1 0 38548 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__351__A
timestamp 1586364061
transform 1 0 38640 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _351_
timestamp 1586364061
transform 1 0 38824 0 1 11424
box -38 -48 866 592
use scs8hd_fill_2  FILLER_17_419
timestamp 1586364061
transform 1 0 39652 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_428
timestamp 1586364061
transform 1 0 40480 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_423
timestamp 1586364061
transform 1 0 40020 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40204 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_316
timestamp 1586364061
transform 1 0 40388 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42964 0 1 11424
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41216 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42780 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42228 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41032 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40664 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_432
timestamp 1586364061
transform 1 0 40848 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_445
timestamp 1586364061
transform 1 0 42044 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_449
timestamp 1586364061
transform 1 0 42412 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44528 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44988 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43976 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_464
timestamp 1586364061
transform 1 0 43792 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_468
timestamp 1586364061
transform 1 0 44160 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_475
timestamp 1586364061
transform 1 0 44804 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_479
timestamp 1586364061
transform 1 0 45172 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_317
timestamp 1586364061
transform 1 0 46000 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_487
timestamp 1586364061
transform 1 0 45908 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_489
timestamp 1586364061
transform 1 0 46092 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_501
timestamp 1586364061
transform 1 0 47196 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 48852 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_513
timestamp 1586364061
transform 1 0 48300 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_318
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_54
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_319
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_18_114
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_118
timestamp 1586364061
transform 1 0 11960 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_8  _607_
timestamp 1586364061
transform 1 0 15364 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_320
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_147
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__601__B
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_164
timestamp 1586364061
transform 1 0 16192 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_168
timestamp 1586364061
transform 1 0 16560 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_180
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_321
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22908 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_236
timestamp 1586364061
transform 1 0 22816 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25760 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_250
timestamp 1586364061
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_254
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_265
timestamp 1586364061
transform 1 0 25484 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _375_
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_322
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__364__B
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_270
timestamp 1586364061
transform 1 0 25944 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_285
timestamp 1586364061
transform 1 0 27324 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_290
timestamp 1586364061
transform 1 0 27784 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 28612 0 -1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30360 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_298
timestamp 1586364061
transform 1 0 28520 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_310
timestamp 1586364061
transform 1 0 29624 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_314
timestamp 1586364061
transform 1 0 29992 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_323
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31464 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_327
timestamp 1586364061
transform 1 0 31188 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_332
timestamp 1586364061
transform 1 0 31648 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_346
timestamp 1586364061
transform 1 0 32936 0 -1 12512
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__332__A
timestamp 1586364061
transform 1 0 35236 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_358
timestamp 1586364061
transform 1 0 34040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_369
timestamp 1586364061
transform 1 0 35052 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_4  FILLER_18_382
timestamp 1586364061
transform 1 0 36248 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_379
timestamp 1586364061
transform 1 0 35972 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36064 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_393
timestamp 1586364061
transform 1 0 37260 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_389
timestamp 1586364061
transform 1 0 36892 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36616 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_401
timestamp 1586364061
transform 1 0 37996 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_324
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 39652 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__352__B
timestamp 1586364061
transform 1 0 38824 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_409
timestamp 1586364061
transform 1 0 38732 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_412
timestamp 1586364061
transform 1 0 39008 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_418
timestamp 1586364061
transform 1 0 39560 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41400 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40848 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41216 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_430
timestamp 1586364061
transform 1 0 40664 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_434
timestamp 1586364061
transform 1 0 41032 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_447
timestamp 1586364061
transform 1 0 42228 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_455
timestamp 1586364061
transform 1 0 42964 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_325
timestamp 1586364061
transform 1 0 43240 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_468
timestamp 1586364061
transform 1 0 44160 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_480
timestamp 1586364061
transform 1 0 45264 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_492
timestamp 1586364061
transform 1 0 46368 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_504
timestamp 1586364061
transform 1 0 47472 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 48852 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_37
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 4508 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_334
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_50
timestamp 1586364061
transform 1 0 5704 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_19_45
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_41
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 4692 0 -1 13600
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_58
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_326
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_72
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_76
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_89
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_100
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_96
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__306__A
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_335
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 866 592
use scs8hd_buf_1  _306_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_103
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_106
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_327
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_134
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_151
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__606__A
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_336
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_8  _606_
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_158
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_171
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_162
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__601__A
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _601_
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_176
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_328
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1050 592
use scs8hd_conb_1  _637_
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_191
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__575__A
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__576__A
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _575_
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__575__B
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_337
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_225
timestamp 1586364061
transform 1 0 21804 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_226
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_222
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_218
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_237
timestamp 1586364061
transform 1 0 22908 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23184 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_253
timestamp 1586364061
transform 1 0 24380 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_329
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_264
timestamp 1586364061
transform 1 0 25392 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_260
timestamp 1586364061
transform 1 0 25024 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_265
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 590 592
use scs8hd_decap_3  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24748 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 1050 592
use scs8hd_nor2_4  _364_
timestamp 1586364061
transform 1 0 27600 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_338
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__364__A
timestamp 1586364061
transform 1 0 27416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_279
timestamp 1586364061
transform 1 0 26772 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_283
timestamp 1586364061
transform 1 0 27140 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_272
timestamp 1586364061
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_287
timestamp 1586364061
transform 1 0 27508 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_303
timestamp 1586364061
transform 1 0 28980 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_299
timestamp 1586364061
transform 1 0 28612 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_302
timestamp 1586364061
transform 1 0 28888 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_297
timestamp 1586364061
transform 1 0 28428 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29164 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28704 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_330
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28704 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_307
timestamp 1586364061
transform 1 0 29348 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29532 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29532 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29992 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_317
timestamp 1586364061
transform 1 0 30268 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_322
timestamp 1586364061
transform 1 0 30728 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30544 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_328
timestamp 1586364061
transform 1 0 31280 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_327
timestamp 1586364061
transform 1 0 31188 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31464 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31004 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_332
timestamp 1586364061
transform 1 0 31648 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_339
timestamp 1586364061
transform 1 0 32292 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32476 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_339
timestamp 1586364061
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_346
timestamp 1586364061
transform 1 0 32936 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_347
timestamp 1586364061
transform 1 0 33028 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_343
timestamp 1586364061
transform 1 0 32660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32844 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_350
timestamp 1586364061
transform 1 0 33304 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_358
timestamp 1586364061
transform 1 0 34040 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__335__A
timestamp 1586364061
transform 1 0 33580 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _335_
timestamp 1586364061
transform 1 0 33856 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_365
timestamp 1586364061
transform 1 0 34684 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_362
timestamp 1586364061
transform 1 0 34408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__332__B
timestamp 1586364061
transform 1 0 34868 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__335__B
timestamp 1586364061
transform 1 0 34592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_331
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _332_
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_369
timestamp 1586364061
transform 1 0 35052 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35236 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_379
timestamp 1586364061
transform 1 0 35972 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_382
timestamp 1586364061
transform 1 0 36248 0 1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_376
timestamp 1586364061
transform 1 0 35696 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36064 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_393
timestamp 1586364061
transform 1 0 37260 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_389
timestamp 1586364061
transform 1 0 36892 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36616 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36800 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_401
timestamp 1586364061
transform 1 0 37996 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_401
timestamp 1586364061
transform 1 0 37996 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_397
timestamp 1586364061
transform 1 0 37628 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37812 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_340
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_405
timestamp 1586364061
transform 1 0 38364 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_19_407
timestamp 1586364061
transform 1 0 38548 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__352__A
timestamp 1586364061
transform 1 0 38640 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _352_
timestamp 1586364061
transform 1 0 38824 0 1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_417
timestamp 1586364061
transform 1 0 39468 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_428
timestamp 1586364061
transform 1 0 40480 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_423
timestamp 1586364061
transform 1 0 40020 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_419
timestamp 1586364061
transform 1 0 39652 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_332
timestamp 1586364061
transform 1 0 40388 0 1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 39560 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_20_429
timestamp 1586364061
transform 1 0 40572 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_437
timestamp 1586364061
transform 1 0 41308 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_433
timestamp 1586364061
transform 1 0 40940 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40756 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40756 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41400 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_447
timestamp 1586364061
transform 1 0 42228 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_6  FILLER_19_448
timestamp 1586364061
transform 1 0 42320 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_444
timestamp 1586364061
transform 1 0 41952 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_440
timestamp 1586364061
transform 1 0 41584 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42136 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41768 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_455
timestamp 1586364061
transform 1 0 42964 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42872 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43056 0 1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_20_462
timestamp 1586364061
transform 1 0 43608 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_469
timestamp 1586364061
transform 1 0 44252 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_465
timestamp 1586364061
transform 1 0 43884 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44068 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_341
timestamp 1586364061
transform 1 0 43240 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_474
timestamp 1586364061
transform 1 0 44712 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_480
timestamp 1586364061
transform 1 0 45264 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_476
timestamp 1586364061
transform 1 0 44896 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45080 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44620 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_333
timestamp 1586364061
transform 1 0 46000 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_489
timestamp 1586364061
transform 1 0 46092 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_501
timestamp 1586364061
transform 1 0 47196 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_486
timestamp 1586364061
transform 1 0 45816 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_498
timestamp 1586364061
transform 1 0 46920 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 48852 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 48852 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_513
timestamp 1586364061
transform 1 0 48300 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_510
timestamp 1586364061
transform 1 0 48024 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_29
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_33
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_48
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_54
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_342
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_88
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_106
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_343
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_130
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_126
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_137
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_141
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_158
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _605_
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_344
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__605__A
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__604__A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_162
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_190
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__577__B
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__577__A
timestamp 1586364061
transform 1 0 18768 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _577_
timestamp 1586364061
transform 1 0 18952 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_207
timestamp 1586364061
transform 1 0 20148 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_203
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__576__B
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_214
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_218
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_225
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_229
timestamp 1586364061
transform 1 0 22172 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_345
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_252
timestamp 1586364061
transform 1 0 24288 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_256
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_273
timestamp 1586364061
transform 1 0 26220 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__376__A
timestamp 1586364061
transform 1 0 26036 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _376_
timestamp 1586364061
transform 1 0 26588 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_286
timestamp 1586364061
transform 1 0 27416 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__365__A
timestamp 1586364061
transform 1 0 27600 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_290
timestamp 1586364061
transform 1 0 27784 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__365__B
timestamp 1586364061
transform 1 0 27968 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_301
timestamp 1586364061
transform 1 0 28796 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_297
timestamp 1586364061
transform 1 0 28428 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_346
timestamp 1586364061
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_319
timestamp 1586364061
transform 1 0 30452 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_315
timestamp 1586364061
transform 1 0 30084 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30636 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30268 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31464 0 1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33028 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31004 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_323
timestamp 1586364061
transform 1 0 30820 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_327
timestamp 1586364061
transform 1 0 31188 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_339
timestamp 1586364061
transform 1 0 32292 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_343
timestamp 1586364061
transform 1 0 32660 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 34868 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_347
timestamp 1586364061
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 34592 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_356
timestamp 1586364061
transform 1 0 33856 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_362
timestamp 1586364061
transform 1 0 34408 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36616 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36064 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36432 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37996 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37628 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_378
timestamp 1586364061
transform 1 0 35880 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_382
timestamp 1586364061
transform 1 0 36248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_395
timestamp 1586364061
transform 1 0 37444 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_399
timestamp 1586364061
transform 1 0 37812 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_412
timestamp 1586364061
transform 1 0 39008 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38180 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_420
timestamp 1586364061
transform 1 0 39744 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_416
timestamp 1586364061
transform 1 0 39376 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39928 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39192 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 39560 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_424
timestamp 1586364061
transform 1 0 40112 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_348
timestamp 1586364061
transform 1 0 40388 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_435
timestamp 1586364061
transform 1 0 41124 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_431
timestamp 1586364061
transform 1 0 40756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41308 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41492 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_448
timestamp 1586364061
transform 1 0 42320 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_452
timestamp 1586364061
transform 1 0 42688 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42872 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42504 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43056 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43516 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43884 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_459
timestamp 1586364061
transform 1 0 43332 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_463
timestamp 1586364061
transform 1 0 43700 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_467
timestamp 1586364061
transform 1 0 44068 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_479
timestamp 1586364061
transform 1 0 45172 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_349
timestamp 1586364061
transform 1 0 46000 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_487
timestamp 1586364061
transform 1 0 45908 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_489
timestamp 1586364061
transform 1 0 46092 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_501
timestamp 1586364061
transform 1 0 47196 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 48852 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_513
timestamp 1586364061
transform 1 0 48300 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_350
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_47
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  FILLER_22_59
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_351
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_86
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_4  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_99
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_118
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_352
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_157
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_161
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_8  _604_
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__600__A
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_167
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_180
timestamp 1586364061
transform 1 0 17664 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _576_
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_353
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_194
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_204
timestamp 1586364061
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_208
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_232
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24840 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_243
timestamp 1586364061
transform 1 0 23460 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_4  FILLER_22_253
timestamp 1586364061
transform 1 0 24380 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_257
timestamp 1586364061
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_261
timestamp 1586364061
transform 1 0 25116 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_265
timestamp 1586364061
transform 1 0 25484 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _365_
timestamp 1586364061
transform 1 0 27508 0 -1 14688
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_354
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__376__B
timestamp 1586364061
transform 1 0 26956 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27324 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_273
timestamp 1586364061
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_279
timestamp 1586364061
transform 1 0 26772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_283
timestamp 1586364061
transform 1 0 27140 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29072 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_296
timestamp 1586364061
transform 1 0 28336 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_313
timestamp 1586364061
transform 1 0 29900 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 14688
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_355
timestamp 1586364061
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31464 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_328
timestamp 1586364061
transform 1 0 31280 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_332
timestamp 1586364061
transform 1 0 31648 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_346
timestamp 1586364061
transform 1 0 32936 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34224 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35236 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_369
timestamp 1586364061
transform 1 0 35052 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_373
timestamp 1586364061
transform 1 0 35420 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_356
timestamp 1586364061
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_379
timestamp 1586364061
transform 1 0 35972 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_389
timestamp 1586364061
transform 1 0 36892 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_398
timestamp 1586364061
transform 1 0 37720 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 39560 0 -1 14688
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38548 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__353__B
timestamp 1586364061
transform 1 0 39008 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_406
timestamp 1586364061
transform 1 0 38456 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_410
timestamp 1586364061
transform 1 0 38824 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_414
timestamp 1586364061
transform 1 0 39192 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_429
timestamp 1586364061
transform 1 0 40572 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41492 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40848 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41308 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_434
timestamp 1586364061
transform 1 0 41032 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_448
timestamp 1586364061
transform 1 0 42320 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_456
timestamp 1586364061
transform 1 0 43056 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_357
timestamp 1586364061
transform 1 0 43240 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43792 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_462
timestamp 1586364061
transform 1 0 43608 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_466
timestamp 1586364061
transform 1 0 43976 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_478
timestamp 1586364061
transform 1 0 45080 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_490
timestamp 1586364061
transform 1 0 46184 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_502
timestamp 1586364061
transform 1 0 47288 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 48852 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_514
timestamp 1586364061
transform 1 0 48392 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__534__B
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__534__A
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_28
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_47
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_55
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_65
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_358
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_23_69
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 590 592
use scs8hd_decap_3  FILLER_23_78
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_96
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_100
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_359
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_140
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_23_157
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_161
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _600_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_360
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__547__B
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_187
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__573__A
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__547__A
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__573__B
timestamp 1586364061
transform 1 0 18952 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_191
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_200
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_215
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 774 592
use scs8hd_decap_4  FILLER_23_225
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_234
timestamp 1586364061
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_238
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_248
timestamp 1586364061
transform 1 0 23920 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_242
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_361
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_256
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_252
timestamp 1586364061
transform 1 0 24288 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26680 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26128 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27692 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28244 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_270
timestamp 1586364061
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_274
timestamp 1586364061
transform 1 0 26312 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_287
timestamp 1586364061
transform 1 0 27508 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_291
timestamp 1586364061
transform 1 0 27876 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29256 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_362
timestamp 1586364061
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30452 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_297
timestamp 1586364061
transform 1 0 28428 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_301
timestamp 1586364061
transform 1 0 28796 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_317
timestamp 1586364061
transform 1 0 30268 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_321
timestamp 1586364061
transform 1 0 30636 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31004 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_327
timestamp 1586364061
transform 1 0 31188 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31372 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_332
timestamp 1586364061
transform 1 0 31648 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_336
timestamp 1586364061
transform 1 0 32016 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31832 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32200 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32384 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_343
timestamp 1586364061
transform 1 0 32660 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_347
timestamp 1586364061
transform 1 0 33028 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _322_
timestamp 1586364061
transform 1 0 33396 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_363
timestamp 1586364061
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34132 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__322__A
timestamp 1586364061
transform 1 0 33212 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_354
timestamp 1586364061
transform 1 0 33672 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_358
timestamp 1586364061
transform 1 0 34040 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_361
timestamp 1586364061
transform 1 0 34316 0 1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_383
timestamp 1586364061
transform 1 0 36340 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_380
timestamp 1586364061
transform 1 0 36064 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_376
timestamp 1586364061
transform 1 0 35696 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36156 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_23_393
timestamp 1586364061
transform 1 0 37260 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_401
timestamp 1586364061
transform 1 0 37996 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_397
timestamp 1586364061
transform 1 0 37628 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__355__B
timestamp 1586364061
transform 1 0 37812 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_405
timestamp 1586364061
transform 1 0 38364 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__355__A
timestamp 1586364061
transform 1 0 38180 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__353__A
timestamp 1586364061
transform 1 0 38548 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _353_
timestamp 1586364061
transform 1 0 38732 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  FILLER_23_418
timestamp 1586364061
transform 1 0 39560 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__348__A
timestamp 1586364061
transform 1 0 39836 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_423
timestamp 1586364061
transform 1 0 40020 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_364
timestamp 1586364061
transform 1 0 40388 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 14688
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42044 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42504 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42872 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41492 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_437
timestamp 1586364061
transform 1 0 41308 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_441
timestamp 1586364061
transform 1 0 41676 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_448
timestamp 1586364061
transform 1 0 42320 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_452
timestamp 1586364061
transform 1 0 42688 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_456
timestamp 1586364061
transform 1 0 43056 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44988 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43424 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45448 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44804 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43240 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44436 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_469
timestamp 1586364061
transform 1 0 44252 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_473
timestamp 1586364061
transform 1 0 44620 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_480
timestamp 1586364061
transform 1 0 45264 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_365
timestamp 1586364061
transform 1 0 46000 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_484
timestamp 1586364061
transform 1 0 45632 0 1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_23_489
timestamp 1586364061
transform 1 0 46092 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_501
timestamp 1586364061
transform 1 0 47196 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 48852 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_513
timestamp 1586364061
transform 1 0 48300 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_nor2_4  _534_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_366
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_45
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_73
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_79
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_367
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_85
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_114
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_118
timestamp 1586364061
transform 1 0 11960 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_122
timestamp 1586364061
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_368
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_4  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_158
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use scs8hd_or2_4  _547_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 682 592
use scs8hd_decap_12  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_24_180
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 314 592
use scs8hd_or2_4  _573_
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_369
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__308__A
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_194
timestamp 1586364061
transform 1 0 18952 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_205
timestamp 1586364061
transform 1 0 19964 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_213
timestamp 1586364061
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21620 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_6  FILLER_24_226
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25208 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_243
timestamp 1586364061
transform 1 0 23460 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_247
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_260
timestamp 1586364061
transform 1 0 25024 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_264
timestamp 1586364061
transform 1 0 25392 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_370
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25944 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_272
timestamp 1586364061
transform 1 0 26128 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_287
timestamp 1586364061
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29072 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__360__A
timestamp 1586364061
transform 1 0 28796 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_299
timestamp 1586364061
transform 1 0 28612 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_303
timestamp 1586364061
transform 1 0 28980 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_313
timestamp 1586364061
transform 1 0 29900 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_371
timestamp 1586364061
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_328
timestamp 1586364061
transform 1 0 31280 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_3  FILLER_24_346
timestamp 1586364061
transform 1 0 32936 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34132 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35144 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__341__A
timestamp 1586364061
transform 1 0 33212 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34868 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_351
timestamp 1586364061
transform 1 0 33396 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_4  FILLER_24_362
timestamp 1586364061
transform 1 0 34408 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_366
timestamp 1586364061
transform 1 0 34776 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_369
timestamp 1586364061
transform 1 0 35052 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_373
timestamp 1586364061
transform 1 0 35420 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36156 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_384
timestamp 1586364061
transform 1 0 36432 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36616 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_388
timestamp 1586364061
transform 1 0 36800 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36984 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_392
timestamp 1586364061
transform 1 0 37168 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_398
timestamp 1586364061
transform 1 0 37720 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_372
timestamp 1586364061
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_402
timestamp 1586364061
transform 1 0 38088 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37904 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  _348_
timestamp 1586364061
transform 1 0 39836 0 -1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _355_
timestamp 1586364061
transform 1 0 38272 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40480 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_413
timestamp 1586364061
transform 1 0 39100 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_4  FILLER_24_424
timestamp 1586364061
transform 1 0 40112 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40848 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 42228 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_430
timestamp 1586364061
transform 1 0 40664 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_441
timestamp 1586364061
transform 1 0 41676 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_6  FILLER_24_449
timestamp 1586364061
transform 1 0 42412 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_455
timestamp 1586364061
transform 1 0 42964 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44896 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_373
timestamp 1586364061
transform 1 0 43240 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_468
timestamp 1586364061
transform 1 0 44160 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_472
timestamp 1586364061
transform 1 0 44528 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_479
timestamp 1586364061
transform 1 0 45172 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_491
timestamp 1586364061
transform 1 0 46276 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_503
timestamp 1586364061
transform 1 0 47380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 48852 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_515
timestamp 1586364061
transform 1 0 48484 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__535__A
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__535__B
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_16
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_20
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__531__A
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__533__A
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__531__B
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_30
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_50
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_374
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__533__B
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_54
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_58
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_81
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_88
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_103
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_107
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_375
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_139
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_154
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 1142 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_376
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__527__A
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__307__A
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__527__B
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_or2_4  _308_
timestamp 1586364061
transform 1 0 18768 0 1 15776
box -38 -48 682 592
use scs8hd_buf_1  _574_
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__308__B
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__574__A
timestamp 1586364061
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_189
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_199
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_203
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__619__A
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_218
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_224
timestamp 1586364061
transform 1 0 21712 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_377
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_254
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_266
timestamp 1586364061
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__379__A
timestamp 1586364061
transform 1 0 27140 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__379__B
timestamp 1586364061
transform 1 0 27508 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_281
timestamp 1586364061
transform 1 0 26956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_285
timestamp 1586364061
transform 1 0 27324 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_289
timestamp 1586364061
transform 1 0 27692 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_293
timestamp 1586364061
transform 1 0 28060 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_301
timestamp 1586364061
transform 1 0 28796 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_297
timestamp 1586364061
transform 1 0 28428 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__368__A
timestamp 1586364061
transform 1 0 28980 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_378
timestamp 1586364061
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _368_
timestamp 1586364061
transform 1 0 29256 0 1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_25_319
timestamp 1586364061
transform 1 0 30452 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_315
timestamp 1586364061
transform 1 0 30084 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30636 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31372 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__341__B
timestamp 1586364061
transform 1 0 33028 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31188 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32384 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_323
timestamp 1586364061
transform 1 0 30820 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_338
timestamp 1586364061
transform 1 0 32200 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_342
timestamp 1586364061
transform 1 0 32568 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_346
timestamp 1586364061
transform 1 0 32936 0 1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _341_
timestamp 1586364061
transform 1 0 33212 0 1 15776
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_379
timestamp 1586364061
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 34224 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35236 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_358
timestamp 1586364061
transform 1 0 34040 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_362
timestamp 1586364061
transform 1 0 34408 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_367
timestamp 1586364061
transform 1 0 34868 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_380
timestamp 1586364061
transform 1 0 36064 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_376
timestamp 1586364061
transform 1 0 35696 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36248 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_25_393
timestamp 1586364061
transform 1 0 37260 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37444 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_401
timestamp 1586364061
transform 1 0 37996 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_397
timestamp 1586364061
transform 1 0 37628 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38088 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 38640 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_380
timestamp 1586364061
transform 1 0 40388 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 38456 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__347__A
timestamp 1586364061
transform 1 0 39836 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_404
timestamp 1586364061
transform 1 0 38272 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_419
timestamp 1586364061
transform 1 0 39652 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_423
timestamp 1586364061
transform 1 0 40020 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_428
timestamp 1586364061
transform 1 0 40480 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 42228 0 1 15776
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40664 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 42044 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_439
timestamp 1586364061
transform 1 0 41492 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_443
timestamp 1586364061
transform 1 0 41860 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43976 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44988 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43792 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43424 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_458
timestamp 1586364061
transform 1 0 43240 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_462
timestamp 1586364061
transform 1 0 43608 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_475
timestamp 1586364061
transform 1 0 44804 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_479
timestamp 1586364061
transform 1 0 45172 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_381
timestamp 1586364061
transform 1 0 46000 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_487
timestamp 1586364061
transform 1 0 45908 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_489
timestamp 1586364061
transform 1 0 46092 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_501
timestamp 1586364061
transform 1 0 47196 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 48852 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_513
timestamp 1586364061
transform 1 0 48300 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_26_11
timestamp 1586364061
transform 1 0 2116 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_25
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__532__B
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _535_
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_29
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__532__A
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__530__A
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_382
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _531_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _530_
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_46
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_42
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__530__B
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _533_
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 866 592
use scs8hd_buf_1  _529_
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_58
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__529__A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__544__B
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__543__A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_390
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _543_
timestamp 1586364061
transform 1 0 6900 0 1 16864
box -38 -48 866 592
use scs8hd_decap_6  FILLER_27_76
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_72
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_67
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__544__A
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__545__B
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_82
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_85
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_383
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__546__A
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__546__B
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _546_
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 866 592
use scs8hd_decap_6  FILLER_26_82
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_102
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__545__A
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_109
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_114
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__537__B
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__537__A
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_127
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__538__B
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__538__A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_391
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _538_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_143
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_137
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_137
timestamp 1586364061
transform 1 0 13708 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__540__B
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__536__A
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__540__A
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_1  _536_
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_384
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_159
timestamp 1586364061
transform 1 0 15732 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15916 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_168
timestamp 1586364061
transform 1 0 16560 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_164
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__554__A
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_179
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_171
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__528__A
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _528_
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 314 592
use scs8hd_or2_4  _527_
timestamp 1586364061
transform 1 0 16928 0 -1 16864
box -38 -48 682 592
use scs8hd_fill_1  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_183
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__599__A
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__B
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_392
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_or2_4  _599_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 682 592
use scs8hd_inv_8  _307_
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_195
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_191
timestamp 1586364061
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_196
timestamp 1586364061
transform 1 0 19136 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__599__B
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_206
timestamp 1586364061
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_202
timestamp 1586364061
transform 1 0 19688 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_201
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__579__B
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__579__A
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_209
timestamp 1586364061
transform 1 0 20332 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_385
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _619_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_233
timestamp 1586364061
transform 1 0 22540 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_227
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_233
timestamp 1586364061
transform 1 0 22540 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_229
timestamp 1586364061
transform 1 0 22172 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 22632 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_241
timestamp 1586364061
transform 1 0 23276 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_237
timestamp 1586364061
transform 1 0 22908 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_236
timestamp 1586364061
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23000 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_3  FILLER_27_249
timestamp 1586364061
transform 1 0 24012 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_247
timestamp 1586364061
transform 1 0 23828 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__552__C
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__552__B
timestamp 1586364061
transform 1 0 23828 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_393
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_259
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_258
timestamp 1586364061
transform 1 0 24840 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_254
timestamp 1586364061
transform 1 0 24472 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__227__B
timestamp 1586364061
transform 1 0 24288 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 314 592
use scs8hd_or2_4  _227_
timestamp 1586364061
transform 1 0 24288 0 1 16864
box -38 -48 682 592
use scs8hd_decap_4  FILLER_27_267
timestamp 1586364061
transform 1 0 25668 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_263
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_266
timestamp 1586364061
transform 1 0 25576 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__345__A
timestamp 1586364061
transform 1 0 25484 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_271
timestamp 1586364061
transform 1 0 26036 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_271
timestamp 1586364061
transform 1 0 26036 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__378__B
timestamp 1586364061
transform 1 0 25852 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__378__A
timestamp 1586364061
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__317__A
timestamp 1586364061
transform 1 0 26128 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_386
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _379_
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _378_
timestamp 1586364061
transform 1 0 26312 0 1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_287
timestamp 1586364061
transform 1 0 27508 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_283
timestamp 1586364061
transform 1 0 27140 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_285
timestamp 1586364061
transform 1 0 27324 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__346__D
timestamp 1586364061
transform 1 0 27600 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__317__B
timestamp 1586364061
transform 1 0 27324 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_291
timestamp 1586364061
transform 1 0 27876 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_290
timestamp 1586364061
transform 1 0 27784 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__359__A
timestamp 1586364061
transform 1 0 28152 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__315__A
timestamp 1586364061
transform 1 0 27968 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _359_
timestamp 1586364061
transform 1 0 28152 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__320__C
timestamp 1586364061
transform 1 0 28612 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_296
timestamp 1586364061
transform 1 0 28336 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_300
timestamp 1586364061
transform 1 0 28704 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_297
timestamp 1586364061
transform 1 0 28428 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _360_
timestamp 1586364061
transform 1 0 28796 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__320__D
timestamp 1586364061
transform 1 0 28980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_304
timestamp 1586364061
transform 1 0 29072 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_301
timestamp 1586364061
transform 1 0 28796 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_394
timestamp 1586364061
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__368__B
timestamp 1586364061
transform 1 0 29256 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_306
timestamp 1586364061
transform 1 0 29256 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_311
timestamp 1586364061
transform 1 0 29716 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_312
timestamp 1586364061
transform 1 0 29808 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_308
timestamp 1586364061
transform 1 0 29440 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__367__B
timestamp 1586364061
transform 1 0 29624 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__367__A
timestamp 1586364061
transform 1 0 29532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 29900 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 30084 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 30176 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_27_326
timestamp 1586364061
transform 1 0 31096 0 1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_26_331
timestamp 1586364061
transform 1 0 31556 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_327
timestamp 1586364061
transform 1 0 31188 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31372 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31648 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_387
timestamp 1586364061
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31832 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_347
timestamp 1586364061
transform 1 0 33028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_343
timestamp 1586364061
transform 1 0 32660 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_346
timestamp 1586364061
transform 1 0 32936 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__321__A
timestamp 1586364061
transform 1 0 32844 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_358
timestamp 1586364061
transform 1 0 34040 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_354
timestamp 1586364061
transform 1 0 33672 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_356
timestamp 1586364061
transform 1 0 33856 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_352
timestamp 1586364061
transform 1 0 33488 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__344__A
timestamp 1586364061
transform 1 0 33304 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__344__B
timestamp 1586364061
transform 1 0 33212 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33856 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33396 0 1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 33948 0 -1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_371
timestamp 1586364061
transform 1 0 35236 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_367
timestamp 1586364061
transform 1 0 34868 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_368
timestamp 1586364061
transform 1 0 34960 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__402__B
timestamp 1586364061
transform 1 0 34592 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__402__A
timestamp 1586364061
transform 1 0 35052 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_395
timestamp 1586364061
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35420 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_380
timestamp 1586364061
transform 1 0 36064 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_376
timestamp 1586364061
transform 1 0 35696 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_387
timestamp 1586364061
transform 1 0 36708 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35880 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36248 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 35696 0 -1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_397
timestamp 1586364061
transform 1 0 37628 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_393
timestamp 1586364061
transform 1 0 37260 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_391
timestamp 1586364061
transform 1 0 37076 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37812 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36892 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_388
timestamp 1586364061
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37996 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_410
timestamp 1586364061
transform 1 0 38824 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_407
timestamp 1586364061
transform 1 0 38548 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_418
timestamp 1586364061
transform 1 0 39560 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_414
timestamp 1586364061
transform 1 0 39192 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_418
timestamp 1586364061
transform 1 0 39560 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__390__B
timestamp 1586364061
transform 1 0 39744 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__356__B
timestamp 1586364061
transform 1 0 39376 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__356__A
timestamp 1586364061
transform 1 0 39008 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _347_
timestamp 1586364061
transform 1 0 39284 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_426
timestamp 1586364061
transform 1 0 40296 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_422
timestamp 1586364061
transform 1 0 39928 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_427
timestamp 1586364061
transform 1 0 40388 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_424
timestamp 1586364061
transform 1 0 40112 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40204 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40572 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__390__A
timestamp 1586364061
transform 1 0 40112 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_396
timestamp 1586364061
transform 1 0 40388 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_442
timestamp 1586364061
transform 1 0 41768 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_435
timestamp 1586364061
transform 1 0 41124 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_431
timestamp 1586364061
transform 1 0 40756 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_440
timestamp 1586364061
transform 1 0 41584 0 -1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40756 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41492 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_27_450
timestamp 1586364061
transform 1 0 42504 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_446
timestamp 1586364061
transform 1 0 42136 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_452
timestamp 1586364061
transform 1 0 42688 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42320 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41952 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43056 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44896 0 -1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_389
timestamp 1586364061
transform 1 0 43240 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43516 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_468
timestamp 1586364061
transform 1 0 44160 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_26_479
timestamp 1586364061
transform 1 0 45172 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_459
timestamp 1586364061
transform 1 0 43332 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_463
timestamp 1586364061
transform 1 0 43700 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_475
timestamp 1586364061
transform 1 0 44804 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_397
timestamp 1586364061
transform 1 0 46000 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_491
timestamp 1586364061
transform 1 0 46276 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_503
timestamp 1586364061
transform 1 0 47380 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_487
timestamp 1586364061
transform 1 0 45908 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_489
timestamp 1586364061
transform 1 0 46092 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_501
timestamp 1586364061
transform 1 0 47196 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 48852 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 48852 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_515
timestamp 1586364061
transform 1 0 48484 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_513
timestamp 1586364061
transform 1 0 48300 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_nor2_4  _532_
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_398
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__556__B
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _544_
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__543__B
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_60
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_78
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _545_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_399
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_83
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _537_
timestamp 1586364061
transform 1 0 11684 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__539__B
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_114
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_124
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_134
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _540_
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_400
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__541__B
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_144
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_148
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_or2_4  _232_
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 682 592
use scs8hd_buf_1  _554_
timestamp 1586364061
transform 1 0 17020 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_165
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_176
timestamp 1586364061
transform 1 0 17296 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_180
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 406 592
use scs8hd_or2_4  _579_
timestamp 1586364061
transform 1 0 19412 0 -1 17952
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_401
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_191
timestamp 1586364061
transform 1 0 18676 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_8  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use scs8hd_buf_1  _228_
timestamp 1586364061
transform 1 0 22632 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__552__A
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_232
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_237
timestamp 1586364061
transform 1 0 22908 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_241
timestamp 1586364061
transform 1 0 23276 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_1  _345_
timestamp 1586364061
transform 1 0 25392 0 -1 17952
box -38 -48 314 592
use scs8hd_or4_4  _552_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23644 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__231__B
timestamp 1586364061
transform 1 0 25208 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__526__C
timestamp 1586364061
transform 1 0 24656 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__552__D
timestamp 1586364061
transform 1 0 23460 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_254
timestamp 1586364061
transform 1 0 24472 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_258
timestamp 1586364061
transform 1 0 24840 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__369__D
timestamp 1586364061
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__319__A
timestamp 1586364061
transform 1 0 25852 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_402
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_or2_4  _317_
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 682 592
use scs8hd_fill_1  FILLER_28_287
timestamp 1586364061
transform 1 0 27508 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_283
timestamp 1586364061
transform 1 0 27140 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__346__B
timestamp 1586364061
transform 1 0 27600 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_290
timestamp 1586364061
transform 1 0 27784 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_8  _315_
timestamp 1586364061
transform 1 0 27968 0 -1 17952
box -38 -48 866 592
use scs8hd_nor2_4  _367_
timestamp 1586364061
transform 1 0 29532 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__358__B
timestamp 1586364061
transform 1 0 29256 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30544 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_301
timestamp 1586364061
transform 1 0 28796 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_305
timestamp 1586364061
transform 1 0 29164 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_308
timestamp 1586364061
transform 1 0 29440 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_318
timestamp 1586364061
transform 1 0 30360 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_322
timestamp 1586364061
transform 1 0 30728 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_326
timestamp 1586364061
transform 1 0 31096 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30912 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_331
timestamp 1586364061
transform 1 0 31556 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__399__A
timestamp 1586364061
transform 1 0 31372 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_335
timestamp 1586364061
transform 1 0 31924 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__399__B
timestamp 1586364061
transform 1 0 31740 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_403
timestamp 1586364061
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_337
timestamp 1586364061
transform 1 0 32108 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_1  _321_
timestamp 1586364061
transform 1 0 32292 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_346
timestamp 1586364061
transform 1 0 32936 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_342
timestamp 1586364061
transform 1 0 32568 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__400__B
timestamp 1586364061
transform 1 0 32752 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _344_
timestamp 1586364061
transform 1 0 33304 0 -1 17952
box -38 -48 866 592
use scs8hd_nor2_4  _402_
timestamp 1586364061
transform 1 0 34868 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_359
timestamp 1586364061
transform 1 0 34132 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_4  FILLER_28_380
timestamp 1586364061
transform 1 0 36064 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_376
timestamp 1586364061
transform 1 0 35696 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 35880 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_387
timestamp 1586364061
transform 1 0 36708 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36892 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_28_391
timestamp 1586364061
transform 1 0 37076 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_4  FILLER_28_402
timestamp 1586364061
transform 1 0 38088 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_398
timestamp 1586364061
transform 1 0 37720 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37904 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_404
timestamp 1586364061
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _356_
timestamp 1586364061
transform 1 0 38548 0 -1 17952
box -38 -48 866 592
use scs8hd_nor2_4  _390_
timestamp 1586364061
transform 1 0 40112 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_1  FILLER_28_406
timestamp 1586364061
transform 1 0 38456 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_416
timestamp 1586364061
transform 1 0 39376 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41676 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41124 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42228 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42596 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_433
timestamp 1586364061
transform 1 0 40940 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_437
timestamp 1586364061
transform 1 0 41308 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  FILLER_28_444
timestamp 1586364061
transform 1 0 41952 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_449
timestamp 1586364061
transform 1 0 42412 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_453
timestamp 1586364061
transform 1 0 42780 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_405
timestamp 1586364061
transform 1 0 43240 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_457
timestamp 1586364061
transform 1 0 43148 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_459
timestamp 1586364061
transform 1 0 43332 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_471
timestamp 1586364061
transform 1 0 44436 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_483
timestamp 1586364061
transform 1 0 45540 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_495
timestamp 1586364061
transform 1 0 46644 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_507
timestamp 1586364061
transform 1 0 47748 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 48852 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_515
timestamp 1586364061
transform 1 0 48484 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_nor2_4  _556_
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__556__A
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__559__A
timestamp 1586364061
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__559__B
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_43
timestamp 1586364061
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_406
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 866 592
use scs8hd_nor2_4  _572_
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__572__A
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__572__B
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_85
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_89
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_102
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_106
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__539__A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_407
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _539_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _541_
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 866 592
use scs8hd_nor2_4  _542_
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__408__A
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__541__A
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__542__A
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_153
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 590 592
use scs8hd_or2_4  _553_
timestamp 1586364061
transform 1 0 18124 0 1 17952
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_408
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__553__B
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_178
timestamp 1586364061
transform 1 0 17480 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_192
timestamp 1586364061
transform 1 0 18768 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__553__A
timestamp 1586364061
transform 1 0 18952 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_204
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_200
timestamp 1586364061
transform 1 0 19504 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__618__A
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use scs8hd_inv_8  _618_
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_29_221
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_225
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__578__C
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_or4_4  _231_
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 866 592
use scs8hd_or4_4  _578_
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_409
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__578__A
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__526__B
timestamp 1586364061
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_254
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use scs8hd_or4_4  _346_
timestamp 1586364061
transform 1 0 27600 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__369__A
timestamp 1586364061
transform 1 0 26588 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__346__A
timestamp 1586364061
transform 1 0 27416 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__D
timestamp 1586364061
transform 1 0 26220 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__369__B
timestamp 1586364061
transform 1 0 26956 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_271
timestamp 1586364061
transform 1 0 26036 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_275
timestamp 1586364061
transform 1 0 26404 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_279
timestamp 1586364061
transform 1 0 26772 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_283
timestamp 1586364061
transform 1 0 27140 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_301
timestamp 1586364061
transform 1 0 28796 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_297
timestamp 1586364061
transform 1 0 28428 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__320__A
timestamp 1586364061
transform 1 0 28612 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__358__A
timestamp 1586364061
transform 1 0 28980 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_410
timestamp 1586364061
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use scs8hd_or4_4  _358_
timestamp 1586364061
transform 1 0 29256 0 1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_29_319
timestamp 1586364061
transform 1 0 30452 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_315
timestamp 1586364061
transform 1 0 30084 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__358__D
timestamp 1586364061
transform 1 0 30636 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30268 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _399_
timestamp 1586364061
transform 1 0 31372 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31004 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__400__A
timestamp 1586364061
transform 1 0 32384 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__403__A
timestamp 1586364061
transform 1 0 33028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_323
timestamp 1586364061
transform 1 0 30820 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_327
timestamp 1586364061
transform 1 0 31188 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_338
timestamp 1586364061
transform 1 0 32200 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_342
timestamp 1586364061
transform 1 0 32568 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_346
timestamp 1586364061
transform 1 0 32936 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_358
timestamp 1586364061
transform 1 0 34040 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__401__A
timestamp 1586364061
transform 1 0 34224 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _403_
timestamp 1586364061
transform 1 0 33212 0 1 17952
box -38 -48 866 592
use scs8hd_decap_4  FILLER_29_367
timestamp 1586364061
transform 1 0 34868 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_362
timestamp 1586364061
transform 1 0 34408 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__401__B
timestamp 1586364061
transform 1 0 34592 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 35236 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_411
timestamp 1586364061
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_373
timestamp 1586364061
transform 1 0 35420 0 1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 35512 0 1 17952
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37260 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37720 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37076 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36708 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_385
timestamp 1586364061
transform 1 0 36524 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_389
timestamp 1586364061
transform 1 0 36892 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_396
timestamp 1586364061
transform 1 0 37536 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_400
timestamp 1586364061
transform 1 0 37904 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_406
timestamp 1586364061
transform 1 0 38456 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__388__B
timestamp 1586364061
transform 1 0 38272 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__388__A
timestamp 1586364061
transform 1 0 38640 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _388_
timestamp 1586364061
transform 1 0 38824 0 1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_29_423
timestamp 1586364061
transform 1 0 40020 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_419
timestamp 1586364061
transform 1 0 39652 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_412
timestamp 1586364061
transform 1 0 40388 0 1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 40480 0 1 17952
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42228 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__398__A
timestamp 1586364061
transform 1 0 41952 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_439
timestamp 1586364061
transform 1 0 41492 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_443
timestamp 1586364061
transform 1 0 41860 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_446
timestamp 1586364061
transform 1 0 42136 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_456
timestamp 1586364061
transform 1 0 43056 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43700 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_461
timestamp 1586364061
transform 1 0 43516 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_465
timestamp 1586364061
transform 1 0 43884 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_477
timestamp 1586364061
transform 1 0 44988 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_413
timestamp 1586364061
transform 1 0 46000 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_485
timestamp 1586364061
transform 1 0 45724 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_489
timestamp 1586364061
transform 1 0 46092 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_501
timestamp 1586364061
transform 1 0 47196 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 48852 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_513
timestamp 1586364061
transform 1 0 48300 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__558__B
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_20
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _559_
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_414
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 4324 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_28
timestamp 1586364061
transform 1 0 3680 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_37
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_54
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_58
timestamp 1586364061
transform 1 0 6440 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_61
timestamp 1586364061
transform 1 0 6716 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_73
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_415
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__571__A
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_98
timestamp 1586364061
transform 1 0 10120 0 -1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12236 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_113
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_30_132
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_1  _408_
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_416
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__542__B
timestamp 1586364061
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_136
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_159
timestamp 1586364061
transform 1 0 15732 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 19040
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18124 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_30_183
timestamp 1586364061
transform 1 0 17940 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_187
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_417
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_8  _229_
timestamp 1586364061
transform 1 0 22264 0 -1 19040
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__578__D
timestamp 1586364061
transform 1 0 23276 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_218
timestamp 1586364061
transform 1 0 21160 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_222
timestamp 1586364061
transform 1 0 21528 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_1  _319_
timestamp 1586364061
transform 1 0 25392 0 -1 19040
box -38 -48 314 592
use scs8hd_or4_4  _526_
timestamp 1586364061
transform 1 0 23828 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__578__B
timestamp 1586364061
transform 1 0 23644 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__C
timestamp 1586364061
transform 1 0 25208 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__526__D
timestamp 1586364061
transform 1 0 24840 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_243
timestamp 1586364061
transform 1 0 23460 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_256
timestamp 1586364061
transform 1 0 24656 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_260
timestamp 1586364061
transform 1 0 25024 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_267
timestamp 1586364061
transform 1 0 25668 0 -1 19040
box -38 -48 590 592
use scs8hd_or4_4  _320_
timestamp 1586364061
transform 1 0 28152 0 -1 19040
box -38 -48 866 592
use scs8hd_or4_4  _369_
timestamp 1586364061
transform 1 0 26588 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_418
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__320__B
timestamp 1586364061
transform 1 0 27968 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__346__C
timestamp 1586364061
transform 1 0 27600 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__369__C
timestamp 1586364061
transform 1 0 26220 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_286
timestamp 1586364061
transform 1 0 27416 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_290
timestamp 1586364061
transform 1 0 27784 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29716 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__438__D
timestamp 1586364061
transform 1 0 29256 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__358__C
timestamp 1586364061
transform 1 0 30176 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__B
timestamp 1586364061
transform 1 0 30544 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_303
timestamp 1586364061
transform 1 0 28980 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_308
timestamp 1586364061
transform 1 0 29440 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_314
timestamp 1586364061
transform 1 0 29992 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_318
timestamp 1586364061
transform 1 0 30360 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_322
timestamp 1586364061
transform 1 0 30728 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _400_
timestamp 1586364061
transform 1 0 32108 0 -1 19040
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_419
timestamp 1586364061
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__438__C
timestamp 1586364061
transform 1 0 31464 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31832 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_328
timestamp 1586364061
transform 1 0 31280 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_332
timestamp 1586364061
transform 1 0 31648 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_346
timestamp 1586364061
transform 1 0 32936 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _401_
timestamp 1586364061
transform 1 0 33672 0 -1 19040
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 35236 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__403__B
timestamp 1586364061
transform 1 0 33212 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35052 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34684 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_351
timestamp 1586364061
transform 1 0 33396 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_363
timestamp 1586364061
transform 1 0 34500 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_367
timestamp 1586364061
transform 1 0 34868 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_420
timestamp 1586364061
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36800 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36432 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_382
timestamp 1586364061
transform 1 0 36248 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_386
timestamp 1586364061
transform 1 0 36616 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_390
timestamp 1586364061
transform 1 0 36984 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_396
timestamp 1586364061
transform 1 0 37536 0 -1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 40204 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__393__B
timestamp 1586364061
transform 1 0 39284 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__391__B
timestamp 1586364061
transform 1 0 38824 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40020 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_407
timestamp 1586364061
transform 1 0 38548 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_412
timestamp 1586364061
transform 1 0 39008 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_30_417
timestamp 1586364061
transform 1 0 39468 0 -1 19040
box -38 -48 590 592
use scs8hd_buf_1  _398_
timestamp 1586364061
transform 1 0 41952 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 42412 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41584 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_436
timestamp 1586364061
transform 1 0 41216 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_442
timestamp 1586364061
transform 1 0 41768 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_447
timestamp 1586364061
transform 1 0 42228 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_451
timestamp 1586364061
transform 1 0 42596 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_421
timestamp 1586364061
transform 1 0 43240 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_457
timestamp 1586364061
transform 1 0 43148 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_468
timestamp 1586364061
transform 1 0 44160 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_480
timestamp 1586364061
transform 1 0 45264 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_492
timestamp 1586364061
transform 1 0 46368 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_504
timestamp 1586364061
transform 1 0 47472 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 48852 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _558_
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__558__A
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_46
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_50
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_54
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_422
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__555__A
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 866 592
use scs8hd_nor2_4  _571_
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__269__A
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_88
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_92
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_109
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__564__B
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__564__A
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_423
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_153
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_424
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_166
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_170
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_31_176
timestamp 1586364061
transform 1 0 17296 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_180
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__617__A
timestamp 1586364061
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_214
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__318__B
timestamp 1586364061
transform 1 0 22724 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__318__A
timestamp 1586364061
transform 1 0 23092 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_227
timestamp 1586364061
transform 1 0 21988 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_237
timestamp 1586364061
transform 1 0 22908 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_241
timestamp 1586364061
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use scs8hd_inv_8  _316_
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_425
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__316__A
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__381__A
timestamp 1586364061
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__526__A
timestamp 1586364061
transform 1 0 23828 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_249
timestamp 1586364061
transform 1 0 24012 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_264
timestamp 1586364061
transform 1 0 25392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_268
timestamp 1586364061
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__357__B
timestamp 1586364061
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use scs8hd_or2_4  _357_
timestamp 1586364061
transform 1 0 26128 0 1 19040
box -38 -48 682 592
use scs8hd_fill_2  FILLER_31_283
timestamp 1586364061
transform 1 0 27140 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_279
timestamp 1586364061
transform 1 0 26772 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__357__A
timestamp 1586364061
transform 1 0 26956 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_290
timestamp 1586364061
transform 1 0 27784 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__328__A
timestamp 1586364061
transform 1 0 27324 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _331_
timestamp 1586364061
transform 1 0 27508 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_294
timestamp 1586364061
transform 1 0 28152 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__383__A
timestamp 1586364061
transform 1 0 27968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_302
timestamp 1586364061
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_298
timestamp 1586364061
transform 1 0 28520 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__383__B
timestamp 1586364061
transform 1 0 28336 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__438__B
timestamp 1586364061
transform 1 0 28980 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_426
timestamp 1586364061
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_306
timestamp 1586364061
transform 1 0 29256 0 1 19040
box -38 -48 130 592
use scs8hd_or4_4  _396_
timestamp 1586364061
transform 1 0 29348 0 1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_31_320
timestamp 1586364061
transform 1 0 30544 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_316
timestamp 1586364061
transform 1 0 30176 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__D
timestamp 1586364061
transform 1 0 30360 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30728 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 31924 0 1 19040
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30912 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 31740 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 31372 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33120 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_327
timestamp 1586364061
transform 1 0 31188 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_331
timestamp 1586364061
transform 1 0 31556 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_346
timestamp 1586364061
transform 1 0 32936 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_357
timestamp 1586364061
transform 1 0 33948 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_350
timestamp 1586364061
transform 1 0 33304 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33488 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34132 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33672 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_367
timestamp 1586364061
transform 1 0 34868 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_361
timestamp 1586364061
transform 1 0 34316 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 34592 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_427
timestamp 1586364061
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 35052 0 1 19040
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36800 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37812 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36616 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_380
timestamp 1586364061
transform 1 0 36064 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_384
timestamp 1586364061
transform 1 0 36432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_397
timestamp 1586364061
transform 1 0 37628 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_401
timestamp 1586364061
transform 1 0 37996 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_405
timestamp 1586364061
transform 1 0 38364 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38180 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__391__A
timestamp 1586364061
transform 1 0 38640 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _391_
timestamp 1586364061
transform 1 0 38824 0 1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_31_423
timestamp 1586364061
transform 1 0 40020 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_419
timestamp 1586364061
transform 1 0 39652 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__393__A
timestamp 1586364061
transform 1 0 39836 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_428
timestamp 1586364061
transform 1 0 40388 0 1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 40480 0 1 19040
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 42412 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 42228 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_439
timestamp 1586364061
transform 1 0 41492 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_443
timestamp 1586364061
transform 1 0 41860 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44988 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43608 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43976 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_460
timestamp 1586364061
transform 1 0 43424 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_464
timestamp 1586364061
transform 1 0 43792 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_468
timestamp 1586364061
transform 1 0 44160 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_476
timestamp 1586364061
transform 1 0 44896 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_479
timestamp 1586364061
transform 1 0 45172 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_429
timestamp 1586364061
transform 1 0 46000 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_487
timestamp 1586364061
transform 1 0 45908 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_489
timestamp 1586364061
transform 1 0 46092 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_501
timestamp 1586364061
transform 1 0 47196 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 48852 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_513
timestamp 1586364061
transform 1 0 48300 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__557__B
timestamp 1586364061
transform 1 0 2668 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 4324 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_430
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_46
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_1  _555_
timestamp 1586364061
transform 1 0 8096 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__570__A
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_54
timestamp 1586364061
transform 1 0 6072 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_74
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_79
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_87
timestamp 1586364061
transform 1 0 9108 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_431
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_buf_1  _269_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_96
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__571__B
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_100
timestamp 1586364061
transform 1 0 10304 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 314 592
use scs8hd_nor2_4  _564_
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__563__B
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_109
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_432
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18124 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_164
timestamp 1586364061
transform 1 0 16192 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_183
timestamp 1586364061
transform 1 0 17940 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_187
timestamp 1586364061
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_433
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_200
timestamp 1586364061
transform 1 0 19504 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_204
timestamp 1586364061
transform 1 0 19872 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_208
timestamp 1586364061
transform 1 0 20240 0 -1 20128
box -38 -48 590 592
use scs8hd_nand2_4  _318_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22724 0 -1 20128
box -38 -48 866 592
use scs8hd_inv_8  _617_
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_224
timestamp 1586364061
transform 1 0 21712 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_232
timestamp 1586364061
transform 1 0 22448 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_8  _381_
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__504__D
timestamp 1586364061
transform 1 0 24656 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__504__A
timestamp 1586364061
transform 1 0 24288 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_244
timestamp 1586364061
transform 1 0 23552 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_254
timestamp 1586364061
transform 1 0 24472 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_267
timestamp 1586364061
transform 1 0 25668 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_271
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__482__B
timestamp 1586364061
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__482__D
timestamp 1586364061
transform 1 0 25852 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_434
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_buf_1  _328_
timestamp 1586364061
transform 1 0 26680 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_285
timestamp 1586364061
transform 1 0 27324 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_281
timestamp 1586364061
transform 1 0 26956 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__B
timestamp 1586364061
transform 1 0 27140 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__331__A
timestamp 1586364061
transform 1 0 27508 0 -1 20128
box -38 -48 222 592
use scs8hd_nand2_4  _383_
timestamp 1586364061
transform 1 0 27692 0 -1 20128
box -38 -48 866 592
use scs8hd_or4_4  _438_
timestamp 1586364061
transform 1 0 29256 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__449__D
timestamp 1586364061
transform 1 0 29072 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__438__A
timestamp 1586364061
transform 1 0 28704 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__A
timestamp 1586364061
transform 1 0 30268 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__449__C
timestamp 1586364061
transform 1 0 30636 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_298
timestamp 1586364061
transform 1 0 28520 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_302
timestamp 1586364061
transform 1 0 28888 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_315
timestamp 1586364061
transform 1 0 30084 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_319
timestamp 1586364061
transform 1 0 30452 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 32200 0 -1 20128
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30820 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_435
timestamp 1586364061
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__385__B
timestamp 1586364061
transform 1 0 31280 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__C
timestamp 1586364061
transform 1 0 31648 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_326
timestamp 1586364061
transform 1 0 31096 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_330
timestamp 1586364061
transform 1 0 31464 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_334
timestamp 1586364061
transform 1 0 31832 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_337
timestamp 1586364061
transform 1 0 32108 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33948 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33396 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35052 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33764 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_349
timestamp 1586364061
transform 1 0 33212 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_353
timestamp 1586364061
transform 1 0 33580 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_366
timestamp 1586364061
transform 1 0 34776 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_371
timestamp 1586364061
transform 1 0 35236 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_436
timestamp 1586364061
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_379
timestamp 1586364061
transform 1 0 35972 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_389
timestamp 1586364061
transform 1 0 36892 0 -1 20128
box -38 -48 774 592
use scs8hd_nor2_4  _393_
timestamp 1586364061
transform 1 0 39284 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40480 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_407
timestamp 1586364061
transform 1 0 38548 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_32_424
timestamp 1586364061
transform 1 0 40112 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41584 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41216 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40848 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_430
timestamp 1586364061
transform 1 0 40664 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_434
timestamp 1586364061
transform 1 0 41032 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_438
timestamp 1586364061
transform 1 0 41400 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_449
timestamp 1586364061
transform 1 0 42412 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44988 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43424 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_437
timestamp 1586364061
transform 1 0 43240 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_457
timestamp 1586364061
transform 1 0 43148 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_459
timestamp 1586364061
transform 1 0 43332 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_469
timestamp 1586364061
transform 1 0 44252 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_480
timestamp 1586364061
transform 1 0 45264 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_492
timestamp 1586364061
transform 1 0 46368 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_504
timestamp 1586364061
transform 1 0 47472 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 48852 0 -1 20128
box -38 -48 314 592
use scs8hd_nor2_4  _557_
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__557__A
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_26
timestamp 1586364061
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_30
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__560__A
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_446
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 1050 592
use scs8hd_nor2_4  _560_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_50
timestamp 1586364061
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_46
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  FILLER_34_41
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_49
timestamp 1586364061
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_45
timestamp 1586364061
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__560__B
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_62
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_54
timestamp 1586364061
transform 1 0 6072 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6900 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_438
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_69
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_65
timestamp 1586364061
transform 1 0 7084 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_68
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__570__B
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__569__A
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _570_
timestamp 1586364061
transform 1 0 7728 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _569_
timestamp 1586364061
transform 1 0 7728 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_89
timestamp 1586364061
transform 1 0 9292 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_81
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_85
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__569__B
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_447
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_34_104
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_104
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_100
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_115
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_111
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_121
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__562__A
timestamp 1586364061
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_439
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_buf_1  _562_
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_134
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_130
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__563__A
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _563_
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_144
timestamp 1586364061
transform 1 0 14352 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_138
timestamp 1586364061
transform 1 0 13800 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_33_149
timestamp 1586364061
transform 1 0 14812 0 1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_34_148
timestamp 1586364061
transform 1 0 14720 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_448
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_153
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_156
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_157
timestamp 1586364061
transform 1 0 15548 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_161
timestamp 1586364061
transform 1 0 15916 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_165
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_164
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_173
timestamp 1586364061
transform 1 0 17020 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_180
timestamp 1586364061
transform 1 0 17664 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_176
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_187
timestamp 1586364061
transform 1 0 18308 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_183
timestamp 1586364061
transform 1 0 17940 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18124 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_440
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_197
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_193
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__614__A
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_inv_8  _614_
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_204
timestamp 1586364061
transform 1 0 19872 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_200
timestamp 1586364061
transform 1 0 19504 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__489__B
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 866 592
use scs8hd_decap_6  FILLER_33_210
timestamp 1586364061
transform 1 0 20424 0 1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_449
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_220
timestamp 1586364061
transform 1 0 21344 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__616__A
timestamp 1586364061
transform 1 0 21160 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__492__B
timestamp 1586364061
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use scs8hd_inv_8  _616_
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _492_
timestamp 1586364061
transform 1 0 21620 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_232
timestamp 1586364061
transform 1 0 22448 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_6  FILLER_33_231
timestamp 1586364061
transform 1 0 22356 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_227
timestamp 1586364061
transform 1 0 21988 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__492__A
timestamp 1586364061
transform 1 0 22172 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_236
timestamp 1586364061
transform 1 0 22816 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_240
timestamp 1586364061
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_237
timestamp 1586364061
transform 1 0 22908 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22908 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__483__A
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  _483_
timestamp 1586364061
transform 1 0 23184 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_247
timestamp 1586364061
transform 1 0 23828 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_243
timestamp 1586364061
transform 1 0 23460 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_441
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_or2_4  _230_
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 682 592
use scs8hd_fill_2  FILLER_34_254
timestamp 1586364061
transform 1 0 24472 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_260
timestamp 1586364061
transform 1 0 25024 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_256
timestamp 1586364061
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_252
timestamp 1586364061
transform 1 0 24288 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__504__B
timestamp 1586364061
transform 1 0 24656 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__504__C
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__B
timestamp 1586364061
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use scs8hd_or4_4  _504_
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_267
timestamp 1586364061
transform 1 0 25668 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__482__C
timestamp 1586364061
transform 1 0 25300 0 1 20128
box -38 -48 222 592
use scs8hd_or4_4  _482_
timestamp 1586364061
transform 1 0 25484 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_271
timestamp 1586364061
transform 1 0 26036 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_278
timestamp 1586364061
transform 1 0 26680 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_274
timestamp 1586364061
transform 1 0 26312 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__494__A
timestamp 1586364061
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__482__A
timestamp 1586364061
transform 1 0 25852 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__C
timestamp 1586364061
transform 1 0 26496 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_450
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_or4_4  _493_
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_285
timestamp 1586364061
transform 1 0 27324 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_285
timestamp 1586364061
transform 1 0 27324 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__A
timestamp 1586364061
transform 1 0 27508 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__460__D
timestamp 1586364061
transform 1 0 27508 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__D
timestamp 1586364061
transform 1 0 26864 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  _494_
timestamp 1586364061
transform 1 0 27048 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_289
timestamp 1586364061
transform 1 0 27692 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_289
timestamp 1586364061
transform 1 0 27692 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__471__C
timestamp 1586364061
transform 1 0 27876 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27968 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28060 0 -1 21216
box -38 -48 314 592
use scs8hd_buf_1  _226_
timestamp 1586364061
transform 1 0 28152 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 28612 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__471__D
timestamp 1586364061
transform 1 0 28520 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_297
timestamp 1586364061
transform 1 0 28428 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_296
timestamp 1586364061
transform 1 0 28336 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_300
timestamp 1586364061
transform 1 0 28704 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_442
timestamp 1586364061
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__449__B
timestamp 1586364061
transform 1 0 28980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__449__A
timestamp 1586364061
transform 1 0 28888 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_301
timestamp 1586364061
transform 1 0 28796 0 1 20128
box -38 -48 222 592
use scs8hd_or4_4  _449_
timestamp 1586364061
transform 1 0 29072 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_313
timestamp 1586364061
transform 1 0 29900 0 -1 21216
box -38 -48 222 592
use scs8hd_or4_4  _427_
timestamp 1586364061
transform 1 0 29256 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_317
timestamp 1586364061
transform 1 0 30268 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_319
timestamp 1586364061
transform 1 0 30452 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_315
timestamp 1586364061
transform 1 0 30084 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__427__B
timestamp 1586364061
transform 1 0 30452 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__427__D
timestamp 1586364061
transform 1 0 30084 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__385__D
timestamp 1586364061
transform 1 0 30268 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__380__A
timestamp 1586364061
transform 1 0 30636 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  _380_
timestamp 1586364061
transform 1 0 30636 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_332
timestamp 1586364061
transform 1 0 31648 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_328
timestamp 1586364061
transform 1 0 31280 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_324
timestamp 1586364061
transform 1 0 30912 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_332
timestamp 1586364061
transform 1 0 31648 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__385__C
timestamp 1586364061
transform 1 0 31464 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__385__A
timestamp 1586364061
transform 1 0 31096 0 -1 21216
box -38 -48 222 592
use scs8hd_or4_4  _385_
timestamp 1586364061
transform 1 0 30820 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_451
timestamp 1586364061
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__427__C
timestamp 1586364061
transform 1 0 31832 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__427__A
timestamp 1586364061
transform 1 0 32200 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_336
timestamp 1586364061
transform 1 0 32016 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_337
timestamp 1586364061
transform 1 0 32108 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__404__B
timestamp 1586364061
transform 1 0 32292 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_340
timestamp 1586364061
transform 1 0 32384 0 1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_34_341
timestamp 1586364061
transform 1 0 32476 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 32844 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_344
timestamp 1586364061
transform 1 0 32752 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_345
timestamp 1586364061
transform 1 0 32844 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33028 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 32936 0 -1 21216
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_34_357
timestamp 1586364061
transform 1 0 33948 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_356
timestamp 1586364061
transform 1 0 33856 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_365
timestamp 1586364061
transform 1 0 34684 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_33_360
timestamp 1586364061
transform 1 0 34224 0 1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34040 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_443
timestamp 1586364061
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_371
timestamp 1586364061
transform 1 0 35236 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_371
timestamp 1586364061
transform 1 0 35236 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_367
timestamp 1586364061
transform 1 0 34868 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35512 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35052 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34960 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_383
timestamp 1586364061
transform 1 0 36340 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_379
timestamp 1586364061
transform 1 0 35972 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36524 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36156 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35972 0 -1 21216
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35696 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_392
timestamp 1586364061
transform 1 0 37168 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_388
timestamp 1586364061
transform 1 0 36800 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_392
timestamp 1586364061
transform 1 0 37168 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_387
timestamp 1586364061
transform 1 0 36708 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36984 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37352 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36892 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_398
timestamp 1586364061
transform 1 0 37720 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_396
timestamp 1586364061
transform 1 0 37536 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_396
timestamp 1586364061
transform 1 0 37536 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__384__A
timestamp 1586364061
transform 1 0 37720 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_452
timestamp 1586364061
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_1  _384_
timestamp 1586364061
transform 1 0 37904 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38548 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38548 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_403
timestamp 1586364061
transform 1 0 38180 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_406
timestamp 1586364061
transform 1 0 38456 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__392__B
timestamp 1586364061
transform 1 0 39008 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_409
timestamp 1586364061
transform 1 0 38732 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_410
timestamp 1586364061
transform 1 0 38824 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39192 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_413
timestamp 1586364061
transform 1 0 39100 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_414
timestamp 1586364061
transform 1 0 39192 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_423
timestamp 1586364061
transform 1 0 40020 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_419
timestamp 1586364061
transform 1 0 39652 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40204 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39376 0 1 20128
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 39560 0 -1 21216
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_34_429
timestamp 1586364061
transform 1 0 40572 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_428
timestamp 1586364061
transform 1 0 40480 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_444
timestamp 1586364061
transform 1 0 40388 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_432
timestamp 1586364061
transform 1 0 40848 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40664 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41124 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41032 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41216 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41308 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_12  FILLER_34_446
timestamp 1586364061
transform 1 0 42136 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_452
timestamp 1586364061
transform 1 0 42688 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_449
timestamp 1586364061
transform 1 0 42412 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_445
timestamp 1586364061
transform 1 0 42044 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42504 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42872 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_456
timestamp 1586364061
transform 1 0 43056 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_468
timestamp 1586364061
transform 1 0 44160 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_469
timestamp 1586364061
transform 1 0 44252 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43240 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_453
timestamp 1586364061
transform 1 0 43240 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43424 0 1 20128
box -38 -48 866 592
use scs8hd_decap_12  FILLER_34_479
timestamp 1586364061
transform 1 0 45172 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_480
timestamp 1586364061
transform 1 0 45264 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_473
timestamp 1586364061
transform 1 0 44620 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44436 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44896 0 -1 21216
box -38 -48 314 592
use scs8hd_conb_1  _651_
timestamp 1586364061
transform 1 0 44988 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45448 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_445
timestamp 1586364061
transform 1 0 46000 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_484
timestamp 1586364061
transform 1 0 45632 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_33_489
timestamp 1586364061
transform 1 0 46092 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_501
timestamp 1586364061
transform 1 0 47196 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_491
timestamp 1586364061
transform 1 0 46276 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_503
timestamp 1586364061
transform 1 0 47380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 48852 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 48852 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_513
timestamp 1586364061
transform 1 0 48300 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_515
timestamp 1586364061
transform 1 0 48484 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_35_12
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_9
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _245_
timestamp 1586364061
transform 1 0 2300 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_20
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_16
timestamp 1586364061
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__245__A
timestamp 1586364061
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_24
timestamp 1586364061
transform 1 0 3312 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__265__A
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_30
timestamp 1586364061
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_49
timestamp 1586364061
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_454
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_76
timestamp 1586364061
transform 1 0 8096 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__300__A
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__252__A
timestamp 1586364061
transform 1 0 8280 0 1 21216
box -38 -48 222 592
use scs8hd_or2_4  _252_
timestamp 1586364061
transform 1 0 8464 0 1 21216
box -38 -48 682 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__252__B
timestamp 1586364061
transform 1 0 9292 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__253__A
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_91
timestamp 1586364061
transform 1 0 9476 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_101
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__339__A
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_455
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_126
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_130
timestamp 1586364061
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__565__A
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_134
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__565__B
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 13892 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_150
timestamp 1586364061
transform 1 0 14904 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_154
timestamp 1586364061
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_456
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_167
timestamp 1586364061
transform 1 0 16468 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _489_
timestamp 1586364061
transform 1 0 19688 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__489__A
timestamp 1586364061
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_193
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_198
timestamp 1586364061
transform 1 0 19320 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21804 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_217
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_221
timestamp 1586364061
transform 1 0 21436 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_236
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_240
timestamp 1586364061
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use scs8hd_or4_4  _515_
timestamp 1586364061
transform 1 0 25208 0 1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_457
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__515__C
timestamp 1586364061
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__515__D
timestamp 1586364061
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_254
timestamp 1586364061
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_258
timestamp 1586364061
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use scs8hd_or4_4  _460_
timestamp 1586364061
transform 1 0 27508 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__460__B
timestamp 1586364061
transform 1 0 27324 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__334__A
timestamp 1586364061
transform 1 0 26956 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__515__A
timestamp 1586364061
transform 1 0 26220 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__460__A
timestamp 1586364061
transform 1 0 26588 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_271
timestamp 1586364061
transform 1 0 26036 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_275
timestamp 1586364061
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_279
timestamp 1586364061
transform 1 0 26772 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_283
timestamp 1586364061
transform 1 0 27140 0 1 21216
box -38 -48 222 592
use scs8hd_or4_4  _409_
timestamp 1586364061
transform 1 0 29256 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_458
timestamp 1586364061
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__471__B
timestamp 1586364061
transform 1 0 28520 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__409__D
timestamp 1586364061
transform 1 0 28980 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__406__A
timestamp 1586364061
transform 1 0 30452 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_296
timestamp 1586364061
transform 1 0 28336 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_300
timestamp 1586364061
transform 1 0 28704 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_315
timestamp 1586364061
transform 1 0 30084 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_321
timestamp 1586364061
transform 1 0 30636 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _382_
timestamp 1586364061
transform 1 0 30820 0 1 21216
box -38 -48 314 592
use scs8hd_nor2_4  _404_
timestamp 1586364061
transform 1 0 32108 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33120 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__404__A
timestamp 1586364061
transform 1 0 31924 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__382__A
timestamp 1586364061
transform 1 0 31280 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_326
timestamp 1586364061
transform 1 0 31096 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_330
timestamp 1586364061
transform 1 0 31464 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_334
timestamp 1586364061
transform 1 0 31832 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_346
timestamp 1586364061
transform 1 0 32936 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_357
timestamp 1586364061
transform 1 0 33948 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_350
timestamp 1586364061
transform 1 0 33304 0 1 21216
box -38 -48 406 592
use scs8hd_conb_1  _650_
timestamp 1586364061
transform 1 0 33672 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_367
timestamp 1586364061
transform 1 0 34868 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_365
timestamp 1586364061
transform 1 0 34684 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_361
timestamp 1586364061
transform 1 0 34316 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34500 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34132 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_459
timestamp 1586364061
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35052 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35236 0 1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36800 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37812 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36616 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_380
timestamp 1586364061
transform 1 0 36064 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_384
timestamp 1586364061
transform 1 0 36432 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_397
timestamp 1586364061
transform 1 0 37628 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_401
timestamp 1586364061
transform 1 0 37996 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_406
timestamp 1586364061
transform 1 0 38456 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__392__A
timestamp 1586364061
transform 1 0 38272 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__389__A
timestamp 1586364061
transform 1 0 38640 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _389_
timestamp 1586364061
transform 1 0 38824 0 1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_35_423
timestamp 1586364061
transform 1 0 40020 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_419
timestamp 1586364061
transform 1 0 39652 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__389__B
timestamp 1586364061
transform 1 0 39836 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_460
timestamp 1586364061
transform 1 0 40388 0 1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 40480 0 1 21216
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42228 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42044 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_439
timestamp 1586364061
transform 1 0 41492 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_443
timestamp 1586364061
transform 1 0 41860 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_456
timestamp 1586364061
transform 1 0 43056 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43792 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43332 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__397__A
timestamp 1586364061
transform 1 0 44804 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_461
timestamp 1586364061
transform 1 0 43516 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_473
timestamp 1586364061
transform 1 0 44620 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_477
timestamp 1586364061
transform 1 0 44988 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_461
timestamp 1586364061
transform 1 0 46000 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_485
timestamp 1586364061
transform 1 0 45724 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_489
timestamp 1586364061
transform 1 0 46092 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_501
timestamp 1586364061
transform 1 0 47196 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 48852 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_513
timestamp 1586364061
transform 1 0 48300 0 1 21216
box -38 -48 314 592
use scs8hd_inv_8  _240_
timestamp 1586364061
transform 1 0 2024 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_9
timestamp 1586364061
transform 1 0 1932 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_19
timestamp 1586364061
transform 1 0 2852 0 -1 22304
box -38 -48 1142 592
use scs8hd_buf_1  _265_
timestamp 1586364061
transform 1 0 4140 0 -1 22304
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_462
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__561__A
timestamp 1586364061
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_36
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_40
timestamp 1586364061
transform 1 0 4784 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_1  _300_
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__305__A
timestamp 1586364061
transform 1 0 8188 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__296__D
timestamp 1586364061
transform 1 0 6348 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_55
timestamp 1586364061
transform 1 0 6164 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_59
timestamp 1586364061
transform 1 0 6532 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_36_72
timestamp 1586364061
transform 1 0 7728 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_76
timestamp 1586364061
transform 1 0 8096 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_79
timestamp 1586364061
transform 1 0 8372 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_1  _253_
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_463
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__270__A
timestamp 1586364061
transform 1 0 10580 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__270__B
timestamp 1586364061
transform 1 0 10948 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_83
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_91
timestamp 1586364061
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_96
timestamp 1586364061
transform 1 0 9936 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_1  _339_
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 314 592
use scs8hd_nor2_4  _565_
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_4  FILLER_36_109
timestamp 1586364061
transform 1 0 11132 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_116
timestamp 1586364061
transform 1 0 11776 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_124
timestamp 1586364061
transform 1 0 12512 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_134
timestamp 1586364061
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_464
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__566__B
timestamp 1586364061
transform 1 0 13616 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_138
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_12  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_175
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_465
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_194
timestamp 1586364061
transform 1 0 18952 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_36_201
timestamp 1586364061
transform 1 0 19596 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_205
timestamp 1586364061
transform 1 0 19964 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_208
timestamp 1586364061
transform 1 0 20240 0 -1 22304
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22908 0 -1 22304
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__491__B
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__484__A
timestamp 1586364061
transform 1 0 22356 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_224
timestamp 1586364061
transform 1 0 21712 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_229
timestamp 1586364061
transform 1 0 22172 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_233
timestamp 1586364061
transform 1 0 22540 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__515__B
timestamp 1586364061
transform 1 0 25668 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_248
timestamp 1586364061
transform 1 0 23920 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_265
timestamp 1586364061
transform 1 0 25484 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_269
timestamp 1586364061
transform 1 0 25852 0 -1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__503__A
timestamp 1586364061
transform 1 0 26680 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_466
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_285
timestamp 1586364061
transform 1 0 27324 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_280
timestamp 1586364061
transform 1 0 26864 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__460__C
timestamp 1586364061
transform 1 0 27508 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_1  _334_
timestamp 1586364061
transform 1 0 27048 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_289
timestamp 1586364061
transform 1 0 27692 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__471__A
timestamp 1586364061
transform 1 0 27876 0 -1 22304
box -38 -48 222 592
use scs8hd_or4_4  _471_
timestamp 1586364061
transform 1 0 28060 0 -1 22304
box -38 -48 866 592
use scs8hd_nor2_4  _406_
timestamp 1586364061
transform 1 0 30452 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__409__B
timestamp 1586364061
transform 1 0 29256 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__409__C
timestamp 1586364061
transform 1 0 29624 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__406__B
timestamp 1586364061
transform 1 0 30268 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_302
timestamp 1586364061
transform 1 0 28888 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_308
timestamp 1586364061
transform 1 0 29440 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_312
timestamp 1586364061
transform 1 0 29808 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_316
timestamp 1586364061
transform 1 0 30176 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32752 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_467
timestamp 1586364061
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32292 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_328
timestamp 1586364061
transform 1 0 31280 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_337
timestamp 1586364061
transform 1 0 32108 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_341
timestamp 1586364061
transform 1 0 32476 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_347
timestamp 1586364061
transform 1 0 33028 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33764 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35236 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_364
timestamp 1586364061
transform 1 0 34592 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_370
timestamp 1586364061
transform 1 0 35144 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_373
timestamp 1586364061
transform 1 0 35420 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_468
timestamp 1586364061
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_377
timestamp 1586364061
transform 1 0 35788 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_389
timestamp 1586364061
transform 1 0 36892 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_4  FILLER_36_401
timestamp 1586364061
transform 1 0 37996 0 -1 22304
box -38 -48 406 592
use scs8hd_nor2_4  _392_
timestamp 1586364061
transform 1 0 38732 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__395__A
timestamp 1586364061
transform 1 0 38364 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40480 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_407
timestamp 1586364061
transform 1 0 38548 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_418
timestamp 1586364061
transform 1 0 39560 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_426
timestamp 1586364061
transform 1 0 40296 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41216 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42228 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_430
timestamp 1586364061
transform 1 0 40664 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_445
timestamp 1586364061
transform 1 0 42044 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_449
timestamp 1586364061
transform 1 0 42412 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_455
timestamp 1586364061
transform 1 0 42964 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_1  _397_
timestamp 1586364061
transform 1 0 44344 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_469
timestamp 1586364061
transform 1 0 43240 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43792 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44160 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_462
timestamp 1586364061
transform 1 0 43608 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_466
timestamp 1586364061
transform 1 0 43976 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_473
timestamp 1586364061
transform 1 0 44620 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_485
timestamp 1586364061
transform 1 0 45724 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_497
timestamp 1586364061
transform 1 0 46828 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_509
timestamp 1586364061
transform 1 0 47932 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 48852 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_515
timestamp 1586364061
transform 1 0 48484 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_8  _237_
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__258__A
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__561__B
timestamp 1586364061
transform 1 0 3496 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_37_20
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_24
timestamp 1586364061
transform 1 0 3312 0 1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _561_
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__296__C
timestamp 1586364061
transform 1 0 5612 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__264__A
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__296__B
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__264__B
timestamp 1586364061
transform 1 0 3864 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_28
timestamp 1586364061
transform 1 0 3680 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_32
timestamp 1586364061
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_45
timestamp 1586364061
transform 1 0 5244 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_55
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__296__A
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_470
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_buf_1  _297_
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_65
timestamp 1586364061
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__336__A
timestamp 1586364061
transform 1 0 7268 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_69
timestamp 1586364061
transform 1 0 7452 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__268__A
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__305__B
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_79
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use scs8hd_or2_4  _268_
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 682 592
use scs8hd_or2_4  _270_
timestamp 1586364061
transform 1 0 10580 0 1 22304
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__268__B
timestamp 1586364061
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__254__A
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__254__B
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_88
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_96
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_100
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__271__B
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__271__A
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_129
timestamp 1586364061
transform 1 0 12972 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__566__A
timestamp 1586364061
transform 1 0 12788 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_471
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 13340 0 1 22304
box -38 -48 1050 592
use scs8hd_buf_1  _272_
timestamp 1586364061
transform 1 0 15088 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__272__A
timestamp 1586364061
transform 1 0 15548 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_144
timestamp 1586364061
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_148
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_155
timestamp 1586364061
transform 1 0 15364 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_169
timestamp 1586364061
transform 1 0 16652 0 1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_37_163
timestamp 1586364061
transform 1 0 16100 0 1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_472
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_inv_8  _615_
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20056 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19872 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_193
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_197
timestamp 1586364061
transform 1 0 19228 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_203
timestamp 1586364061
transform 1 0 19780 0 1 22304
box -38 -48 130 592
use scs8hd_nor2_4  _491_
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__491__A
timestamp 1586364061
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_217
timestamp 1586364061
transform 1 0 21068 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_221
timestamp 1586364061
transform 1 0 21436 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_473
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_buf_1  _343_
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_248
timestamp 1586364061
transform 1 0 23920 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_252
timestamp 1586364061
transform 1 0 24288 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__343__A
timestamp 1586364061
transform 1 0 24104 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  _337_
timestamp 1586364061
transform 1 0 24656 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_259
timestamp 1586364061
transform 1 0 24932 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_263
timestamp 1586364061
transform 1 0 25300 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__337__A
timestamp 1586364061
transform 1 0 25116 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  _314_
timestamp 1586364061
transform 1 0 25668 0 1 22304
box -38 -48 314 592
use scs8hd_nor2_4  _503_
timestamp 1586364061
transform 1 0 26680 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 27968 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__314__A
timestamp 1586364061
transform 1 0 26128 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__325__A
timestamp 1586364061
transform 1 0 26496 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_270
timestamp 1586364061
transform 1 0 25944 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_274
timestamp 1586364061
transform 1 0 26312 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_287
timestamp 1586364061
transform 1 0 27508 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_291
timestamp 1586364061
transform 1 0 27876 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_294
timestamp 1586364061
transform 1 0 28152 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_302
timestamp 1586364061
transform 1 0 28888 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_298
timestamp 1586364061
transform 1 0 28520 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28336 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__409__A
timestamp 1586364061
transform 1 0 28980 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_474
timestamp 1586364061
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_309
timestamp 1586364061
transform 1 0 29532 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__405__B
timestamp 1586364061
transform 1 0 29900 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  _472_
timestamp 1586364061
transform 1 0 29256 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_315
timestamp 1586364061
transform 1 0 30084 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30268 0 1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _405_
timestamp 1586364061
transform 1 0 30452 0 1 22304
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 32016 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 31832 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 31464 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_328
timestamp 1586364061
transform 1 0 31280 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_332
timestamp 1586364061
transform 1 0 31648 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_347
timestamp 1586364061
transform 1 0 33028 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_351
timestamp 1586364061
transform 1 0 33396 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33212 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33580 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_358
timestamp 1586364061
transform 1 0 34040 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_362
timestamp 1586364061
transform 1 0 34408 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_475
timestamp 1586364061
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_370
timestamp 1586364061
transform 1 0 35144 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_374
timestamp 1586364061
transform 1 0 35512 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_378
timestamp 1586364061
transform 1 0 35880 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35696 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36064 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36248 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_385
timestamp 1586364061
transform 1 0 36524 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36708 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_389
timestamp 1586364061
transform 1 0 36892 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__394__B
timestamp 1586364061
transform 1 0 37076 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37260 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_396
timestamp 1586364061
transform 1 0 37536 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37720 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_400
timestamp 1586364061
transform 1 0 37904 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__394__A
timestamp 1586364061
transform 1 0 38088 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_404
timestamp 1586364061
transform 1 0 38272 0 1 22304
box -38 -48 130 592
use scs8hd_nor2_4  _395_
timestamp 1586364061
transform 1 0 38364 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  FILLER_37_422
timestamp 1586364061
transform 1 0 39928 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_418
timestamp 1586364061
transform 1 0 39560 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_414
timestamp 1586364061
transform 1 0 39192 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39744 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 39376 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40204 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_476
timestamp 1586364061
transform 1 0 40388 0 1 22304
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_435
timestamp 1586364061
transform 1 0 41124 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_431
timestamp 1586364061
transform 1 0 40756 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41308 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41492 0 1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_37_446
timestamp 1586364061
transform 1 0 42136 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_442
timestamp 1586364061
transform 1 0 41768 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41952 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_452
timestamp 1586364061
transform 1 0 42688 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42504 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42872 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43056 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44896 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44068 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_465
timestamp 1586364061
transform 1 0 43884 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_469
timestamp 1586364061
transform 1 0 44252 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_475
timestamp 1586364061
transform 1 0 44804 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_478
timestamp 1586364061
transform 1 0 45080 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_477
timestamp 1586364061
transform 1 0 46000 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_486
timestamp 1586364061
transform 1 0 45816 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_489
timestamp 1586364061
transform 1 0 46092 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_501
timestamp 1586364061
transform 1 0 47196 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 48852 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_513
timestamp 1586364061
transform 1 0 48300 0 1 22304
box -38 -48 314 592
use scs8hd_buf_1  _258_
timestamp 1586364061
transform 1 0 2300 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__246__B
timestamp 1586364061
transform 1 0 2944 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__C
timestamp 1586364061
transform 1 0 3312 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_11
timestamp 1586364061
transform 1 0 2116 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_16
timestamp 1586364061
transform 1 0 2576 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_22
timestamp 1586364061
transform 1 0 3128 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_26
timestamp 1586364061
transform 1 0 3496 0 -1 23392
box -38 -48 314 592
use scs8hd_or2_4  _264_
timestamp 1586364061
transform 1 0 4232 0 -1 23392
box -38 -48 682 592
use scs8hd_or4_4  _296_
timestamp 1586364061
transform 1 0 5612 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_478
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__263__B
timestamp 1586364061
transform 1 0 5060 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__B
timestamp 1586364061
transform 1 0 5428 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__249__C
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_41
timestamp 1586364061
transform 1 0 4876 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_45
timestamp 1586364061
transform 1 0 5244 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_58
timestamp 1586364061
transform 1 0 6440 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__263__A
timestamp 1586364061
transform 1 0 6624 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_69
timestamp 1586364061
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_62
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__297__A
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_1  _336_
timestamp 1586364061
transform 1 0 7176 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_73
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__255__B
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__299__A
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 222 592
use scs8hd_or2_4  _305_
timestamp 1586364061
transform 1 0 8188 0 -1 23392
box -38 -48 682 592
use scs8hd_or2_4  _254_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_479
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__282__B
timestamp 1586364061
transform 1 0 9108 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__274__A
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_89
timestamp 1586364061
transform 1 0 9292 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_100
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_106
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 222 592
use scs8hd_or2_4  _271_
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 682 592
use scs8hd_nor2_4  _566_
timestamp 1586364061
transform 1 0 13156 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__283__B
timestamp 1586364061
transform 1 0 12236 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_115
timestamp 1586364061
transform 1 0 11684 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_8  FILLER_38_123
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_480
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__287__B
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_144
timestamp 1586364061
transform 1 0 14352 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_152
timestamp 1586364061
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_158
timestamp 1586364061
transform 1 0 15640 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__615__A
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_4  FILLER_38_180
timestamp 1586364061
transform 1 0 17664 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_186
timestamp 1586364061
transform 1 0 18216 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_481
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_197
timestamp 1586364061
transform 1 0 19228 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_38_209
timestamp 1586364061
transform 1 0 20332 0 -1 23392
box -38 -48 314 592
use scs8hd_buf_1  _484_
timestamp 1586364061
transform 1 0 21896 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22908 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_218
timestamp 1586364061
transform 1 0 21160 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_222
timestamp 1586364061
transform 1 0 21528 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_229
timestamp 1586364061
transform 1 0 22172 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_246
timestamp 1586364061
transform 1 0 23736 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_1  _325_
timestamp 1586364061
transform 1 0 26680 0 -1 23392
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 27968 0 -1 23392
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_482
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__503__B
timestamp 1586364061
transform 1 0 27140 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_281
timestamp 1586364061
transform 1 0 26956 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_285
timestamp 1586364061
transform 1 0 27324 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_291
timestamp 1586364061
transform 1 0 27876 0 -1 23392
box -38 -48 130 592
use scs8hd_buf_1  _495_
timestamp 1586364061
transform 1 0 29716 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__405__A
timestamp 1586364061
transform 1 0 30452 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__472__A
timestamp 1586364061
transform 1 0 29256 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_303
timestamp 1586364061
transform 1 0 28980 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_308
timestamp 1586364061
transform 1 0 29440 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_314
timestamp 1586364061
transform 1 0 29992 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_318
timestamp 1586364061
transform 1 0 30360 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_321
timestamp 1586364061
transform 1 0 30636 0 -1 23392
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 23392
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30820 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_483
timestamp 1586364061
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31280 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_326
timestamp 1586364061
transform 1 0 31096 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_330
timestamp 1586364061
transform 1 0 31464 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_38_348
timestamp 1586364061
transform 1 0 33120 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34868 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35236 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35604 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_352
timestamp 1586364061
transform 1 0 33488 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_365
timestamp 1586364061
transform 1 0 34684 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_369
timestamp 1586364061
transform 1 0 35052 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_373
timestamp 1586364061
transform 1 0 35420 0 -1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _394_
timestamp 1586364061
transform 1 0 37812 0 -1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_484
timestamp 1586364061
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_377
timestamp 1586364061
transform 1 0 35788 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_389
timestamp 1586364061
transform 1 0 36892 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_393
timestamp 1586364061
transform 1 0 37260 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_398
timestamp 1586364061
transform 1 0 37720 0 -1 23392
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 39376 0 -1 23392
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__395__B
timestamp 1586364061
transform 1 0 38824 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_408
timestamp 1586364061
transform 1 0 38640 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_412
timestamp 1586364061
transform 1 0 39008 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_6  FILLER_38_427
timestamp 1586364061
transform 1 0 40388 0 -1 23392
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41124 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40940 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_444
timestamp 1586364061
transform 1 0 41952 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44896 0 -1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_485
timestamp 1586364061
transform 1 0 43240 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_468
timestamp 1586364061
transform 1 0 44160 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_479
timestamp 1586364061
transform 1 0 45172 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_491
timestamp 1586364061
transform 1 0 46276 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_503
timestamp 1586364061
transform 1 0 47380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 48852 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_515
timestamp 1586364061
transform 1 0 48484 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_inv_8  _238_
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 866 592
use scs8hd_buf_1  _236_
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_16
timestamp 1586364061
transform 1 0 2576 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_16
timestamp 1586364061
transform 1 0 2576 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_12
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__A
timestamp 1586364061
transform 1 0 2760 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_26
timestamp 1586364061
transform 1 0 3496 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_22
timestamp 1586364061
transform 1 0 3128 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__247__A
timestamp 1586364061
transform 1 0 3312 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__D
timestamp 1586364061
transform 1 0 2944 0 -1 24480
box -38 -48 222 592
use scs8hd_or4_4  _246_
timestamp 1586364061
transform 1 0 2944 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_29
timestamp 1586364061
transform 1 0 3772 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__259__A
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__249__A
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__249__D
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_494
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_or4_4  _249_
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_45
timestamp 1586364061
transform 1 0 5244 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_41
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_38
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__263__C
timestamp 1586364061
transform 1 0 5060 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__249__B
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use scs8hd_or3_4  _263_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__C
timestamp 1586364061
transform 1 0 5428 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_or3_4  _241_
timestamp 1586364061
transform 1 0 5612 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_62
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_58
timestamp 1586364061
transform 1 0 6440 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_55
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__595__B
timestamp 1586364061
transform 1 0 6624 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__255__A
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_486
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_73
timestamp 1586364061
transform 1 0 7820 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__595__A
timestamp 1586364061
transform 1 0 6992 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__299__C
timestamp 1586364061
transform 1 0 6992 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__299__B
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_or4_4  _299_
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 866 592
use scs8hd_or2_4  _255_
timestamp 1586364061
transform 1 0 7176 0 -1 24480
box -38 -48 682 592
use scs8hd_decap_4  FILLER_40_77
timestamp 1586364061
transform 1 0 8188 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_79
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__299__D
timestamp 1586364061
transform 1 0 8004 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_89
timestamp 1586364061
transform 1 0 9292 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_83
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__333__A
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__282__C
timestamp 1586364061
transform 1 0 9108 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__282__A
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use scs8hd_buf_1  _333_
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 314 592
use scs8hd_or3_4  _282_
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_98
timestamp 1586364061
transform 1 0 10120 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_100
timestamp 1586364061
transform 1 0 10304 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_96
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__303__A
timestamp 1586364061
transform 1 0 10304 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__275__B
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_495
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_1  _303_
timestamp 1586364061
transform 1 0 9844 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_102
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__274__B
timestamp 1586364061
transform 1 0 10488 0 1 23392
box -38 -48 222 592
use scs8hd_or2_4  _275_
timestamp 1586364061
transform 1 0 10856 0 -1 24480
box -38 -48 682 592
use scs8hd_or2_4  _274_
timestamp 1586364061
transform 1 0 10672 0 1 23392
box -38 -48 682 592
use scs8hd_decap_8  FILLER_40_113
timestamp 1586364061
transform 1 0 11500 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__275__A
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_119
timestamp 1586364061
transform 1 0 12052 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__283__A
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_487
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_buf_1  _342_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 314 592
use scs8hd_or2_4  _283_
timestamp 1586364061
transform 1 0 12236 0 -1 24480
box -38 -48 682 592
use scs8hd_fill_2  FILLER_40_132
timestamp 1586364061
transform 1 0 13248 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_128
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_130
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_126
timestamp 1586364061
transform 1 0 12696 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__567__B
timestamp 1586364061
transform 1 0 13064 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__342__A
timestamp 1586364061
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__292__B
timestamp 1586364061
transform 1 0 13432 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__287__A
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_143
timestamp 1586364061
transform 1 0 14260 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_145
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__567__A
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _567_
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 866 592
use scs8hd_or2_4  _287_
timestamp 1586364061
transform 1 0 13616 0 -1 24480
box -38 -48 682 592
use scs8hd_fill_2  FILLER_40_151
timestamp 1586364061
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_147
timestamp 1586364061
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_149
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__568__B
timestamp 1586364061
transform 1 0 14812 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14996 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_496
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15180 0 1 23392
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_40_165
timestamp 1586364061
transform 1 0 16284 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_168
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_164
timestamp 1586364061
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_174
timestamp 1586364061
transform 1 0 17112 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_171
timestamp 1586364061
transform 1 0 16836 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__612__A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 -1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 23392
box -38 -48 314 592
use scs8hd_inv_8  _612_
timestamp 1586364061
transform 1 0 17296 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_185
timestamp 1586364061
transform 1 0 18124 0 -1 24480
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__613__A
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_488
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_inv_8  _613_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_40_196
timestamp 1586364061
transform 1 0 19136 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_197
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__327__A
timestamp 1586364061
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use scs8hd_buf_1  _327_
timestamp 1586364061
transform 1 0 18860 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_206
timestamp 1586364061
transform 1 0 20056 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_204
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 20056 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__486__B
timestamp 1586364061
transform 1 0 19872 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__487__A
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 19596 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_497
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 866 592
use scs8hd_fill_1  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_221
timestamp 1586364061
transform 1 0 21436 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_233
timestamp 1586364061
transform 1 0 22540 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_225
timestamp 1586364061
transform 1 0 21804 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_6  FILLER_39_225
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_240
timestamp 1586364061
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_236
timestamp 1586364061
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_4  FILLER_40_248
timestamp 1586364061
transform 1 0 23920 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_244
timestamp 1586364061
transform 1 0 23552 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_250
timestamp 1586364061
transform 1 0 24104 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23736 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_489
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_252
timestamp 1586364061
transform 1 0 24288 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_264
timestamp 1586364061
transform 1 0 25392 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_267
timestamp 1586364061
transform 1 0 25668 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_279
timestamp 1586364061
transform 1 0 26772 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_272
timestamp 1586364061
transform 1 0 26128 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_271
timestamp 1586364061
transform 1 0 26036 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__340__A
timestamp 1586364061
transform 1 0 26128 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__502__A
timestamp 1586364061
transform 1 0 26496 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_498
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_nor2_4  _502_
timestamp 1586364061
transform 1 0 26680 0 1 23392
box -38 -48 866 592
use scs8hd_buf_1  _340_
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_290
timestamp 1586364061
transform 1 0 27784 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_287
timestamp 1586364061
transform 1 0 27508 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_283
timestamp 1586364061
transform 1 0 27140 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_291
timestamp 1586364061
transform 1 0 27876 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_287
timestamp 1586364061
transform 1 0 27508 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27600 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__502__B
timestamp 1586364061
transform 1 0 26956 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 27968 0 1 23392
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 27968 0 -1 24480
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_39_294
timestamp 1586364061
transform 1 0 28152 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_303
timestamp 1586364061
transform 1 0 28980 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_39_304
timestamp 1586364061
transform 1 0 29072 0 1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_39_298
timestamp 1586364061
transform 1 0 28520 0 1 23392
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28336 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_490
timestamp 1586364061
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_312
timestamp 1586364061
transform 1 0 29808 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_308
timestamp 1586364061
transform 1 0 29440 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_313
timestamp 1586364061
transform 1 0 29900 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_39_310
timestamp 1586364061
transform 1 0 29624 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_306
timestamp 1586364061
transform 1 0 29256 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29624 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29256 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__495__A
timestamp 1586364061
transform 1 0 29716 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_318
timestamp 1586364061
transform 1 0 30360 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_319
timestamp 1586364061
transform 1 0 30452 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30636 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 24480
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30176 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_328
timestamp 1586364061
transform 1 0 31280 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_323
timestamp 1586364061
transform 1 0 30820 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31464 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31004 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31188 0 1 23392
box -38 -48 866 592
use scs8hd_decap_3  FILLER_40_337
timestamp 1586364061
transform 1 0 32108 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_332
timestamp 1586364061
transform 1 0 31648 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_340
timestamp 1586364061
transform 1 0 32384 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_336
timestamp 1586364061
transform 1 0 32016 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32200 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32384 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_499
timestamp 1586364061
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_347
timestamp 1586364061
transform 1 0 33028 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_342
timestamp 1586364061
transform 1 0 32568 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_346
timestamp 1586364061
transform 1 0 32936 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32752 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32752 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_40_358
timestamp 1586364061
transform 1 0 34040 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_4  FILLER_40_351
timestamp 1586364061
transform 1 0 33396 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_358
timestamp 1586364061
transform 1 0 34040 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 -1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_362
timestamp 1586364061
transform 1 0 34408 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_491
timestamp 1586364061
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34776 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_375
timestamp 1586364061
transform 1 0 35604 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_380
timestamp 1586364061
transform 1 0 36064 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_376
timestamp 1586364061
transform 1 0 35696 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36248 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36340 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_40_390
timestamp 1586364061
transform 1 0 36984 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_386
timestamp 1586364061
transform 1 0 36616 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_393
timestamp 1586364061
transform 1 0 37260 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36800 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_401
timestamp 1586364061
transform 1 0 37996 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_396
timestamp 1586364061
transform 1 0 37536 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_400
timestamp 1586364061
transform 1 0 37904 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_397
timestamp 1586364061
transform 1 0 37628 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37720 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_500
timestamp 1586364061
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37996 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_413
timestamp 1586364061
transform 1 0 39100 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_409
timestamp 1586364061
transform 1 0 38732 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_405
timestamp 1586364061
transform 1 0 38364 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_410
timestamp 1586364061
transform 1 0 38824 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38548 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38180 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 39192 0 1 23392
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 39192 0 -1 24480
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_40_425
timestamp 1586364061
transform 1 0 40204 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_424
timestamp 1586364061
transform 1 0 40112 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_420
timestamp 1586364061
transform 1 0 39744 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_416
timestamp 1586364061
transform 1 0 39376 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39560 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_428
timestamp 1586364061
transform 1 0 40480 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_492
timestamp 1586364061
transform 1 0 40388 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40756 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40940 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40940 0 1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_448
timestamp 1586364061
transform 1 0 42320 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_40_442
timestamp 1586364061
transform 1 0 41768 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_446
timestamp 1586364061
transform 1 0 42136 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_442
timestamp 1586364061
transform 1 0 41768 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41952 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42136 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_456
timestamp 1586364061
transform 1 0 43056 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_452
timestamp 1586364061
transform 1 0 42688 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42504 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42872 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43056 0 1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_468
timestamp 1586364061
transform 1 0 44160 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_469
timestamp 1586364061
transform 1 0 44252 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_465
timestamp 1586364061
transform 1 0 43884 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44068 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_501
timestamp 1586364061
transform 1 0 43240 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_12  FILLER_40_479
timestamp 1586364061
transform 1 0 45172 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_480
timestamp 1586364061
transform 1 0 45264 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_476
timestamp 1586364061
transform 1 0 44896 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45080 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44620 0 1 23392
box -38 -48 314 592
use scs8hd_buf_1  _410_
timestamp 1586364061
transform 1 0 44896 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__410__A
timestamp 1586364061
transform 1 0 45448 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_493
timestamp 1586364061
transform 1 0 46000 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_484
timestamp 1586364061
transform 1 0 45632 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_39_489
timestamp 1586364061
transform 1 0 46092 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_501
timestamp 1586364061
transform 1 0 47196 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_491
timestamp 1586364061
transform 1 0 46276 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_503
timestamp 1586364061
transform 1 0 47380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 48852 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 48852 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_513
timestamp 1586364061
transform 1 0 48300 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_515
timestamp 1586364061
transform 1 0 48484 0 -1 24480
box -38 -48 130 592
use scs8hd_inv_8  _235_
timestamp 1586364061
transform 1 0 2392 0 1 24480
box -38 -48 866 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 2208 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__259__B
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 1840 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_7
timestamp 1586364061
transform 1 0 1748 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_10
timestamp 1586364061
transform 1 0 2024 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_23
timestamp 1586364061
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__260__A
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 222 592
use scs8hd_or3_4  _259_
timestamp 1586364061
transform 1 0 3956 0 1 24480
box -38 -48 866 592
use scs8hd_decap_3  FILLER_41_44
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_40
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__259__C
timestamp 1586364061
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_49
timestamp 1586364061
transform 1 0 5612 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 5428 0 1 24480
box -38 -48 222 592
use scs8hd_buf_1  _256_
timestamp 1586364061
transform 1 0 5704 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__256__A
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__B
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_502
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__293__B
timestamp 1586364061
transform 1 0 7084 0 1 24480
box -38 -48 222 592
use scs8hd_or2_4  _293_
timestamp 1586364061
transform 1 0 7268 0 1 24480
box -38 -48 682 592
use scs8hd_fill_2  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__286__B
timestamp 1586364061
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_78
timestamp 1586364061
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__286__C
timestamp 1586364061
transform 1 0 8464 0 1 24480
box -38 -48 222 592
use scs8hd_or3_4  _286_
timestamp 1586364061
transform 1 0 8648 0 1 24480
box -38 -48 866 592
use scs8hd_or2_4  _302_
timestamp 1586364061
transform 1 0 10396 0 1 24480
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__302__A
timestamp 1586364061
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__598__A
timestamp 1586364061
transform 1 0 9660 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_91
timestamp 1586364061
transform 1 0 9476 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_95
timestamp 1586364061
transform 1 0 9844 0 1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_41_112
timestamp 1586364061
transform 1 0 11408 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_108
timestamp 1586364061
transform 1 0 11040 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__302__B
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__279__A
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__279__B
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_503
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__290__A
timestamp 1586364061
transform 1 0 12604 0 1 24480
box -38 -48 222 592
use scs8hd_or2_4  _290_
timestamp 1586364061
transform 1 0 12788 0 1 24480
box -38 -48 682 592
use scs8hd_fill_2  FILLER_41_134
timestamp 1586364061
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use scs8hd_buf_1  _330_
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 314 592
use scs8hd_nor2_4  _568_
timestamp 1586364061
transform 1 0 14168 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__330__A
timestamp 1586364061
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__290__B
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__292__A
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__288__A
timestamp 1586364061
transform 1 0 15180 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_138
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_151
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_155
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_162
timestamp 1586364061
transform 1 0 16008 0 1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_41_169
timestamp 1586364061
transform 1 0 16652 0 1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_41_166
timestamp 1586364061
transform 1 0 16376 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 16468 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_180
timestamp 1586364061
transform 1 0 17664 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__313__A
timestamp 1586364061
transform 1 0 17480 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_504
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_buf_1  _324_
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_187
timestamp 1586364061
transform 1 0 18308 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_195
timestamp 1586364061
transform 1 0 19044 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_191
timestamp 1586364061
transform 1 0 18676 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__487__B
timestamp 1586364061
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__486__A
timestamp 1586364061
transform 1 0 19228 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__324__A
timestamp 1586364061
transform 1 0 18492 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_199
timestamp 1586364061
transform 1 0 19412 0 1 24480
box -38 -48 130 592
use scs8hd_nor2_4  _487_
timestamp 1586364061
transform 1 0 19504 0 1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_41_213
timestamp 1586364061
transform 1 0 20700 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_209
timestamp 1586364061
transform 1 0 20332 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_226
timestamp 1586364061
transform 1 0 21896 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_230
timestamp 1586364061
transform 1 0 22264 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_234
timestamp 1586364061
transform 1 0 22632 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_240
timestamp 1586364061
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_505
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_254
timestamp 1586364061
transform 1 0 24472 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_258
timestamp 1586364061
transform 1 0 24840 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_262
timestamp 1586364061
transform 1 0 25208 0 1 24480
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26588 0 1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 27232 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_273
timestamp 1586364061
transform 1 0 26220 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_280
timestamp 1586364061
transform 1 0 26864 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_286
timestamp 1586364061
transform 1 0 27416 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_301
timestamp 1586364061
transform 1 0 28796 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_297
timestamp 1586364061
transform 1 0 28428 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28980 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_506
timestamp 1586364061
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_41_319
timestamp 1586364061
transform 1 0 30452 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_315
timestamp 1586364061
transform 1 0 30084 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30268 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30636 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30820 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_332
timestamp 1586364061
transform 1 0 31648 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_336
timestamp 1586364061
transform 1 0 32016 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_339
timestamp 1586364061
transform 1 0 32292 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_41_357
timestamp 1586364061
transform 1 0 33948 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_353
timestamp 1586364061
transform 1 0 33580 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_349
timestamp 1586364061
transform 1 0 33212 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33764 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33396 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_362
timestamp 1586364061
transform 1 0 34408 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_507
timestamp 1586364061
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 24480
box -38 -48 866 592
use scs8hd_buf_1  _386_
timestamp 1586364061
transform 1 0 37996 0 1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36248 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35880 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_376
timestamp 1586364061
transform 1 0 35696 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_380
timestamp 1586364061
transform 1 0 36064 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_393
timestamp 1586364061
transform 1 0 37260 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_397
timestamp 1586364061
transform 1 0 37628 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_404
timestamp 1586364061
transform 1 0 38272 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__386__A
timestamp 1586364061
transform 1 0 38456 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_408
timestamp 1586364061
transform 1 0 38640 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__387__A
timestamp 1586364061
transform 1 0 38824 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_412
timestamp 1586364061
transform 1 0 39008 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39192 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39376 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_419
timestamp 1586364061
transform 1 0 39652 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_423
timestamp 1586364061
transform 1 0 40020 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_428
timestamp 1586364061
transform 1 0 40480 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_508
timestamp 1586364061
transform 1 0 40388 0 1 24480
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42780 0 1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40940 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41952 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42596 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40756 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_442
timestamp 1586364061
transform 1 0 41768 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_446
timestamp 1586364061
transform 1 0 42136 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_450
timestamp 1586364061
transform 1 0 42504 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_41_456
timestamp 1586364061
transform 1 0 43056 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_461
timestamp 1586364061
transform 1 0 43516 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43332 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_467
timestamp 1586364061
transform 1 0 44068 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44252 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43792 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_471
timestamp 1586364061
transform 1 0 44436 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__428__A
timestamp 1586364061
transform 1 0 44620 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44804 0 1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_41_482
timestamp 1586364061
transform 1 0 45448 0 1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_41_478
timestamp 1586364061
transform 1 0 45080 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45264 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_509
timestamp 1586364061
transform 1 0 46000 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_489
timestamp 1586364061
transform 1 0 46092 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_501
timestamp 1586364061
transform 1 0 47196 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 48852 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_513
timestamp 1586364061
transform 1 0 48300 0 1 24480
box -38 -48 314 592
use scs8hd_buf_1  _239_
timestamp 1586364061
transform 1 0 1932 0 -1 25568
box -38 -48 314 592
use scs8hd_buf_1  _247_
timestamp 1586364061
transform 1 0 2944 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_8  FILLER_42_12
timestamp 1586364061
transform 1 0 2208 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_8  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 774 592
use scs8hd_or2_4  _242_
timestamp 1586364061
transform 1 0 5428 0 -1 25568
box -38 -48 682 592
use scs8hd_or2_4  _260_
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_510
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__260__B
timestamp 1586364061
transform 1 0 4876 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_39
timestamp 1586364061
transform 1 0 4692 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_43
timestamp 1586364061
transform 1 0 5060 0 -1 25568
box -38 -48 406 592
use scs8hd_nor2_4  _595_
timestamp 1586364061
transform 1 0 7452 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__295__A
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__293__A
timestamp 1586364061
transform 1 0 7268 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_54
timestamp 1586364061
transform 1 0 6072 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_60
timestamp 1586364061
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_64
timestamp 1586364061
transform 1 0 6992 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_78
timestamp 1586364061
transform 1 0 8280 0 -1 25568
box -38 -48 406 592
use scs8hd_nor2_4  _598_
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_511
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__286__A
timestamp 1586364061
transform 1 0 8648 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__598__B
timestamp 1586364061
transform 1 0 9384 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_84
timestamp 1586364061
transform 1 0 8832 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_42_102
timestamp 1586364061
transform 1 0 10488 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 774 592
use scs8hd_or2_4  _279_
timestamp 1586364061
transform 1 0 11776 0 -1 25568
box -38 -48 682 592
use scs8hd_nor2_4  _292_
timestamp 1586364061
transform 1 0 13432 0 -1 25568
box -38 -48 866 592
use scs8hd_fill_2  FILLER_42_114
timestamp 1586364061
transform 1 0 11592 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_123
timestamp 1586364061
transform 1 0 12420 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_131
timestamp 1586364061
transform 1 0 13156 0 -1 25568
box -38 -48 314 592
use scs8hd_buf_1  _288_
timestamp 1586364061
transform 1 0 15272 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_512
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__568__A
timestamp 1586364061
transform 1 0 14444 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_143
timestamp 1586364061
transform 1 0 14260 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_147
timestamp 1586364061
transform 1 0 14628 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_8  FILLER_42_157
timestamp 1586364061
transform 1 0 15548 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_1  _233_
timestamp 1586364061
transform 1 0 16468 0 -1 25568
box -38 -48 314 592
use scs8hd_buf_1  _313_
timestamp 1586364061
transform 1 0 17480 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__635__A
timestamp 1586364061
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_165
timestamp 1586364061
transform 1 0 16284 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_170
timestamp 1586364061
transform 1 0 16744 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_181
timestamp 1586364061
transform 1 0 17756 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_186
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 774 592
use scs8hd_nor2_4  _486_
timestamp 1586364061
transform 1 0 19228 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_513
timestamp 1586364061
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_194
timestamp 1586364061
transform 1 0 18952 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_206
timestamp 1586364061
transform 1 0 20056 0 -1 25568
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_226
timestamp 1586364061
transform 1 0 21896 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 25568
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24564 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_247
timestamp 1586364061
transform 1 0 23828 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_42_252
timestamp 1586364061
transform 1 0 24288 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_264
timestamp 1586364061
transform 1 0 25392 0 -1 25568
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 27232 0 -1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_514
timestamp 1586364061
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27048 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_272
timestamp 1586364061
transform 1 0 26128 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_276
timestamp 1586364061
transform 1 0 26496 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_42_295
timestamp 1586364061
transform 1 0 28244 0 -1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30728 0 -1 25568
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28980 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28428 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_299
timestamp 1586364061
transform 1 0 28612 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_8  FILLER_42_312
timestamp 1586364061
transform 1 0 29808 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_320
timestamp 1586364061
transform 1 0 30544 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_325
timestamp 1586364061
transform 1 0 31004 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_329
timestamp 1586364061
transform 1 0 31372 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31556 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31188 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_333
timestamp 1586364061
transform 1 0 31740 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_515
timestamp 1586364061
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_340
timestamp 1586364061
transform 1 0 32384 0 -1 25568
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_346
timestamp 1586364061
transform 1 0 32936 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32752 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 -1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 -1 25568
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33304 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34684 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_359
timestamp 1586364061
transform 1 0 34132 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_42_382
timestamp 1586364061
transform 1 0 36248 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_376
timestamp 1586364061
transform 1 0 35696 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 36064 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_387
timestamp 1586364061
transform 1 0 36708 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36892 0 -1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_391
timestamp 1586364061
transform 1 0 37076 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_42_402
timestamp 1586364061
transform 1 0 38088 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_398
timestamp 1586364061
transform 1 0 37720 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37904 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_516
timestamp 1586364061
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use scs8hd_buf_1  _387_
timestamp 1586364061
transform 1 0 38548 0 -1 25568
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39560 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38272 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_406
timestamp 1586364061
transform 1 0 38456 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_410
timestamp 1586364061
transform 1 0 38824 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_6  FILLER_42_427
timestamp 1586364061
transform 1 0 40388 0 -1 25568
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42136 0 -1 25568
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41124 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41584 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41952 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40940 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_438
timestamp 1586364061
transform 1 0 41400 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_442
timestamp 1586364061
transform 1 0 41768 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_449
timestamp 1586364061
transform 1 0 42412 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_1  _428_
timestamp 1586364061
transform 1 0 44344 0 -1 25568
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_517
timestamp 1586364061
transform 1 0 43240 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_457
timestamp 1586364061
transform 1 0 43148 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_462
timestamp 1586364061
transform 1 0 43608 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_12  FILLER_42_473
timestamp 1586364061
transform 1 0 44620 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_485
timestamp 1586364061
transform 1 0 45724 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_497
timestamp 1586364061
transform 1 0 46828 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_509
timestamp 1586364061
transform 1 0 47932 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 48852 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_515
timestamp 1586364061
transform 1 0 48484 0 -1 25568
box -38 -48 130 592
use scs8hd_buf_1  _250_
timestamp 1586364061
transform 1 0 3128 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_43_21
timestamp 1586364061
transform 1 0 3036 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_25
timestamp 1586364061
transform 1 0 3404 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_29
timestamp 1586364061
transform 1 0 3772 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__250__A
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__266__B
timestamp 1586364061
transform 1 0 3956 0 1 25568
box -38 -48 222 592
use scs8hd_buf_1  _261_
timestamp 1586364061
transform 1 0 4140 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_36
timestamp 1586364061
transform 1 0 4416 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__266__A
timestamp 1586364061
transform 1 0 4600 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_40
timestamp 1586364061
transform 1 0 4784 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__261__A
timestamp 1586364061
transform 1 0 4968 0 1 25568
box -38 -48 222 592
use scs8hd_buf_1  _243_
timestamp 1586364061
transform 1 0 5152 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_47
timestamp 1586364061
transform 1 0 5428 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 5612 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 5980 0 1 25568
box -38 -48 222 592
use scs8hd_buf_1  _294_
timestamp 1586364061
transform 1 0 8372 0 1 25568
box -38 -48 314 592
use scs8hd_nor2_4  _295_
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_518
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__294__A
timestamp 1586364061
transform 1 0 8188 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__295__B
timestamp 1586364061
transform 1 0 7820 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_55
timestamp 1586364061
transform 1 0 6164 0 1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_43_71
timestamp 1586364061
transform 1 0 7636 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_75
timestamp 1586364061
transform 1 0 8004 0 1 25568
box -38 -48 222 592
use scs8hd_nor2_4  _304_
timestamp 1586364061
transform 1 0 9476 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__304__A
timestamp 1586364061
transform 1 0 9292 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__276__A
timestamp 1586364061
transform 1 0 8832 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__304__B
timestamp 1586364061
transform 1 0 10856 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_82
timestamp 1586364061
transform 1 0 8648 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_86
timestamp 1586364061
transform 1 0 9016 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_100
timestamp 1586364061
transform 1 0 10304 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_104
timestamp 1586364061
transform 1 0 10672 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_108
timestamp 1586364061
transform 1 0 11040 0 1 25568
box -38 -48 314 592
use scs8hd_buf_1  _267_
timestamp 1586364061
transform 1 0 11316 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_114
timestamp 1586364061
transform 1 0 11592 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_118
timestamp 1586364061
transform 1 0 11960 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__267__A
timestamp 1586364061
transform 1 0 11776 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__291__A
timestamp 1586364061
transform 1 0 12144 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_519
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 222 592
use scs8hd_buf_1  _284_
timestamp 1586364061
transform 1 0 12604 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_128
timestamp 1586364061
transform 1 0 12880 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__284__A
timestamp 1586364061
transform 1 0 13064 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_132
timestamp 1586364061
transform 1 0 13248 0 1 25568
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 14260 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__289__A
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_137
timestamp 1586364061
transform 1 0 13708 0 1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_43_154
timestamp 1586364061
transform 1 0 15272 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_158
timestamp 1586364061
transform 1 0 15640 0 1 25568
box -38 -48 222 592
use scs8hd_buf_1  _580_
timestamp 1586364061
transform 1 0 16928 0 1 25568
box -38 -48 314 592
use scs8hd_inv_8  _635_
timestamp 1586364061
transform 1 0 18032 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_520
timestamp 1586364061
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__580__A
timestamp 1586364061
transform 1 0 17756 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_162
timestamp 1586364061
transform 1 0 16008 0 1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_43_175
timestamp 1586364061
transform 1 0 17204 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_179
timestamp 1586364061
transform 1 0 17572 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 19872 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 19688 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__634__A
timestamp 1586364061
transform 1 0 19044 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_193
timestamp 1586364061
transform 1 0 18860 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_197
timestamp 1586364061
transform 1 0 19228 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_201
timestamp 1586364061
transform 1 0 19596 0 1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_43_222
timestamp 1586364061
transform 1 0 21528 0 1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_43_219
timestamp 1586364061
transform 1 0 21252 0 1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_43_215
timestamp 1586364061
transform 1 0 20884 0 1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 1 25568
box -38 -48 866 592
use scs8hd_fill_2  FILLER_43_232
timestamp 1586364061
transform 1 0 22448 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_240
timestamp 1586364061
transform 1 0 23184 0 1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_43_236
timestamp 1586364061
transform 1 0 22816 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_521
timestamp 1586364061
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_245
timestamp 1586364061
transform 1 0 23644 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_259
timestamp 1586364061
transform 1 0 24932 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_263
timestamp 1586364061
transform 1 0 25300 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_267
timestamp 1586364061
transform 1 0 25668 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_271
timestamp 1586364061
transform 1 0 26036 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__501__B
timestamp 1586364061
transform 1 0 25852 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__501__A
timestamp 1586364061
transform 1 0 26220 0 1 25568
box -38 -48 222 592
use scs8hd_nor2_4  _501_
timestamp 1586364061
transform 1 0 26404 0 1 25568
box -38 -48 866 592
use scs8hd_fill_2  FILLER_43_288
timestamp 1586364061
transform 1 0 27600 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_284
timestamp 1586364061
transform 1 0 27232 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 27416 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_295
timestamp 1586364061
transform 1 0 28244 0 1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27784 0 1 25568
box -38 -48 222 592
use scs8hd_conb_1  _642_
timestamp 1586364061
transform 1 0 27968 0 1 25568
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30176 0 1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_522
timestamp 1586364061
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30636 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28980 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_301
timestamp 1586364061
transform 1 0 28796 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_306
timestamp 1586364061
transform 1 0 29256 0 1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_43_314
timestamp 1586364061
transform 1 0 29992 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_319
timestamp 1586364061
transform 1 0 30452 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32752 0 1 25568
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31188 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32200 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31004 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32568 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_323
timestamp 1586364061
transform 1 0 30820 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_336
timestamp 1586364061
transform 1 0 32016 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_340
timestamp 1586364061
transform 1 0 32384 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_353
timestamp 1586364061
transform 1 0 33580 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_357
timestamp 1586364061
transform 1 0 33948 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33764 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_361
timestamp 1586364061
transform 1 0 34316 0 1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34132 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_365
timestamp 1586364061
transform 1 0 34684 0 1 25568
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_523
timestamp 1586364061
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_370
timestamp 1586364061
transform 1 0 35144 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_374
timestamp 1586364061
transform 1 0 35512 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 36064 0 1 25568
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37904 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35696 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 37260 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37720 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_378
timestamp 1586364061
transform 1 0 35880 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_391
timestamp 1586364061
transform 1 0 37076 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_395
timestamp 1586364061
transform 1 0 37444 0 1 25568
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_524
timestamp 1586364061
transform 1 0 40388 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39468 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38916 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39836 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_409
timestamp 1586364061
transform 1 0 38732 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_413
timestamp 1586364061
transform 1 0 39100 0 1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_43_419
timestamp 1586364061
transform 1 0 39652 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_423
timestamp 1586364061
transform 1 0 40020 0 1 25568
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41584 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41400 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42596 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_431
timestamp 1586364061
transform 1 0 40756 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_435
timestamp 1586364061
transform 1 0 41124 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_449
timestamp 1586364061
transform 1 0 42412 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_453
timestamp 1586364061
transform 1 0 42780 0 1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44160 0 1 25568
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43148 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44620 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43608 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43976 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_460
timestamp 1586364061
transform 1 0 43424 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_464
timestamp 1586364061
transform 1 0 43792 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_471
timestamp 1586364061
transform 1 0 44436 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_475
timestamp 1586364061
transform 1 0 44804 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_525
timestamp 1586364061
transform 1 0 46000 0 1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_43_487
timestamp 1586364061
transform 1 0 45908 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_489
timestamp 1586364061
transform 1 0 46092 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_501
timestamp 1586364061
transform 1 0 47196 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 48852 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_513
timestamp 1586364061
transform 1 0 48300 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_buf_1  _234_
timestamp 1586364061
transform 1 0 5612 0 -1 26656
box -38 -48 314 592
use scs8hd_nor2_4  _266_
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_526
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_41
timestamp 1586364061
transform 1 0 4876 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_8  FILLER_44_52
timestamp 1586364061
transform 1 0 5888 0 -1 26656
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 26656
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_44_71
timestamp 1586364061
transform 1 0 7636 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_44_79
timestamp 1586364061
transform 1 0 8372 0 -1 26656
box -38 -48 222 592
use scs8hd_buf_1  _276_
timestamp 1586364061
transform 1 0 8556 0 -1 26656
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10212 0 -1 26656
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_527
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__301__A
timestamp 1586364061
transform 1 0 9844 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_84
timestamp 1586364061
transform 1 0 8832 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_97
timestamp 1586364061
transform 1 0 10028 0 -1 26656
box -38 -48 222 592
use scs8hd_buf_1  _291_
timestamp 1586364061
transform 1 0 12512 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__281__B
timestamp 1586364061
transform 1 0 12144 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__289__B
timestamp 1586364061
transform 1 0 13340 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_110
timestamp 1586364061
transform 1 0 11224 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_44_118
timestamp 1586364061
transform 1 0 11960 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_122
timestamp 1586364061
transform 1 0 12328 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_127
timestamp 1586364061
transform 1 0 12788 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_131
timestamp 1586364061
transform 1 0 13156 0 -1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _289_
timestamp 1586364061
transform 1 0 13524 0 -1 26656
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_528
timestamp 1586364061
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_144
timestamp 1586364061
transform 1 0 14352 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_148
timestamp 1586364061
transform 1 0 14720 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_44_152
timestamp 1586364061
transform 1 0 15088 0 -1 26656
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17388 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_163
timestamp 1586364061
transform 1 0 16100 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_4  FILLER_44_173
timestamp 1586364061
transform 1 0 17020 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_44_186
timestamp 1586364061
transform 1 0 18216 0 -1 26656
box -38 -48 222 592
use scs8hd_inv_8  _634_
timestamp 1586364061
transform 1 0 18952 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_529
timestamp 1586364061
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_190
timestamp 1586364061
transform 1 0 18584 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_44_203
timestamp 1586364061
transform 1 0 19780 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_207
timestamp 1586364061
transform 1 0 20148 0 -1 26656
box -38 -48 590 592
use scs8hd_fill_1  FILLER_44_213
timestamp 1586364061
transform 1 0 20700 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_223
timestamp 1586364061
transform 1 0 21620 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_219
timestamp 1586364061
transform 1 0 21252 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_215
timestamp 1586364061
transform 1 0 20884 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_227
timestamp 1586364061
transform 1 0 21988 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22172 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 -1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22356 0 -1 26656
box -38 -48 866 592
use scs8hd_decap_8  FILLER_44_240
timestamp 1586364061
transform 1 0 23184 0 -1 26656
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_250
timestamp 1586364061
transform 1 0 24104 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_263
timestamp 1586364061
transform 1 0 25300 0 -1 26656
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 26864 0 -1 26656
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_530
timestamp 1586364061
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__497__B
timestamp 1586364061
transform 1 0 28060 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_276
timestamp 1586364061
transform 1 0 26496 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_44_291
timestamp 1586364061
transform 1 0 27876 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_295
timestamp 1586364061
transform 1 0 28244 0 -1 26656
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28612 0 -1 26656
box -38 -48 866 592
use scs8hd_decap_12  FILLER_44_308
timestamp 1586364061
transform 1 0 29440 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_44_320
timestamp 1586364061
transform 1 0 30544 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_326
timestamp 1586364061
transform 1 0 31096 0 -1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30820 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_4  FILLER_44_330
timestamp 1586364061
transform 1 0 31464 0 -1 26656
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31280 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_531
timestamp 1586364061
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_341
timestamp 1586364061
transform 1 0 32476 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_337
timestamp 1586364061
transform 1 0 32108 0 -1 26656
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32200 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_4  FILLER_44_345
timestamp 1586364061
transform 1 0 32844 0 -1 26656
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32660 0 -1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34776 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__437__A
timestamp 1586364061
transform 1 0 35236 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__437__B
timestamp 1586364061
transform 1 0 35604 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_358
timestamp 1586364061
transform 1 0 34040 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_44_369
timestamp 1586364061
transform 1 0 35052 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_373
timestamp 1586364061
transform 1 0 35420 0 -1 26656
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 35880 0 -1 26656
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37904 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_532
timestamp 1586364061
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_1  FILLER_44_377
timestamp 1586364061
transform 1 0 35788 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_8  FILLER_44_389
timestamp 1586364061
transform 1 0 36892 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_44_398
timestamp 1586364061
transform 1 0 37720 0 -1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39468 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38916 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39284 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_409
timestamp 1586364061
transform 1 0 38732 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_413
timestamp 1586364061
transform 1 0 39100 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_426
timestamp 1586364061
transform 1 0 40296 0 -1 26656
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_438
timestamp 1586364061
transform 1 0 41400 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_8  FILLER_44_450
timestamp 1586364061
transform 1 0 42504 0 -1 26656
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_533
timestamp 1586364061
transform 1 0 43240 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_468
timestamp 1586364061
transform 1 0 44160 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_480
timestamp 1586364061
transform 1 0 45264 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_492
timestamp 1586364061
transform 1 0 46368 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_504
timestamp 1586364061
transform 1 0 47472 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 48852 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 774 592
use scs8hd_fill_1  FILLER_45_23
timestamp 1586364061
transform 1 0 3220 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_26
timestamp 1586364061
transform 1 0 3496 0 1 26656
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 4232 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__298__A
timestamp 1586364061
transform 1 0 5888 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__298__B
timestamp 1586364061
transform 1 0 5520 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_30
timestamp 1586364061
transform 1 0 3864 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_45
timestamp 1586364061
transform 1 0 5244 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_50
timestamp 1586364061
transform 1 0 5704 0 1 26656
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_534
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_54
timestamp 1586364061
transform 1 0 6072 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_58
timestamp 1586364061
transform 1 0 6440 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_73
timestamp 1586364061
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_77
timestamp 1586364061
transform 1 0 8188 0 1 26656
box -38 -48 222 592
use scs8hd_buf_1  _278_
timestamp 1586364061
transform 1 0 8556 0 1 26656
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9844 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__278__A
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_84
timestamp 1586364061
transform 1 0 8832 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_88
timestamp 1586364061
transform 1 0 9200 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_92
timestamp 1586364061
transform 1 0 9568 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_106
timestamp 1586364061
transform 1 0 10856 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_114
timestamp 1586364061
transform 1 0 11592 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_110
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__301__B
timestamp 1586364061
transform 1 0 11040 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__281__A
timestamp 1586364061
transform 1 0 11776 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_118
timestamp 1586364061
transform 1 0 11960 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_535
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 866 592
use scs8hd_decap_4  FILLER_45_132
timestamp 1586364061
transform 1 0 13248 0 1 26656
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15916 0 1 26656
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14168 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__280__A
timestamp 1586364061
transform 1 0 13616 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_138
timestamp 1586364061
transform 1 0 13800 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_153
timestamp 1586364061
transform 1 0 15180 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_157
timestamp 1586364061
transform 1 0 15548 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_168
timestamp 1586364061
transform 1 0 16560 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_164
timestamp 1586364061
transform 1 0 16192 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_179
timestamp 1586364061
transform 1 0 17572 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_175
timestamp 1586364061
transform 1 0 17204 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_536
timestamp 1586364061
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 26656
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20516 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_193
timestamp 1586364061
transform 1 0 18860 0 1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_45_197
timestamp 1586364061
transform 1 0 19228 0 1 26656
box -38 -48 590 592
use scs8hd_decap_4  FILLER_45_205
timestamp 1586364061
transform 1 0 19964 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_214
timestamp 1586364061
transform 1 0 20792 0 1 26656
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 21528 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 21344 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_218
timestamp 1586364061
transform 1 0 21160 0 1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_45_233
timestamp 1586364061
transform 1 0 22540 0 1 26656
box -38 -48 774 592
use scs8hd_fill_1  FILLER_45_241
timestamp 1586364061
transform 1 0 23276 0 1 26656
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 23644 0 1 26656
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_537
timestamp 1586364061
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__496__B
timestamp 1586364061
transform 1 0 25760 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_256
timestamp 1586364061
transform 1 0 24656 0 1 26656
box -38 -48 1142 592
use scs8hd_nor2_4  _496_
timestamp 1586364061
transform 1 0 26312 0 1 26656
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27876 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27324 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__496__A
timestamp 1586364061
transform 1 0 26128 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__497__A
timestamp 1586364061
transform 1 0 27692 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_270
timestamp 1586364061
transform 1 0 25944 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_283
timestamp 1586364061
transform 1 0 27140 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_287
timestamp 1586364061
transform 1 0 27508 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_294
timestamp 1586364061
transform 1 0 28152 0 1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_45_302
timestamp 1586364061
transform 1 0 28888 0 1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_45_298
timestamp 1586364061
transform 1 0 28520 0 1 26656
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28980 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28336 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_538
timestamp 1586364061
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_313
timestamp 1586364061
transform 1 0 29900 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_309
timestamp 1586364061
transform 1 0 29532 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 29716 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_317
timestamp 1586364061
transform 1 0 30268 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30544 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30084 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30728 0 1 26656
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32292 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32108 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31740 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_331
timestamp 1586364061
transform 1 0 31556 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_335
timestamp 1586364061
transform 1 0 31924 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_348
timestamp 1586364061
transform 1 0 33120 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_356
timestamp 1586364061
transform 1 0 33856 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_352
timestamp 1586364061
transform 1 0 33488 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33672 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_367
timestamp 1586364061
transform 1 0 34868 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_362
timestamp 1586364061
transform 1 0 34408 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__436__B
timestamp 1586364061
transform 1 0 34224 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__436__A
timestamp 1586364061
transform 1 0 34592 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_539
timestamp 1586364061
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use scs8hd_nor2_4  _436_
timestamp 1586364061
transform 1 0 35144 0 1 26656
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 36708 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 36524 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38088 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36156 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_379
timestamp 1586364061
transform 1 0 35972 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_383
timestamp 1586364061
transform 1 0 36340 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_398
timestamp 1586364061
transform 1 0 37720 0 1 26656
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38456 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_540
timestamp 1586364061
transform 1 0 40388 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39652 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40020 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_404
timestamp 1586364061
transform 1 0 38272 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_415
timestamp 1586364061
transform 1 0 39284 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_421
timestamp 1586364061
transform 1 0 39836 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_425
timestamp 1586364061
transform 1 0 40204 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_428
timestamp 1586364061
transform 1 0 40480 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_437
timestamp 1586364061
transform 1 0 41308 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_433
timestamp 1586364061
transform 1 0 40940 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41492 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41124 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40664 0 1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_45_454
timestamp 1586364061
transform 1 0 42872 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_450
timestamp 1586364061
transform 1 0 42504 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42688 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43240 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43700 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44068 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_461
timestamp 1586364061
transform 1 0 43516 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_465
timestamp 1586364061
transform 1 0 43884 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_469
timestamp 1586364061
transform 1 0 44252 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_45_481
timestamp 1586364061
transform 1 0 45356 0 1 26656
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_541
timestamp 1586364061
transform 1 0 46000 0 1 26656
box -38 -48 130 592
use scs8hd_fill_1  FILLER_45_487
timestamp 1586364061
transform 1 0 45908 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_489
timestamp 1586364061
transform 1 0 46092 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_501
timestamp 1586364061
transform 1 0 47196 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 48852 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_513
timestamp 1586364061
transform 1 0 48300 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_47_23
timestamp 1586364061
transform 1 0 3220 0 1 27744
box -38 -48 130 592
use scs8hd_decap_8  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  FILLER_46_23
timestamp 1586364061
transform 1 0 3220 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__262__A
timestamp 1586364061
transform 1 0 3312 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__262__B
timestamp 1586364061
transform 1 0 3496 0 -1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _262_
timestamp 1586364061
transform 1 0 3496 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_35
timestamp 1586364061
transform 1 0 4324 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_28
timestamp 1586364061
transform 1 0 3680 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_542
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_47_49
timestamp 1586364061
transform 1 0 5612 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_43
timestamp 1586364061
transform 1 0 5060 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 406 592
use scs8hd_decap_8  FILLER_46_43
timestamp 1586364061
transform 1 0 5060 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 1 27744
box -38 -48 314 592
use scs8hd_decap_4  FILLER_47_53
timestamp 1586364061
transform 1 0 5980 0 1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_46_51
timestamp 1586364061
transform 1 0 5796 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _298_
timestamp 1586364061
transform 1 0 5888 0 -1 27744
box -38 -48 866 592
use scs8hd_decap_3  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_59
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_61
timestamp 1586364061
transform 1 0 6716 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6900 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_550
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_72
timestamp 1586364061
transform 1 0 7728 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_68
timestamp 1586364061
transform 1 0 7360 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_73
timestamp 1586364061
transform 1 0 7820 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_69
timestamp 1586364061
transform 1 0 7452 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_65
timestamp 1586364061
transform 1 0 7084 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_90
timestamp 1586364061
transform 1 0 9384 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_85
timestamp 1586364061
transform 1 0 8924 0 1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_46_84
timestamp 1586364061
transform 1 0 8832 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 9568 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_543
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_nor2_4  _301_
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_101
timestamp 1586364061
transform 1 0 10396 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_97
timestamp 1586364061
transform 1 0 10028 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_102
timestamp 1586364061
transform 1 0 10488 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 27744
box -38 -48 866 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 9752 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_107
timestamp 1586364061
transform 1 0 10948 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_118
timestamp 1586364061
transform 1 0 11960 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_114
timestamp 1586364061
transform 1 0 11592 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_119
timestamp 1586364061
transform 1 0 12052 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_129
timestamp 1586364061
transform 1 0 12972 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_551
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 12788 0 1 27744
box -38 -48 1050 592
use scs8hd_nor2_4  _281_
timestamp 1586364061
transform 1 0 12144 0 -1 27744
box -38 -48 866 592
use scs8hd_decap_4  FILLER_46_133
timestamp 1586364061
transform 1 0 13340 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_142
timestamp 1586364061
transform 1 0 14168 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_138
timestamp 1586364061
transform 1 0 13800 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_144
timestamp 1586364061
transform 1 0 14352 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_140
timestamp 1586364061
transform 1 0 13984 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 27744
box -38 -48 222 592
use scs8hd_buf_1  _280_
timestamp 1586364061
transform 1 0 13708 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_151
timestamp 1586364061
transform 1 0 14996 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_146
timestamp 1586364061
transform 1 0 14536 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_46_152
timestamp 1586364061
transform 1 0 15088 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_544
timestamp 1586364061
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_1  FILLER_47_168
timestamp 1586364061
transform 1 0 16560 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_164
timestamp 1586364061
transform 1 0 16192 0 1 27744
box -38 -48 406 592
use scs8hd_decap_6  FILLER_46_163
timestamp 1586364061
transform 1 0 16100 0 -1 27744
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_179
timestamp 1586364061
transform 1 0 17572 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_175
timestamp 1586364061
transform 1 0 17204 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_171
timestamp 1586364061
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_180
timestamp 1586364061
transform 1 0 17664 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 17388 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 27744
box -38 -48 866 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 16928 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_47_184
timestamp 1586364061
transform 1 0 18032 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_46_187
timestamp 1586364061
transform 1 0 18308 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_184
timestamp 1586364061
transform 1 0 18032 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__633__A
timestamp 1586364061
transform 1 0 18124 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_552
timestamp 1586364061
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use scs8hd_inv_8  _633_
timestamp 1586364061
transform 1 0 18124 0 1 27744
box -38 -48 866 592
use scs8hd_decap_3  FILLER_47_194
timestamp 1586364061
transform 1 0 18952 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_46_196
timestamp 1586364061
transform 1 0 19136 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_192
timestamp 1586364061
transform 1 0 18768 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__525__B
timestamp 1586364061
transform 1 0 19228 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__525__A
timestamp 1586364061
transform 1 0 19228 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18492 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_47_203
timestamp 1586364061
transform 1 0 19780 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_199
timestamp 1586364061
transform 1 0 19412 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_46_206
timestamp 1586364061
transform 1 0 20056 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_199
timestamp 1586364061
transform 1 0 19412 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__488__A
timestamp 1586364061
transform 1 0 19872 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 27744
box -38 -48 314 592
use scs8hd_nor2_4  _488_
timestamp 1586364061
transform 1 0 20056 0 1 27744
box -38 -48 866 592
use scs8hd_decap_4  FILLER_46_210
timestamp 1586364061
transform 1 0 20424 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__488__B
timestamp 1586364061
transform 1 0 20240 0 -1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_545
timestamp 1586364061
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_1  FILLER_47_223
timestamp 1586364061
transform 1 0 21620 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_219
timestamp 1586364061
transform 1 0 21252 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_215
timestamp 1586364061
transform 1 0 20884 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_226
timestamp 1586364061
transform 1 0 21896 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__485__B
timestamp 1586364061
transform 1 0 21436 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__485__A
timestamp 1586364061
transform 1 0 21068 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 1 27744
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 27744
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_47_237
timestamp 1586364061
transform 1 0 22908 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_233
timestamp 1586364061
transform 1 0 22540 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_234
timestamp 1586364061
transform 1 0 22632 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_46_230
timestamp 1586364061
transform 1 0 22264 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__490__A
timestamp 1586364061
transform 1 0 22724 0 1 27744
box -38 -48 222 592
use scs8hd_conb_1  _643_
timestamp 1586364061
transform 1 0 22908 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  FILLER_47_241
timestamp 1586364061
transform 1 0 23276 0 1 27744
box -38 -48 314 592
use scs8hd_decap_4  FILLER_46_240
timestamp 1586364061
transform 1 0 23184 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__490__B
timestamp 1586364061
transform 1 0 23092 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_249
timestamp 1586364061
transform 1 0 24012 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_245
timestamp 1586364061
transform 1 0 23644 0 1 27744
box -38 -48 130 592
use scs8hd_fill_1  FILLER_46_247
timestamp 1586364061
transform 1 0 23828 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_1  FILLER_46_244
timestamp 1586364061
transform 1 0 23552 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23644 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24196 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_553
timestamp 1586364061
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 -1 27744
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23736 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_253
timestamp 1586364061
transform 1 0 24380 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_261
timestamp 1586364061
transform 1 0 25116 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_257
timestamp 1586364061
transform 1 0 24748 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__514__A
timestamp 1586364061
transform 1 0 24932 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__513__A
timestamp 1586364061
transform 1 0 24564 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _514_
timestamp 1586364061
transform 1 0 24748 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_266
timestamp 1586364061
transform 1 0 25576 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_265
timestamp 1586364061
transform 1 0 25484 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__513__B
timestamp 1586364061
transform 1 0 25300 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__514__B
timestamp 1586364061
transform 1 0 25760 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_274
timestamp 1586364061
transform 1 0 26312 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_270
timestamp 1586364061
transform 1 0 25944 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_46_273
timestamp 1586364061
transform 1 0 26220 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26404 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_546
timestamp 1586364061
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 27744
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26588 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_284
timestamp 1586364061
transform 1 0 27232 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_280
timestamp 1586364061
transform 1 0 26864 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_287
timestamp 1586364061
transform 1 0 27508 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_8  FILLER_46_279
timestamp 1586364061
transform 1 0 26772 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__500__A
timestamp 1586364061
transform 1 0 27600 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__498__A
timestamp 1586364061
transform 1 0 27416 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27048 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _500_
timestamp 1586364061
transform 1 0 27600 0 1 27744
box -38 -48 866 592
use scs8hd_nor2_4  _497_
timestamp 1586364061
transform 1 0 27784 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_306
timestamp 1586364061
transform 1 0 29256 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_301
timestamp 1586364061
transform 1 0 28796 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_297
timestamp 1586364061
transform 1 0 28428 0 1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_46_299
timestamp 1586364061
transform 1 0 28612 0 -1 27744
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29164 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__500__B
timestamp 1586364061
transform 1 0 28612 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_554
timestamp 1586364061
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 29348 0 -1 27744
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_46_318
timestamp 1586364061
transform 1 0 30360 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 29440 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 29624 0 1 27744
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_47_321
timestamp 1586364061
transform 1 0 30636 0 1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30728 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_47_327
timestamp 1586364061
transform 1 0 31188 0 1 27744
box -38 -48 590 592
use scs8hd_decap_12  FILLER_46_324
timestamp 1586364061
transform 1 0 30912 0 -1 27744
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__516__A
timestamp 1586364061
transform 1 0 31004 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_335
timestamp 1586364061
transform 1 0 31924 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_346
timestamp 1586364061
transform 1 0 32936 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_547
timestamp 1586364061
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 27744
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 32292 0 1 27744
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_47_358
timestamp 1586364061
transform 1 0 34040 0 1 27744
box -38 -48 590 592
use scs8hd_fill_2  FILLER_47_354
timestamp 1586364061
transform 1 0 33672 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_350
timestamp 1586364061
transform 1 0 33304 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33488 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33672 0 -1 27744
box -38 -48 866 592
use scs8hd_decap_8  FILLER_46_363
timestamp 1586364061
transform 1 0 34500 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__423__A
timestamp 1586364061
transform 1 0 34592 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_555
timestamp 1586364061
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_374
timestamp 1586364061
transform 1 0 35512 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_370
timestamp 1586364061
transform 1 0 35144 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _437_
timestamp 1586364061
transform 1 0 35236 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_378
timestamp 1586364061
transform 1 0 35880 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_384
timestamp 1586364061
transform 1 0 36432 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_380
timestamp 1586364061
transform 1 0 36064 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36616 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__430__B
timestamp 1586364061
transform 1 0 36248 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__430__A
timestamp 1586364061
transform 1 0 35696 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 36064 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 36248 0 1 27744
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_47_393
timestamp 1586364061
transform 1 0 37260 0 1 27744
box -38 -48 774 592
use scs8hd_decap_4  FILLER_46_398
timestamp 1586364061
transform 1 0 37720 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_46_396
timestamp 1586364061
transform 1 0 37536 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_8  FILLER_46_388
timestamp 1586364061
transform 1 0 36800 0 -1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_548
timestamp 1586364061
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38088 0 -1 27744
box -38 -48 866 592
use scs8hd_conb_1  _648_
timestamp 1586364061
transform 1 0 37996 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_412
timestamp 1586364061
transform 1 0 39008 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_408
timestamp 1586364061
transform 1 0 38640 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_404
timestamp 1586364061
transform 1 0 38272 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_411
timestamp 1586364061
transform 1 0 38916 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38824 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 38456 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_421
timestamp 1586364061
transform 1 0 39836 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_417
timestamp 1586364061
transform 1 0 39468 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_415
timestamp 1586364061
transform 1 0 39284 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39100 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39652 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39652 0 -1 27744
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39192 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_47_426
timestamp 1586364061
transform 1 0 40296 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_46_428
timestamp 1586364061
transform 1 0 40480 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40112 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_556
timestamp 1586364061
transform 1 0 40388 0 1 27744
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_47_439
timestamp 1586364061
transform 1 0 41492 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_435
timestamp 1586364061
transform 1 0 41124 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_431
timestamp 1586364061
transform 1 0 40756 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_438
timestamp 1586364061
transform 1 0 41400 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_6  FILLER_46_432
timestamp 1586364061
transform 1 0 40848 0 -1 27744
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40664 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41584 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41768 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_455
timestamp 1586364061
transform 1 0 42964 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_451
timestamp 1586364061
transform 1 0 42596 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_450
timestamp 1586364061
transform 1 0 42504 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42780 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_466
timestamp 1586364061
transform 1 0 43976 0 1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_462
timestamp 1586364061
transform 1 0 43608 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_462
timestamp 1586364061
transform 1 0 43608 0 -1 27744
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43148 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43792 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_549
timestamp 1586364061
transform 1 0 43240 0 -1 27744
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 1 27744
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_47_478
timestamp 1586364061
transform 1 0 45080 0 1 27744
box -38 -48 774 592
use scs8hd_decap_12  FILLER_46_474
timestamp 1586364061
transform 1 0 44712 0 -1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_557
timestamp 1586364061
transform 1 0 46000 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_486
timestamp 1586364061
transform 1 0 45816 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_498
timestamp 1586364061
transform 1 0 46920 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_486
timestamp 1586364061
transform 1 0 45816 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_489
timestamp 1586364061
transform 1 0 46092 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_501
timestamp 1586364061
transform 1 0 47196 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 48852 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 48852 0 1 27744
box -38 -48 314 592
use scs8hd_decap_6  FILLER_46_510
timestamp 1586364061
transform 1 0 48024 0 -1 27744
box -38 -48 590 592
use scs8hd_decap_3  FILLER_47_513
timestamp 1586364061
transform 1 0 48300 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__244__B
timestamp 1586364061
transform 1 0 2668 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_48_19
timestamp 1586364061
transform 1 0 2852 0 -1 28832
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 28832
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_558
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4784 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_38
timestamp 1586364061
transform 1 0 4600 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_42
timestamp 1586364061
transform 1 0 4968 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_8  FILLER_48_49
timestamp 1586364061
transform 1 0 5612 0 -1 28832
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7912 0 -1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_66
timestamp 1586364061
transform 1 0 7176 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_48_77
timestamp 1586364061
transform 1 0 8188 0 -1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_559
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_81
timestamp 1586364061
transform 1 0 8556 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_85
timestamp 1586364061
transform 1 0 8924 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_88
timestamp 1586364061
transform 1 0 9200 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_8  FILLER_48_102
timestamp 1586364061
transform 1 0 10488 0 -1 28832
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_110
timestamp 1586364061
transform 1 0 11224 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_121
timestamp 1586364061
transform 1 0 12236 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_125
timestamp 1586364061
transform 1 0 12604 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_129
timestamp 1586364061
transform 1 0 12972 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_133
timestamp 1586364061
transform 1 0 13340 0 -1 28832
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_560
timestamp 1586364061
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_145
timestamp 1586364061
transform 1 0 14444 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_48_157
timestamp 1586364061
transform 1 0 15548 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_161
timestamp 1586364061
transform 1 0 15916 0 -1 28832
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16652 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_48_165
timestamp 1586364061
transform 1 0 16284 0 -1 28832
box -38 -48 130 592
use scs8hd_fill_1  FILLER_48_168
timestamp 1586364061
transform 1 0 16560 0 -1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_48_178
timestamp 1586364061
transform 1 0 17480 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_182
timestamp 1586364061
transform 1 0 17848 0 -1 28832
box -38 -48 406 592
use scs8hd_nor2_4  _525_
timestamp 1586364061
transform 1 0 19228 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_561
timestamp 1586364061
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_189
timestamp 1586364061
transform 1 0 18492 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_8  FILLER_48_206
timestamp 1586364061
transform 1 0 20056 0 -1 28832
box -38 -48 774 592
use scs8hd_nor2_4  _485_
timestamp 1586364061
transform 1 0 20884 0 -1 28832
box -38 -48 866 592
use scs8hd_nor2_4  _490_
timestamp 1586364061
transform 1 0 22448 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__507__B
timestamp 1586364061
transform 1 0 21988 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_224
timestamp 1586364061
transform 1 0 21712 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_48_229
timestamp 1586364061
transform 1 0 22172 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_241
timestamp 1586364061
transform 1 0 23276 0 -1 28832
box -38 -48 1142 592
use scs8hd_nor2_4  _513_
timestamp 1586364061
transform 1 0 24840 0 -1 28832
box -38 -48 866 592
use scs8hd_decap_4  FILLER_48_253
timestamp 1586364061
transform 1 0 24380 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_257
timestamp 1586364061
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_6  FILLER_48_267
timestamp 1586364061
transform 1 0 25668 0 -1 28832
box -38 -48 590 592
use scs8hd_nor2_4  _498_
timestamp 1586364061
transform 1 0 27692 0 -1 28832
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_562
timestamp 1586364061
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__498__B
timestamp 1586364061
transform 1 0 27508 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27140 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_279
timestamp 1586364061
transform 1 0 26772 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_48_285
timestamp 1586364061
transform 1 0 27324 0 -1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 29256 0 -1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30452 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_298
timestamp 1586364061
transform 1 0 28520 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_48_317
timestamp 1586364061
transform 1 0 30268 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_321
timestamp 1586364061
transform 1 0 30636 0 -1 28832
box -38 -48 406 592
use scs8hd_buf_1  _516_
timestamp 1586364061
transform 1 0 31004 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_328
timestamp 1586364061
transform 1 0 31280 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31464 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_332
timestamp 1586364061
transform 1 0 31648 0 -1 28832
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_563
timestamp 1586364061
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_48_341
timestamp 1586364061
transform 1 0 32476 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_48_337
timestamp 1586364061
transform 1 0 32108 0 -1 28832
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32200 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_4  FILLER_48_345
timestamp 1586364061
transform 1 0 32844 0 -1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32660 0 -1 28832
box -38 -48 222 592
use scs8hd_buf_1  _423_
timestamp 1586364061
transform 1 0 34776 0 -1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__435__A
timestamp 1586364061
transform 1 0 35236 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_358
timestamp 1586364061
transform 1 0 34040 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_48_369
timestamp 1586364061
transform 1 0 35052 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_373
timestamp 1586364061
transform 1 0 35420 0 -1 28832
box -38 -48 406 592
use scs8hd_nor2_4  _430_
timestamp 1586364061
transform 1 0 35880 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_564
timestamp 1586364061
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__433__A
timestamp 1586364061
transform 1 0 36892 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38088 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_48_377
timestamp 1586364061
transform 1 0 35788 0 -1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_48_387
timestamp 1586364061
transform 1 0 36708 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_48_391
timestamp 1586364061
transform 1 0 37076 0 -1 28832
box -38 -48 590 592
use scs8hd_decap_4  FILLER_48_398
timestamp 1586364061
transform 1 0 37720 0 -1 28832
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 38364 0 -1 28832
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40112 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39928 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_48_404
timestamp 1586364061
transform 1 0 38272 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_6  FILLER_48_416
timestamp 1586364061
transform 1 0 39376 0 -1 28832
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41124 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_433
timestamp 1586364061
transform 1 0 40940 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_437
timestamp 1586364061
transform 1 0 41308 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_8  FILLER_48_450
timestamp 1586364061
transform 1 0 42504 0 -1 28832
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_565
timestamp 1586364061
transform 1 0 43240 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_459
timestamp 1586364061
transform 1 0 43332 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_471
timestamp 1586364061
transform 1 0 44436 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_483
timestamp 1586364061
transform 1 0 45540 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_495
timestamp 1586364061
transform 1 0 46644 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_48_507
timestamp 1586364061
transform 1 0 47748 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 48852 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_48_515
timestamp 1586364061
transform 1 0 48484 0 -1 28832
box -38 -48 130 592
use scs8hd_nor2_4  _244_
timestamp 1586364061
transform 1 0 2668 0 1 28832
box -38 -48 866 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__244__A
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_49_26
timestamp 1586364061
transform 1 0 3496 0 1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 4232 0 1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__257__A
timestamp 1586364061
transform 1 0 5796 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_30
timestamp 1586364061
transform 1 0 3864 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_45
timestamp 1586364061
transform 1 0 5244 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_49
timestamp 1586364061
transform 1 0 5612 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_53
timestamp 1586364061
transform 1 0 5980 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_57
timestamp 1586364061
transform 1 0 6348 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__257__B
timestamp 1586364061
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_566
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 866 592
use scs8hd_fill_2  FILLER_49_71
timestamp 1586364061
transform 1 0 7636 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_79
timestamp 1586364061
transform 1 0 8372 0 1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_49_75
timestamp 1586364061
transform 1 0 8004 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 28832
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9016 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__273__A
timestamp 1586364061
transform 1 0 10764 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_83
timestamp 1586364061
transform 1 0 8740 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_95
timestamp 1586364061
transform 1 0 9844 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_99
timestamp 1586364061
transform 1 0 10212 0 1 28832
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_567
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__273__B
timestamp 1586364061
transform 1 0 11408 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_110
timestamp 1586364061
transform 1 0 11224 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_114
timestamp 1586364061
transform 1 0 11592 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_118
timestamp 1586364061
transform 1 0 11960 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_132
timestamp 1586364061
transform 1 0 13248 0 1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_49_139
timestamp 1586364061
transform 1 0 13892 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_136
timestamp 1586364061
transform 1 0 13616 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13708 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 866 592
use scs8hd_fill_2  FILLER_49_152
timestamp 1586364061
transform 1 0 15088 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_160
timestamp 1586364061
transform 1 0 15824 0 1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_49_156
timestamp 1586364061
transform 1 0 15456 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 28832
box -38 -48 222 592
use scs8hd_inv_8  _632_
timestamp 1586364061
transform 1 0 18216 0 1 28832
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_568
timestamp 1586364061
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__519__B
timestamp 1586364061
transform 1 0 17756 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_175
timestamp 1586364061
transform 1 0 17204 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_179
timestamp 1586364061
transform 1 0 17572 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_184
timestamp 1586364061
transform 1 0 18032 0 1 28832
box -38 -48 222 592
use scs8hd_nor2_4  _524_
timestamp 1586364061
transform 1 0 19872 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__519__A
timestamp 1586364061
transform 1 0 19228 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__524__A
timestamp 1586364061
transform 1 0 19688 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_195
timestamp 1586364061
transform 1 0 19044 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_199
timestamp 1586364061
transform 1 0 19412 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_213
timestamp 1586364061
transform 1 0 20700 0 1 28832
box -38 -48 314 592
use scs8hd_nor2_4  _507_
timestamp 1586364061
transform 1 0 21988 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__507__A
timestamp 1586364061
transform 1 0 21804 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__508__A
timestamp 1586364061
transform 1 0 20976 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__508__B
timestamp 1586364061
transform 1 0 21344 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_218
timestamp 1586364061
transform 1 0 21160 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_222
timestamp 1586364061
transform 1 0 21528 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_236
timestamp 1586364061
transform 1 0 22816 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_240
timestamp 1586364061
transform 1 0 23184 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_249
timestamp 1586364061
transform 1 0 24012 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_245
timestamp 1586364061
transform 1 0 23644 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23828 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23368 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__506__A
timestamp 1586364061
transform 1 0 24196 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_569
timestamp 1586364061
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use scs8hd_buf_1  _506_
timestamp 1586364061
transform 1 0 24380 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_260
timestamp 1586364061
transform 1 0 25024 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_256
timestamp 1586364061
transform 1 0 24656 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 25208 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 24840 0 1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 25392 0 1 28832
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 27140 0 1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 26956 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_275
timestamp 1586364061
transform 1 0 26404 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_279
timestamp 1586364061
transform 1 0 26772 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_294
timestamp 1586364061
transform 1 0 28152 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_298
timestamp 1586364061
transform 1 0 28520 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__499__B
timestamp 1586364061
transform 1 0 28704 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__499__A
timestamp 1586364061
transform 1 0 28336 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_302
timestamp 1586364061
transform 1 0 28888 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_309
timestamp 1586364061
transform 1 0 29532 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_570
timestamp 1586364061
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use scs8hd_buf_1  _505_
timestamp 1586364061
transform 1 0 29256 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_313
timestamp 1586364061
transform 1 0 29900 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__505__A
timestamp 1586364061
transform 1 0 29716 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_317
timestamp 1586364061
transform 1 0 30268 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__475__B
timestamp 1586364061
transform 1 0 30084 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__475__A
timestamp 1586364061
transform 1 0 30452 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_321
timestamp 1586364061
transform 1 0 30636 0 1 28832
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 31188 0 1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 31004 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__478__A
timestamp 1586364061
transform 1 0 32384 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__478__B
timestamp 1586364061
transform 1 0 32752 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_338
timestamp 1586364061
transform 1 0 32200 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_342
timestamp 1586364061
transform 1 0 32568 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_346
timestamp 1586364061
transform 1 0 32936 0 1 28832
box -38 -48 590 592
use scs8hd_fill_2  FILLER_49_356
timestamp 1586364061
transform 1 0 33856 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_352
timestamp 1586364061
transform 1 0 33488 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34040 0 1 28832
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33580 0 1 28832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_49_367
timestamp 1586364061
transform 1 0 34868 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_364
timestamp 1586364061
transform 1 0 34592 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_360
timestamp 1586364061
transform 1 0 34224 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34408 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_571
timestamp 1586364061
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use scs8hd_nor2_4  _435_
timestamp 1586364061
transform 1 0 34960 0 1 28832
box -38 -48 866 592
use scs8hd_nor2_4  _433_
timestamp 1586364061
transform 1 0 36524 0 1 28832
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 38088 0 1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 37904 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__431__A
timestamp 1586364061
transform 1 0 36064 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__433__B
timestamp 1586364061
transform 1 0 37536 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_377
timestamp 1586364061
transform 1 0 35788 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_382
timestamp 1586364061
transform 1 0 36248 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_394
timestamp 1586364061
transform 1 0 37352 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_398
timestamp 1586364061
transform 1 0 37720 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_572
timestamp 1586364061
transform 1 0 40388 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 39284 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39652 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_413
timestamp 1586364061
transform 1 0 39100 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_417
timestamp 1586364061
transform 1 0 39468 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_421
timestamp 1586364061
transform 1 0 39836 0 1 28832
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42044 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41860 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41492 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_437
timestamp 1586364061
transform 1 0 41308 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_441
timestamp 1586364061
transform 1 0 41676 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_454
timestamp 1586364061
transform 1 0 42872 0 1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43700 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_458
timestamp 1586364061
transform 1 0 43240 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_461
timestamp 1586364061
transform 1 0 43516 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_465
timestamp 1586364061
transform 1 0 43884 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_477
timestamp 1586364061
transform 1 0 44988 0 1 28832
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_573
timestamp 1586364061
transform 1 0 46000 0 1 28832
box -38 -48 130 592
use scs8hd_decap_3  FILLER_49_485
timestamp 1586364061
transform 1 0 45724 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_489
timestamp 1586364061
transform 1 0 46092 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_501
timestamp 1586364061
transform 1 0 47196 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 48852 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_513
timestamp 1586364061
transform 1 0 48300 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__248__B
timestamp 1586364061
transform 1 0 3220 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_4  FILLER_50_25
timestamp 1586364061
transform 1 0 3404 0 -1 29920
box -38 -48 406 592
use scs8hd_nor2_4  _257_
timestamp 1586364061
transform 1 0 5796 0 -1 29920
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_574
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__251__B
timestamp 1586364061
transform 1 0 5244 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_43
timestamp 1586364061
transform 1 0 5060 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_47
timestamp 1586364061
transform 1 0 5428 0 -1 29920
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_60
timestamp 1586364061
transform 1 0 6624 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_64
timestamp 1586364061
transform 1 0 6992 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_50_77
timestamp 1586364061
transform 1 0 8188 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_87
timestamp 1586364061
transform 1 0 9108 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_4  FILLER_50_81
timestamp 1586364061
transform 1 0 8556 0 -1 29920
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_97
timestamp 1586364061
transform 1 0 10028 0 -1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 130 592
use scs8hd_fill_1  FILLER_50_91
timestamp 1586364061
transform 1 0 9476 0 -1 29920
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_575
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _273_
timestamp 1586364061
transform 1 0 10764 0 -1 29920
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12328 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__285__B
timestamp 1586364061
transform 1 0 13340 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_114
timestamp 1586364061
transform 1 0 11592 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_118
timestamp 1586364061
transform 1 0 11960 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_50_131
timestamp 1586364061
transform 1 0 13156 0 -1 29920
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13892 0 -1 29920
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_576
timestamp 1586364061
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14352 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13708 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_135
timestamp 1586364061
transform 1 0 13524 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_142
timestamp 1586364061
transform 1 0 14168 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_146
timestamp 1586364061
transform 1 0 14536 0 -1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_50_152
timestamp 1586364061
transform 1 0 15088 0 -1 29920
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__632__A
timestamp 1586364061
transform 1 0 18216 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_163
timestamp 1586364061
transform 1 0 16100 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_6  FILLER_50_180
timestamp 1586364061
transform 1 0 17664 0 -1 29920
box -38 -48 590 592
use scs8hd_nor2_4  _519_
timestamp 1586364061
transform 1 0 18400 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_577
timestamp 1586364061
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__524__B
timestamp 1586364061
transform 1 0 19872 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_197
timestamp 1586364061
transform 1 0 19228 0 -1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_50_203
timestamp 1586364061
transform 1 0 19780 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_206
timestamp 1586364061
transform 1 0 20056 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_50_212
timestamp 1586364061
transform 1 0 20608 0 -1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _508_
timestamp 1586364061
transform 1 0 20976 0 -1 29920
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 22540 0 -1 29920
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_50_215
timestamp 1586364061
transform 1 0 20884 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_50_225
timestamp 1586364061
transform 1 0 21804 0 -1 29920
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 24288 0 -1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25484 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23736 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_244
timestamp 1586364061
transform 1 0 23552 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_248
timestamp 1586364061
transform 1 0 23920 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_263
timestamp 1586364061
transform 1 0 25300 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_267
timestamp 1586364061
transform 1 0 25668 0 -1 29920
box -38 -48 590 592
use scs8hd_nor2_4  _499_
timestamp 1586364061
transform 1 0 28152 0 -1 29920
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_578
timestamp 1586364061
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_285
timestamp 1586364061
transform 1 0 27324 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_1  FILLER_50_293
timestamp 1586364061
transform 1 0 28060 0 -1 29920
box -38 -48 130 592
use scs8hd_nor2_4  _475_
timestamp 1586364061
transform 1 0 30452 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__477__B
timestamp 1586364061
transform 1 0 29900 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_303
timestamp 1586364061
transform 1 0 28980 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_50_311
timestamp 1586364061
transform 1 0 29716 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_315
timestamp 1586364061
transform 1 0 30084 0 -1 29920
box -38 -48 406 592
use scs8hd_nor2_4  _478_
timestamp 1586364061
transform 1 0 32108 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_579
timestamp 1586364061
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_328
timestamp 1586364061
transform 1 0 31280 0 -1 29920
box -38 -48 590 592
use scs8hd_decap_8  FILLER_50_346
timestamp 1586364061
transform 1 0 32936 0 -1 29920
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33672 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_357
timestamp 1586364061
transform 1 0 33948 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34132 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_361
timestamp 1586364061
transform 1 0 34316 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34500 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_368
timestamp 1586364061
transform 1 0 34960 0 -1 29920
box -38 -48 222 592
use scs8hd_buf_1  _421_
timestamp 1586364061
transform 1 0 34684 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__421__A
timestamp 1586364061
transform 1 0 35144 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_372
timestamp 1586364061
transform 1 0 35328 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__435__B
timestamp 1586364061
transform 1 0 35512 0 -1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _431_
timestamp 1586364061
transform 1 0 36064 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_580
timestamp 1586364061
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__431__B
timestamp 1586364061
transform 1 0 35880 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_376
timestamp 1586364061
transform 1 0 35696 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_389
timestamp 1586364061
transform 1 0 36892 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_8  FILLER_50_398
timestamp 1586364061
transform 1 0 37720 0 -1 29920
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 38640 0 -1 29920
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40388 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40204 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_406
timestamp 1586364061
transform 1 0 38456 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_419
timestamp 1586364061
transform 1 0 39652 0 -1 29920
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41952 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41400 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42412 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_436
timestamp 1586364061
transform 1 0 41216 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_440
timestamp 1586364061
transform 1 0 41584 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_50_447
timestamp 1586364061
transform 1 0 42228 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_451
timestamp 1586364061
transform 1 0 42596 0 -1 29920
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_581
timestamp 1586364061
transform 1 0 43240 0 -1 29920
box -38 -48 130 592
use scs8hd_fill_1  FILLER_50_457
timestamp 1586364061
transform 1 0 43148 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_468
timestamp 1586364061
transform 1 0 44160 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_480
timestamp 1586364061
transform 1 0 45264 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_492
timestamp 1586364061
transform 1 0 46368 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_504
timestamp 1586364061
transform 1 0 47472 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 48852 0 -1 29920
box -38 -48 314 592
use scs8hd_nor2_4  _248_
timestamp 1586364061
transform 1 0 3220 0 1 29920
box -38 -48 866 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__248__A
timestamp 1586364061
transform 1 0 3036 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 590 592
use scs8hd_nor2_4  _251_
timestamp 1586364061
transform 1 0 4784 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__251__A
timestamp 1586364061
transform 1 0 4600 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_32
timestamp 1586364061
transform 1 0 4048 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_36
timestamp 1586364061
transform 1 0 4416 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_49
timestamp 1586364061
transform 1 0 5612 0 1 29920
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_582
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_55
timestamp 1586364061
transform 1 0 6164 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_77
timestamp 1586364061
transform 1 0 8188 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 29920
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 10580 0 1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_81
timestamp 1586364061
transform 1 0 8556 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_94
timestamp 1586364061
transform 1 0 9752 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_98
timestamp 1586364061
transform 1 0 10120 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_114
timestamp 1586364061
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_118
timestamp 1586364061
transform 1 0 11960 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_583
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_128
timestamp 1586364061
transform 1 0 12880 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__285__A
timestamp 1586364061
transform 1 0 13064 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_132
timestamp 1586364061
transform 1 0 13248 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 29920
box -38 -48 222 592
use scs8hd_inv_8  _631_
timestamp 1586364061
transform 1 0 15640 0 1 29920
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 13616 0 1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__629__A
timestamp 1586364061
transform 1 0 15364 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__631__A
timestamp 1586364061
transform 1 0 14996 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_147
timestamp 1586364061
transform 1 0 14628 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_153
timestamp 1586364061
transform 1 0 15180 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_157
timestamp 1586364061
transform 1 0 15548 0 1 29920
box -38 -48 130 592
use scs8hd_nor2_4  _518_
timestamp 1586364061
transform 1 0 18308 0 1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_584
timestamp 1586364061
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__518__B
timestamp 1586364061
transform 1 0 17756 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__630__A
timestamp 1586364061
transform 1 0 16928 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_167
timestamp 1586364061
transform 1 0 16468 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_171
timestamp 1586364061
transform 1 0 16836 0 1 29920
box -38 -48 130 592
use scs8hd_decap_6  FILLER_51_174
timestamp 1586364061
transform 1 0 17112 0 1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_51_180
timestamp 1586364061
transform 1 0 17664 0 1 29920
box -38 -48 130 592
use scs8hd_decap_3  FILLER_51_184
timestamp 1586364061
transform 1 0 18032 0 1 29920
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20424 0 1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 19320 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20240 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19688 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_196
timestamp 1586364061
transform 1 0 19136 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_200
timestamp 1586364061
transform 1 0 19504 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_204
timestamp 1586364061
transform 1 0 19872 0 1 29920
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__517__A
timestamp 1586364061
transform 1 0 21620 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_221
timestamp 1586364061
transform 1 0 21436 0 1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_51_225
timestamp 1586364061
transform 1 0 21804 0 1 29920
box -38 -48 590 592
use scs8hd_fill_2  FILLER_51_236
timestamp 1586364061
transform 1 0 22816 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_240
timestamp 1586364061
transform 1 0 23184 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_245
timestamp 1586364061
transform 1 0 23644 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_585
timestamp 1586364061
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23736 0 1 29920
box -38 -48 866 592
use scs8hd_decap_4  FILLER_51_259
timestamp 1586364061
transform 1 0 24932 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_255
timestamp 1586364061
transform 1 0 24564 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24748 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_267
timestamp 1586364061
transform 1 0 25668 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_263
timestamp 1586364061
transform 1 0 25300 0 1 29920
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_271
timestamp 1586364061
transform 1 0 26036 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26220 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26404 0 1 29920
box -38 -48 866 592
use scs8hd_fill_2  FILLER_51_288
timestamp 1586364061
transform 1 0 27600 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_284
timestamp 1586364061
transform 1 0 27232 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_295
timestamp 1586364061
transform 1 0 28244 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27784 0 1 29920
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27968 0 1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_51_304
timestamp 1586364061
transform 1 0 29072 0 1 29920
box -38 -48 130 592
use scs8hd_decap_3  FILLER_51_299
timestamp 1586364061
transform 1 0 28612 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__473__A
timestamp 1586364061
transform 1 0 28888 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28428 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_586
timestamp 1586364061
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use scs8hd_buf_1  _417_
timestamp 1586364061
transform 1 0 29256 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_317
timestamp 1586364061
transform 1 0 30268 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_313
timestamp 1586364061
transform 1 0 29900 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_309
timestamp 1586364061
transform 1 0 29532 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__477__A
timestamp 1586364061
transform 1 0 30084 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__417__A
timestamp 1586364061
transform 1 0 29716 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 30452 0 1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 30636 0 1 29920
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 33028 0 1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 32844 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32476 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32108 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_332
timestamp 1586364061
transform 1 0 31648 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_336
timestamp 1586364061
transform 1 0 32016 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_339
timestamp 1586364061
transform 1 0 32292 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_343
timestamp 1586364061
transform 1 0 32660 0 1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _434_
timestamp 1586364061
transform 1 0 34960 0 1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_587
timestamp 1586364061
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__434__A
timestamp 1586364061
transform 1 0 34592 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__434__B
timestamp 1586364061
transform 1 0 34224 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_358
timestamp 1586364061
transform 1 0 34040 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_362
timestamp 1586364061
transform 1 0 34408 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_367
timestamp 1586364061
transform 1 0 34868 0 1 29920
box -38 -48 130 592
use scs8hd_nor2_4  _432_
timestamp 1586364061
transform 1 0 36524 0 1 29920
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38088 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__425__A
timestamp 1586364061
transform 1 0 37720 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__432__A
timestamp 1586364061
transform 1 0 36340 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__432__B
timestamp 1586364061
transform 1 0 35972 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_377
timestamp 1586364061
transform 1 0 35788 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_381
timestamp 1586364061
transform 1 0 36156 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_394
timestamp 1586364061
transform 1 0 37352 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_400
timestamp 1586364061
transform 1 0 37904 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_405
timestamp 1586364061
transform 1 0 38364 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38548 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_409
timestamp 1586364061
transform 1 0 38732 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__407__A
timestamp 1586364061
transform 1 0 38916 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_416
timestamp 1586364061
transform 1 0 39376 0 1 29920
box -38 -48 406 592
use scs8hd_buf_1  _429_
timestamp 1586364061
transform 1 0 39100 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__415__A
timestamp 1586364061
transform 1 0 39744 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_426
timestamp 1586364061
transform 1 0 40296 0 1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_51_422
timestamp 1586364061
transform 1 0 39928 0 1 29920
box -38 -48 406 592
use scs8hd_decap_3  FILLER_51_428
timestamp 1586364061
transform 1 0 40480 0 1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_588
timestamp 1586364061
transform 1 0 40388 0 1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 40940 0 1 29920
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42688 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 40756 0 1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_51_444
timestamp 1586364061
transform 1 0 41952 0 1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_51_455
timestamp 1586364061
transform 1 0 42964 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43148 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_459
timestamp 1586364061
transform 1 0 43332 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_471
timestamp 1586364061
transform 1 0 44436 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_51_483
timestamp 1586364061
transform 1 0 45540 0 1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_589
timestamp 1586364061
transform 1 0 46000 0 1 29920
box -38 -48 130 592
use scs8hd_fill_1  FILLER_51_487
timestamp 1586364061
transform 1 0 45908 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_489
timestamp 1586364061
transform 1 0 46092 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_501
timestamp 1586364061
transform 1 0 47196 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 48852 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_513
timestamp 1586364061
transform 1 0 48300 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_34
timestamp 1586364061
transform 1 0 4232 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_31
timestamp 1586364061
transform 1 0 3956 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__586__A
timestamp 1586364061
transform 1 0 4048 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_590
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 4232 0 -1 31008
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 1 31008
box -38 -48 314 592
use scs8hd_decap_4  FILLER_53_50
timestamp 1586364061
transform 1 0 5704 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_43
timestamp 1586364061
transform 1 0 5060 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_45
timestamp 1586364061
transform 1 0 5244 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5612 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__586__B
timestamp 1586364061
transform 1 0 4876 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_52_51
timestamp 1586364061
transform 1 0 5796 0 -1 31008
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 31008
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_53_57
timestamp 1586364061
transform 1 0 6348 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_54
timestamp 1586364061
transform 1 0 6072 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__596__A
timestamp 1586364061
transform 1 0 6164 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_598
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_71
timestamp 1586364061
transform 1 0 7636 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_64
timestamp 1586364061
transform 1 0 6992 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__596__B
timestamp 1586364061
transform 1 0 7176 0 -1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_79
timestamp 1586364061
transform 1 0 8372 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_75
timestamp 1586364061
transform 1 0 8004 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_92
timestamp 1586364061
transform 1 0 9568 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_91
timestamp 1586364061
transform 1 0 9476 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_6  FILLER_52_85
timestamp 1586364061
transform 1 0 8924 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_2  FILLER_52_81
timestamp 1586364061
transform 1 0 8556 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_591
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 31008
box -38 -48 866 592
use scs8hd_decap_3  FILLER_53_100
timestamp 1586364061
transform 1 0 10304 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_96
timestamp 1586364061
transform 1 0 9936 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_99
timestamp 1586364061
transform 1 0 10212 0 -1 31008
box -38 -48 590 592
use scs8hd_decap_3  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__597__B
timestamp 1586364061
transform 1 0 10120 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__597__A
timestamp 1586364061
transform 1 0 9752 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__277__A
timestamp 1586364061
transform 1 0 10580 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__277__B
timestamp 1586364061
transform 1 0 10764 0 -1 31008
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 10948 0 -1 31008
box -38 -48 1050 592
use scs8hd_nor2_4  _277_
timestamp 1586364061
transform 1 0 10764 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_114
timestamp 1586364061
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__589__A
timestamp 1586364061
transform 1 0 11776 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_118
timestamp 1586364061
transform 1 0 11960 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_126
timestamp 1586364061
transform 1 0 12696 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_2  FILLER_52_122
timestamp 1586364061
transform 1 0 12328 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_118
timestamp 1586364061
transform 1 0 11960 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__589__B
timestamp 1586364061
transform 1 0 12144 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_599
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_132
timestamp 1586364061
transform 1 0 13248 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__588__A
timestamp 1586364061
transform 1 0 13432 0 1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _285_
timestamp 1586364061
transform 1 0 13248 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_1  FILLER_53_144
timestamp 1586364061
transform 1 0 14352 0 1 31008
box -38 -48 130 592
use scs8hd_decap_8  FILLER_53_136
timestamp 1586364061
transform 1 0 13616 0 1 31008
box -38 -48 774 592
use scs8hd_decap_12  FILLER_52_141
timestamp 1586364061
transform 1 0 14076 0 -1 31008
box -38 -48 1142 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 14444 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_152
timestamp 1586364061
transform 1 0 15088 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_148
timestamp 1586364061
transform 1 0 14720 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_154
timestamp 1586364061
transform 1 0 15272 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__628__A
timestamp 1586364061
transform 1 0 15272 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 14904 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_592
timestamp 1586364061
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use scs8hd_inv_8  _629_
timestamp 1586364061
transform 1 0 15364 0 -1 31008
box -38 -48 866 592
use scs8hd_inv_8  _628_
timestamp 1586364061
transform 1 0 15456 0 1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_53_169
timestamp 1586364061
transform 1 0 16652 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_165
timestamp 1586364061
transform 1 0 16284 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_164
timestamp 1586364061
transform 1 0 16192 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16468 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_179
timestamp 1586364061
transform 1 0 17572 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_175
timestamp 1586364061
transform 1 0 17204 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__521__B
timestamp 1586364061
transform 1 0 17388 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__521__A
timestamp 1586364061
transform 1 0 17020 0 1 31008
box -38 -48 222 592
use scs8hd_inv_8  _630_
timestamp 1586364061
transform 1 0 16928 0 -1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_53_184
timestamp 1586364061
transform 1 0 18032 0 1 31008
box -38 -48 406 592
use scs8hd_decap_6  FILLER_52_181
timestamp 1586364061
transform 1 0 17756 0 -1 31008
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__518__A
timestamp 1586364061
transform 1 0 18308 0 -1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_600
timestamp 1586364061
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_190
timestamp 1586364061
transform 1 0 18584 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_189
timestamp 1586364061
transform 1 0 18492 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 18768 0 1 31008
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 18860 0 -1 31008
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 18952 0 1 31008
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_53_209
timestamp 1586364061
transform 1 0 20332 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_205
timestamp 1586364061
transform 1 0 19964 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_204
timestamp 1586364061
transform 1 0 19872 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_212
timestamp 1586364061
transform 1 0 20608 0 -1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_593
timestamp 1586364061
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 20700 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_224
timestamp 1586364061
transform 1 0 21712 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_220
timestamp 1586364061
transform 1 0 21344 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_216
timestamp 1586364061
transform 1 0 20976 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_218
timestamp 1586364061
transform 1 0 21160 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 21160 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 31008
box -38 -48 222 592
use scs8hd_buf_1  _517_
timestamp 1586364061
transform 1 0 20884 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_232
timestamp 1586364061
transform 1 0 22448 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_228
timestamp 1586364061
transform 1 0 22080 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__510__A
timestamp 1586364061
transform 1 0 21896 0 -1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 -1 31008
box -38 -48 314 592
use scs8hd_nor2_4  _510_
timestamp 1586364061
transform 1 0 21896 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_239
timestamp 1586364061
transform 1 0 23092 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_235
timestamp 1586364061
transform 1 0 22724 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_236
timestamp 1586364061
transform 1 0 22816 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23276 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 22908 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_249
timestamp 1586364061
transform 1 0 24012 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_245
timestamp 1586364061
transform 1 0 23644 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_243
timestamp 1586364061
transform 1 0 23460 0 1 31008
box -38 -48 130 592
use scs8hd_fill_1  FILLER_52_244
timestamp 1586364061
transform 1 0 23552 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__512__A
timestamp 1586364061
transform 1 0 24104 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_601
timestamp 1586364061
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_261
timestamp 1586364061
transform 1 0 25116 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_258
timestamp 1586364061
transform 1 0 24840 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_254
timestamp 1586364061
transform 1 0 24472 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__512__B
timestamp 1586364061
transform 1 0 24656 0 -1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _512_
timestamp 1586364061
transform 1 0 24288 0 1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_53_265
timestamp 1586364061
transform 1 0 25484 0 1 31008
box -38 -48 406 592
use scs8hd_decap_6  FILLER_52_267
timestamp 1586364061
transform 1 0 25668 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_2  FILLER_52_262
timestamp 1586364061
transform 1 0 25208 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25300 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_275
timestamp 1586364061
transform 1 0 26404 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_271
timestamp 1586364061
transform 1 0 26036 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25852 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26220 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26588 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_594
timestamp 1586364061
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26772 0 1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 31008
box -38 -48 866 592
use scs8hd_decap_8  FILLER_53_292
timestamp 1586364061
transform 1 0 27968 0 1 31008
box -38 -48 774 592
use scs8hd_fill_2  FILLER_53_288
timestamp 1586364061
transform 1 0 27600 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_285
timestamp 1586364061
transform 1 0 27324 0 -1 31008
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27784 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_300
timestamp 1586364061
transform 1 0 28704 0 1 31008
box -38 -48 314 592
use scs8hd_decap_4  FILLER_52_305
timestamp 1586364061
transform 1 0 29164 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_52_301
timestamp 1586364061
transform 1 0 28796 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_297
timestamp 1586364061
transform 1 0 28428 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__479__A
timestamp 1586364061
transform 1 0 28980 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_602
timestamp 1586364061
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use scs8hd_buf_1  _473_
timestamp 1586364061
transform 1 0 28888 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_52_311
timestamp 1586364061
transform 1 0 29716 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29532 0 -1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _479_
timestamp 1586364061
transform 1 0 29256 0 1 31008
box -38 -48 866 592
use scs8hd_nor2_4  _477_
timestamp 1586364061
transform 1 0 29900 0 -1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_53_319
timestamp 1586364061
transform 1 0 30452 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_315
timestamp 1586364061
transform 1 0 30084 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_322
timestamp 1586364061
transform 1 0 30728 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_330
timestamp 1586364061
transform 1 0 31464 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_326
timestamp 1586364061
transform 1 0 31096 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_326
timestamp 1586364061
transform 1 0 31096 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30912 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__419__A
timestamp 1586364061
transform 1 0 31280 0 1 31008
box -38 -48 222 592
use scs8hd_buf_1  _419_
timestamp 1586364061
transform 1 0 30820 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_337
timestamp 1586364061
transform 1 0 32108 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31648 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_595
timestamp 1586364061
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32200 0 -1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31832 0 1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_53_347
timestamp 1586364061
transform 1 0 33028 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_343
timestamp 1586364061
transform 1 0 32660 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_52_347
timestamp 1586364061
transform 1 0 33028 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32844 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_356
timestamp 1586364061
transform 1 0 33856 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_352
timestamp 1586364061
transform 1 0 33488 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33672 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33396 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34040 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 31008
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33580 0 1 31008
box -38 -48 314 592
use scs8hd_decap_4  FILLER_53_360
timestamp 1586364061
transform 1 0 34224 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_52_365
timestamp 1586364061
transform 1 0 34684 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__424__A
timestamp 1586364061
transform 1 0 34868 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__424__B
timestamp 1586364061
transform 1 0 34592 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_603
timestamp 1586364061
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use scs8hd_nor2_4  _424_
timestamp 1586364061
transform 1 0 34868 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_52_369
timestamp 1586364061
transform 1 0 35052 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35236 0 -1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35420 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_380
timestamp 1586364061
transform 1 0 36064 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_376
timestamp 1586364061
transform 1 0 35696 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_382
timestamp 1586364061
transform 1 0 36248 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__416__A
timestamp 1586364061
transform 1 0 36432 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__416__B
timestamp 1586364061
transform 1 0 36248 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__426__B
timestamp 1586364061
transform 1 0 35880 0 1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _416_
timestamp 1586364061
transform 1 0 36432 0 1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_53_393
timestamp 1586364061
transform 1 0 37260 0 1 31008
box -38 -48 406 592
use scs8hd_decap_3  FILLER_52_394
timestamp 1586364061
transform 1 0 37352 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_8  FILLER_52_386
timestamp 1586364061
transform 1 0 36616 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_3  FILLER_53_400
timestamp 1586364061
transform 1 0 37904 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_53_397
timestamp 1586364061
transform 1 0 37628 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_52_401
timestamp 1586364061
transform 1 0 37996 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 37720 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_596
timestamp 1586364061
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use scs8hd_buf_1  _425_
timestamp 1586364061
transform 1 0 37720 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_410
timestamp 1586364061
transform 1 0 38824 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_406
timestamp 1586364061
transform 1 0 38456 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_405
timestamp 1586364061
transform 1 0 38364 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38180 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38640 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38180 0 1 31008
box -38 -48 314 592
use scs8hd_buf_1  _407_
timestamp 1586364061
transform 1 0 38732 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_417
timestamp 1586364061
transform 1 0 39468 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_416
timestamp 1586364061
transform 1 0 39376 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_52_412
timestamp 1586364061
transform 1 0 39008 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39008 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__429__A
timestamp 1586364061
transform 1 0 39192 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 39652 0 1 31008
box -38 -48 222 592
use scs8hd_buf_1  _415_
timestamp 1586364061
transform 1 0 39744 0 -1 31008
box -38 -48 314 592
use scs8hd_buf_1  _413_
timestamp 1586364061
transform 1 0 39192 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_425
timestamp 1586364061
transform 1 0 40204 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_421
timestamp 1586364061
transform 1 0 39836 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_423
timestamp 1586364061
transform 1 0 40020 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__413__A
timestamp 1586364061
transform 1 0 40020 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_604
timestamp 1586364061
transform 1 0 40388 0 1 31008
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_441
timestamp 1586364061
transform 1 0 41676 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_435
timestamp 1586364061
transform 1 0 41124 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_431
timestamp 1586364061
transform 1 0 40756 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_438
timestamp 1586364061
transform 1 0 41400 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_52_431
timestamp 1586364061
transform 1 0 40756 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40940 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 41492 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41124 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_454
timestamp 1586364061
transform 1 0 42872 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_450
timestamp 1586364061
transform 1 0 42504 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_445
timestamp 1586364061
transform 1 0 42044 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_450
timestamp 1586364061
transform 1 0 42504 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41860 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42688 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42228 0 1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_469
timestamp 1586364061
transform 1 0 44252 0 1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_465
timestamp 1586364061
transform 1 0 43884 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_461
timestamp 1586364061
transform 1 0 43516 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_459
timestamp 1586364061
transform 1 0 43332 0 -1 31008
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44068 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43700 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_597
timestamp 1586364061
transform 1 0 43240 0 -1 31008
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43240 0 1 31008
box -38 -48 314 592
use scs8hd_decap_6  FILLER_53_481
timestamp 1586364061
transform 1 0 45356 0 1 31008
box -38 -48 590 592
use scs8hd_decap_12  FILLER_52_471
timestamp 1586364061
transform 1 0 44436 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_483
timestamp 1586364061
transform 1 0 45540 0 -1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_605
timestamp 1586364061
transform 1 0 46000 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_495
timestamp 1586364061
transform 1 0 46644 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_52_507
timestamp 1586364061
transform 1 0 47748 0 -1 31008
box -38 -48 774 592
use scs8hd_fill_1  FILLER_53_487
timestamp 1586364061
transform 1 0 45908 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_53_489
timestamp 1586364061
transform 1 0 46092 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_501
timestamp 1586364061
transform 1 0 47196 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 48852 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 48852 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_515
timestamp 1586364061
transform 1 0 48484 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_513
timestamp 1586364061
transform 1 0 48300 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_nor2_4  _586_
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_606
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5428 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_6  FILLER_54_41
timestamp 1586364061
transform 1 0 4876 0 -1 32096
box -38 -48 590 592
use scs8hd_fill_2  FILLER_54_52
timestamp 1586364061
transform 1 0 5888 0 -1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _596_
timestamp 1586364061
transform 1 0 6900 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7912 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_54_56
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 590 592
use scs8hd_fill_1  FILLER_54_62
timestamp 1586364061
transform 1 0 6808 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_72
timestamp 1586364061
transform 1 0 7728 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_76
timestamp 1586364061
transform 1 0 8096 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 130 592
use scs8hd_nor2_4  _597_
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_607
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_54_84
timestamp 1586364061
transform 1 0 8832 0 -1 32096
box -38 -48 590 592
use scs8hd_decap_8  FILLER_54_102
timestamp 1586364061
transform 1 0 10488 0 -1 32096
box -38 -48 774 592
use scs8hd_buf_1  _588_
timestamp 1586364061
transform 1 0 13432 0 -1 32096
box -38 -48 314 592
use scs8hd_nor2_4  _589_
timestamp 1586364061
transform 1 0 11316 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__591__B
timestamp 1586364061
transform 1 0 13156 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__590__B
timestamp 1586364061
transform 1 0 12420 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_110
timestamp 1586364061
transform 1 0 11224 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  FILLER_54_120
timestamp 1586364061
transform 1 0 12144 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_6  FILLER_54_125
timestamp 1586364061
transform 1 0 12604 0 -1 32096
box -38 -48 590 592
use scs8hd_fill_1  FILLER_54_133
timestamp 1586364061
transform 1 0 13340 0 -1 32096
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_608
timestamp 1586364061
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__594__A
timestamp 1586364061
transform 1 0 15640 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__593__B
timestamp 1586364061
transform 1 0 14076 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_137
timestamp 1586364061
transform 1 0 13708 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_8  FILLER_54_143
timestamp 1586364061
transform 1 0 14260 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_2  FILLER_54_151
timestamp 1586364061
transform 1 0 14996 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_154
timestamp 1586364061
transform 1 0 15272 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_160
timestamp 1586364061
transform 1 0 15824 0 -1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _521_
timestamp 1586364061
transform 1 0 17020 0 -1 32096
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16008 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__520__B
timestamp 1586364061
transform 1 0 18032 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_165
timestamp 1586364061
transform 1 0 16284 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_2  FILLER_54_182
timestamp 1586364061
transform 1 0 17848 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_186
timestamp 1586364061
transform 1 0 18216 0 -1 32096
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_609
timestamp 1586364061
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_196
timestamp 1586364061
transform 1 0 19136 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_206
timestamp 1586364061
transform 1 0 20056 0 -1 32096
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 22632 0 -1 32096
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__510__B
timestamp 1586364061
transform 1 0 21988 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_215
timestamp 1586364061
transform 1 0 20884 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_221
timestamp 1586364061
transform 1 0 21436 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_225
timestamp 1586364061
transform 1 0 21804 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_229
timestamp 1586364061
transform 1 0 22172 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_233
timestamp 1586364061
transform 1 0 22540 0 -1 32096
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_245
timestamp 1586364061
transform 1 0 23644 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_249
timestamp 1586364061
transform 1 0 24012 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_262
timestamp 1586364061
transform 1 0 25208 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_266
timestamp 1586364061
transform 1 0 25576 0 -1 32096
box -38 -48 774 592
use scs8hd_conb_1  _641_
timestamp 1586364061
transform 1 0 28060 0 -1 32096
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_610
timestamp 1586364061
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27508 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_274
timestamp 1586364061
transform 1 0 26312 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_285
timestamp 1586364061
transform 1 0 27324 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_289
timestamp 1586364061
transform 1 0 27692 0 -1 32096
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 29532 0 -1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__479__B
timestamp 1586364061
transform 1 0 29256 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30728 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_296
timestamp 1586364061
transform 1 0 28336 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_2  FILLER_54_304
timestamp 1586364061
transform 1 0 29072 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_308
timestamp 1586364061
transform 1 0 29440 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_320
timestamp 1586364061
transform 1 0 30544 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_54_324
timestamp 1586364061
transform 1 0 30912 0 -1 32096
box -38 -48 590 592
use scs8hd_decap_3  FILLER_54_333
timestamp 1586364061
transform 1 0 31740 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_54_330
timestamp 1586364061
transform 1 0 31464 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__476__B
timestamp 1586364061
transform 1 0 31556 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_341
timestamp 1586364061
transform 1 0 32476 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_337
timestamp 1586364061
transform 1 0 32108 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32292 0 -1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_611
timestamp 1586364061
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_348
timestamp 1586364061
transform 1 0 33120 0 -1 32096
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32844 0 -1 32096
box -38 -48 314 592
use scs8hd_nor2_4  _426_
timestamp 1586364061
transform 1 0 35512 0 -1 32096
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__426__A
timestamp 1586364061
transform 1 0 35328 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33672 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_352
timestamp 1586364061
transform 1 0 33488 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_54_365
timestamp 1586364061
transform 1 0 34684 0 -1 32096
box -38 -48 590 592
use scs8hd_fill_1  FILLER_54_371
timestamp 1586364061
transform 1 0 35236 0 -1 32096
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_612
timestamp 1586364061
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37352 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_383
timestamp 1586364061
transform 1 0 36340 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  FILLER_54_391
timestamp 1586364061
transform 1 0 37076 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_54_396
timestamp 1586364061
transform 1 0 37536 0 -1 32096
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 39468 0 -1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38916 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_409
timestamp 1586364061
transform 1 0 38732 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_413
timestamp 1586364061
transform 1 0 39100 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_428
timestamp 1586364061
transform 1 0 40480 0 -1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 41492 0 -1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40664 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41032 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_432
timestamp 1586364061
transform 1 0 40848 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_54_436
timestamp 1586364061
transform 1 0 41216 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_8  FILLER_54_450
timestamp 1586364061
transform 1 0 42504 0 -1 32096
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_613
timestamp 1586364061
transform 1 0 43240 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_468
timestamp 1586364061
transform 1 0 44160 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_480
timestamp 1586364061
transform 1 0 45264 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_492
timestamp 1586364061
transform 1 0 46368 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_504
timestamp 1586364061
transform 1 0 47472 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 48852 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__583__A
timestamp 1586364061
transform 1 0 3496 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__583__B
timestamp 1586364061
transform 1 0 3128 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 590 592
use scs8hd_fill_1  FILLER_55_21
timestamp 1586364061
transform 1 0 3036 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_24
timestamp 1586364061
transform 1 0 3312 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _582_
timestamp 1586364061
transform 1 0 4048 0 1 32096
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__582__A
timestamp 1586364061
transform 1 0 3864 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__585__B
timestamp 1586364061
transform 1 0 5520 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__582__B
timestamp 1586364061
transform 1 0 5060 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_28
timestamp 1586364061
transform 1 0 3680 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_41
timestamp 1586364061
transform 1 0 4876 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_45
timestamp 1586364061
transform 1 0 5244 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_53
timestamp 1586364061
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_65
timestamp 1586364061
transform 1 0 7084 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_57
timestamp 1586364061
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__581__A
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__585__A
timestamp 1586364061
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_614
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_buf_1  _581_
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_70
timestamp 1586364061
transform 1 0 7544 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7360 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_85
timestamp 1586364061
transform 1 0 8924 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_89
timestamp 1586364061
transform 1 0 9292 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_104
timestamp 1586364061
transform 1 0 10672 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_114
timestamp 1586364061
transform 1 0 11592 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_108
timestamp 1586364061
transform 1 0 11040 0 1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_118
timestamp 1586364061
transform 1 0 11960 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__590__A
timestamp 1586364061
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_615
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_nor2_4  _590_
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 866 592
use scs8hd_fill_2  FILLER_55_132
timestamp 1586364061
transform 1 0 13248 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__591__A
timestamp 1586364061
transform 1 0 13432 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _593_
timestamp 1586364061
transform 1 0 14076 0 1 32096
box -38 -48 866 592
use scs8hd_nor2_4  _594_
timestamp 1586364061
transform 1 0 15640 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__593__A
timestamp 1586364061
transform 1 0 13892 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_136
timestamp 1586364061
transform 1 0 13616 0 1 32096
box -38 -48 314 592
use scs8hd_decap_4  FILLER_55_150
timestamp 1586364061
transform 1 0 14904 0 1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_55_156
timestamp 1586364061
transform 1 0 15456 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_167
timestamp 1586364061
transform 1 0 16468 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__594__B
timestamp 1586364061
transform 1 0 16652 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_179
timestamp 1586364061
transform 1 0 17572 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_175
timestamp 1586364061
transform 1 0 17204 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_171
timestamp 1586364061
transform 1 0 16836 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__520__A
timestamp 1586364061
transform 1 0 17756 0 1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_616
timestamp 1586364061
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use scs8hd_nor2_4  _520_
timestamp 1586364061
transform 1 0 18032 0 1 32096
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20700 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_193
timestamp 1586364061
transform 1 0 18860 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_198
timestamp 1586364061
transform 1 0 19320 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_211
timestamp 1586364061
transform 1 0 20516 0 1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 23184 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__509__A
timestamp 1586364061
transform 1 0 22264 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__509__B
timestamp 1586364061
transform 1 0 21068 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22816 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_215
timestamp 1586364061
transform 1 0 20884 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_228
timestamp 1586364061
transform 1 0 22080 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_232
timestamp 1586364061
transform 1 0 22448 0 1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_55_238
timestamp 1586364061
transform 1 0 23000 0 1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 25208 0 1 32096
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_617
timestamp 1586364061
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 25024 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_242
timestamp 1586364061
transform 1 0 23368 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_254
timestamp 1586364061
transform 1 0 24472 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_258
timestamp 1586364061
transform 1 0 24840 0 1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26956 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26496 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27968 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_273
timestamp 1586364061
transform 1 0 26220 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_278
timestamp 1586364061
transform 1 0 26680 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_290
timestamp 1586364061
transform 1 0 27784 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_294
timestamp 1586364061
transform 1 0 28152 0 1 32096
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 29808 0 1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_618
timestamp 1586364061
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 29624 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__474__A
timestamp 1586364061
transform 1 0 28888 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__474__B
timestamp 1586364061
transform 1 0 28520 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_300
timestamp 1586364061
transform 1 0 28704 0 1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_55_304
timestamp 1586364061
transform 1 0 29072 0 1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_55_306
timestamp 1586364061
transform 1 0 29256 0 1 32096
box -38 -48 406 592
use scs8hd_nor2_4  _476_
timestamp 1586364061
transform 1 0 31556 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 32568 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__476__A
timestamp 1586364061
transform 1 0 31372 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33028 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31004 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_323
timestamp 1586364061
transform 1 0 30820 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_327
timestamp 1586364061
transform 1 0 31188 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_340
timestamp 1586364061
transform 1 0 32384 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_344
timestamp 1586364061
transform 1 0 32752 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_358
timestamp 1586364061
transform 1 0 34040 0 1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 32096
box -38 -48 866 592
use scs8hd_decap_4  FILLER_55_367
timestamp 1586364061
transform 1 0 34868 0 1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_55_362
timestamp 1586364061
transform 1 0 34408 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_619
timestamp 1586364061
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_373
timestamp 1586364061
transform 1 0 35420 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__412__B
timestamp 1586364061
transform 1 0 35236 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__412__A
timestamp 1586364061
transform 1 0 35604 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _412_
timestamp 1586364061
transform 1 0 35788 0 1 32096
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 37352 0 1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 37168 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36800 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_386
timestamp 1586364061
transform 1 0 36616 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_390
timestamp 1586364061
transform 1 0 36984 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_409
timestamp 1586364061
transform 1 0 38732 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_405
timestamp 1586364061
transform 1 0 38364 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38916 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__411__A
timestamp 1586364061
transform 1 0 38548 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_419
timestamp 1586364061
transform 1 0 39652 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_413
timestamp 1586364061
transform 1 0 39100 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 32096
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39376 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_423
timestamp 1586364061
transform 1 0 40020 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_620
timestamp 1586364061
transform 1 0 40388 0 1 32096
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 32096
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42044 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41860 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_437
timestamp 1586364061
transform 1 0 41308 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_441
timestamp 1586364061
transform 1 0 41676 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_454
timestamp 1586364061
transform 1 0 42872 0 1 32096
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43608 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43332 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44620 0 1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_55_458
timestamp 1586364061
transform 1 0 43240 0 1 32096
box -38 -48 130 592
use scs8hd_fill_1  FILLER_55_461
timestamp 1586364061
transform 1 0 43516 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_471
timestamp 1586364061
transform 1 0 44436 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_475
timestamp 1586364061
transform 1 0 44804 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_621
timestamp 1586364061
transform 1 0 46000 0 1 32096
box -38 -48 130 592
use scs8hd_fill_1  FILLER_55_487
timestamp 1586364061
transform 1 0 45908 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_489
timestamp 1586364061
transform 1 0 46092 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_501
timestamp 1586364061
transform 1 0 47196 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 48852 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_513
timestamp 1586364061
transform 1 0 48300 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__584__B
timestamp 1586364061
transform 1 0 3404 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_56_23
timestamp 1586364061
transform 1 0 3220 0 -1 33184
box -38 -48 222 592
use scs8hd_nor2_4  _583_
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 866 592
use scs8hd_nor2_4  _585_
timestamp 1586364061
transform 1 0 5796 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_622
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__587__B
timestamp 1586364061
transform 1 0 5060 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_56_41
timestamp 1586364061
transform 1 0 4876 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_45
timestamp 1586364061
transform 1 0 5244 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_49
timestamp 1586364061
transform 1 0 5612 0 -1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_60
timestamp 1586364061
transform 1 0 6624 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_64
timestamp 1586364061
transform 1 0 6992 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_623
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_104
timestamp 1586364061
transform 1 0 10672 0 -1 33184
box -38 -48 774 592
use scs8hd_nor2_4  _591_
timestamp 1586364061
transform 1 0 13156 0 -1 33184
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__592__B
timestamp 1586364061
transform 1 0 12880 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_123
timestamp 1586364061
transform 1 0 12420 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_127
timestamp 1586364061
transform 1 0 12788 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_1  FILLER_56_130
timestamp 1586364061
transform 1 0 13064 0 -1 33184
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_624
timestamp 1586364061
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_140
timestamp 1586364061
transform 1 0 13984 0 -1 33184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_56_146
timestamp 1586364061
transform 1 0 14536 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_149
timestamp 1586364061
transform 1 0 14812 0 -1 33184
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 17388 0 -1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17204 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_165
timestamp 1586364061
transform 1 0 16284 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_56_173
timestamp 1586364061
transform 1 0 17020 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_192
timestamp 1586364061
transform 1 0 18768 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_188
timestamp 1586364061
transform 1 0 18400 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18952 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 33184
box -38 -48 866 592
use scs8hd_fill_2  FILLER_56_205
timestamp 1586364061
transform 1 0 19964 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_213
timestamp 1586364061
transform 1 0 20700 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_209
timestamp 1586364061
transform 1 0 20332 0 -1 33184
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_625
timestamp 1586364061
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use scs8hd_nor2_4  _509_
timestamp 1586364061
transform 1 0 21620 0 -1 33184
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 23184 0 -1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_215
timestamp 1586364061
transform 1 0 20884 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_219
timestamp 1586364061
transform 1 0 21252 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_1  FILLER_56_222
timestamp 1586364061
transform 1 0 21528 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_232
timestamp 1586364061
transform 1 0 22448 0 -1 33184
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25208 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_251
timestamp 1586364061
transform 1 0 24196 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_3  FILLER_56_259
timestamp 1586364061
transform 1 0 24932 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_56_267
timestamp 1586364061
transform 1 0 25668 0 -1 33184
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 33184
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27508 0 -1 33184
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_626
timestamp 1586364061
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26956 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27324 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_279
timestamp 1586364061
transform 1 0 26772 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_283
timestamp 1586364061
transform 1 0 27140 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_290
timestamp 1586364061
transform 1 0 27784 0 -1 33184
box -38 -48 774 592
use scs8hd_nor2_4  _474_
timestamp 1586364061
transform 1 0 28888 0 -1 33184
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__480__B
timestamp 1586364061
transform 1 0 28520 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29900 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_300
timestamp 1586364061
transform 1 0 28704 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_311
timestamp 1586364061
transform 1 0 29716 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_315
timestamp 1586364061
transform 1 0 30084 0 -1 33184
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_627
timestamp 1586364061
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_328
timestamp 1586364061
transform 1 0 31280 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_8  FILLER_56_348
timestamp 1586364061
transform 1 0 33120 0 -1 33184
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 33184
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35420 0 -1 33184
box -38 -48 866 592
use scs8hd_decap_8  FILLER_56_365
timestamp 1586364061
transform 1 0 34684 0 -1 33184
box -38 -48 774 592
use scs8hd_buf_1  _411_
timestamp 1586364061
transform 1 0 37720 0 -1 33184
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_628
timestamp 1586364061
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__414__B
timestamp 1586364061
transform 1 0 36432 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__418__A
timestamp 1586364061
transform 1 0 36800 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_382
timestamp 1586364061
transform 1 0 36248 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_386
timestamp 1586364061
transform 1 0 36616 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_390
timestamp 1586364061
transform 1 0 36984 0 -1 33184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_56_396
timestamp 1586364061
transform 1 0 37536 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_401
timestamp 1586364061
transform 1 0 37996 0 -1 33184
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40388 0 -1 33184
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38824 0 -1 33184
box -38 -48 866 592
use scs8hd_fill_1  FILLER_56_409
timestamp 1586364061
transform 1 0 38732 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_419
timestamp 1586364061
transform 1 0 39652 0 -1 33184
box -38 -48 774 592
use scs8hd_conb_1  _649_
timestamp 1586364061
transform 1 0 42228 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42688 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42044 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_436
timestamp 1586364061
transform 1 0 41216 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_1  FILLER_56_444
timestamp 1586364061
transform 1 0 41952 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_56_450
timestamp 1586364061
transform 1 0 42504 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_454
timestamp 1586364061
transform 1 0 42872 0 -1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 33184
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_629
timestamp 1586364061
transform 1 0 43240 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43792 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44160 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_462
timestamp 1586364061
transform 1 0 43608 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_466
timestamp 1586364061
transform 1 0 43976 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_56_470
timestamp 1586364061
transform 1 0 44344 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_482
timestamp 1586364061
transform 1 0 45448 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_494
timestamp 1586364061
transform 1 0 46552 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_56_506
timestamp 1586364061
transform 1 0 47656 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 48852 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_56_514
timestamp 1586364061
transform 1 0 48392 0 -1 33184
box -38 -48 222 592
use scs8hd_nor2_4  _584_
timestamp 1586364061
transform 1 0 3404 0 1 33184
box -38 -48 866 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__584__A
timestamp 1586364061
transform 1 0 3220 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 4968 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__587__A
timestamp 1586364061
transform 1 0 4416 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_34
timestamp 1586364061
transform 1 0 4232 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_38
timestamp 1586364061
transform 1 0 4600 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_53
timestamp 1586364061
transform 1 0 5980 0 1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_630
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_57
timestamp 1586364061
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_73
timestamp 1586364061
transform 1 0 7820 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_77
timestamp 1586364061
transform 1 0 8188 0 1 33184
box -38 -48 406 592
use scs8hd_decap_3  FILLER_57_83
timestamp 1586364061
transform 1 0 8740 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9200 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_91
timestamp 1586364061
transform 1 0 9476 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_95
timestamp 1586364061
transform 1 0 9844 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_102
timestamp 1586364061
transform 1 0 10488 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_106
timestamp 1586364061
transform 1 0 10856 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_114
timestamp 1586364061
transform 1 0 11592 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_118
timestamp 1586364061
transform 1 0 11960 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__592__A
timestamp 1586364061
transform 1 0 12696 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_631
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_nor2_4  _592_
timestamp 1586364061
transform 1 0 12880 0 1 33184
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14628 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__621__A
timestamp 1586364061
transform 1 0 15824 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_137
timestamp 1586364061
transform 1 0 13708 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_141
timestamp 1586364061
transform 1 0 14076 0 1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_57_158
timestamp 1586364061
transform 1 0 15640 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_162
timestamp 1586364061
transform 1 0 16008 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16192 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_169
timestamp 1586364061
transform 1 0 16652 0 1 33184
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 1 33184
box -38 -48 314 592
use scs8hd_fill_1  FILLER_57_173
timestamp 1586364061
transform 1 0 17020 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__522__A
timestamp 1586364061
transform 1 0 17112 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_180
timestamp 1586364061
transform 1 0 17664 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_176
timestamp 1586364061
transform 1 0 17296 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__522__B
timestamp 1586364061
transform 1 0 17480 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_184
timestamp 1586364061
transform 1 0 18032 0 1 33184
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_632
timestamp 1586364061
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18584 0 1 33184
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20332 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18400 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20792 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_201
timestamp 1586364061
transform 1 0 19596 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_205
timestamp 1586364061
transform 1 0 19964 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_212
timestamp 1586364061
transform 1 0 20608 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_216
timestamp 1586364061
transform 1 0 20976 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_229
timestamp 1586364061
transform 1 0 22172 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_234
timestamp 1586364061
transform 1 0 22632 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_238
timestamp 1586364061
transform 1 0 23000 0 1 33184
box -38 -48 406 592
use scs8hd_nor2_4  _511_
timestamp 1586364061
transform 1 0 23644 0 1 33184
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 33184
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_633
timestamp 1586364061
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__511__A
timestamp 1586364061
transform 1 0 23368 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_254
timestamp 1586364061
transform 1 0 24472 0 1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_57_258
timestamp 1586364061
transform 1 0 24840 0 1 33184
box -38 -48 590 592
use scs8hd_fill_2  FILLER_57_273
timestamp 1586364061
transform 1 0 26220 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_269
timestamp 1586364061
transform 1 0 25852 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26404 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26588 0 1 33184
box -38 -48 866 592
use scs8hd_fill_2  FILLER_57_286
timestamp 1586364061
transform 1 0 27416 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27600 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_290
timestamp 1586364061
transform 1 0 27784 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27968 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_301
timestamp 1586364061
transform 1 0 28796 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_297
timestamp 1586364061
transform 1 0 28428 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__480__A
timestamp 1586364061
transform 1 0 28980 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_634
timestamp 1586364061
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_313
timestamp 1586364061
transform 1 0 29900 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_309
timestamp 1586364061
transform 1 0 29532 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_317
timestamp 1586364061
transform 1 0 30268 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30084 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30452 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30636 0 1 33184
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31740 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_330
timestamp 1586364061
transform 1 0 31464 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_335
timestamp 1586364061
transform 1 0 31924 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_339
timestamp 1586364061
transform 1 0 32292 0 1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_57_353
timestamp 1586364061
transform 1 0 33580 0 1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_57_349
timestamp 1586364061
transform 1 0 33212 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33396 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_364
timestamp 1586364061
transform 1 0 34592 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_361
timestamp 1586364061
transform 1 0 34316 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34408 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_635
timestamp 1586364061
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_57_374
timestamp 1586364061
transform 1 0 35512 0 1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_57_370
timestamp 1586364061
transform 1 0 35144 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 33184
box -38 -48 314 592
use scs8hd_nor2_4  _418_
timestamp 1586364061
transform 1 0 36156 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 37720 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__418__B
timestamp 1586364061
transform 1 0 35972 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__414__A
timestamp 1586364061
transform 1 0 37168 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38088 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_378
timestamp 1586364061
transform 1 0 35880 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_390
timestamp 1586364061
transform 1 0 36984 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_394
timestamp 1586364061
transform 1 0 37352 0 1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_57_400
timestamp 1586364061
transform 1 0 37904 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 33184
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38732 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_636
timestamp 1586364061
transform 1 0 40388 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39836 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38548 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_404
timestamp 1586364061
transform 1 0 38272 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_418
timestamp 1586364061
transform 1 0 39560 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_423
timestamp 1586364061
transform 1 0 40020 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42596 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42228 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41860 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_437
timestamp 1586364061
transform 1 0 41308 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_441
timestamp 1586364061
transform 1 0 41676 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_445
timestamp 1586364061
transform 1 0 42044 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_449
timestamp 1586364061
transform 1 0 42412 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44160 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43976 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43608 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_460
timestamp 1586364061
transform 1 0 43424 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_464
timestamp 1586364061
transform 1 0 43792 0 1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_57_477
timestamp 1586364061
transform 1 0 44988 0 1 33184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_637
timestamp 1586364061
transform 1 0 46000 0 1 33184
box -38 -48 130 592
use scs8hd_decap_3  FILLER_57_485
timestamp 1586364061
transform 1 0 45724 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_489
timestamp 1586364061
transform 1 0 46092 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_501
timestamp 1586364061
transform 1 0 47196 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 48852 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_513
timestamp 1586364061
transform 1 0 48300 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_nor2_4  _587_
timestamp 1586364061
transform 1 0 4416 0 -1 34272
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5980 0 -1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_638
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_45
timestamp 1586364061
transform 1 0 5244 0 -1 34272
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7176 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 774 592
use scs8hd_fill_2  FILLER_58_64
timestamp 1586364061
transform 1 0 6992 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_73
timestamp 1586364061
transform 1 0 7820 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_58_79
timestamp 1586364061
transform 1 0 8372 0 -1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 34272
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_639
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_58_84
timestamp 1586364061
transform 1 0 8832 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_8  FILLER_58_102
timestamp 1586364061
transform 1 0 10488 0 -1 34272
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13340 0 -1 34272
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 34272
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_58_110
timestamp 1586364061
transform 1 0 11224 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_122
timestamp 1586364061
transform 1 0 12328 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_4  FILLER_58_128
timestamp 1586364061
transform 1 0 12880 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_132
timestamp 1586364061
transform 1 0 13248 0 -1 34272
box -38 -48 130 592
use scs8hd_inv_8  _621_
timestamp 1586364061
transform 1 0 15548 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_640
timestamp 1586364061
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_136
timestamp 1586364061
transform 1 0 13616 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_58_140
timestamp 1586364061
transform 1 0 13984 0 -1 34272
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_58_152
timestamp 1586364061
transform 1 0 15088 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  FILLER_58_154
timestamp 1586364061
transform 1 0 15272 0 -1 34272
box -38 -48 314 592
use scs8hd_nor2_4  _522_
timestamp 1586364061
transform 1 0 17112 0 -1 34272
box -38 -48 866 592
use scs8hd_decap_8  FILLER_58_166
timestamp 1586364061
transform 1 0 16376 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_4  FILLER_58_183
timestamp 1586364061
transform 1 0 17940 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_187
timestamp 1586364061
transform 1 0 18308 0 -1 34272
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_641
timestamp 1586364061
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18400 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_190
timestamp 1586364061
transform 1 0 18584 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_194
timestamp 1586364061
transform 1 0 18952 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_58_206
timestamp 1586364061
transform 1 0 20056 0 -1 34272
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 34272
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_224
timestamp 1586364061
transform 1 0 21712 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_228
timestamp 1586364061
transform 1 0 22080 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_8  FILLER_58_235
timestamp 1586364061
transform 1 0 22724 0 -1 34272
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 34272
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__511__B
timestamp 1586364061
transform 1 0 23644 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_243
timestamp 1586364061
transform 1 0 23460 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_250
timestamp 1586364061
transform 1 0 24104 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_254
timestamp 1586364061
transform 1 0 24472 0 -1 34272
box -38 -48 774 592
use scs8hd_fill_2  FILLER_58_262
timestamp 1586364061
transform 1 0 25208 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_267
timestamp 1586364061
transform 1 0 25668 0 -1 34272
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26680 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_642
timestamp 1586364061
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_276
timestamp 1586364061
transform 1 0 26496 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_287
timestamp 1586364061
transform 1 0 27508 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_3  FILLER_58_295
timestamp 1586364061
transform 1 0 28244 0 -1 34272
box -38 -48 314 592
use scs8hd_nor2_4  _480_
timestamp 1586364061
transform 1 0 28520 0 -1 34272
box -38 -48 866 592
use scs8hd_conb_1  _644_
timestamp 1586364061
transform 1 0 30360 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29532 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_307
timestamp 1586364061
transform 1 0 29348 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_311
timestamp 1586364061
transform 1 0 29716 0 -1 34272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_58_317
timestamp 1586364061
transform 1 0 30268 0 -1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_58_321
timestamp 1586364061
transform 1 0 30636 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_325
timestamp 1586364061
transform 1 0 31004 0 -1 34272
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30820 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_333
timestamp 1586364061
transform 1 0 31740 0 -1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_643
timestamp 1586364061
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_3  FILLER_58_348
timestamp 1586364061
transform 1 0 33120 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_58_344
timestamp 1586364061
transform 1 0 32752 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_340
timestamp 1586364061
transform 1 0 32384 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32936 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32568 0 -1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33396 0 -1 34272
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34408 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_58_354
timestamp 1586364061
transform 1 0 33672 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_58_365
timestamp 1586364061
transform 1 0 34684 0 -1 34272
box -38 -48 1142 592
use scs8hd_nor2_4  _414_
timestamp 1586364061
transform 1 0 36064 0 -1 34272
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 34272
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_644
timestamp 1586364061
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  FILLER_58_377
timestamp 1586364061
transform 1 0 35788 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_58_389
timestamp 1586364061
transform 1 0 36892 0 -1 34272
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40388 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39008 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39376 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_409
timestamp 1586364061
transform 1 0 38732 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_58_414
timestamp 1586364061
transform 1 0 39192 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_418
timestamp 1586364061
transform 1 0 39560 0 -1 34272
box -38 -48 774 592
use scs8hd_fill_1  FILLER_58_426
timestamp 1586364061
transform 1 0 40296 0 -1 34272
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42228 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42688 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41676 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_436
timestamp 1586364061
transform 1 0 41216 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_440
timestamp 1586364061
transform 1 0 41584 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_443
timestamp 1586364061
transform 1 0 41860 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_58_450
timestamp 1586364061
transform 1 0 42504 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_454
timestamp 1586364061
transform 1 0 42872 0 -1 34272
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_645
timestamp 1586364061
transform 1 0 43240 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_468
timestamp 1586364061
transform 1 0 44160 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_480
timestamp 1586364061
transform 1 0 45264 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_492
timestamp 1586364061
transform 1 0 46368 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_504
timestamp 1586364061
transform 1 0 47472 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 48852 0 -1 34272
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_32
timestamp 1586364061
transform 1 0 4048 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_28
timestamp 1586364061
transform 1 0 3680 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 3864 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_654
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 4324 0 -1 35360
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 4416 0 1 34272
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_60_46
timestamp 1586364061
transform 1 0 5336 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_47
timestamp 1586364061
transform 1 0 5428 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_60_65
timestamp 1586364061
transform 1 0 7084 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_60
timestamp 1586364061
transform 1 0 6624 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_56
timestamp 1586364061
transform 1 0 6256 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_646
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 6072 0 -1 35360
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_60_69
timestamp 1586364061
transform 1 0 7452 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_75
timestamp 1586364061
transform 1 0 8004 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_69
timestamp 1586364061
transform 1 0 7452 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 34272
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7176 0 1 34272
box -38 -48 314 592
use scs8hd_decap_6  FILLER_60_86
timestamp 1586364061
transform 1 0 9016 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_2  FILLER_60_82
timestamp 1586364061
transform 1 0 8648 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_90
timestamp 1586364061
transform 1 0 9384 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_86
timestamp 1586364061
transform 1 0 9016 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_655
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 34272
box -38 -48 866 592
use scs8hd_decap_6  FILLER_60_107
timestamp 1586364061
transform 1 0 10948 0 -1 35360
box -38 -48 590 592
use scs8hd_decap_3  FILLER_60_102
timestamp 1586364061
transform 1 0 10488 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_107
timestamp 1586364061
transform 1 0 10948 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_103
timestamp 1586364061
transform 1 0 10580 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_116
timestamp 1586364061
transform 1 0 11776 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_118
timestamp 1586364061
transform 1 0 11960 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_114
timestamp 1586364061
transform 1 0 11592 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 34272
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_124
timestamp 1586364061
transform 1 0 12512 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_128
timestamp 1586364061
transform 1 0 12880 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 13064 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_647
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 35360
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 13248 0 1 34272
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_60_141
timestamp 1586364061
transform 1 0 14076 0 -1 35360
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_60_137
timestamp 1586364061
transform 1 0 13708 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_143
timestamp 1586364061
transform 1 0 14260 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_154
timestamp 1586364061
transform 1 0 15272 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_153
timestamp 1586364061
transform 1 0 15180 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_149
timestamp 1586364061
transform 1 0 14812 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_656
timestamp 1586364061
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 34272
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_164
timestamp 1586364061
transform 1 0 16192 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_170
timestamp 1586364061
transform 1 0 16744 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_166
timestamp 1586364061
transform 1 0 16376 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_175
timestamp 1586364061
transform 1 0 17204 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_59_180
timestamp 1586364061
transform 1 0 17664 0 1 34272
box -38 -48 130 592
use scs8hd_decap_6  FILLER_59_174
timestamp 1586364061
transform 1 0 17112 0 1 34272
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17572 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_186
timestamp 1586364061
transform 1 0 18216 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_60_181
timestamp 1586364061
transform 1 0 17756 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__523__B
timestamp 1586364061
transform 1 0 18032 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__523__A
timestamp 1586364061
transform 1 0 17756 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_648
timestamp 1586364061
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use scs8hd_nor2_4  _523_
timestamp 1586364061
transform 1 0 18032 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_60_199
timestamp 1586364061
transform 1 0 19412 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_197
timestamp 1586364061
transform 1 0 19228 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_193
timestamp 1586364061
transform 1 0 18860 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18400 0 -1 35360
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_60_211
timestamp 1586364061
transform 1 0 20516 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_60_203
timestamp 1586364061
transform 1 0 19780 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_209
timestamp 1586364061
transform 1 0 20332 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_205
timestamp 1586364061
transform 1 0 19964 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_201
timestamp 1586364061
transform 1 0 19596 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20516 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_657
timestamp 1586364061
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20700 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_226
timestamp 1586364061
transform 1 0 21896 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_220
timestamp 1586364061
transform 1 0 21344 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_216
timestamp 1586364061
transform 1 0 20976 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21160 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 1 34272
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 35360
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_60_237
timestamp 1586364061
transform 1 0 22908 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_4  FILLER_60_230
timestamp 1586364061
transform 1 0 22264 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_4  FILLER_59_237
timestamp 1586364061
transform 1 0 22908 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_233
timestamp 1586364061
transform 1 0 22540 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22632 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_1  FILLER_59_241
timestamp 1586364061
transform 1 0 23276 0 1 34272
box -38 -48 130 592
use scs8hd_decap_3  FILLER_60_247
timestamp 1586364061
transform 1 0 23828 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23644 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_649
timestamp 1586364061
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 35360
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 23644 0 1 34272
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_60_259
timestamp 1586364061
transform 1 0 24932 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_59_260
timestamp 1586364061
transform 1 0 25024 0 1 34272
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_256
timestamp 1586364061
transform 1 0 24656 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_271
timestamp 1586364061
transform 1 0 26036 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_273
timestamp 1586364061
transform 1 0 26220 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_269
timestamp 1586364061
transform 1 0 25852 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26404 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_658
timestamp 1586364061
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26588 0 1 34272
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_285
timestamp 1586364061
transform 1 0 27324 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_286
timestamp 1586364061
transform 1 0 27416 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27600 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_60_293
timestamp 1586364061
transform 1 0 28060 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_290
timestamp 1586364061
transform 1 0 27784 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27968 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 34272
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28336 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__481__B
timestamp 1586364061
transform 1 0 28796 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_297
timestamp 1586364061
transform 1 0 28428 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_301
timestamp 1586364061
transform 1 0 28796 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_60_299
timestamp 1586364061
transform 1 0 28612 0 -1 35360
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_650
timestamp 1586364061
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28980 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_303
timestamp 1586364061
transform 1 0 28980 0 -1 35360
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 29348 0 -1 35360
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_60_318
timestamp 1586364061
transform 1 0 30360 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_313
timestamp 1586364061
transform 1 0 29900 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_309
timestamp 1586364061
transform 1 0 29532 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30084 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 29716 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30268 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_60_322
timestamp 1586364061
transform 1 0 30728 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30544 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_60_326
timestamp 1586364061
transform 1 0 31096 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_1  FILLER_59_330
timestamp 1586364061
transform 1 0 31464 0 1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_59_326
timestamp 1586364061
transform 1 0 31096 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30912 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31556 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_60_334
timestamp 1586364061
transform 1 0 31832 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_333
timestamp 1586364061
transform 1 0 31740 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31648 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31924 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_659
timestamp 1586364061
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 1 34272
box -38 -48 866 592
use scs8hd_decap_3  FILLER_60_346
timestamp 1586364061
transform 1 0 32936 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_346
timestamp 1586364061
transform 1 0 32936 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_60_351
timestamp 1586364061
transform 1 0 33396 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_357
timestamp 1586364061
transform 1 0 33948 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_350
timestamp 1586364061
transform 1 0 33304 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33488 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33212 0 -1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33672 0 -1 35360
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33672 0 1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_60_363
timestamp 1586364061
transform 1 0 34500 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_1  FILLER_59_365
timestamp 1586364061
transform 1 0 34684 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_361
timestamp 1586364061
transform 1 0 34316 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34500 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34132 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_651
timestamp 1586364061
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_374
timestamp 1586364061
transform 1 0 35512 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_370
timestamp 1586364061
transform 1 0 35144 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35236 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_384
timestamp 1586364061
transform 1 0 36432 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_60_380
timestamp 1586364061
transform 1 0 36064 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_386
timestamp 1586364061
transform 1 0 36616 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_382
timestamp 1586364061
transform 1 0 36248 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_378
timestamp 1586364061
transform 1 0 35880 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36064 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36432 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35696 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__422__A
timestamp 1586364061
transform 1 0 36248 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_60_398
timestamp 1586364061
transform 1 0 37720 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_395
timestamp 1586364061
transform 1 0 37444 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_392
timestamp 1586364061
transform 1 0 37168 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37260 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 36800 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_660
timestamp 1586364061
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 36984 0 1 34272
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_59_401
timestamp 1586364061
transform 1 0 37996 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37996 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_1  FILLER_60_411
timestamp 1586364061
transform 1 0 38916 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_1  FILLER_60_408
timestamp 1586364061
transform 1 0 38640 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_4  FILLER_60_404
timestamp 1586364061
transform 1 0 38272 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_405
timestamp 1586364061
transform 1 0 38364 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38732 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38548 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38180 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38732 0 1 34272
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39008 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_421
timestamp 1586364061
transform 1 0 39836 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_4  FILLER_59_422
timestamp 1586364061
transform 1 0 39928 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_418
timestamp 1586364061
transform 1 0 39560 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39744 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_426
timestamp 1586364061
transform 1 0 40296 0 1 34272
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_652
timestamp 1586364061
transform 1 0 40388 0 1 34272
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 34272
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40572 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_60_438
timestamp 1586364061
transform 1 0 41400 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_4  FILLER_60_432
timestamp 1586364061
transform 1 0 40848 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_439
timestamp 1586364061
transform 1 0 41492 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_435
timestamp 1586364061
transform 1 0 41124 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_431
timestamp 1586364061
transform 1 0 40756 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41216 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41308 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_443
timestamp 1586364061
transform 1 0 41860 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42228 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42412 0 1 34272
box -38 -48 866 592
use scs8hd_decap_4  FILLER_60_454
timestamp 1586364061
transform 1 0 42872 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_60_450
timestamp 1586364061
transform 1 0 42504 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42688 0 -1 35360
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 35360
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_661
timestamp 1586364061
transform 1 0 43240 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43424 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_458
timestamp 1586364061
transform 1 0 43240 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_462
timestamp 1586364061
transform 1 0 43608 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_474
timestamp 1586364061
transform 1 0 44712 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_462
timestamp 1586364061
transform 1 0 43608 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_474
timestamp 1586364061
transform 1 0 44712 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_653
timestamp 1586364061
transform 1 0 46000 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_486
timestamp 1586364061
transform 1 0 45816 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_489
timestamp 1586364061
transform 1 0 46092 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_501
timestamp 1586364061
transform 1 0 47196 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_486
timestamp 1586364061
transform 1 0 45816 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_498
timestamp 1586364061
transform 1 0 46920 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 48852 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 48852 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_59_513
timestamp 1586364061
transform 1 0 48300 0 1 34272
box -38 -48 314 592
use scs8hd_decap_6  FILLER_60_510
timestamp 1586364061
transform 1 0 48024 0 -1 35360
box -38 -48 590 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 4600 0 1 35360
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5888 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_30
timestamp 1586364061
transform 1 0 3864 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_34
timestamp 1586364061
transform 1 0 4232 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_49
timestamp 1586364061
transform 1 0 5612 0 1 35360
box -38 -48 314 592
use scs8hd_fill_1  FILLER_61_58
timestamp 1586364061
transform 1 0 6440 0 1 35360
box -38 -48 130 592
use scs8hd_decap_4  FILLER_61_54
timestamp 1586364061
transform 1 0 6072 0 1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_662
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 866 592
use scs8hd_decap_12  FILLER_61_79
timestamp 1586364061
transform 1 0 8372 0 1 35360
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_61_75
timestamp 1586364061
transform 1 0 8004 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_71
timestamp 1586364061
transform 1 0 7636 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_91
timestamp 1586364061
transform 1 0 9476 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_95
timestamp 1586364061
transform 1 0 9844 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_99
timestamp 1586364061
transform 1 0 10212 0 1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_61_114
timestamp 1586364061
transform 1 0 11592 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_118
timestamp 1586364061
transform 1 0 11960 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_663
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_fill_1  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_127
timestamp 1586364061
transform 1 0 12788 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_131
timestamp 1586364061
transform 1 0 13156 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_144
timestamp 1586364061
transform 1 0 14352 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_148
timestamp 1586364061
transform 1 0 14720 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_161
timestamp 1586364061
transform 1 0 15916 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_165
timestamp 1586364061
transform 1 0 16284 0 1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__620__A
timestamp 1586364061
transform 1 0 16100 0 1 35360
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 16652 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_172
timestamp 1586364061
transform 1 0 16928 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 17112 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_176
timestamp 1586364061
transform 1 0 17296 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17572 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_184
timestamp 1586364061
transform 1 0 18032 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_181
timestamp 1586364061
transform 1 0 17756 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_664
timestamp 1586364061
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use scs8hd_conb_1  _640_
timestamp 1586364061
transform 1 0 18308 0 1 35360
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19320 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_190
timestamp 1586364061
transform 1 0 18584 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_194
timestamp 1586364061
transform 1 0 18952 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_207
timestamp 1586364061
transform 1 0 20148 0 1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_61_211
timestamp 1586364061
transform 1 0 20516 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_214
timestamp 1586364061
transform 1 0 20792 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_227
timestamp 1586364061
transform 1 0 21988 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_231
timestamp 1586364061
transform 1 0 22356 0 1 35360
box -38 -48 406 592
use scs8hd_decap_4  FILLER_61_237
timestamp 1586364061
transform 1 0 22908 0 1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_61_241
timestamp 1586364061
transform 1 0 23276 0 1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_665
timestamp 1586364061
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25208 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_245
timestamp 1586364061
transform 1 0 23644 0 1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_61_260
timestamp 1586364061
transform 1 0 25024 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_264
timestamp 1586364061
transform 1 0 25392 0 1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_61_268
timestamp 1586364061
transform 1 0 25760 0 1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26404 0 1 35360
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__481__A
timestamp 1586364061
transform 1 0 27968 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26220 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25852 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27416 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_271
timestamp 1586364061
transform 1 0 26036 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_284
timestamp 1586364061
transform 1 0 27232 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_288
timestamp 1586364061
transform 1 0 27600 0 1 35360
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 29256 0 1 35360
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_666
timestamp 1586364061
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_297
timestamp 1586364061
transform 1 0 28428 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_301
timestamp 1586364061
transform 1 0 28796 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_317
timestamp 1586364061
transform 1 0 30268 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_321
timestamp 1586364061
transform 1 0 30636 0 1 35360
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31648 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__459__A
timestamp 1586364061
transform 1 0 32660 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__459__B
timestamp 1586364061
transform 1 0 31464 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33028 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31096 0 1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_61_325
timestamp 1586364061
transform 1 0 31004 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_328
timestamp 1586364061
transform 1 0 31280 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_341
timestamp 1586364061
transform 1 0 32476 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_345
timestamp 1586364061
transform 1 0 32844 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_667
timestamp 1586364061
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__420__B
timestamp 1586364061
transform 1 0 35512 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__439__A
timestamp 1586364061
transform 1 0 35052 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_358
timestamp 1586364061
transform 1 0 34040 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_362
timestamp 1586364061
transform 1 0 34408 0 1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_61_367
timestamp 1586364061
transform 1 0 34868 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_371
timestamp 1586364061
transform 1 0 35236 0 1 35360
box -38 -48 314 592
use scs8hd_nor2_4  _420_
timestamp 1586364061
transform 1 0 35696 0 1 35360
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 37260 0 1 35360
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 37076 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__422__B
timestamp 1586364061
transform 1 0 36708 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_385
timestamp 1586364061
transform 1 0 36524 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_389
timestamp 1586364061
transform 1 0 36892 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_404
timestamp 1586364061
transform 1 0 38272 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__440__A
timestamp 1586364061
transform 1 0 38456 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_408
timestamp 1586364061
transform 1 0 38640 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38824 0 1 35360
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39008 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_415
timestamp 1586364061
transform 1 0 39284 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39468 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_419
timestamp 1586364061
transform 1 0 39652 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39836 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_423
timestamp 1586364061
transform 1 0 40020 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40204 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_428
timestamp 1586364061
transform 1 0 40480 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_668
timestamp 1586364061
transform 1 0 40388 0 1 35360
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 41216 0 1 35360
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42964 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42412 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 41032 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42780 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40664 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_432
timestamp 1586364061
transform 1 0 40848 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_447
timestamp 1586364061
transform 1 0 42228 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_451
timestamp 1586364061
transform 1 0 42596 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43976 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_464
timestamp 1586364061
transform 1 0 43792 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_468
timestamp 1586364061
transform 1 0 44160 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_480
timestamp 1586364061
transform 1 0 45264 0 1 35360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_669
timestamp 1586364061
transform 1 0 46000 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_489
timestamp 1586364061
transform 1 0 46092 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_501
timestamp 1586364061
transform 1 0 47196 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 48852 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_513
timestamp 1586364061
transform 1 0 48300 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 590 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_670
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_62_40
timestamp 1586364061
transform 1 0 4784 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 -1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_4  FILLER_62_48
timestamp 1586364061
transform 1 0 5520 0 -1 36448
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_61
timestamp 1586364061
transform 1 0 6716 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_62_67
timestamp 1586364061
transform 1 0 7268 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_62_78
timestamp 1586364061
transform 1 0 8280 0 -1 36448
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_671
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_90
timestamp 1586364061
transform 1 0 9384 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_62_106
timestamp 1586364061
transform 1 0 10856 0 -1 36448
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_123
timestamp 1586364061
transform 1 0 12420 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_6  FILLER_62_129
timestamp 1586364061
transform 1 0 12972 0 -1 36448
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 -1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_672
timestamp 1586364061
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_62_137
timestamp 1586364061
transform 1 0 13708 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_141
timestamp 1586364061
transform 1 0 14076 0 -1 36448
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_62_154
timestamp 1586364061
transform 1 0 15272 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_158
timestamp 1586364061
transform 1 0 15640 0 -1 36448
box -38 -48 406 592
use scs8hd_inv_8  _620_
timestamp 1586364061
transform 1 0 16008 0 -1 36448
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17572 0 -1 36448
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_62_171
timestamp 1586364061
transform 1 0 16836 0 -1 36448
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_673
timestamp 1586364061
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_62_190
timestamp 1586364061
transform 1 0 18584 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_62_195
timestamp 1586364061
transform 1 0 19044 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_62_201
timestamp 1586364061
transform 1 0 19596 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_62_205
timestamp 1586364061
transform 1 0 19964 0 -1 36448
box -38 -48 774 592
use scs8hd_fill_1  FILLER_62_213
timestamp 1586364061
transform 1 0 20700 0 -1 36448
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22724 0 -1 36448
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_62_215
timestamp 1586364061
transform 1 0 20884 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_62_227
timestamp 1586364061
transform 1 0 21988 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_231
timestamp 1586364061
transform 1 0 22356 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_8  FILLER_62_238
timestamp 1586364061
transform 1 0 23000 0 -1 36448
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__469__B
timestamp 1586364061
transform 1 0 25116 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_246
timestamp 1586364061
transform 1 0 23736 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_259
timestamp 1586364061
transform 1 0 24932 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_62_263
timestamp 1586364061
transform 1 0 25300 0 -1 36448
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_674
timestamp 1586364061
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__463__B
timestamp 1586364061
transform 1 0 27508 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_285
timestamp 1586364061
transform 1 0 27324 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_62_289
timestamp 1586364061
transform 1 0 27692 0 -1 36448
box -38 -48 774 592
use scs8hd_nor2_4  _481_
timestamp 1586364061
transform 1 0 28612 0 -1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30360 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__452__B
timestamp 1586364061
transform 1 0 29624 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29992 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_297
timestamp 1586364061
transform 1 0 28428 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_308
timestamp 1586364061
transform 1 0 29440 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_312
timestamp 1586364061
transform 1 0 29808 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_316
timestamp 1586364061
transform 1 0 30176 0 -1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _459_
timestamp 1586364061
transform 1 0 32108 0 -1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_675
timestamp 1586364061
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__458__B
timestamp 1586364061
transform 1 0 31648 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33120 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_327
timestamp 1586364061
transform 1 0 31188 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_331
timestamp 1586364061
transform 1 0 31556 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_62_334
timestamp 1586364061
transform 1 0 31832 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_346
timestamp 1586364061
transform 1 0 32936 0 -1 36448
box -38 -48 222 592
use scs8hd_buf_1  _439_
timestamp 1586364061
transform 1 0 34684 0 -1 36448
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33672 0 -1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__447__B
timestamp 1586364061
transform 1 0 35328 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_350
timestamp 1586364061
transform 1 0 33304 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_8  FILLER_62_357
timestamp 1586364061
transform 1 0 33948 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_4  FILLER_62_368
timestamp 1586364061
transform 1 0 34960 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_62_374
timestamp 1586364061
transform 1 0 35512 0 -1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _422_
timestamp 1586364061
transform 1 0 36064 0 -1 36448
box -38 -48 866 592
use scs8hd_buf_1  _440_
timestamp 1586364061
transform 1 0 37720 0 -1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_676
timestamp 1586364061
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__420__A
timestamp 1586364061
transform 1 0 35696 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_378
timestamp 1586364061
transform 1 0 35880 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_62_389
timestamp 1586364061
transform 1 0 36892 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_8  FILLER_62_401
timestamp 1586364061
transform 1 0 37996 0 -1 36448
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40572 0 -1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39008 0 -1 36448
box -38 -48 866 592
use scs8hd_decap_3  FILLER_62_409
timestamp 1586364061
transform 1 0 38732 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_8  FILLER_62_421
timestamp 1586364061
transform 1 0 39836 0 -1 36448
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42136 0 -1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_62_438
timestamp 1586364061
transform 1 0 41400 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_6  FILLER_62_449
timestamp 1586364061
transform 1 0 42412 0 -1 36448
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_677
timestamp 1586364061
transform 1 0 43240 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_1  FILLER_62_457
timestamp 1586364061
transform 1 0 43148 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_462
timestamp 1586364061
transform 1 0 43608 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_474
timestamp 1586364061
transform 1 0 44712 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_486
timestamp 1586364061
transform 1 0 45816 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_498
timestamp 1586364061
transform 1 0 46920 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 48852 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_6  FILLER_62_510
timestamp 1586364061
transform 1 0 48024 0 -1 36448
box -38 -48 590 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5428 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  FILLER_63_52
timestamp 1586364061
transform 1 0 5888 0 1 36448
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_678
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_57
timestamp 1586364061
transform 1 0 6348 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 222 592
use scs8hd_decap_6  FILLER_63_78
timestamp 1586364061
transform 1 0 8280 0 1 36448
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_90
timestamp 1586364061
transform 1 0 9384 0 1 36448
box -38 -48 222 592
use scs8hd_decap_6  FILLER_63_103
timestamp 1586364061
transform 1 0 10580 0 1 36448
box -38 -48 590 592
use scs8hd_fill_2  FILLER_63_112
timestamp 1586364061
transform 1 0 11408 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_109
timestamp 1586364061
transform 1 0 11132 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 222 592
use scs8hd_decap_6  FILLER_63_116
timestamp 1586364061
transform 1 0 11776 0 1 36448
box -38 -48 590 592
use scs8hd_decap_4  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_679
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_63_129
timestamp 1586364061
transform 1 0 12972 0 1 36448
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13892 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 222 592
use scs8hd_decap_6  FILLER_63_148
timestamp 1586364061
transform 1 0 14720 0 1 36448
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_680
timestamp 1586364061
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__623__A
timestamp 1586364061
transform 1 0 16468 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_165
timestamp 1586364061
transform 1 0 16284 0 1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_63_169
timestamp 1586364061
transform 1 0 16652 0 1 36448
box -38 -48 774 592
use scs8hd_fill_2  FILLER_63_179
timestamp 1586364061
transform 1 0 17572 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_184
timestamp 1586364061
transform 1 0 18032 0 1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_195
timestamp 1586364061
transform 1 0 19044 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_199
timestamp 1586364061
transform 1 0 19412 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_212
timestamp 1586364061
transform 1 0 20608 0 1 36448
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21804 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_216
timestamp 1586364061
transform 1 0 20976 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_219
timestamp 1586364061
transform 1 0 21252 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_223
timestamp 1586364061
transform 1 0 21620 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_234
timestamp 1586364061
transform 1 0 22632 0 1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_63_240
timestamp 1586364061
transform 1 0 23184 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_248
timestamp 1586364061
transform 1 0 23920 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23368 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 24104 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_681
timestamp 1586364061
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_256
timestamp 1586364061
transform 1 0 24656 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_252
timestamp 1586364061
transform 1 0 24288 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__469__A
timestamp 1586364061
transform 1 0 24932 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _469_
timestamp 1586364061
transform 1 0 25116 0 1 36448
box -38 -48 866 592
use scs8hd_nor2_4  _468_
timestamp 1586364061
transform 1 0 26680 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__463__A
timestamp 1586364061
transform 1 0 26496 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__468__A
timestamp 1586364061
transform 1 0 26128 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__468__B
timestamp 1586364061
transform 1 0 27692 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_270
timestamp 1586364061
transform 1 0 25944 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_274
timestamp 1586364061
transform 1 0 26312 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_287
timestamp 1586364061
transform 1 0 27508 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_291
timestamp 1586364061
transform 1 0 27876 0 1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_63_295
timestamp 1586364061
transform 1 0 28244 0 1 36448
box -38 -48 130 592
use scs8hd_nor2_4  _470_
timestamp 1586364061
transform 1 0 29256 0 1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_682
timestamp 1586364061
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__452__A
timestamp 1586364061
transform 1 0 30268 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__470__A
timestamp 1586364061
transform 1 0 28980 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__461__A
timestamp 1586364061
transform 1 0 28336 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_298
timestamp 1586364061
transform 1 0 28520 0 1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_63_302
timestamp 1586364061
transform 1 0 28888 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_315
timestamp 1586364061
transform 1 0 30084 0 1 36448
box -38 -48 222 592
use scs8hd_decap_6  FILLER_63_319
timestamp 1586364061
transform 1 0 30452 0 1 36448
box -38 -48 590 592
use scs8hd_nor2_4  _458_
timestamp 1586364061
transform 1 0 31648 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 32844 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31004 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__458__A
timestamp 1586364061
transform 1 0 31464 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_327
timestamp 1586364061
transform 1 0 31188 0 1 36448
box -38 -48 314 592
use scs8hd_decap_4  FILLER_63_341
timestamp 1586364061
transform 1 0 32476 0 1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_63_347
timestamp 1586364061
transform 1 0 33028 0 1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _447_
timestamp 1586364061
transform 1 0 35420 0 1 36448
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33212 0 1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_683
timestamp 1586364061
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33672 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__447__A
timestamp 1586364061
transform 1 0 35236 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__448__A
timestamp 1586364061
transform 1 0 34592 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_352
timestamp 1586364061
transform 1 0 33488 0 1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_63_356
timestamp 1586364061
transform 1 0 33856 0 1 36448
box -38 -48 774 592
use scs8hd_decap_4  FILLER_63_367
timestamp 1586364061
transform 1 0 34868 0 1 36448
box -38 -48 406 592
use scs8hd_nor2_4  _441_
timestamp 1586364061
transform 1 0 36984 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__441__A
timestamp 1586364061
transform 1 0 36800 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__448__B
timestamp 1586364061
transform 1 0 36432 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_382
timestamp 1586364061
transform 1 0 36248 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_386
timestamp 1586364061
transform 1 0 36616 0 1 36448
box -38 -48 222 592
use scs8hd_decap_6  FILLER_63_399
timestamp 1586364061
transform 1 0 37812 0 1 36448
box -38 -48 590 592
use scs8hd_fill_2  FILLER_63_411
timestamp 1586364061
transform 1 0 38916 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_405
timestamp 1586364061
transform 1 0 38364 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38456 0 1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38640 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_419
timestamp 1586364061
transform 1 0 39652 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_415
timestamp 1586364061
transform 1 0 39284 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39836 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39468 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 39100 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_423
timestamp 1586364061
transform 1 0 40020 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40204 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_684
timestamp 1586364061
transform 1 0 40388 0 1 36448
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42044 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 41492 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41860 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_437
timestamp 1586364061
transform 1 0 41308 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_441
timestamp 1586364061
transform 1 0 41676 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_454
timestamp 1586364061
transform 1 0 42872 0 1 36448
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43332 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_458
timestamp 1586364061
transform 1 0 43240 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_461
timestamp 1586364061
transform 1 0 43516 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_473
timestamp 1586364061
transform 1 0 44620 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_685
timestamp 1586364061
transform 1 0 46000 0 1 36448
box -38 -48 130 592
use scs8hd_decap_3  FILLER_63_485
timestamp 1586364061
transform 1 0 45724 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_489
timestamp 1586364061
transform 1 0 46092 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_501
timestamp 1586364061
transform 1 0 47196 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 48852 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_513
timestamp 1586364061
transform 1 0 48300 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_686
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 866 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_71
timestamp 1586364061
transform 1 0 7636 0 -1 37536
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_687
timestamp 1586364061
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_83
timestamp 1586364061
transform 1 0 8740 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_3  FILLER_64_89
timestamp 1586364061
transform 1 0 9292 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_3  FILLER_64_102
timestamp 1586364061
transform 1 0 10488 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_3  FILLER_64_107
timestamp 1586364061
transform 1 0 10948 0 -1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 37536
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 37536
box -38 -48 866 592
use scs8hd_decap_8  FILLER_64_119
timestamp 1586364061
transform 1 0 12052 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_8  FILLER_64_144
timestamp 1586364061
transform 1 0 14352 0 -1 37536
box -38 -48 774 592
use scs8hd_fill_2  FILLER_64_140
timestamp 1586364061
transform 1 0 13984 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_136
timestamp 1586364061
transform 1 0 13616 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__626__A
timestamp 1586364061
transform 1 0 13800 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_1  FILLER_64_152
timestamp 1586364061
transform 1 0 15088 0 -1 37536
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_688
timestamp 1586364061
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use scs8hd_fill_1  FILLER_64_158
timestamp 1586364061
transform 1 0 15640 0 -1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_64_154
timestamp 1586364061
transform 1 0 15272 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 37536
box -38 -48 222 592
use scs8hd_inv_8  _623_
timestamp 1586364061
transform 1 0 15732 0 -1 37536
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17848 0 -1 37536
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_64_168
timestamp 1586364061
transform 1 0 16560 0 -1 37536
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_64_180
timestamp 1586364061
transform 1 0 17664 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_185
timestamp 1586364061
transform 1 0 18124 0 -1 37536
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_689
timestamp 1586364061
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_189
timestamp 1586364061
transform 1 0 18492 0 -1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_64_202
timestamp 1586364061
transform 1 0 19688 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_206
timestamp 1586364061
transform 1 0 20056 0 -1 37536
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23000 0 -1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22724 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_215
timestamp 1586364061
transform 1 0 20884 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_4  FILLER_64_230
timestamp 1586364061
transform 1 0 22264 0 -1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_64_234
timestamp 1586364061
transform 1 0 22632 0 -1 37536
box -38 -48 130 592
use scs8hd_fill_1  FILLER_64_237
timestamp 1586364061
transform 1 0 22908 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_8  FILLER_64_241
timestamp 1586364061
transform 1 0 23276 0 -1 37536
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 24104 0 -1 37536
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_64_249
timestamp 1586364061
transform 1 0 24012 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_261
timestamp 1586364061
transform 1 0 25116 0 -1 37536
box -38 -48 1142 592
use scs8hd_nor2_4  _463_
timestamp 1586364061
transform 1 0 26772 0 -1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_690
timestamp 1586364061
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_64_273
timestamp 1586364061
transform 1 0 26220 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_64_276
timestamp 1586364061
transform 1 0 26496 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_8  FILLER_64_288
timestamp 1586364061
transform 1 0 27600 0 -1 37536
box -38 -48 774 592
use scs8hd_nor2_4  _452_
timestamp 1586364061
transform 1 0 29440 0 -1 37536
box -38 -48 866 592
use scs8hd_buf_1  _461_
timestamp 1586364061
transform 1 0 28336 0 -1 37536
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__470__B
timestamp 1586364061
transform 1 0 29256 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_6  FILLER_64_299
timestamp 1586364061
transform 1 0 28612 0 -1 37536
box -38 -48 590 592
use scs8hd_fill_1  FILLER_64_305
timestamp 1586364061
transform 1 0 29164 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_8  FILLER_64_317
timestamp 1586364061
transform 1 0 30268 0 -1 37536
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 32844 0 -1 37536
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_691
timestamp 1586364061
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32476 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_328
timestamp 1586364061
transform 1 0 31280 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_4  FILLER_64_337
timestamp 1586364061
transform 1 0 32108 0 -1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_64_343
timestamp 1586364061
transform 1 0 32660 0 -1 37536
box -38 -48 222 592
use scs8hd_nor2_4  _448_
timestamp 1586364061
transform 1 0 35420 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_356
timestamp 1586364061
transform 1 0 33856 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  FILLER_64_364
timestamp 1586364061
transform 1 0 34592 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_4  FILLER_64_369
timestamp 1586364061
transform 1 0 35052 0 -1 37536
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_692
timestamp 1586364061
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__441__B
timestamp 1586364061
transform 1 0 36984 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37904 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37352 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_382
timestamp 1586364061
transform 1 0 36248 0 -1 37536
box -38 -48 774 592
use scs8hd_fill_2  FILLER_64_392
timestamp 1586364061
transform 1 0 37168 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_1  FILLER_64_396
timestamp 1586364061
transform 1 0 37536 0 -1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_64_398
timestamp 1586364061
transform 1 0 37720 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_6  FILLER_64_402
timestamp 1586364061
transform 1 0 38088 0 -1 37536
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 38640 0 -1 37536
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40480 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_419
timestamp 1586364061
transform 1 0 39652 0 -1 37536
box -38 -48 774 592
use scs8hd_fill_1  FILLER_64_427
timestamp 1586364061
transform 1 0 40388 0 -1 37536
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 40756 0 -1 37536
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41952 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42320 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_1  FILLER_64_430
timestamp 1586364061
transform 1 0 40664 0 -1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_64_442
timestamp 1586364061
transform 1 0 41768 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_446
timestamp 1586364061
transform 1 0 42136 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_450
timestamp 1586364061
transform 1 0 42504 0 -1 37536
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_693
timestamp 1586364061
transform 1 0 43240 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_462
timestamp 1586364061
transform 1 0 43608 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_474
timestamp 1586364061
transform 1 0 44712 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_486
timestamp 1586364061
transform 1 0 45816 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_498
timestamp 1586364061
transform 1 0 46920 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 48852 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_6  FILLER_64_510
timestamp 1586364061
transform 1 0 48024 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_3  PHY_130
timestamp 1586364061
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_65_3
timestamp 1586364061
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_15
timestamp 1586364061
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_27
timestamp 1586364061
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_39
timestamp 1586364061
transform 1 0 4692 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_65_51
timestamp 1586364061
transform 1 0 5796 0 1 37536
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_694
timestamp 1586364061
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_59
timestamp 1586364061
transform 1 0 6532 0 1 37536
box -38 -48 222 592
use scs8hd_decap_6  FILLER_65_62
timestamp 1586364061
transform 1 0 6808 0 1 37536
box -38 -48 590 592
use scs8hd_decap_6  FILLER_65_79
timestamp 1586364061
transform 1 0 8372 0 1 37536
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 37536
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_96
timestamp 1586364061
transform 1 0 9936 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_65_100
timestamp 1586364061
transform 1 0 10304 0 1 37536
box -38 -48 314 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 12420 0 1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_695
timestamp 1586364061
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 12880 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__625__A
timestamp 1586364061
transform 1 0 11776 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_114
timestamp 1586364061
transform 1 0 11592 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_118
timestamp 1586364061
transform 1 0 11960 0 1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_65_126
timestamp 1586364061
transform 1 0 12696 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_130
timestamp 1586364061
transform 1 0 13064 0 1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_65_134
timestamp 1586364061
transform 1 0 13432 0 1 37536
box -38 -48 130 592
use scs8hd_inv_8  _622_
timestamp 1586364061
transform 1 0 15272 0 1 37536
box -38 -48 866 592
use scs8hd_inv_8  _626_
timestamp 1586364061
transform 1 0 13708 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__622__A
timestamp 1586364061
transform 1 0 14720 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_146
timestamp 1586364061
transform 1 0 14536 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_150
timestamp 1586364061
transform 1 0 14904 0 1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_65_163
timestamp 1586364061
transform 1 0 16100 0 1 37536
box -38 -48 774 592
use scs8hd_fill_2  FILLER_65_178
timestamp 1586364061
transform 1 0 17480 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_174
timestamp 1586364061
transform 1 0 17112 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 17296 0 1 37536
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 16836 0 1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_65_187
timestamp 1586364061
transform 1 0 18308 0 1 37536
box -38 -48 222 592
use scs8hd_fill_1  FILLER_65_182
timestamp 1586364061
transform 1 0 17848 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17664 0 1 37536
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_696
timestamp 1586364061
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19412 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_191
timestamp 1586364061
transform 1 0 18676 0 1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_65_197
timestamp 1586364061
transform 1 0 19228 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_65_208
timestamp 1586364061
transform 1 0 20240 0 1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_65_213
timestamp 1586364061
transform 1 0 20700 0 1 37536
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_65_217
timestamp 1586364061
transform 1 0 21068 0 1 37536
box -38 -48 314 592
use scs8hd_decap_4  FILLER_65_231
timestamp 1586364061
transform 1 0 22356 0 1 37536
box -38 -48 406 592
use scs8hd_decap_4  FILLER_65_237
timestamp 1586364061
transform 1 0 22908 0 1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_65_241
timestamp 1586364061
transform 1 0 23276 0 1 37536
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 24196 0 1 37536
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_697
timestamp 1586364061
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 24012 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25392 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_245
timestamp 1586364061
transform 1 0 23644 0 1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_65_262
timestamp 1586364061
transform 1 0 25208 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_266
timestamp 1586364061
transform 1 0 25576 0 1 37536
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 26496 0 1 37536
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 26312 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25944 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27692 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_272
timestamp 1586364061
transform 1 0 26128 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_287
timestamp 1586364061
transform 1 0 27508 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_291
timestamp 1586364061
transform 1 0 27876 0 1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_65_295
timestamp 1586364061
transform 1 0 28244 0 1 37536
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 30084 0 1 37536
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_698
timestamp 1586364061
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 29900 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__455__A
timestamp 1586364061
transform 1 0 28980 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__455__B
timestamp 1586364061
transform 1 0 29440 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_306
timestamp 1586364061
transform 1 0 29256 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_65_310
timestamp 1586364061
transform 1 0 29624 0 1 37536
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 32476 0 1 37536
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 32292 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__462__A
timestamp 1586364061
transform 1 0 31280 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_326
timestamp 1586364061
transform 1 0 31096 0 1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_65_330
timestamp 1586364061
transform 1 0 31464 0 1 37536
box -38 -48 774 592
use scs8hd_fill_1  FILLER_65_338
timestamp 1586364061
transform 1 0 32200 0 1 37536
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_699
timestamp 1586364061
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33672 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34040 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_352
timestamp 1586364061
transform 1 0 33488 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_356
timestamp 1586364061
transform 1 0 33856 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_360
timestamp 1586364061
transform 1 0 34224 0 1 37536
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 37168 0 1 37536
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 36984 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__446__A
timestamp 1586364061
transform 1 0 36064 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__446__B
timestamp 1586364061
transform 1 0 36432 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_376
timestamp 1586364061
transform 1 0 35696 0 1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_65_382
timestamp 1586364061
transform 1 0 36248 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_386
timestamp 1586364061
transform 1 0 36616 0 1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_65_407
timestamp 1586364061
transform 1 0 38548 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_403
timestamp 1586364061
transform 1 0 38180 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 38364 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38732 0 1 37536
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38916 0 1 37536
box -38 -48 314 592
use scs8hd_decap_3  FILLER_65_414
timestamp 1586364061
transform 1 0 39192 0 1 37536
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 39468 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_419
timestamp 1586364061
transform 1 0 39652 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39836 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_423
timestamp 1586364061
transform 1 0 40020 0 1 37536
box -38 -48 406 592
use scs8hd_decap_3  FILLER_65_428
timestamp 1586364061
transform 1 0 40480 0 1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_700
timestamp 1586364061
transform 1 0 40388 0 1 37536
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40756 0 1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41768 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41216 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41584 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_434
timestamp 1586364061
transform 1 0 41032 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_438
timestamp 1586364061
transform 1 0 41400 0 1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_65_451
timestamp 1586364061
transform 1 0 42596 0 1 37536
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 1 37536
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43792 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44160 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_462
timestamp 1586364061
transform 1 0 43608 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_466
timestamp 1586364061
transform 1 0 43976 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_470
timestamp 1586364061
transform 1 0 44344 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_65_482
timestamp 1586364061
transform 1 0 45448 0 1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_701
timestamp 1586364061
transform 1 0 46000 0 1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_65_489
timestamp 1586364061
transform 1 0 46092 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_501
timestamp 1586364061
transform 1 0 47196 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_3  PHY_131
timestamp 1586364061
transform -1 0 48852 0 1 37536
box -38 -48 314 592
use scs8hd_decap_3  FILLER_65_513
timestamp 1586364061
transform 1 0 48300 0 1 37536
box -38 -48 314 592
use scs8hd_decap_3  PHY_132
timestamp 1586364061
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_134
timestamp 1586364061
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_66_3
timestamp 1586364061
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_15
timestamp 1586364061
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_3
timestamp 1586364061
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_15
timestamp 1586364061
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_702
timestamp 1586364061
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_27
timestamp 1586364061
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use scs8hd_decap_12  FILLER_66_32
timestamp 1586364061
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_44
timestamp 1586364061
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_27
timestamp 1586364061
transform 1 0 3588 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_39
timestamp 1586364061
transform 1 0 4692 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_67_51
timestamp 1586364061
transform 1 0 5796 0 1 38624
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_710
timestamp 1586364061
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_66_56
timestamp 1586364061
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_66_68
timestamp 1586364061
transform 1 0 7360 0 -1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_66_72
timestamp 1586364061
transform 1 0 7728 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_67_59
timestamp 1586364061
transform 1 0 6532 0 1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_67_62
timestamp 1586364061
transform 1 0 6808 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_74
timestamp 1586364061
transform 1 0 7912 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_86
timestamp 1586364061
transform 1 0 9016 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_66_84
timestamp 1586364061
transform 1 0 8832 0 -1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_703
timestamp 1586364061
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_1  FILLER_67_102
timestamp 1586364061
transform 1 0 10488 0 1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_67_98
timestamp 1586364061
transform 1 0 10120 0 1 38624
box -38 -48 406 592
use scs8hd_decap_3  FILLER_66_102
timestamp 1586364061
transform 1 0 10488 0 -1 38624
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 38624
box -38 -48 866 592
use scs8hd_decap_3  FILLER_66_107
timestamp 1586364061
transform 1 0 10948 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_4  FILLER_67_118
timestamp 1586364061
transform 1 0 11960 0 1 38624
box -38 -48 406 592
use scs8hd_fill_2  FILLER_67_114
timestamp 1586364061
transform 1 0 11592 0 1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_66_119
timestamp 1586364061
transform 1 0 12052 0 -1 38624
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__624__A
timestamp 1586364061
transform 1 0 11776 0 1 38624
box -38 -48 222 592
use scs8hd_inv_8  _625_
timestamp 1586364061
transform 1 0 11224 0 -1 38624
box -38 -48 866 592
use scs8hd_decap_4  FILLER_67_130
timestamp 1586364061
transform 1 0 13064 0 1 38624
box -38 -48 406 592
use scs8hd_fill_2  FILLER_67_126
timestamp 1586364061
transform 1 0 12696 0 1 38624
box -38 -48 222 592
use scs8hd_decap_4  FILLER_66_131
timestamp 1586364061
transform 1 0 13156 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_711
timestamp 1586364061
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 38624
box -38 -48 314 592
use scs8hd_fill_1  FILLER_67_134
timestamp 1586364061
transform 1 0 13432 0 1 38624
box -38 -48 130 592
use scs8hd_fill_1  FILLER_66_135
timestamp 1586364061
transform 1 0 13524 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__627__A
timestamp 1586364061
transform 1 0 13524 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 38624
box -38 -48 866 592
use scs8hd_inv_8  _627_
timestamp 1586364061
transform 1 0 13708 0 1 38624
box -38 -48 866 592
use scs8hd_decap_4  FILLER_67_150
timestamp 1586364061
transform 1 0 14904 0 1 38624
box -38 -48 406 592
use scs8hd_fill_2  FILLER_67_146
timestamp 1586364061
transform 1 0 14536 0 1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_145
timestamp 1586364061
transform 1 0 14444 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 14720 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_704
timestamp 1586364061
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_67_161
timestamp 1586364061
transform 1 0 15916 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_157
timestamp 1586364061
transform 1 0 15548 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15732 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 38624
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 1 38624
box -38 -48 314 592
use scs8hd_decap_8  FILLER_67_172
timestamp 1586364061
transform 1 0 16928 0 1 38624
box -38 -48 774 592
use scs8hd_fill_2  FILLER_67_168
timestamp 1586364061
transform 1 0 16560 0 1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_163
timestamp 1586364061
transform 1 0 16100 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16100 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 38624
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 38624
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 1 38624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_67_184
timestamp 1586364061
transform 1 0 18032 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_67_180
timestamp 1586364061
transform 1 0 17664 0 1 38624
box -38 -48 314 592
use scs8hd_decap_8  FILLER_66_186
timestamp 1586364061
transform 1 0 18216 0 -1 38624
box -38 -48 774 592
use scs8hd_decap_12  FILLER_66_174
timestamp 1586364061
transform 1 0 17112 0 -1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_712
timestamp 1586364061
transform 1 0 17940 0 1 38624
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 38624
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 -1 38624
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_705
timestamp 1586364061
transform 1 0 20792 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_194
timestamp 1586364061
transform 1 0 18952 0 -1 38624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_66_198
timestamp 1586364061
transform 1 0 19320 0 -1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_66_202
timestamp 1586364061
transform 1 0 19688 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_196
timestamp 1586364061
transform 1 0 19136 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_67_208
timestamp 1586364061
transform 1 0 20240 0 1 38624
box -38 -48 406 592
use scs8hd_fill_2  FILLER_67_219
timestamp 1586364061
transform 1 0 21252 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_215
timestamp 1586364061
transform 1 0 20884 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_224
timestamp 1586364061
transform 1 0 21712 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21436 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 38624
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21620 0 1 38624
box -38 -48 314 592
use scs8hd_decap_4  FILLER_67_234
timestamp 1586364061
transform 1 0 22632 0 1 38624
box -38 -48 406 592
use scs8hd_fill_2  FILLER_67_230
timestamp 1586364061
transform 1 0 22264 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_226
timestamp 1586364061
transform 1 0 21896 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_234
timestamp 1586364061
transform 1 0 22632 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_6  FILLER_66_228
timestamp 1586364061
transform 1 0 22080 0 -1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 22080 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_240
timestamp 1586364061
transform 1 0 23184 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22724 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_66_248
timestamp 1586364061
transform 1 0 23920 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_244
timestamp 1586364061
transform 1 0 23552 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23736 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_713
timestamp 1586364061
transform 1 0 23552 0 1 38624
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 38624
box -38 -48 866 592
use scs8hd_decap_3  FILLER_67_258
timestamp 1586364061
transform 1 0 24840 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_254
timestamp 1586364061
transform 1 0 24472 0 1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_66_261
timestamp 1586364061
transform 1 0 25116 0 -1 38624
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_1  FILLER_67_263
timestamp 1586364061
transform 1 0 25300 0 1 38624
box -38 -48 130 592
use scs8hd_decap_6  FILLER_66_266
timestamp 1586364061
transform 1 0 25576 0 -1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25392 0 -1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25392 0 1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_278
timestamp 1586364061
transform 1 0 26680 0 1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_67_273
timestamp 1586364061
transform 1 0 26220 0 1 38624
box -38 -48 314 592
use scs8hd_fill_1  FILLER_66_272
timestamp 1586364061
transform 1 0 26128 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26864 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_706
timestamp 1586364061
transform 1 0 26404 0 -1 38624
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_282
timestamp 1586364061
transform 1 0 27048 0 1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_285
timestamp 1586364061
transform 1 0 27324 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 27232 0 1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 27416 0 1 38624
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_66_295
timestamp 1586364061
transform 1 0 28244 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__466__B
timestamp 1586364061
transform 1 0 28060 0 -1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_67_306
timestamp 1586364061
transform 1 0 29256 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_301
timestamp 1586364061
transform 1 0 28796 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_297
timestamp 1586364061
transform 1 0 28428 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28980 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__466__A
timestamp 1586364061
transform 1 0 28612 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_714
timestamp 1586364061
transform 1 0 29164 0 1 38624
box -38 -48 130 592
use scs8hd_nor2_4  _455_
timestamp 1586364061
transform 1 0 28980 0 -1 38624
box -38 -48 866 592
use scs8hd_decap_3  FILLER_66_317
timestamp 1586364061
transform 1 0 30268 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  FILLER_66_312
timestamp 1586364061
transform 1 0 29808 0 -1 38624
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30084 0 -1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 29532 0 1 38624
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_67_320
timestamp 1586364061
transform 1 0 30544 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30728 0 1 38624
box -38 -48 222 592
use scs8hd_buf_1  _462_
timestamp 1586364061
transform 1 0 30544 0 -1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_324
timestamp 1586364061
transform 1 0 30912 0 1 38624
box -38 -48 222 592
use scs8hd_decap_6  FILLER_66_330
timestamp 1586364061
transform 1 0 31464 0 -1 38624
box -38 -48 590 592
use scs8hd_fill_1  FILLER_66_327
timestamp 1586364061
transform 1 0 31188 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_323
timestamp 1586364061
transform 1 0 30820 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31280 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31096 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31280 0 1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_341
timestamp 1586364061
transform 1 0 32476 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_337
timestamp 1586364061
transform 1 0 32108 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_341
timestamp 1586364061
transform 1 0 32476 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_337
timestamp 1586364061
transform 1 0 32108 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 32292 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_707
timestamp 1586364061
transform 1 0 32016 0 -1 38624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_67_345
timestamp 1586364061
transform 1 0 32844 0 1 38624
box -38 -48 222 592
use scs8hd_decap_4  FILLER_66_345
timestamp 1586364061
transform 1 0 32844 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32660 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33028 0 1 38624
box -38 -48 222 592
use scs8hd_conb_1  _646_
timestamp 1586364061
transform 1 0 32568 0 -1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_358
timestamp 1586364061
transform 1 0 34040 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_351
timestamp 1586364061
transform 1 0 33396 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 -1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 38624
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33580 0 -1 38624
box -38 -48 866 592
use scs8hd_decap_3  FILLER_67_367
timestamp 1586364061
transform 1 0 34868 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_362
timestamp 1586364061
transform 1 0 34408 0 1 38624
box -38 -48 222 592
use scs8hd_decap_4  FILLER_66_366
timestamp 1586364061
transform 1 0 34776 0 -1 38624
box -38 -48 406 592
use scs8hd_fill_2  FILLER_66_362
timestamp 1586364061
transform 1 0 34408 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__444__B
timestamp 1586364061
transform 1 0 34592 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_715
timestamp 1586364061
transform 1 0 34776 0 1 38624
box -38 -48 130 592
use scs8hd_decap_6  FILLER_66_372
timestamp 1586364061
transform 1 0 35328 0 -1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__444__A
timestamp 1586364061
transform 1 0 35144 0 -1 38624
box -38 -48 222 592
use scs8hd_nor2_4  _444_
timestamp 1586364061
transform 1 0 35144 0 1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_383
timestamp 1586364061
transform 1 0 36340 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_379
timestamp 1586364061
transform 1 0 35972 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__442__B
timestamp 1586364061
transform 1 0 35880 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__442__A
timestamp 1586364061
transform 1 0 36156 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 36524 0 1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 36708 0 1 38624
box -38 -48 1050 592
use scs8hd_nor2_4  _446_
timestamp 1586364061
transform 1 0 36064 0 -1 38624
box -38 -48 866 592
use scs8hd_decap_4  FILLER_67_398
timestamp 1586364061
transform 1 0 37720 0 1 38624
box -38 -48 406 592
use scs8hd_decap_4  FILLER_66_393
timestamp 1586364061
transform 1 0 37260 0 -1 38624
box -38 -48 406 592
use scs8hd_fill_2  FILLER_66_389
timestamp 1586364061
transform 1 0 36892 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37076 0 -1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_708
timestamp 1586364061
transform 1 0 37628 0 -1 38624
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 38624
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38088 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_404
timestamp 1586364061
transform 1 0 38272 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_413
timestamp 1586364061
transform 1 0 39100 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_409
timestamp 1586364061
transform 1 0 38732 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38916 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38456 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38640 0 1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_425
timestamp 1586364061
transform 1 0 40204 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_421
timestamp 1586364061
transform 1 0 39836 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_417
timestamp 1586364061
transform 1 0 39468 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39284 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39652 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40020 0 1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 39468 0 -1 38624
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_67_428
timestamp 1586364061
transform 1 0 40480 0 1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_428
timestamp 1586364061
transform 1 0 40480 0 -1 38624
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_716
timestamp 1586364061
transform 1 0 40388 0 1 38624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_67_437
timestamp 1586364061
transform 1 0 41308 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_433
timestamp 1586364061
transform 1 0 40940 0 1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_66_436
timestamp 1586364061
transform 1 0 41216 0 -1 38624
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41492 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41124 0 1 38624
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40664 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_66_448
timestamp 1586364061
transform 1 0 42320 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_444
timestamp 1586364061
transform 1 0 41952 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42136 0 -1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 1 38624
box -38 -48 866 592
use scs8hd_conb_1  _647_
timestamp 1586364061
transform 1 0 41676 0 -1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_454
timestamp 1586364061
transform 1 0 42872 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_450
timestamp 1586364061
transform 1 0 42504 0 1 38624
box -38 -48 222 592
use scs8hd_decap_6  FILLER_66_452
timestamp 1586364061
transform 1 0 42688 0 -1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42504 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42688 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43056 0 1 38624
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 38624
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43240 0 1 38624
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_709
timestamp 1586364061
transform 1 0 43240 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44252 0 1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_66_462
timestamp 1586364061
transform 1 0 43608 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_474
timestamp 1586364061
transform 1 0 44712 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_67_467
timestamp 1586364061
transform 1 0 44068 0 1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_67_471
timestamp 1586364061
transform 1 0 44436 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_67_483
timestamp 1586364061
transform 1 0 45540 0 1 38624
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_717
timestamp 1586364061
transform 1 0 46000 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_486
timestamp 1586364061
transform 1 0 45816 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_498
timestamp 1586364061
transform 1 0 46920 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_67_487
timestamp 1586364061
transform 1 0 45908 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_67_489
timestamp 1586364061
transform 1 0 46092 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_501
timestamp 1586364061
transform 1 0 47196 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_3  PHY_133
timestamp 1586364061
transform -1 0 48852 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_135
timestamp 1586364061
transform -1 0 48852 0 1 38624
box -38 -48 314 592
use scs8hd_decap_6  FILLER_66_510
timestamp 1586364061
transform 1 0 48024 0 -1 38624
box -38 -48 590 592
use scs8hd_decap_3  FILLER_67_513
timestamp 1586364061
transform 1 0 48300 0 1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_136
timestamp 1586364061
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_68_3
timestamp 1586364061
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_15
timestamp 1586364061
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_718
timestamp 1586364061
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_68_27
timestamp 1586364061
transform 1 0 3588 0 -1 39712
box -38 -48 406 592
use scs8hd_decap_12  FILLER_68_32
timestamp 1586364061
transform 1 0 4048 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_44
timestamp 1586364061
transform 1 0 5152 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_56
timestamp 1586364061
transform 1 0 6256 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_68
timestamp 1586364061
transform 1 0 7360 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_80
timestamp 1586364061
transform 1 0 8464 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_719
timestamp 1586364061
transform 1 0 9568 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_93
timestamp 1586364061
transform 1 0 9660 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_68_105
timestamp 1586364061
transform 1 0 10764 0 -1 39712
box -38 -48 774 592
use scs8hd_inv_8  _624_
timestamp 1586364061
transform 1 0 11592 0 -1 39712
box -38 -48 866 592
use scs8hd_fill_1  FILLER_68_113
timestamp 1586364061
transform 1 0 11500 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_123
timestamp 1586364061
transform 1 0 12420 0 -1 39712
box -38 -48 1142 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 13984 0 -1 39712
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 39712
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_720
timestamp 1586364061
transform 1 0 15180 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_68_135
timestamp 1586364061
transform 1 0 13524 0 -1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_68_139
timestamp 1586364061
transform 1 0 13892 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_8  FILLER_68_143
timestamp 1586364061
transform 1 0 14260 0 -1 39712
box -38 -48 774 592
use scs8hd_fill_2  FILLER_68_151
timestamp 1586364061
transform 1 0 14996 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_68_157
timestamp 1586364061
transform 1 0 15548 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_169
timestamp 1586364061
transform 1 0 16652 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_181
timestamp 1586364061
transform 1 0 17756 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_721
timestamp 1586364061
transform 1 0 20792 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_193
timestamp 1586364061
transform 1 0 18860 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_68_205
timestamp 1586364061
transform 1 0 19964 0 -1 39712
box -38 -48 774 592
use scs8hd_fill_1  FILLER_68_213
timestamp 1586364061
transform 1 0 20700 0 -1 39712
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 21804 0 -1 39712
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_68_215
timestamp 1586364061
transform 1 0 20884 0 -1 39712
box -38 -48 774 592
use scs8hd_fill_2  FILLER_68_223
timestamp 1586364061
transform 1 0 21620 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_236
timestamp 1586364061
transform 1 0 22816 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_68_240
timestamp 1586364061
transform 1 0 23184 0 -1 39712
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25116 0 -1 39712
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23552 0 -1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25576 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_68_253
timestamp 1586364061
transform 1 0 24380 0 -1 39712
box -38 -48 774 592
use scs8hd_fill_2  FILLER_68_264
timestamp 1586364061
transform 1 0 25392 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_68_268
timestamp 1586364061
transform 1 0 25760 0 -1 39712
box -38 -48 590 592
use scs8hd_nor2_4  _466_
timestamp 1586364061
transform 1 0 28060 0 -1 39712
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 39712
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_722
timestamp 1586364061
transform 1 0 26404 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__465__B
timestamp 1586364061
transform 1 0 27508 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_68_274
timestamp 1586364061
transform 1 0 26312 0 -1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_68_285
timestamp 1586364061
transform 1 0 27324 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_68_289
timestamp 1586364061
transform 1 0 27692 0 -1 39712
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 29532 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29992 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_68_302
timestamp 1586364061
transform 1 0 28888 0 -1 39712
box -38 -48 590 592
use scs8hd_fill_1  FILLER_68_308
timestamp 1586364061
transform 1 0 29440 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_3  FILLER_68_311
timestamp 1586364061
transform 1 0 29716 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_3  FILLER_68_316
timestamp 1586364061
transform 1 0 30176 0 -1 39712
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 39712
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_723
timestamp 1586364061
transform 1 0 32016 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31464 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_328
timestamp 1586364061
transform 1 0 31280 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_68_332
timestamp 1586364061
transform 1 0 31648 0 -1 39712
box -38 -48 406 592
use scs8hd_fill_2  FILLER_68_348
timestamp 1586364061
transform 1 0 33120 0 -1 39712
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__443__A
timestamp 1586364061
transform 1 0 35236 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33672 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_352
timestamp 1586364061
transform 1 0 33488 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_68_365
timestamp 1586364061
transform 1 0 34684 0 -1 39712
box -38 -48 590 592
use scs8hd_decap_3  FILLER_68_373
timestamp 1586364061
transform 1 0 35420 0 -1 39712
box -38 -48 314 592
use scs8hd_nor2_4  _442_
timestamp 1586364061
transform 1 0 35880 0 -1 39712
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_724
timestamp 1586364061
transform 1 0 37628 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__445__B
timestamp 1586364061
transform 1 0 35696 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36892 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_387
timestamp 1586364061
transform 1 0 36708 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_68_391
timestamp 1586364061
transform 1 0 37076 0 -1 39712
box -38 -48 590 592
use scs8hd_decap_8  FILLER_68_398
timestamp 1586364061
transform 1 0 37720 0 -1 39712
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40020 0 -1 39712
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38456 0 -1 39712
box -38 -48 866 592
use scs8hd_decap_8  FILLER_68_415
timestamp 1586364061
transform 1 0 39284 0 -1 39712
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_68_432
timestamp 1586364061
transform 1 0 40848 0 -1 39712
box -38 -48 590 592
use scs8hd_fill_1  FILLER_68_438
timestamp 1586364061
transform 1 0 41400 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_8  FILLER_68_450
timestamp 1586364061
transform 1 0 42504 0 -1 39712
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 39712
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_725
timestamp 1586364061
transform 1 0 43240 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_462
timestamp 1586364061
transform 1 0 43608 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_474
timestamp 1586364061
transform 1 0 44712 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_486
timestamp 1586364061
transform 1 0 45816 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_498
timestamp 1586364061
transform 1 0 46920 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_137
timestamp 1586364061
transform -1 0 48852 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_6  FILLER_68_510
timestamp 1586364061
transform 1 0 48024 0 -1 39712
box -38 -48 590 592
use scs8hd_decap_3  PHY_138
timestamp 1586364061
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_69_3
timestamp 1586364061
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_15
timestamp 1586364061
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_27
timestamp 1586364061
transform 1 0 3588 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_39
timestamp 1586364061
transform 1 0 4692 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_69_51
timestamp 1586364061
transform 1 0 5796 0 1 39712
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_726
timestamp 1586364061
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_59
timestamp 1586364061
transform 1 0 6532 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_62
timestamp 1586364061
transform 1 0 6808 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_74
timestamp 1586364061
transform 1 0 7912 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_86
timestamp 1586364061
transform 1 0 9016 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_98
timestamp 1586364061
transform 1 0 10120 0 1 39712
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 39712
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_727
timestamp 1586364061
transform 1 0 12328 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_110
timestamp 1586364061
transform 1 0 11224 0 1 39712
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_69_126
timestamp 1586364061
transform 1 0 12696 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_130
timestamp 1586364061
transform 1 0 13064 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_142
timestamp 1586364061
transform 1 0 14168 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_154
timestamp 1586364061
transform 1 0 15272 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_728
timestamp 1586364061
transform 1 0 17940 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_166
timestamp 1586364061
transform 1 0 16376 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_69_178
timestamp 1586364061
transform 1 0 17480 0 1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_69_182
timestamp 1586364061
transform 1 0 17848 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_184
timestamp 1586364061
transform 1 0 18032 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_196
timestamp 1586364061
transform 1 0 19136 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_69_208
timestamp 1586364061
transform 1 0 20240 0 1 39712
box -38 -48 774 592
use scs8hd_decap_3  FILLER_69_216
timestamp 1586364061
transform 1 0 20976 0 1 39712
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21252 0 1 39712
box -38 -48 314 592
use scs8hd_fill_2  FILLER_69_222
timestamp 1586364061
transform 1 0 21528 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21712 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_226
timestamp 1586364061
transform 1 0 21896 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22080 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_233
timestamp 1586364061
transform 1 0 22540 0 1 39712
box -38 -48 222 592
use scs8hd_conb_1  _645_
timestamp 1586364061
transform 1 0 22264 0 1 39712
box -38 -48 314 592
use scs8hd_decap_4  FILLER_69_237
timestamp 1586364061
transform 1 0 22908 0 1 39712
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22724 0 1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_69_241
timestamp 1586364061
transform 1 0 23276 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_248
timestamp 1586364061
transform 1 0 23920 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 39712
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_729
timestamp 1586364061
transform 1 0 23552 0 1 39712
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 39712
box -38 -48 314 592
use scs8hd_fill_2  FILLER_69_260
timestamp 1586364061
transform 1 0 25024 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_256
timestamp 1586364061
transform 1 0 24656 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_252
timestamp 1586364061
transform 1 0 24288 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25208 0 1 39712
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25392 0 1 39712
box -38 -48 866 592
use scs8hd_nor2_4  _465_
timestamp 1586364061
transform 1 0 27232 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__464__A
timestamp 1586364061
transform 1 0 27048 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__465__A
timestamp 1586364061
transform 1 0 26680 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__464__B
timestamp 1586364061
transform 1 0 28244 0 1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_69_273
timestamp 1586364061
transform 1 0 26220 0 1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_69_277
timestamp 1586364061
transform 1 0 26588 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_280
timestamp 1586364061
transform 1 0 26864 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_293
timestamp 1586364061
transform 1 0 28060 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_301
timestamp 1586364061
transform 1 0 28796 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_297
timestamp 1586364061
transform 1 0 28428 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__450__A
timestamp 1586364061
transform 1 0 28612 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__453__A
timestamp 1586364061
transform 1 0 28980 0 1 39712
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_730
timestamp 1586364061
transform 1 0 29164 0 1 39712
box -38 -48 130 592
use scs8hd_nor2_4  _453_
timestamp 1586364061
transform 1 0 29256 0 1 39712
box -38 -48 866 592
use scs8hd_fill_2  FILLER_69_319
timestamp 1586364061
transform 1 0 30452 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_315
timestamp 1586364061
transform 1 0 30084 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__457__A
timestamp 1586364061
transform 1 0 30636 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 39712
box -38 -48 222 592
use scs8hd_nor2_4  _457_
timestamp 1586364061
transform 1 0 30820 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__451__A
timestamp 1586364061
transform 1 0 32108 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33028 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32660 0 1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_69_332
timestamp 1586364061
transform 1 0 31648 0 1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_69_336
timestamp 1586364061
transform 1 0 32016 0 1 39712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_69_339
timestamp 1586364061
transform 1 0 32292 0 1 39712
box -38 -48 406 592
use scs8hd_fill_2  FILLER_69_345
timestamp 1586364061
transform 1 0 32844 0 1 39712
box -38 -48 222 592
use scs8hd_nor2_4  _443_
timestamp 1586364061
transform 1 0 35236 0 1 39712
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 39712
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_731
timestamp 1586364061
transform 1 0 34776 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35052 0 1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_69_358
timestamp 1586364061
transform 1 0 34040 0 1 39712
box -38 -48 774 592
use scs8hd_fill_2  FILLER_69_367
timestamp 1586364061
transform 1 0 34868 0 1 39712
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 36800 0 1 39712
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 36616 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38088 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__445__A
timestamp 1586364061
transform 1 0 36248 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_380
timestamp 1586364061
transform 1 0 36064 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_384
timestamp 1586364061
transform 1 0 36432 0 1 39712
box -38 -48 222 592
use scs8hd_decap_3  FILLER_69_399
timestamp 1586364061
transform 1 0 37812 0 1 39712
box -38 -48 314 592
use scs8hd_decap_3  FILLER_69_404
timestamp 1586364061
transform 1 0 38272 0 1 39712
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38548 0 1 39712
box -38 -48 866 592
use scs8hd_fill_2  FILLER_69_420
timestamp 1586364061
transform 1 0 39744 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_416
timestamp 1586364061
transform 1 0 39376 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39560 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39928 0 1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_69_428
timestamp 1586364061
transform 1 0 40480 0 1 39712
box -38 -48 130 592
use scs8hd_decap_3  FILLER_69_424
timestamp 1586364061
transform 1 0 40112 0 1 39712
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_732
timestamp 1586364061
transform 1 0 40388 0 1 39712
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40572 0 1 39712
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41584 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41032 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42964 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41400 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42596 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_432
timestamp 1586364061
transform 1 0 40848 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_436
timestamp 1586364061
transform 1 0 41216 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_449
timestamp 1586364061
transform 1 0 42412 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_453
timestamp 1586364061
transform 1 0 42780 0 1 39712
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43148 0 1 39712
box -38 -48 866 592
use scs8hd_decap_12  FILLER_69_466
timestamp 1586364061
transform 1 0 43976 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_69_478
timestamp 1586364061
transform 1 0 45080 0 1 39712
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_733
timestamp 1586364061
transform 1 0 46000 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_486
timestamp 1586364061
transform 1 0 45816 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_489
timestamp 1586364061
transform 1 0 46092 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_501
timestamp 1586364061
transform 1 0 47196 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_139
timestamp 1586364061
transform -1 0 48852 0 1 39712
box -38 -48 314 592
use scs8hd_decap_3  FILLER_69_513
timestamp 1586364061
transform 1 0 48300 0 1 39712
box -38 -48 314 592
use scs8hd_decap_3  PHY_140
timestamp 1586364061
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_70_3
timestamp 1586364061
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_15
timestamp 1586364061
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_734
timestamp 1586364061
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_4  FILLER_70_27
timestamp 1586364061
transform 1 0 3588 0 -1 40800
box -38 -48 406 592
use scs8hd_decap_12  FILLER_70_32
timestamp 1586364061
transform 1 0 4048 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_44
timestamp 1586364061
transform 1 0 5152 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_56
timestamp 1586364061
transform 1 0 6256 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_68
timestamp 1586364061
transform 1 0 7360 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_80
timestamp 1586364061
transform 1 0 8464 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_735
timestamp 1586364061
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_93
timestamp 1586364061
transform 1 0 9660 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_105
timestamp 1586364061
transform 1 0 10764 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_117
timestamp 1586364061
transform 1 0 11868 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_129
timestamp 1586364061
transform 1 0 12972 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_736
timestamp 1586364061
transform 1 0 15180 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_141
timestamp 1586364061
transform 1 0 14076 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_154
timestamp 1586364061
transform 1 0 15272 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_166
timestamp 1586364061
transform 1 0 16376 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_178
timestamp 1586364061
transform 1 0 17480 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_737
timestamp 1586364061
transform 1 0 20792 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_190
timestamp 1586364061
transform 1 0 18584 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_202
timestamp 1586364061
transform 1 0 19688 0 -1 40800
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 -1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22356 0 -1 40800
box -38 -48 866 592
use scs8hd_decap_4  FILLER_70_215
timestamp 1586364061
transform 1 0 20884 0 -1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_70_219
timestamp 1586364061
transform 1 0 21252 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_8  FILLER_70_223
timestamp 1586364061
transform 1 0 21620 0 -1 40800
box -38 -48 774 592
use scs8hd_fill_2  FILLER_70_240
timestamp 1586364061
transform 1 0 23184 0 -1 40800
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 -1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25208 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_70_244
timestamp 1586364061
transform 1 0 23552 0 -1 40800
box -38 -48 406 592
use scs8hd_decap_4  FILLER_70_257
timestamp 1586364061
transform 1 0 24748 0 -1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_70_261
timestamp 1586364061
transform 1 0 25116 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_8  FILLER_70_264
timestamp 1586364061
transform 1 0 25392 0 -1 40800
box -38 -48 774 592
use scs8hd_nor2_4  _464_
timestamp 1586364061
transform 1 0 27324 0 -1 40800
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_738
timestamp 1586364061
transform 1 0 26404 0 -1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26956 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_3  FILLER_70_272
timestamp 1586364061
transform 1 0 26128 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_4  FILLER_70_276
timestamp 1586364061
transform 1 0 26496 0 -1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_70_280
timestamp 1586364061
transform 1 0 26864 0 -1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_70_283
timestamp 1586364061
transform 1 0 27140 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_294
timestamp 1586364061
transform 1 0 28152 0 -1 40800
box -38 -48 774 592
use scs8hd_buf_1  _450_
timestamp 1586364061
transform 1 0 28980 0 -1 40800
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 29992 0 -1 40800
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__453__B
timestamp 1586364061
transform 1 0 29440 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29808 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_1  FILLER_70_302
timestamp 1586364061
transform 1 0 28888 0 -1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_70_306
timestamp 1586364061
transform 1 0 29256 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_310
timestamp 1586364061
transform 1 0 29624 0 -1 40800
box -38 -48 222 592
use scs8hd_buf_1  _451_
timestamp 1586364061
transform 1 0 32108 0 -1 40800
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_739
timestamp 1586364061
transform 1 0 32016 0 -1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__457__B
timestamp 1586364061
transform 1 0 31188 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_325
timestamp 1586364061
transform 1 0 31004 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_70_329
timestamp 1586364061
transform 1 0 31372 0 -1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_70_333
timestamp 1586364061
transform 1 0 31740 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_8  FILLER_70_340
timestamp 1586364061
transform 1 0 32384 0 -1 40800
box -38 -48 774 592
use scs8hd_fill_2  FILLER_70_348
timestamp 1586364061
transform 1 0 33120 0 -1 40800
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 -1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33304 0 -1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__443__B
timestamp 1586364061
transform 1 0 35328 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_359
timestamp 1586364061
transform 1 0 34132 0 -1 40800
box -38 -48 774 592
use scs8hd_fill_2  FILLER_70_370
timestamp 1586364061
transform 1 0 35144 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_374
timestamp 1586364061
transform 1 0 35512 0 -1 40800
box -38 -48 222 592
use scs8hd_nor2_4  _445_
timestamp 1586364061
transform 1 0 35880 0 -1 40800
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38088 0 -1 40800
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_740
timestamp 1586364061
transform 1 0 37628 0 -1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35696 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_387
timestamp 1586364061
transform 1 0 36708 0 -1 40800
box -38 -48 774 592
use scs8hd_fill_2  FILLER_70_395
timestamp 1586364061
transform 1 0 37444 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_70_398
timestamp 1586364061
transform 1 0 37720 0 -1 40800
box -38 -48 406 592
use scs8hd_fill_2  FILLER_70_409
timestamp 1586364061
transform 1 0 38732 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_405
timestamp 1586364061
transform 1 0 38364 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38916 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38548 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_413
timestamp 1586364061
transform 1 0 39100 0 -1 40800
box -38 -48 774 592
use scs8hd_fill_2  FILLER_70_429
timestamp 1586364061
transform 1 0 40572 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_425
timestamp 1586364061
transform 1 0 40204 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_1  FILLER_70_421
timestamp 1586364061
transform 1 0 39836 0 -1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40388 0 -1 40800
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39928 0 -1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41584 0 -1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40756 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41400 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_70_433
timestamp 1586364061
transform 1 0 40940 0 -1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_70_437
timestamp 1586364061
transform 1 0 41308 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_8  FILLER_70_449
timestamp 1586364061
transform 1 0 42412 0 -1 40800
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_741
timestamp 1586364061
transform 1 0 43240 0 -1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43516 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_1  FILLER_70_457
timestamp 1586364061
transform 1 0 43148 0 -1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_70_459
timestamp 1586364061
transform 1 0 43332 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_70_463
timestamp 1586364061
transform 1 0 43700 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_475
timestamp 1586364061
transform 1 0 44804 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_487
timestamp 1586364061
transform 1 0 45908 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_499
timestamp 1586364061
transform 1 0 47012 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_141
timestamp 1586364061
transform -1 0 48852 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_4  FILLER_70_511
timestamp 1586364061
transform 1 0 48116 0 -1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_70_515
timestamp 1586364061
transform 1 0 48484 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_3  PHY_142
timestamp 1586364061
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_71_3
timestamp 1586364061
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_15
timestamp 1586364061
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_27
timestamp 1586364061
transform 1 0 3588 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_39
timestamp 1586364061
transform 1 0 4692 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_71_51
timestamp 1586364061
transform 1 0 5796 0 1 40800
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_742
timestamp 1586364061
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_59
timestamp 1586364061
transform 1 0 6532 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_62
timestamp 1586364061
transform 1 0 6808 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_74
timestamp 1586364061
transform 1 0 7912 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_86
timestamp 1586364061
transform 1 0 9016 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_98
timestamp 1586364061
transform 1 0 10120 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_743
timestamp 1586364061
transform 1 0 12328 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_110
timestamp 1586364061
transform 1 0 11224 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_123
timestamp 1586364061
transform 1 0 12420 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_135
timestamp 1586364061
transform 1 0 13524 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_147
timestamp 1586364061
transform 1 0 14628 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_159
timestamp 1586364061
transform 1 0 15732 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_744
timestamp 1586364061
transform 1 0 17940 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_171
timestamp 1586364061
transform 1 0 16836 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_184
timestamp 1586364061
transform 1 0 18032 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_196
timestamp 1586364061
transform 1 0 19136 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_208
timestamp 1586364061
transform 1 0 20240 0 1 40800
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21804 0 1 40800
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22264 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23184 0 1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_71_220
timestamp 1586364061
transform 1 0 21344 0 1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_71_224
timestamp 1586364061
transform 1 0 21712 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_228
timestamp 1586364061
transform 1 0 22080 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_232
timestamp 1586364061
transform 1 0 22448 0 1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_71_236
timestamp 1586364061
transform 1 0 22816 0 1 40800
box -38 -48 406 592
use scs8hd_decap_4  FILLER_71_252
timestamp 1586364061
transform 1 0 24288 0 1 40800
box -38 -48 406 592
use scs8hd_fill_2  FILLER_71_248
timestamp 1586364061
transform 1 0 23920 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_242
timestamp 1586364061
transform 1 0 23368 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 40800
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_745
timestamp 1586364061
transform 1 0 23552 0 1 40800
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 40800
box -38 -48 314 592
use scs8hd_fill_2  FILLER_71_258
timestamp 1586364061
transform 1 0 24840 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 25024 0 1 40800
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 25208 0 1 40800
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 26956 0 1 40800
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 26772 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26404 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28152 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_273
timestamp 1586364061
transform 1 0 26220 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_277
timestamp 1586364061
transform 1 0 26588 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_292
timestamp 1586364061
transform 1 0 27968 0 1 40800
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 30084 0 1 40800
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_746
timestamp 1586364061
transform 1 0 29164 0 1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 29900 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__454__A
timestamp 1586364061
transform 1 0 28888 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__454__B
timestamp 1586364061
transform 1 0 29440 0 1 40800
box -38 -48 222 592
use scs8hd_decap_6  FILLER_71_296
timestamp 1586364061
transform 1 0 28336 0 1 40800
box -38 -48 590 592
use scs8hd_fill_1  FILLER_71_304
timestamp 1586364061
transform 1 0 29072 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_306
timestamp 1586364061
transform 1 0 29256 0 1 40800
box -38 -48 222 592
use scs8hd_decap_3  FILLER_71_310
timestamp 1586364061
transform 1 0 29624 0 1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31832 0 1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32844 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31280 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31648 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_326
timestamp 1586364061
transform 1 0 31096 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_330
timestamp 1586364061
transform 1 0 31464 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_343
timestamp 1586364061
transform 1 0 32660 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_347
timestamp 1586364061
transform 1 0 33028 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_358
timestamp 1586364061
transform 1 0 34040 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_354
timestamp 1586364061
transform 1 0 33672 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33212 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33856 0 1 40800
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33396 0 1 40800
box -38 -48 314 592
use scs8hd_fill_2  FILLER_71_362
timestamp 1586364061
transform 1 0 34408 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 40800
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_747
timestamp 1586364061
transform 1 0 34776 0 1 40800
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 40800
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 36616 0 1 40800
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 36432 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37812 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_376
timestamp 1586364061
transform 1 0 35696 0 1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_71_380
timestamp 1586364061
transform 1 0 36064 0 1 40800
box -38 -48 406 592
use scs8hd_fill_2  FILLER_71_397
timestamp 1586364061
transform 1 0 37628 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_401
timestamp 1586364061
transform 1 0 37996 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38180 0 1 40800
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38364 0 1 40800
box -38 -48 866 592
use scs8hd_decap_3  FILLER_71_418
timestamp 1586364061
transform 1 0 39560 0 1 40800
box -38 -48 314 592
use scs8hd_fill_2  FILLER_71_414
timestamp 1586364061
transform 1 0 39192 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39376 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39836 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_423
timestamp 1586364061
transform 1 0 40020 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 40800
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_748
timestamp 1586364061
transform 1 0 40388 0 1 40800
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 40800
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42044 0 1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41768 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_71_437
timestamp 1586364061
transform 1 0 41308 0 1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_71_441
timestamp 1586364061
transform 1 0 41676 0 1 40800
box -38 -48 130 592
use scs8hd_fill_1  FILLER_71_444
timestamp 1586364061
transform 1 0 41952 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_454
timestamp 1586364061
transform 1 0 42872 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_458
timestamp 1586364061
transform 1 0 43240 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_470
timestamp 1586364061
transform 1 0 44344 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_71_482
timestamp 1586364061
transform 1 0 45448 0 1 40800
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_749
timestamp 1586364061
transform 1 0 46000 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_489
timestamp 1586364061
transform 1 0 46092 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_501
timestamp 1586364061
transform 1 0 47196 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_143
timestamp 1586364061
transform -1 0 48852 0 1 40800
box -38 -48 314 592
use scs8hd_decap_3  FILLER_71_513
timestamp 1586364061
transform 1 0 48300 0 1 40800
box -38 -48 314 592
use scs8hd_decap_3  PHY_144
timestamp 1586364061
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_146
timestamp 1586364061
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_72_3
timestamp 1586364061
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_15
timestamp 1586364061
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_3
timestamp 1586364061
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_15
timestamp 1586364061
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_750
timestamp 1586364061
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_27
timestamp 1586364061
transform 1 0 3588 0 -1 41888
box -38 -48 406 592
use scs8hd_decap_12  FILLER_72_32
timestamp 1586364061
transform 1 0 4048 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_44
timestamp 1586364061
transform 1 0 5152 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_27
timestamp 1586364061
transform 1 0 3588 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_39
timestamp 1586364061
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_73_51
timestamp 1586364061
transform 1 0 5796 0 1 41888
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_758
timestamp 1586364061
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_56
timestamp 1586364061
transform 1 0 6256 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_68
timestamp 1586364061
transform 1 0 7360 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_80
timestamp 1586364061
transform 1 0 8464 0 -1 41888
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_73_59
timestamp 1586364061
transform 1 0 6532 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_73_62
timestamp 1586364061
transform 1 0 6808 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_74
timestamp 1586364061
transform 1 0 7912 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_751
timestamp 1586364061
transform 1 0 9568 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_93
timestamp 1586364061
transform 1 0 9660 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_105
timestamp 1586364061
transform 1 0 10764 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_86
timestamp 1586364061
transform 1 0 9016 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_98
timestamp 1586364061
transform 1 0 10120 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_759
timestamp 1586364061
transform 1 0 12328 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_117
timestamp 1586364061
transform 1 0 11868 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_129
timestamp 1586364061
transform 1 0 12972 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_110
timestamp 1586364061
transform 1 0 11224 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_123
timestamp 1586364061
transform 1 0 12420 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_752
timestamp 1586364061
transform 1 0 15180 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_141
timestamp 1586364061
transform 1 0 14076 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_154
timestamp 1586364061
transform 1 0 15272 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_135
timestamp 1586364061
transform 1 0 13524 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_147
timestamp 1586364061
transform 1 0 14628 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_159
timestamp 1586364061
transform 1 0 15732 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_760
timestamp 1586364061
transform 1 0 17940 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_166
timestamp 1586364061
transform 1 0 16376 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_178
timestamp 1586364061
transform 1 0 17480 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_171
timestamp 1586364061
transform 1 0 16836 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_184
timestamp 1586364061
transform 1 0 18032 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_753
timestamp 1586364061
transform 1 0 20792 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_190
timestamp 1586364061
transform 1 0 18584 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_202
timestamp 1586364061
transform 1 0 19688 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_196
timestamp 1586364061
transform 1 0 19136 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_73_208
timestamp 1586364061
transform 1 0 20240 0 1 41888
box -38 -48 774 592
use scs8hd_fill_2  FILLER_73_223
timestamp 1586364061
transform 1 0 21620 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_219
timestamp 1586364061
transform 1 0 21252 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_72_215
timestamp 1586364061
transform 1 0 20884 0 -1 41888
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 41888
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20976 0 1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_240
timestamp 1586364061
transform 1 0 23184 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_236
timestamp 1586364061
transform 1 0 22816 0 1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_232
timestamp 1586364061
transform 1 0 22448 0 -1 41888
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23184 0 -1 41888
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 -1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_72_249
timestamp 1586364061
transform 1 0 24012 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_761
timestamp 1586364061
transform 1 0 23552 0 1 41888
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 41888
box -38 -48 866 592
use scs8hd_decap_4  FILLER_73_258
timestamp 1586364061
transform 1 0 24840 0 1 41888
box -38 -48 406 592
use scs8hd_fill_2  FILLER_73_254
timestamp 1586364061
transform 1 0 24472 0 1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_253
timestamp 1586364061
transform 1 0 24380 0 -1 41888
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 41888
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25116 0 -1 41888
box -38 -48 314 592
use scs8hd_fill_1  FILLER_73_264
timestamp 1586364061
transform 1 0 25392 0 1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_268
timestamp 1586364061
transform 1 0 25760 0 -1 41888
box -38 -48 406 592
use scs8hd_fill_2  FILLER_72_264
timestamp 1586364061
transform 1 0 25392 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25576 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25484 0 1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_73_278
timestamp 1586364061
transform 1 0 26680 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_274
timestamp 1586364061
transform 1 0 26312 0 1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_72_272
timestamp 1586364061
transform 1 0 26128 0 -1 41888
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26864 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_754
timestamp 1586364061
transform 1 0 26404 0 -1 41888
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_73_282
timestamp 1586364061
transform 1 0 27048 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_72_285
timestamp 1586364061
transform 1 0 27324 0 -1 41888
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 27232 0 1 41888
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 27416 0 1 41888
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_73_306
timestamp 1586364061
transform 1 0 29256 0 1 41888
box -38 -48 314 592
use scs8hd_fill_1  FILLER_73_304
timestamp 1586364061
transform 1 0 29072 0 1 41888
box -38 -48 130 592
use scs8hd_fill_1  FILLER_73_301
timestamp 1586364061
transform 1 0 28796 0 1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_73_297
timestamp 1586364061
transform 1 0 28428 0 1 41888
box -38 -48 406 592
use scs8hd_decap_3  FILLER_72_297
timestamp 1586364061
transform 1 0 28428 0 -1 41888
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__456__B
timestamp 1586364061
transform 1 0 28704 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__456__A
timestamp 1586364061
transform 1 0 28888 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_762
timestamp 1586364061
transform 1 0 29164 0 1 41888
box -38 -48 130 592
use scs8hd_nor2_4  _454_
timestamp 1586364061
transform 1 0 28888 0 -1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_72_315
timestamp 1586364061
transform 1 0 30084 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_311
timestamp 1586364061
transform 1 0 29716 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30268 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29900 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 29532 0 1 41888
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29716 0 1 41888
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_73_322
timestamp 1586364061
transform 1 0 30728 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 41888
box -38 -48 866 592
use scs8hd_decap_4  FILLER_73_330
timestamp 1586364061
transform 1 0 31464 0 1 41888
box -38 -48 406 592
use scs8hd_fill_2  FILLER_73_326
timestamp 1586364061
transform 1 0 31096 0 1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_328
timestamp 1586364061
transform 1 0 31280 0 -1 41888
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31280 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30912 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_338
timestamp 1586364061
transform 1 0 32200 0 1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_73_334
timestamp 1586364061
transform 1 0 31832 0 1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_337
timestamp 1586364061
transform 1 0 32108 0 -1 41888
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_755
timestamp 1586364061
transform 1 0 32016 0 -1 41888
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31924 0 1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_342
timestamp 1586364061
transform 1 0 32568 0 1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_345
timestamp 1586364061
transform 1 0 32844 0 -1 41888
box -38 -48 774 592
use scs8hd_fill_1  FILLER_72_341
timestamp 1586364061
transform 1 0 32476 0 -1 41888
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32752 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32384 0 1 41888
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32936 0 1 41888
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32568 0 -1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_357
timestamp 1586364061
transform 1 0 33948 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_353
timestamp 1586364061
transform 1 0 33580 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_349
timestamp 1586364061
transform 1 0 33212 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33764 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33396 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33580 0 -1 41888
box -38 -48 866 592
use scs8hd_decap_3  FILLER_73_361
timestamp 1586364061
transform 1 0 34316 0 1 41888
box -38 -48 314 592
use scs8hd_fill_1  FILLER_72_366
timestamp 1586364061
transform 1 0 34776 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_362
timestamp 1586364061
transform 1 0 34408 0 -1 41888
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34132 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_763
timestamp 1586364061
transform 1 0 34776 0 1 41888
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_374
timestamp 1586364061
transform 1 0 35512 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_370
timestamp 1586364061
transform 1 0 35144 0 1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_72_369
timestamp 1586364061
transform 1 0 35052 0 -1 41888
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35144 0 -1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_73_381
timestamp 1586364061
transform 1 0 36156 0 1 41888
box -38 -48 222 592
use scs8hd_decap_6  FILLER_72_379
timestamp 1586364061
transform 1 0 35972 0 -1 41888
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35696 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36340 0 1 41888
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35880 0 1 41888
box -38 -48 314 592
use scs8hd_fill_1  FILLER_73_393
timestamp 1586364061
transform 1 0 37260 0 1 41888
box -38 -48 130 592
use scs8hd_decap_8  FILLER_73_385
timestamp 1586364061
transform 1 0 36524 0 1 41888
box -38 -48 774 592
use scs8hd_decap_8  FILLER_72_388
timestamp 1586364061
transform 1 0 36800 0 -1 41888
box -38 -48 774 592
use scs8hd_fill_1  FILLER_72_385
timestamp 1586364061
transform 1 0 36524 0 -1 41888
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36616 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_401
timestamp 1586364061
transform 1 0 37996 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_397
timestamp 1586364061
transform 1 0 37628 0 1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_398
timestamp 1586364061
transform 1 0 37720 0 -1 41888
box -38 -48 774 592
use scs8hd_fill_1  FILLER_72_396
timestamp 1586364061
transform 1 0 37536 0 -1 41888
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37812 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_756
timestamp 1586364061
transform 1 0 37628 0 -1 41888
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37352 0 1 41888
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38180 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38456 0 -1 41888
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38364 0 1 41888
box -38 -48 866 592
use scs8hd_decap_3  FILLER_73_418
timestamp 1586364061
transform 1 0 39560 0 1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_414
timestamp 1586364061
transform 1 0 39192 0 1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_415
timestamp 1586364061
transform 1 0 39284 0 -1 41888
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39376 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 41888
box -38 -48 222 592
use scs8hd_decap_4  FILLER_73_423
timestamp 1586364061
transform 1 0 40020 0 1 41888
box -38 -48 406 592
use scs8hd_fill_2  FILLER_72_423
timestamp 1586364061
transform 1 0 40020 0 -1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_764
timestamp 1586364061
transform 1 0 40388 0 1 41888
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40204 0 -1 41888
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 41888
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41768 0 -1 41888
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42228 0 -1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_434
timestamp 1586364061
transform 1 0 41032 0 -1 41888
box -38 -48 774 592
use scs8hd_fill_2  FILLER_72_445
timestamp 1586364061
transform 1 0 42044 0 -1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_449
timestamp 1586364061
transform 1 0 42412 0 -1 41888
box -38 -48 774 592
use scs8hd_fill_2  FILLER_73_431
timestamp 1586364061
transform 1 0 40756 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_73_435
timestamp 1586364061
transform 1 0 41124 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_447
timestamp 1586364061
transform 1 0 42228 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_757
timestamp 1586364061
transform 1 0 43240 0 -1 41888
box -38 -48 130 592
use scs8hd_fill_1  FILLER_72_457
timestamp 1586364061
transform 1 0 43148 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_459
timestamp 1586364061
transform 1 0 43332 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_471
timestamp 1586364061
transform 1 0 44436 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_483
timestamp 1586364061
transform 1 0 45540 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_459
timestamp 1586364061
transform 1 0 43332 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_471
timestamp 1586364061
transform 1 0 44436 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_73_483
timestamp 1586364061
transform 1 0 45540 0 1 41888
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_765
timestamp 1586364061
transform 1 0 46000 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_495
timestamp 1586364061
transform 1 0 46644 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_72_507
timestamp 1586364061
transform 1 0 47748 0 -1 41888
box -38 -48 774 592
use scs8hd_fill_1  FILLER_73_487
timestamp 1586364061
transform 1 0 45908 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_73_489
timestamp 1586364061
transform 1 0 46092 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_501
timestamp 1586364061
transform 1 0 47196 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_3  PHY_145
timestamp 1586364061
transform -1 0 48852 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_147
timestamp 1586364061
transform -1 0 48852 0 1 41888
box -38 -48 314 592
use scs8hd_fill_1  FILLER_72_515
timestamp 1586364061
transform 1 0 48484 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_3  FILLER_73_513
timestamp 1586364061
transform 1 0 48300 0 1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_148
timestamp 1586364061
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_74_3
timestamp 1586364061
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_15
timestamp 1586364061
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_766
timestamp 1586364061
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_74_27
timestamp 1586364061
transform 1 0 3588 0 -1 42976
box -38 -48 406 592
use scs8hd_decap_12  FILLER_74_32
timestamp 1586364061
transform 1 0 4048 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_44
timestamp 1586364061
transform 1 0 5152 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_56
timestamp 1586364061
transform 1 0 6256 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_68
timestamp 1586364061
transform 1 0 7360 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_80
timestamp 1586364061
transform 1 0 8464 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_767
timestamp 1586364061
transform 1 0 9568 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_93
timestamp 1586364061
transform 1 0 9660 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_105
timestamp 1586364061
transform 1 0 10764 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_117
timestamp 1586364061
transform 1 0 11868 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_129
timestamp 1586364061
transform 1 0 12972 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_768
timestamp 1586364061
transform 1 0 15180 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_141
timestamp 1586364061
transform 1 0 14076 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_154
timestamp 1586364061
transform 1 0 15272 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_166
timestamp 1586364061
transform 1 0 16376 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_178
timestamp 1586364061
transform 1 0 17480 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_769
timestamp 1586364061
transform 1 0 20792 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_190
timestamp 1586364061
transform 1 0 18584 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_202
timestamp 1586364061
transform 1 0 19688 0 -1 42976
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22356 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_74_215
timestamp 1586364061
transform 1 0 20884 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_74_227
timestamp 1586364061
transform 1 0 21988 0 -1 42976
box -38 -48 406 592
use scs8hd_decap_8  FILLER_74_234
timestamp 1586364061
transform 1 0 22632 0 -1 42976
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 -1 42976
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23460 0 -1 42976
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 -1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24472 0 -1 42976
box -38 -48 222 592
use scs8hd_fill_1  FILLER_74_242
timestamp 1586364061
transform 1 0 23368 0 -1 42976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_74_252
timestamp 1586364061
transform 1 0 24288 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_6  FILLER_74_256
timestamp 1586364061
transform 1 0 24656 0 -1 42976
box -38 -48 590 592
use scs8hd_fill_2  FILLER_74_265
timestamp 1586364061
transform 1 0 25484 0 -1 42976
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 42976
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_770
timestamp 1586364061
transform 1 0 26404 0 -1 42976
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__467__B
timestamp 1586364061
transform 1 0 27508 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_6  FILLER_74_269
timestamp 1586364061
transform 1 0 25852 0 -1 42976
box -38 -48 590 592
use scs8hd_fill_2  FILLER_74_285
timestamp 1586364061
transform 1 0 27324 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_74_289
timestamp 1586364061
transform 1 0 27692 0 -1 42976
box -38 -48 1142 592
use scs8hd_nor2_4  _456_
timestamp 1586364061
transform 1 0 28888 0 -1 42976
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 42976
box -38 -48 866 592
use scs8hd_fill_1  FILLER_74_301
timestamp 1586364061
transform 1 0 28796 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_8  FILLER_74_311
timestamp 1586364061
transform 1 0 29716 0 -1 42976
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32384 0 -1 42976
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_771
timestamp 1586364061
transform 1 0 32016 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_8  FILLER_74_328
timestamp 1586364061
transform 1 0 31280 0 -1 42976
box -38 -48 774 592
use scs8hd_decap_3  FILLER_74_337
timestamp 1586364061
transform 1 0 32108 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_8  FILLER_74_343
timestamp 1586364061
transform 1 0 32660 0 -1 42976
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34960 0 -1 42976
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33396 0 -1 42976
box -38 -48 866 592
use scs8hd_decap_8  FILLER_74_360
timestamp 1586364061
transform 1 0 34224 0 -1 42976
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38088 0 -1 42976
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_772
timestamp 1586364061
transform 1 0 37628 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_377
timestamp 1586364061
transform 1 0 35788 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_74_389
timestamp 1586364061
transform 1 0 36892 0 -1 42976
box -38 -48 774 592
use scs8hd_decap_4  FILLER_74_398
timestamp 1586364061
transform 1 0 37720 0 -1 42976
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39836 0 -1 42976
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38548 0 -1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_74_405
timestamp 1586364061
transform 1 0 38364 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_74_409
timestamp 1586364061
transform 1 0 38732 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_424
timestamp 1586364061
transform 1 0 40112 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_436
timestamp 1586364061
transform 1 0 41216 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_74_448
timestamp 1586364061
transform 1 0 42320 0 -1 42976
box -38 -48 774 592
use scs8hd_fill_2  FILLER_74_456
timestamp 1586364061
transform 1 0 43056 0 -1 42976
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_773
timestamp 1586364061
transform 1 0 43240 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_459
timestamp 1586364061
transform 1 0 43332 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_471
timestamp 1586364061
transform 1 0 44436 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_483
timestamp 1586364061
transform 1 0 45540 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_495
timestamp 1586364061
transform 1 0 46644 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_74_507
timestamp 1586364061
transform 1 0 47748 0 -1 42976
box -38 -48 774 592
use scs8hd_decap_3  PHY_149
timestamp 1586364061
transform -1 0 48852 0 -1 42976
box -38 -48 314 592
use scs8hd_fill_1  FILLER_74_515
timestamp 1586364061
transform 1 0 48484 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_3  PHY_150
timestamp 1586364061
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_75_3
timestamp 1586364061
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_15
timestamp 1586364061
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_27
timestamp 1586364061
transform 1 0 3588 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_39
timestamp 1586364061
transform 1 0 4692 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_75_51
timestamp 1586364061
transform 1 0 5796 0 1 42976
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_774
timestamp 1586364061
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_75_59
timestamp 1586364061
transform 1 0 6532 0 1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_75_62
timestamp 1586364061
transform 1 0 6808 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_74
timestamp 1586364061
transform 1 0 7912 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_86
timestamp 1586364061
transform 1 0 9016 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_98
timestamp 1586364061
transform 1 0 10120 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_775
timestamp 1586364061
transform 1 0 12328 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_110
timestamp 1586364061
transform 1 0 11224 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_123
timestamp 1586364061
transform 1 0 12420 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_135
timestamp 1586364061
transform 1 0 13524 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_147
timestamp 1586364061
transform 1 0 14628 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_159
timestamp 1586364061
transform 1 0 15732 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_776
timestamp 1586364061
transform 1 0 17940 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_171
timestamp 1586364061
transform 1 0 16836 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_184
timestamp 1586364061
transform 1 0 18032 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_196
timestamp 1586364061
transform 1 0 19136 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_208
timestamp 1586364061
transform 1 0 20240 0 1 42976
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 42976
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23092 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 42976
box -38 -48 222 592
use scs8hd_decap_8  FILLER_75_220
timestamp 1586364061
transform 1 0 21344 0 1 42976
box -38 -48 774 592
use scs8hd_decap_3  FILLER_75_228
timestamp 1586364061
transform 1 0 22080 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  FILLER_75_236
timestamp 1586364061
transform 1 0 22816 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  FILLER_75_241
timestamp 1586364061
transform 1 0 23276 0 1 42976
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25392 0 1 42976
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 42976
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_777
timestamp 1586364061
transform 1 0 23552 0 1 42976
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_254
timestamp 1586364061
transform 1 0 24472 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_258
timestamp 1586364061
transform 1 0 24840 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_262
timestamp 1586364061
transform 1 0 25208 0 1 42976
box -38 -48 222 592
use scs8hd_nor2_4  _467_
timestamp 1586364061
transform 1 0 27508 0 1 42976
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__467__A
timestamp 1586364061
transform 1 0 27324 0 1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_75_273
timestamp 1586364061
transform 1 0 26220 0 1 42976
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_75_304
timestamp 1586364061
transform 1 0 29072 0 1 42976
box -38 -48 130 592
use scs8hd_decap_8  FILLER_75_296
timestamp 1586364061
transform 1 0 28336 0 1 42976
box -38 -48 774 592
use scs8hd_fill_1  FILLER_75_312
timestamp 1586364061
transform 1 0 29808 0 1 42976
box -38 -48 130 592
use scs8hd_decap_6  FILLER_75_306
timestamp 1586364061
transform 1 0 29256 0 1 42976
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_778
timestamp 1586364061
transform 1 0 29164 0 1 42976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_75_320
timestamp 1586364061
transform 1 0 30544 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_316
timestamp 1586364061
transform 1 0 30176 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30360 0 1 42976
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29900 0 1 42976
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30728 0 1 42976
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32476 0 1 42976
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30912 0 1 42976
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32292 0 1 42976
box -38 -48 222 592
use scs8hd_decap_6  FILLER_75_333
timestamp 1586364061
transform 1 0 31740 0 1 42976
box -38 -48 590 592
use scs8hd_decap_8  FILLER_75_358
timestamp 1586364061
transform 1 0 34040 0 1 42976
box -38 -48 774 592
use scs8hd_fill_2  FILLER_75_354
timestamp 1586364061
transform 1 0 33672 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_350
timestamp 1586364061
transform 1 0 33304 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33488 0 1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_75_374
timestamp 1586364061
transform 1 0 35512 0 1 42976
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_75_370
timestamp 1586364061
transform 1 0 35144 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 42976
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_779
timestamp 1586364061
transform 1 0 34776 0 1 42976
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_75_386
timestamp 1586364061
transform 1 0 36616 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_398
timestamp 1586364061
transform 1 0 37720 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_780
timestamp 1586364061
transform 1 0 40388 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_410
timestamp 1586364061
transform 1 0 38824 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_75_422
timestamp 1586364061
transform 1 0 39928 0 1 42976
box -38 -48 406 592
use scs8hd_fill_1  FILLER_75_426
timestamp 1586364061
transform 1 0 40296 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_428
timestamp 1586364061
transform 1 0 40480 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_440
timestamp 1586364061
transform 1 0 41584 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_452
timestamp 1586364061
transform 1 0 42688 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_464
timestamp 1586364061
transform 1 0 43792 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_476
timestamp 1586364061
transform 1 0 44896 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_781
timestamp 1586364061
transform 1 0 46000 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_489
timestamp 1586364061
transform 1 0 46092 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_501
timestamp 1586364061
transform 1 0 47196 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_151
timestamp 1586364061
transform -1 0 48852 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  FILLER_75_513
timestamp 1586364061
transform 1 0 48300 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  PHY_152
timestamp 1586364061
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_76_3
timestamp 1586364061
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_15
timestamp 1586364061
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_782
timestamp 1586364061
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_4  FILLER_76_27
timestamp 1586364061
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use scs8hd_decap_12  FILLER_76_32
timestamp 1586364061
transform 1 0 4048 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_44
timestamp 1586364061
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_56
timestamp 1586364061
transform 1 0 6256 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_68
timestamp 1586364061
transform 1 0 7360 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_80
timestamp 1586364061
transform 1 0 8464 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_783
timestamp 1586364061
transform 1 0 9568 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_93
timestamp 1586364061
transform 1 0 9660 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_105
timestamp 1586364061
transform 1 0 10764 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_117
timestamp 1586364061
transform 1 0 11868 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_129
timestamp 1586364061
transform 1 0 12972 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_784
timestamp 1586364061
transform 1 0 15180 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_141
timestamp 1586364061
transform 1 0 14076 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_154
timestamp 1586364061
transform 1 0 15272 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_166
timestamp 1586364061
transform 1 0 16376 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_178
timestamp 1586364061
transform 1 0 17480 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_785
timestamp 1586364061
transform 1 0 20792 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_190
timestamp 1586364061
transform 1 0 18584 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_202
timestamp 1586364061
transform 1 0 19688 0 -1 44064
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23092 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_76_215
timestamp 1586364061
transform 1 0 20884 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_227
timestamp 1586364061
transform 1 0 21988 0 -1 44064
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_76_247
timestamp 1586364061
transform 1 0 23828 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_3  FILLER_76_242
timestamp 1586364061
transform 1 0 23368 0 -1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23644 0 -1 44064
box -38 -48 222 592
use scs8hd_fill_1  FILLER_76_259
timestamp 1586364061
transform 1 0 24932 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_8  FILLER_76_251
timestamp 1586364061
transform 1 0 24196 0 -1 44064
box -38 -48 774 592
use scs8hd_decap_8  FILLER_76_267
timestamp 1586364061
transform 1 0 25668 0 -1 44064
box -38 -48 774 592
use scs8hd_fill_2  FILLER_76_263
timestamp 1586364061
transform 1 0 25300 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25484 0 -1 44064
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 44064
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_786
timestamp 1586364061
transform 1 0 26404 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_276
timestamp 1586364061
transform 1 0 26496 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_288
timestamp 1586364061
transform 1 0 27600 0 -1 44064
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30360 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_76_300
timestamp 1586364061
transform 1 0 28704 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_76_312
timestamp 1586364061
transform 1 0 29808 0 -1 44064
box -38 -48 590 592
use scs8hd_decap_3  FILLER_76_321
timestamp 1586364061
transform 1 0 30636 0 -1 44064
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_787
timestamp 1586364061
transform 1 0 32016 0 -1 44064
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30912 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31280 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32476 0 -1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_76_326
timestamp 1586364061
transform 1 0 31096 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_6  FILLER_76_330
timestamp 1586364061
transform 1 0 31464 0 -1 44064
box -38 -48 590 592
use scs8hd_decap_4  FILLER_76_337
timestamp 1586364061
transform 1 0 32108 0 -1 44064
box -38 -48 406 592
use scs8hd_decap_6  FILLER_76_343
timestamp 1586364061
transform 1 0 32660 0 -1 44064
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 -1 44064
box -38 -48 866 592
use scs8hd_decap_12  FILLER_76_358
timestamp 1586364061
transform 1 0 34040 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_370
timestamp 1586364061
transform 1 0 35144 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_788
timestamp 1586364061
transform 1 0 37628 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_382
timestamp 1586364061
transform 1 0 36248 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_76_394
timestamp 1586364061
transform 1 0 37352 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_76_398
timestamp 1586364061
transform 1 0 37720 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_410
timestamp 1586364061
transform 1 0 38824 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_422
timestamp 1586364061
transform 1 0 39928 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_434
timestamp 1586364061
transform 1 0 41032 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_446
timestamp 1586364061
transform 1 0 42136 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_789
timestamp 1586364061
transform 1 0 43240 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_459
timestamp 1586364061
transform 1 0 43332 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_471
timestamp 1586364061
transform 1 0 44436 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_483
timestamp 1586364061
transform 1 0 45540 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_495
timestamp 1586364061
transform 1 0 46644 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_76_507
timestamp 1586364061
transform 1 0 47748 0 -1 44064
box -38 -48 774 592
use scs8hd_decap_3  PHY_153
timestamp 1586364061
transform -1 0 48852 0 -1 44064
box -38 -48 314 592
use scs8hd_fill_1  FILLER_76_515
timestamp 1586364061
transform 1 0 48484 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_3  PHY_154
timestamp 1586364061
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_77_3
timestamp 1586364061
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_15
timestamp 1586364061
transform 1 0 2484 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_27
timestamp 1586364061
transform 1 0 3588 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_39
timestamp 1586364061
transform 1 0 4692 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_77_51
timestamp 1586364061
transform 1 0 5796 0 1 44064
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_790
timestamp 1586364061
transform 1 0 6716 0 1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_77_59
timestamp 1586364061
transform 1 0 6532 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_62
timestamp 1586364061
transform 1 0 6808 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_74
timestamp 1586364061
transform 1 0 7912 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_86
timestamp 1586364061
transform 1 0 9016 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_98
timestamp 1586364061
transform 1 0 10120 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_791
timestamp 1586364061
transform 1 0 12328 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_110
timestamp 1586364061
transform 1 0 11224 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_123
timestamp 1586364061
transform 1 0 12420 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_135
timestamp 1586364061
transform 1 0 13524 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_147
timestamp 1586364061
transform 1 0 14628 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_159
timestamp 1586364061
transform 1 0 15732 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_792
timestamp 1586364061
transform 1 0 17940 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_171
timestamp 1586364061
transform 1 0 16836 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_184
timestamp 1586364061
transform 1 0 18032 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_196
timestamp 1586364061
transform 1 0 19136 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_208
timestamp 1586364061
transform 1 0 20240 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_220
timestamp 1586364061
transform 1 0 21344 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_232
timestamp 1586364061
transform 1 0 22448 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_793
timestamp 1586364061
transform 1 0 23552 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_245
timestamp 1586364061
transform 1 0 23644 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_257
timestamp 1586364061
transform 1 0 24748 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_269
timestamp 1586364061
transform 1 0 25852 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_281
timestamp 1586364061
transform 1 0 26956 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_293
timestamp 1586364061
transform 1 0 28060 0 1 44064
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30636 0 1 44064
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_794
timestamp 1586364061
transform 1 0 29164 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_306
timestamp 1586364061
transform 1 0 29256 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_77_318
timestamp 1586364061
transform 1 0 30360 0 1 44064
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33120 0 1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31096 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_324
timestamp 1586364061
transform 1 0 30912 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_328
timestamp 1586364061
transform 1 0 31280 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_77_340
timestamp 1586364061
transform 1 0 32384 0 1 44064
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_795
timestamp 1586364061
transform 1 0 34776 0 1 44064
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33580 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_351
timestamp 1586364061
transform 1 0 33396 0 1 44064
box -38 -48 222 592
use scs8hd_decap_8  FILLER_77_355
timestamp 1586364061
transform 1 0 33764 0 1 44064
box -38 -48 774 592
use scs8hd_decap_3  FILLER_77_363
timestamp 1586364061
transform 1 0 34500 0 1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_77_367
timestamp 1586364061
transform 1 0 34868 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_379
timestamp 1586364061
transform 1 0 35972 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_391
timestamp 1586364061
transform 1 0 37076 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_796
timestamp 1586364061
transform 1 0 40388 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_403
timestamp 1586364061
transform 1 0 38180 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_415
timestamp 1586364061
transform 1 0 39284 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_428
timestamp 1586364061
transform 1 0 40480 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_440
timestamp 1586364061
transform 1 0 41584 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_452
timestamp 1586364061
transform 1 0 42688 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_464
timestamp 1586364061
transform 1 0 43792 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_476
timestamp 1586364061
transform 1 0 44896 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_797
timestamp 1586364061
transform 1 0 46000 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_489
timestamp 1586364061
transform 1 0 46092 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_501
timestamp 1586364061
transform 1 0 47196 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_155
timestamp 1586364061
transform -1 0 48852 0 1 44064
box -38 -48 314 592
use scs8hd_decap_3  FILLER_77_513
timestamp 1586364061
transform 1 0 48300 0 1 44064
box -38 -48 314 592
use scs8hd_decap_3  PHY_156
timestamp 1586364061
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_78_3
timestamp 1586364061
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_15
timestamp 1586364061
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_798
timestamp 1586364061
transform 1 0 3956 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_78_27
timestamp 1586364061
transform 1 0 3588 0 -1 45152
box -38 -48 406 592
use scs8hd_decap_12  FILLER_78_32
timestamp 1586364061
transform 1 0 4048 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_44
timestamp 1586364061
transform 1 0 5152 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_56
timestamp 1586364061
transform 1 0 6256 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_68
timestamp 1586364061
transform 1 0 7360 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_80
timestamp 1586364061
transform 1 0 8464 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_799
timestamp 1586364061
transform 1 0 9568 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_93
timestamp 1586364061
transform 1 0 9660 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_105
timestamp 1586364061
transform 1 0 10764 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_117
timestamp 1586364061
transform 1 0 11868 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_129
timestamp 1586364061
transform 1 0 12972 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_800
timestamp 1586364061
transform 1 0 15180 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_141
timestamp 1586364061
transform 1 0 14076 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_154
timestamp 1586364061
transform 1 0 15272 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_166
timestamp 1586364061
transform 1 0 16376 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_178
timestamp 1586364061
transform 1 0 17480 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_801
timestamp 1586364061
transform 1 0 20792 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_190
timestamp 1586364061
transform 1 0 18584 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_202
timestamp 1586364061
transform 1 0 19688 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_215
timestamp 1586364061
transform 1 0 20884 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_227
timestamp 1586364061
transform 1 0 21988 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_239
timestamp 1586364061
transform 1 0 23092 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_251
timestamp 1586364061
transform 1 0 24196 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_263
timestamp 1586364061
transform 1 0 25300 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_802
timestamp 1586364061
transform 1 0 26404 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_276
timestamp 1586364061
transform 1 0 26496 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_288
timestamp 1586364061
transform 1 0 27600 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_300
timestamp 1586364061
transform 1 0 28704 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_312
timestamp 1586364061
transform 1 0 29808 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_803
timestamp 1586364061
transform 1 0 32016 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_324
timestamp 1586364061
transform 1 0 30912 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_337
timestamp 1586364061
transform 1 0 32108 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_349
timestamp 1586364061
transform 1 0 33212 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_361
timestamp 1586364061
transform 1 0 34316 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_373
timestamp 1586364061
transform 1 0 35420 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_804
timestamp 1586364061
transform 1 0 37628 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_385
timestamp 1586364061
transform 1 0 36524 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_398
timestamp 1586364061
transform 1 0 37720 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_410
timestamp 1586364061
transform 1 0 38824 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_422
timestamp 1586364061
transform 1 0 39928 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_434
timestamp 1586364061
transform 1 0 41032 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_446
timestamp 1586364061
transform 1 0 42136 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_805
timestamp 1586364061
transform 1 0 43240 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_459
timestamp 1586364061
transform 1 0 43332 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_471
timestamp 1586364061
transform 1 0 44436 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_483
timestamp 1586364061
transform 1 0 45540 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_495
timestamp 1586364061
transform 1 0 46644 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_78_507
timestamp 1586364061
transform 1 0 47748 0 -1 45152
box -38 -48 774 592
use scs8hd_decap_3  PHY_157
timestamp 1586364061
transform -1 0 48852 0 -1 45152
box -38 -48 314 592
use scs8hd_fill_1  FILLER_78_515
timestamp 1586364061
transform 1 0 48484 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_3  PHY_158
timestamp 1586364061
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_160
timestamp 1586364061
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_79_3
timestamp 1586364061
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_15
timestamp 1586364061
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_3
timestamp 1586364061
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_15
timestamp 1586364061
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_814
timestamp 1586364061
transform 1 0 3956 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_27
timestamp 1586364061
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_39
timestamp 1586364061
transform 1 0 4692 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_79_51
timestamp 1586364061
transform 1 0 5796 0 1 45152
box -38 -48 774 592
use scs8hd_decap_4  FILLER_80_27
timestamp 1586364061
transform 1 0 3588 0 -1 46240
box -38 -48 406 592
use scs8hd_decap_12  FILLER_80_32
timestamp 1586364061
transform 1 0 4048 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_44
timestamp 1586364061
transform 1 0 5152 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_806
timestamp 1586364061
transform 1 0 6716 0 1 45152
box -38 -48 130 592
use scs8hd_fill_2  FILLER_79_59
timestamp 1586364061
transform 1 0 6532 0 1 45152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_79_62
timestamp 1586364061
transform 1 0 6808 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_74
timestamp 1586364061
transform 1 0 7912 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_56
timestamp 1586364061
transform 1 0 6256 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_68
timestamp 1586364061
transform 1 0 7360 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_80
timestamp 1586364061
transform 1 0 8464 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_815
timestamp 1586364061
transform 1 0 9568 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_86
timestamp 1586364061
transform 1 0 9016 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_98
timestamp 1586364061
transform 1 0 10120 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_93
timestamp 1586364061
transform 1 0 9660 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_105
timestamp 1586364061
transform 1 0 10764 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_807
timestamp 1586364061
transform 1 0 12328 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_110
timestamp 1586364061
transform 1 0 11224 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_123
timestamp 1586364061
transform 1 0 12420 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_117
timestamp 1586364061
transform 1 0 11868 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_129
timestamp 1586364061
transform 1 0 12972 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_816
timestamp 1586364061
transform 1 0 15180 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_135
timestamp 1586364061
transform 1 0 13524 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_147
timestamp 1586364061
transform 1 0 14628 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_159
timestamp 1586364061
transform 1 0 15732 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_141
timestamp 1586364061
transform 1 0 14076 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_154
timestamp 1586364061
transform 1 0 15272 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_808
timestamp 1586364061
transform 1 0 17940 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_171
timestamp 1586364061
transform 1 0 16836 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_184
timestamp 1586364061
transform 1 0 18032 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_166
timestamp 1586364061
transform 1 0 16376 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_178
timestamp 1586364061
transform 1 0 17480 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_817
timestamp 1586364061
transform 1 0 20792 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_196
timestamp 1586364061
transform 1 0 19136 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_208
timestamp 1586364061
transform 1 0 20240 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_190
timestamp 1586364061
transform 1 0 18584 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_202
timestamp 1586364061
transform 1 0 19688 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_220
timestamp 1586364061
transform 1 0 21344 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_232
timestamp 1586364061
transform 1 0 22448 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_215
timestamp 1586364061
transform 1 0 20884 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_227
timestamp 1586364061
transform 1 0 21988 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_239
timestamp 1586364061
transform 1 0 23092 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_809
timestamp 1586364061
transform 1 0 23552 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_245
timestamp 1586364061
transform 1 0 23644 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_257
timestamp 1586364061
transform 1 0 24748 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_251
timestamp 1586364061
transform 1 0 24196 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_263
timestamp 1586364061
transform 1 0 25300 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_818
timestamp 1586364061
transform 1 0 26404 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_269
timestamp 1586364061
transform 1 0 25852 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_281
timestamp 1586364061
transform 1 0 26956 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_293
timestamp 1586364061
transform 1 0 28060 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_276
timestamp 1586364061
transform 1 0 26496 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_288
timestamp 1586364061
transform 1 0 27600 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_810
timestamp 1586364061
transform 1 0 29164 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_306
timestamp 1586364061
transform 1 0 29256 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_318
timestamp 1586364061
transform 1 0 30360 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_300
timestamp 1586364061
transform 1 0 28704 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_312
timestamp 1586364061
transform 1 0 29808 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_819
timestamp 1586364061
transform 1 0 32016 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_330
timestamp 1586364061
transform 1 0 31464 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_342
timestamp 1586364061
transform 1 0 32568 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_324
timestamp 1586364061
transform 1 0 30912 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_337
timestamp 1586364061
transform 1 0 32108 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_811
timestamp 1586364061
transform 1 0 34776 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_354
timestamp 1586364061
transform 1 0 33672 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_367
timestamp 1586364061
transform 1 0 34868 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_349
timestamp 1586364061
transform 1 0 33212 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_361
timestamp 1586364061
transform 1 0 34316 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_373
timestamp 1586364061
transform 1 0 35420 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_820
timestamp 1586364061
transform 1 0 37628 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_379
timestamp 1586364061
transform 1 0 35972 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_391
timestamp 1586364061
transform 1 0 37076 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_385
timestamp 1586364061
transform 1 0 36524 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_398
timestamp 1586364061
transform 1 0 37720 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_812
timestamp 1586364061
transform 1 0 40388 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_403
timestamp 1586364061
transform 1 0 38180 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_415
timestamp 1586364061
transform 1 0 39284 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_428
timestamp 1586364061
transform 1 0 40480 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_410
timestamp 1586364061
transform 1 0 38824 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_422
timestamp 1586364061
transform 1 0 39928 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_440
timestamp 1586364061
transform 1 0 41584 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_452
timestamp 1586364061
transform 1 0 42688 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_434
timestamp 1586364061
transform 1 0 41032 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_446
timestamp 1586364061
transform 1 0 42136 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_821
timestamp 1586364061
transform 1 0 43240 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_464
timestamp 1586364061
transform 1 0 43792 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_476
timestamp 1586364061
transform 1 0 44896 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_459
timestamp 1586364061
transform 1 0 43332 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_471
timestamp 1586364061
transform 1 0 44436 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_483
timestamp 1586364061
transform 1 0 45540 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_813
timestamp 1586364061
transform 1 0 46000 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_489
timestamp 1586364061
transform 1 0 46092 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_501
timestamp 1586364061
transform 1 0 47196 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_495
timestamp 1586364061
transform 1 0 46644 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_80_507
timestamp 1586364061
transform 1 0 47748 0 -1 46240
box -38 -48 774 592
use scs8hd_decap_3  PHY_159
timestamp 1586364061
transform -1 0 48852 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_161
timestamp 1586364061
transform -1 0 48852 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_3  FILLER_79_513
timestamp 1586364061
transform 1 0 48300 0 1 45152
box -38 -48 314 592
use scs8hd_fill_1  FILLER_80_515
timestamp 1586364061
transform 1 0 48484 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_3  PHY_162
timestamp 1586364061
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_81_3
timestamp 1586364061
transform 1 0 1380 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_15
timestamp 1586364061
transform 1 0 2484 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_27
timestamp 1586364061
transform 1 0 3588 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_39
timestamp 1586364061
transform 1 0 4692 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_81_51
timestamp 1586364061
transform 1 0 5796 0 1 46240
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_822
timestamp 1586364061
transform 1 0 6716 0 1 46240
box -38 -48 130 592
use scs8hd_fill_2  FILLER_81_59
timestamp 1586364061
transform 1 0 6532 0 1 46240
box -38 -48 222 592
use scs8hd_decap_12  FILLER_81_62
timestamp 1586364061
transform 1 0 6808 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_74
timestamp 1586364061
transform 1 0 7912 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_86
timestamp 1586364061
transform 1 0 9016 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_98
timestamp 1586364061
transform 1 0 10120 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_823
timestamp 1586364061
transform 1 0 12328 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_110
timestamp 1586364061
transform 1 0 11224 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_123
timestamp 1586364061
transform 1 0 12420 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_135
timestamp 1586364061
transform 1 0 13524 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_147
timestamp 1586364061
transform 1 0 14628 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_159
timestamp 1586364061
transform 1 0 15732 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_824
timestamp 1586364061
transform 1 0 17940 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_171
timestamp 1586364061
transform 1 0 16836 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_184
timestamp 1586364061
transform 1 0 18032 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_196
timestamp 1586364061
transform 1 0 19136 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_208
timestamp 1586364061
transform 1 0 20240 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_220
timestamp 1586364061
transform 1 0 21344 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_232
timestamp 1586364061
transform 1 0 22448 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_825
timestamp 1586364061
transform 1 0 23552 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_245
timestamp 1586364061
transform 1 0 23644 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_257
timestamp 1586364061
transform 1 0 24748 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_269
timestamp 1586364061
transform 1 0 25852 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_281
timestamp 1586364061
transform 1 0 26956 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_293
timestamp 1586364061
transform 1 0 28060 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_826
timestamp 1586364061
transform 1 0 29164 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_306
timestamp 1586364061
transform 1 0 29256 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_318
timestamp 1586364061
transform 1 0 30360 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_330
timestamp 1586364061
transform 1 0 31464 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_342
timestamp 1586364061
transform 1 0 32568 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_827
timestamp 1586364061
transform 1 0 34776 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_354
timestamp 1586364061
transform 1 0 33672 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_367
timestamp 1586364061
transform 1 0 34868 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_379
timestamp 1586364061
transform 1 0 35972 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_391
timestamp 1586364061
transform 1 0 37076 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_828
timestamp 1586364061
transform 1 0 40388 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_403
timestamp 1586364061
transform 1 0 38180 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_415
timestamp 1586364061
transform 1 0 39284 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_428
timestamp 1586364061
transform 1 0 40480 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_440
timestamp 1586364061
transform 1 0 41584 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_452
timestamp 1586364061
transform 1 0 42688 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_464
timestamp 1586364061
transform 1 0 43792 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_476
timestamp 1586364061
transform 1 0 44896 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_829
timestamp 1586364061
transform 1 0 46000 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_489
timestamp 1586364061
transform 1 0 46092 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_501
timestamp 1586364061
transform 1 0 47196 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_3  PHY_163
timestamp 1586364061
transform -1 0 48852 0 1 46240
box -38 -48 314 592
use scs8hd_decap_3  FILLER_81_513
timestamp 1586364061
transform 1 0 48300 0 1 46240
box -38 -48 314 592
use scs8hd_decap_3  PHY_164
timestamp 1586364061
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_82_3
timestamp 1586364061
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_15
timestamp 1586364061
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_830
timestamp 1586364061
transform 1 0 3956 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_4  FILLER_82_27
timestamp 1586364061
transform 1 0 3588 0 -1 47328
box -38 -48 406 592
use scs8hd_decap_12  FILLER_82_32
timestamp 1586364061
transform 1 0 4048 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_44
timestamp 1586364061
transform 1 0 5152 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_831
timestamp 1586364061
transform 1 0 6808 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_56
timestamp 1586364061
transform 1 0 6256 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_63
timestamp 1586364061
transform 1 0 6900 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_75
timestamp 1586364061
transform 1 0 8004 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_832
timestamp 1586364061
transform 1 0 9660 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_87
timestamp 1586364061
transform 1 0 9108 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_94
timestamp 1586364061
transform 1 0 9752 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_106
timestamp 1586364061
transform 1 0 10856 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_833
timestamp 1586364061
transform 1 0 12512 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_118
timestamp 1586364061
transform 1 0 11960 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_125
timestamp 1586364061
transform 1 0 12604 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_834
timestamp 1586364061
transform 1 0 15364 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_137
timestamp 1586364061
transform 1 0 13708 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_149
timestamp 1586364061
transform 1 0 14812 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_156
timestamp 1586364061
transform 1 0 15456 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_835
timestamp 1586364061
transform 1 0 18216 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_168
timestamp 1586364061
transform 1 0 16560 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_180
timestamp 1586364061
transform 1 0 17664 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_187
timestamp 1586364061
transform 1 0 18308 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_199
timestamp 1586364061
transform 1 0 19412 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_211
timestamp 1586364061
transform 1 0 20516 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_836
timestamp 1586364061
transform 1 0 21068 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_218
timestamp 1586364061
transform 1 0 21160 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_230
timestamp 1586364061
transform 1 0 22264 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_837
timestamp 1586364061
transform 1 0 23920 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_242
timestamp 1586364061
transform 1 0 23368 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_249
timestamp 1586364061
transform 1 0 24012 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_261
timestamp 1586364061
transform 1 0 25116 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_838
timestamp 1586364061
transform 1 0 26772 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_273
timestamp 1586364061
transform 1 0 26220 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_280
timestamp 1586364061
transform 1 0 26864 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_292
timestamp 1586364061
transform 1 0 27968 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_839
timestamp 1586364061
transform 1 0 29624 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_304
timestamp 1586364061
transform 1 0 29072 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_311
timestamp 1586364061
transform 1 0 29716 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_840
timestamp 1586364061
transform 1 0 32476 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_323
timestamp 1586364061
transform 1 0 30820 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_335
timestamp 1586364061
transform 1 0 31924 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_342
timestamp 1586364061
transform 1 0 32568 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_841
timestamp 1586364061
transform 1 0 35328 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_354
timestamp 1586364061
transform 1 0 33672 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_366
timestamp 1586364061
transform 1 0 34776 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_373
timestamp 1586364061
transform 1 0 35420 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_385
timestamp 1586364061
transform 1 0 36524 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_397
timestamp 1586364061
transform 1 0 37628 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_842
timestamp 1586364061
transform 1 0 38180 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_404
timestamp 1586364061
transform 1 0 38272 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_416
timestamp 1586364061
transform 1 0 39376 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_428
timestamp 1586364061
transform 1 0 40480 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_843
timestamp 1586364061
transform 1 0 41032 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_435
timestamp 1586364061
transform 1 0 41124 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_447
timestamp 1586364061
transform 1 0 42228 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_844
timestamp 1586364061
transform 1 0 43884 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_459
timestamp 1586364061
transform 1 0 43332 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_466
timestamp 1586364061
transform 1 0 43976 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_478
timestamp 1586364061
transform 1 0 45080 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_845
timestamp 1586364061
transform 1 0 46736 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_490
timestamp 1586364061
transform 1 0 46184 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_497
timestamp 1586364061
transform 1 0 46828 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_509
timestamp 1586364061
transform 1 0 47932 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_3  PHY_165
timestamp 1586364061
transform -1 0 48852 0 -1 47328
box -38 -48 314 592
use scs8hd_fill_1  FILLER_82_515
timestamp 1586364061
transform 1 0 48484 0 -1 47328
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 3544 480 3664 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 10616 480 10736 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 17824 480 17944 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 24896 480 25016 6 address[3]
port 3 nsew default input
rlabel metal2 s 19430 0 19486 480 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 32104 480 32224 6 address[5]
port 5 nsew default input
rlabel metal2 s 24950 0 25006 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 30470 0 30526 480 6 address[7]
port 7 nsew default input
rlabel metal3 s 0 39176 480 39296 6 address[8]
port 8 nsew default input
rlabel metal2 s 36082 0 36138 480 6 address[9]
port 9 nsew default input
rlabel metal2 s 41602 0 41658 480 6 bottom_width_0_height_0__pin_10_
port 10 nsew default tristate
rlabel metal2 s 8298 49520 8354 50000 6 bottom_width_0_height_0__pin_14_
port 11 nsew default input
rlabel metal3 s 49520 24896 50000 25016 6 bottom_width_0_height_0__pin_2_
port 12 nsew default input
rlabel metal2 s 2778 49520 2834 50000 6 bottom_width_0_height_0__pin_6_
port 13 nsew default input
rlabel metal2 s 13818 0 13874 480 6 clk
port 14 nsew default input
rlabel metal3 s 49520 14832 50000 14952 6 data_in
port 15 nsew default input
rlabel metal3 s 49520 4904 50000 5024 6 enable
port 16 nsew default input
rlabel metal2 s 24950 49520 25006 50000 6 left_width_0_height_0__pin_11_
port 17 nsew default tristate
rlabel metal2 s 13818 49520 13874 50000 6 left_width_0_height_0__pin_3_
port 18 nsew default input
rlabel metal2 s 19430 49520 19486 50000 6 left_width_0_height_0__pin_7_
port 19 nsew default input
rlabel metal2 s 8298 0 8354 480 6 reset
port 20 nsew default input
rlabel metal3 s 0 46384 480 46504 6 right_width_0_height_0__pin_13_
port 21 nsew default tristate
rlabel metal2 s 30470 49520 30526 50000 6 right_width_0_height_0__pin_1_
port 22 nsew default input
rlabel metal2 s 36082 49520 36138 50000 6 right_width_0_height_0__pin_5_
port 23 nsew default input
rlabel metal2 s 41602 49520 41658 50000 6 right_width_0_height_0__pin_9_
port 24 nsew default input
rlabel metal2 s 2778 0 2834 480 6 set
port 25 nsew default input
rlabel metal3 s 49520 34824 50000 34944 6 top_width_0_height_0__pin_0_
port 26 nsew default input
rlabel metal2 s 47122 0 47178 480 6 top_width_0_height_0__pin_12_
port 27 nsew default tristate
rlabel metal2 s 47122 49520 47178 50000 6 top_width_0_height_0__pin_4_
port 28 nsew default input
rlabel metal3 s 49520 44888 50000 45008 6 top_width_0_height_0__pin_8_
port 29 nsew default input
rlabel metal4 s 4208 2128 4528 47376 6 vpwr
port 30 nsew default input
rlabel metal4 s 19568 2128 19888 47376 6 vgnd
port 31 nsew default input
<< end >>
