magic
tech EFS8A
magscale 1 2
timestamp 1602269239
<< locali >>
rect 10793 23137 10954 23171
rect 10793 22967 10827 23137
rect 21511 18921 21649 18955
rect 1443 18785 1478 18819
rect 12167 17833 12173 17867
rect 12167 17765 12201 17833
rect 21005 17697 21166 17731
rect 21005 17663 21039 17697
rect 16951 16745 16957 16779
rect 16951 16677 16985 16745
rect 14197 15963 14231 16201
rect 13363 14569 13369 14603
rect 16031 14569 16037 14603
rect 17779 14569 17785 14603
rect 21275 14569 21281 14603
rect 13363 14501 13397 14569
rect 16031 14501 16065 14569
rect 17779 14501 17813 14569
rect 21275 14501 21309 14569
rect 9597 13855 9631 14025
rect 5491 13345 5526 13379
rect 16307 12631 16341 12699
rect 16307 12597 16313 12631
rect 10051 12393 10057 12427
rect 13639 12393 13645 12427
rect 10051 12325 10085 12393
rect 13639 12325 13673 12393
rect 19475 12257 19510 12291
rect 22017 12155 22051 12325
rect 23615 11645 23742 11679
rect 4203 11169 4330 11203
rect 8435 11169 8470 11203
rect 6831 10217 6837 10251
rect 6831 10149 6865 10217
rect 9229 9435 9263 9605
rect 21275 9129 21281 9163
rect 21275 9061 21309 9129
rect 7291 7191 7325 7259
rect 13369 7191 13403 7497
rect 7291 7157 7297 7191
rect 18147 6953 18153 6987
rect 18147 6885 18181 6953
rect 8159 6817 8194 6851
rect 25179 6817 25214 6851
rect 4479 5729 4514 5763
rect 20815 5015 20849 5083
rect 20815 4981 20821 5015
rect 7239 4709 7284 4743
rect 18429 4539 18463 4709
rect 13737 4131 13771 4233
rect 8493 3995 8527 4097
rect 22511 3553 22546 3587
rect 6009 2839 6043 2941
rect 10971 2839 11005 2907
rect 10971 2805 10977 2839
rect 4399 2601 4537 2635
rect 17877 2295 17911 2397
<< viali >>
rect 22820 24225 22854 24259
rect 22891 24021 22925 24055
rect 7021 23817 7055 23851
rect 21925 23817 21959 23851
rect 22845 23817 22879 23851
rect 24225 23817 24259 23851
rect 25237 23817 25271 23851
rect 24823 23749 24857 23783
rect 6837 23613 6871 23647
rect 7389 23613 7423 23647
rect 9204 23613 9238 23647
rect 9597 23613 9631 23647
rect 10333 23613 10367 23647
rect 10885 23613 10919 23647
rect 21741 23613 21775 23647
rect 22293 23613 22327 23647
rect 23724 23613 23758 23647
rect 24752 23613 24786 23647
rect 23811 23545 23845 23579
rect 9275 23477 9309 23511
rect 10517 23477 10551 23511
rect 11023 23273 11057 23307
rect 22820 23137 22854 23171
rect 10793 22933 10827 22967
rect 22891 22933 22925 22967
rect 22845 22729 22879 22763
rect 25145 22729 25179 22763
rect 1409 22525 1443 22559
rect 1961 22525 1995 22559
rect 24644 22525 24678 22559
rect 24731 22457 24765 22491
rect 1593 22389 1627 22423
rect 10977 22389 11011 22423
rect 1593 21641 1627 21675
rect 1409 21437 1443 21471
rect 2053 21301 2087 21335
rect 19809 21097 19843 21131
rect 19625 20961 19659 20995
rect 18751 20485 18785 20519
rect 19625 20485 19659 20519
rect 18680 20349 18714 20383
rect 19073 20349 19107 20383
rect 12608 19873 12642 19907
rect 15336 19873 15370 19907
rect 14013 19805 14047 19839
rect 12679 19669 12713 19703
rect 15439 19669 15473 19703
rect 16037 19669 16071 19703
rect 1593 19465 1627 19499
rect 12265 19465 12299 19499
rect 13737 19465 13771 19499
rect 1409 19261 1443 19295
rect 12817 19261 12851 19295
rect 14968 19261 15002 19295
rect 15393 19261 15427 19295
rect 15945 19261 15979 19295
rect 16497 19261 16531 19295
rect 13461 19193 13495 19227
rect 15761 19193 15795 19227
rect 16681 19193 16715 19227
rect 2053 19125 2087 19159
rect 14749 19125 14783 19159
rect 15071 19125 15105 19159
rect 9965 18921 9999 18955
rect 12817 18921 12851 18955
rect 14197 18921 14231 18955
rect 21649 18921 21683 18955
rect 24777 18921 24811 18955
rect 11805 18853 11839 18887
rect 13277 18853 13311 18887
rect 13369 18853 13403 18887
rect 17049 18853 17083 18887
rect 17141 18853 17175 18887
rect 1409 18785 1443 18819
rect 7849 18785 7883 18819
rect 9781 18785 9815 18819
rect 15393 18785 15427 18819
rect 15853 18785 15887 18819
rect 21440 18785 21474 18819
rect 24593 18785 24627 18819
rect 11713 18717 11747 18751
rect 11989 18717 12023 18751
rect 13737 18717 13771 18751
rect 16129 18717 16163 18751
rect 17693 18717 17727 18751
rect 8033 18649 8067 18683
rect 16773 18649 16807 18683
rect 1547 18581 1581 18615
rect 16405 18581 16439 18615
rect 18061 18581 18095 18615
rect 21925 18581 21959 18615
rect 1869 18377 1903 18411
rect 7941 18377 7975 18411
rect 11805 18377 11839 18411
rect 13645 18377 13679 18411
rect 2237 18241 2271 18275
rect 14289 18241 14323 18275
rect 14565 18241 14599 18275
rect 16221 18241 16255 18275
rect 24593 18241 24627 18275
rect 1460 18173 1494 18207
rect 1547 18173 1581 18207
rect 9648 18173 9682 18207
rect 11396 18173 11430 18207
rect 17877 18173 17911 18207
rect 18061 18173 18095 18207
rect 18521 18173 18555 18207
rect 9735 18105 9769 18139
rect 11483 18105 11517 18139
rect 12725 18105 12759 18139
rect 12817 18105 12851 18139
rect 13369 18105 13403 18139
rect 14105 18105 14139 18139
rect 14381 18105 14415 18139
rect 16313 18105 16347 18139
rect 16865 18105 16899 18139
rect 21373 18105 21407 18139
rect 21925 18105 21959 18139
rect 22017 18105 22051 18139
rect 22569 18105 22603 18139
rect 10057 18037 10091 18071
rect 10517 18037 10551 18071
rect 11161 18037 11195 18071
rect 12265 18037 12299 18071
rect 15393 18037 15427 18071
rect 15853 18037 15887 18071
rect 17141 18037 17175 18071
rect 18153 18037 18187 18071
rect 21649 18037 21683 18071
rect 12173 17833 12207 17867
rect 12725 17833 12759 17867
rect 15945 17833 15979 17867
rect 17233 17833 17267 17867
rect 22109 17833 22143 17867
rect 24777 17833 24811 17867
rect 10333 17765 10367 17799
rect 10425 17765 10459 17799
rect 10977 17765 11011 17799
rect 13829 17765 13863 17799
rect 14381 17765 14415 17799
rect 16313 17765 16347 17799
rect 17877 17765 17911 17799
rect 18429 17765 18463 17799
rect 22569 17765 22603 17799
rect 22661 17765 22695 17799
rect 11713 17697 11747 17731
rect 13369 17697 13403 17731
rect 24593 17697 24627 17731
rect 11805 17629 11839 17663
rect 13737 17629 13771 17663
rect 16221 17629 16255 17663
rect 16865 17629 16899 17663
rect 17785 17629 17819 17663
rect 21005 17629 21039 17663
rect 22845 17629 22879 17663
rect 11253 17493 11287 17527
rect 13001 17493 13035 17527
rect 21235 17493 21269 17527
rect 9597 17289 9631 17323
rect 19073 17289 19107 17323
rect 23029 17289 23063 17323
rect 21097 17221 21131 17255
rect 9919 17153 9953 17187
rect 10885 17153 10919 17187
rect 14381 17153 14415 17187
rect 16313 17153 16347 17187
rect 16957 17153 16991 17187
rect 18429 17153 18463 17187
rect 20545 17153 20579 17187
rect 21465 17153 21499 17187
rect 22109 17153 22143 17187
rect 22385 17153 22419 17187
rect 24731 17153 24765 17187
rect 9832 17085 9866 17119
rect 12633 17085 12667 17119
rect 13553 17085 13587 17119
rect 13921 17085 13955 17119
rect 14289 17085 14323 17119
rect 14473 17085 14507 17119
rect 24644 17085 24678 17119
rect 25421 17085 25455 17119
rect 10977 17017 11011 17051
rect 11529 17017 11563 17051
rect 11897 17017 11931 17051
rect 12265 17017 12299 17051
rect 12995 17017 13029 17051
rect 16129 17017 16163 17051
rect 16405 17017 16439 17051
rect 18153 17017 18187 17051
rect 18245 17017 18279 17051
rect 20361 17017 20395 17051
rect 20637 17017 20671 17051
rect 22201 17017 22235 17051
rect 10241 16949 10275 16983
rect 10701 16949 10735 16983
rect 15761 16949 15795 16983
rect 17417 16949 17451 16983
rect 17785 16949 17819 16983
rect 21925 16949 21959 16983
rect 25053 16949 25087 16983
rect 13737 16745 13771 16779
rect 15669 16745 15703 16779
rect 16129 16745 16163 16779
rect 16957 16745 16991 16779
rect 17509 16745 17543 16779
rect 18429 16745 18463 16779
rect 20545 16745 20579 16779
rect 22477 16745 22511 16779
rect 10609 16677 10643 16711
rect 12909 16677 12943 16711
rect 21281 16677 21315 16711
rect 22753 16677 22787 16711
rect 22845 16677 22879 16711
rect 24409 16677 24443 16711
rect 24961 16677 24995 16711
rect 15485 16609 15519 16643
rect 16589 16609 16623 16643
rect 19073 16609 19107 16643
rect 19257 16609 19291 16643
rect 8585 16541 8619 16575
rect 10517 16541 10551 16575
rect 11161 16541 11195 16575
rect 12817 16541 12851 16575
rect 13461 16541 13495 16575
rect 19533 16541 19567 16575
rect 21189 16541 21223 16575
rect 23029 16541 23063 16575
rect 24317 16541 24351 16575
rect 21741 16473 21775 16507
rect 10241 16405 10275 16439
rect 11805 16405 11839 16439
rect 18153 16405 18187 16439
rect 22109 16405 22143 16439
rect 10149 16201 10183 16235
rect 13921 16201 13955 16235
rect 14197 16201 14231 16235
rect 15577 16201 15611 16235
rect 17417 16201 17451 16235
rect 20729 16201 20763 16235
rect 21097 16201 21131 16235
rect 23121 16201 23155 16235
rect 24685 16201 24719 16235
rect 11713 16133 11747 16167
rect 11069 16065 11103 16099
rect 9356 15997 9390 16031
rect 9781 15997 9815 16031
rect 12817 15997 12851 16031
rect 13185 15997 13219 16031
rect 13369 15997 13403 16031
rect 15117 16133 15151 16167
rect 15853 16133 15887 16167
rect 22845 16133 22879 16167
rect 14565 16065 14599 16099
rect 16405 16065 16439 16099
rect 19809 16065 19843 16099
rect 18061 15997 18095 16031
rect 18613 15997 18647 16031
rect 21557 15997 21591 16031
rect 9459 15929 9493 15963
rect 10425 15929 10459 15963
rect 10517 15929 10551 15963
rect 11437 15929 11471 15963
rect 14197 15929 14231 15963
rect 14657 15929 14691 15963
rect 16129 15929 16163 15963
rect 16221 15929 16255 15963
rect 20171 15929 20205 15963
rect 21878 15929 21912 15963
rect 12173 15861 12207 15895
rect 13185 15861 13219 15895
rect 14289 15861 14323 15895
rect 17049 15861 17083 15895
rect 17877 15861 17911 15895
rect 18153 15861 18187 15895
rect 19073 15861 19107 15895
rect 19717 15861 19751 15895
rect 21373 15861 21407 15895
rect 22477 15861 22511 15895
rect 24225 15861 24259 15895
rect 10057 15657 10091 15691
rect 12817 15657 12851 15691
rect 13829 15657 13863 15691
rect 14565 15657 14599 15691
rect 15393 15657 15427 15691
rect 19257 15657 19291 15691
rect 19809 15657 19843 15691
rect 21189 15657 21223 15691
rect 23121 15657 23155 15691
rect 8217 15589 8251 15623
rect 10425 15589 10459 15623
rect 13271 15589 13305 15623
rect 16726 15589 16760 15623
rect 18337 15589 18371 15623
rect 21741 15589 21775 15623
rect 11964 15521 11998 15555
rect 17325 15521 17359 15555
rect 8125 15453 8159 15487
rect 8401 15453 8435 15487
rect 10333 15453 10367 15487
rect 12909 15453 12943 15487
rect 16405 15453 16439 15487
rect 18245 15453 18279 15487
rect 18521 15453 18555 15487
rect 21649 15453 21683 15487
rect 22293 15453 22327 15487
rect 10885 15385 10919 15419
rect 15945 15385 15979 15419
rect 12035 15317 12069 15351
rect 16221 15317 16255 15351
rect 20453 15317 20487 15351
rect 7849 15113 7883 15147
rect 10701 15113 10735 15147
rect 11069 15113 11103 15147
rect 14105 15113 14139 15147
rect 15485 15113 15519 15147
rect 15853 15113 15887 15147
rect 17509 15113 17543 15147
rect 21649 15113 21683 15147
rect 22247 15113 22281 15147
rect 22661 15113 22695 15147
rect 17049 15045 17083 15079
rect 19073 15045 19107 15079
rect 8309 14977 8343 15011
rect 13185 14977 13219 15011
rect 14749 14977 14783 15011
rect 16497 14977 16531 15011
rect 18153 14977 18187 15011
rect 18429 14977 18463 15011
rect 21925 14977 21959 15011
rect 9505 14909 9539 14943
rect 10425 14909 10459 14943
rect 11396 14909 11430 14943
rect 11897 14909 11931 14943
rect 12265 14909 12299 14943
rect 15301 14909 15335 14943
rect 20361 14909 20395 14943
rect 22176 14909 22210 14943
rect 7113 14841 7147 14875
rect 8033 14841 8067 14875
rect 8125 14841 8159 14875
rect 9827 14841 9861 14875
rect 13506 14841 13540 14875
rect 16589 14841 16623 14875
rect 18245 14841 18279 14875
rect 20682 14841 20716 14875
rect 7481 14773 7515 14807
rect 8953 14773 8987 14807
rect 9413 14773 9447 14807
rect 11483 14773 11517 14807
rect 13001 14773 13035 14807
rect 14473 14773 14507 14807
rect 16221 14773 16255 14807
rect 17877 14773 17911 14807
rect 20269 14773 20303 14807
rect 21281 14773 21315 14807
rect 1593 14569 1627 14603
rect 10609 14569 10643 14603
rect 11529 14569 11563 14603
rect 12541 14569 12575 14603
rect 13369 14569 13403 14603
rect 13921 14569 13955 14603
rect 16037 14569 16071 14603
rect 16865 14569 16899 14603
rect 17233 14569 17267 14603
rect 17785 14569 17819 14603
rect 18337 14569 18371 14603
rect 21281 14569 21315 14603
rect 8769 14501 8803 14535
rect 10010 14501 10044 14535
rect 18613 14501 18647 14535
rect 19901 14501 19935 14535
rect 22845 14501 22879 14535
rect 1409 14433 1443 14467
rect 8125 14433 8159 14467
rect 8585 14433 8619 14467
rect 11437 14433 11471 14467
rect 11897 14433 11931 14467
rect 12817 14433 12851 14467
rect 15577 14433 15611 14467
rect 15669 14433 15703 14467
rect 19165 14433 19199 14467
rect 19625 14433 19659 14467
rect 9689 14365 9723 14399
rect 13001 14365 13035 14399
rect 17417 14365 17451 14399
rect 20913 14365 20947 14399
rect 22753 14365 22787 14399
rect 23029 14365 23063 14399
rect 7205 14229 7239 14263
rect 7941 14229 7975 14263
rect 16589 14229 16623 14263
rect 20177 14229 20211 14263
rect 21833 14229 21867 14263
rect 9597 14025 9631 14059
rect 9781 14025 9815 14059
rect 10057 14025 10091 14059
rect 12265 14025 12299 14059
rect 17785 14025 17819 14059
rect 21097 14025 21131 14059
rect 21833 14025 21867 14059
rect 23029 14025 23063 14059
rect 25421 14025 25455 14059
rect 7849 13889 7883 13923
rect 9413 13889 9447 13923
rect 11437 13957 11471 13991
rect 14289 13957 14323 13991
rect 23489 13957 23523 13991
rect 10241 13889 10275 13923
rect 13921 13889 13955 13923
rect 20177 13889 20211 13923
rect 22753 13889 22787 13923
rect 24041 13889 24075 13923
rect 8585 13821 8619 13855
rect 8769 13821 8803 13855
rect 9137 13821 9171 13855
rect 9597 13821 9631 13855
rect 11161 13821 11195 13855
rect 12725 13821 12759 13855
rect 13093 13821 13127 13855
rect 13277 13821 13311 13855
rect 14657 13821 14691 13855
rect 14841 13821 14875 13855
rect 16313 13821 16347 13855
rect 16681 13821 16715 13855
rect 16865 13821 16899 13855
rect 18429 13821 18463 13855
rect 18613 13821 18647 13855
rect 19165 13821 19199 13855
rect 19349 13821 19383 13855
rect 25237 13821 25271 13855
rect 25789 13821 25823 13855
rect 6653 13753 6687 13787
rect 7205 13753 7239 13787
rect 7297 13753 7331 13787
rect 10603 13753 10637 13787
rect 17141 13753 17175 13787
rect 20539 13753 20573 13787
rect 22109 13753 22143 13787
rect 22201 13753 22235 13787
rect 23765 13753 23799 13787
rect 23857 13753 23891 13787
rect 1685 13685 1719 13719
rect 8125 13685 8159 13719
rect 11805 13685 11839 13719
rect 12909 13685 12943 13719
rect 14473 13685 14507 13719
rect 15761 13685 15795 13719
rect 17417 13685 17451 13719
rect 19625 13685 19659 13719
rect 20085 13685 20119 13719
rect 21373 13685 21407 13719
rect 1593 13481 1627 13515
rect 5595 13481 5629 13515
rect 9413 13481 9447 13515
rect 10609 13481 10643 13515
rect 14381 13481 14415 13515
rect 19165 13481 19199 13515
rect 22569 13481 22603 13515
rect 9827 13413 9861 13447
rect 11345 13413 11379 13447
rect 17233 13413 17267 13447
rect 21234 13413 21268 13447
rect 22845 13413 22879 13447
rect 23397 13413 23431 13447
rect 1409 13345 1443 13379
rect 5457 13345 5491 13379
rect 7056 13345 7090 13379
rect 8309 13345 8343 13379
rect 8493 13345 8527 13379
rect 9724 13345 9758 13379
rect 13093 13345 13127 13379
rect 13369 13345 13403 13379
rect 15761 13345 15795 13379
rect 15945 13345 15979 13379
rect 18889 13345 18923 13379
rect 19349 13345 19383 13379
rect 19901 13345 19935 13379
rect 20913 13345 20947 13379
rect 24276 13345 24310 13379
rect 8769 13277 8803 13311
rect 11253 13277 11287 13311
rect 13461 13277 13495 13311
rect 16129 13277 16163 13311
rect 17141 13277 17175 13311
rect 17785 13277 17819 13311
rect 22753 13277 22787 13311
rect 24363 13277 24397 13311
rect 11805 13209 11839 13243
rect 21833 13209 21867 13243
rect 7159 13141 7193 13175
rect 7941 13141 7975 13175
rect 9137 13141 9171 13175
rect 10149 13141 10183 13175
rect 12725 13141 12759 13175
rect 16497 13141 16531 13175
rect 18613 13141 18647 13175
rect 20637 13141 20671 13175
rect 22201 13141 22235 13175
rect 23673 13141 23707 13175
rect 7067 12937 7101 12971
rect 7389 12937 7423 12971
rect 9045 12937 9079 12971
rect 10517 12937 10551 12971
rect 11897 12937 11931 12971
rect 13645 12937 13679 12971
rect 16865 12937 16899 12971
rect 17233 12937 17267 12971
rect 21833 12937 21867 12971
rect 22523 12937 22557 12971
rect 23213 12937 23247 12971
rect 23811 12937 23845 12971
rect 11207 12869 11241 12903
rect 15485 12869 15519 12903
rect 1685 12801 1719 12835
rect 9597 12801 9631 12835
rect 10057 12801 10091 12835
rect 12725 12801 12759 12835
rect 13001 12801 13035 12835
rect 14565 12801 14599 12835
rect 18429 12801 18463 12835
rect 24823 12801 24857 12835
rect 6653 12733 6687 12767
rect 6964 12733 6998 12767
rect 7849 12733 7883 12767
rect 8217 12733 8251 12767
rect 8401 12733 8435 12767
rect 9321 12733 9355 12767
rect 11136 12733 11170 12767
rect 15945 12733 15979 12767
rect 18981 12733 19015 12767
rect 19441 12733 19475 12767
rect 19717 12733 19751 12767
rect 22452 12733 22486 12767
rect 23740 12733 23774 12767
rect 24736 12733 24770 12767
rect 25145 12733 25179 12767
rect 5549 12665 5583 12699
rect 8677 12665 8711 12699
rect 9689 12665 9723 12699
rect 12817 12665 12851 12699
rect 14289 12665 14323 12699
rect 14381 12665 14415 12699
rect 20913 12665 20947 12699
rect 21005 12665 21039 12699
rect 21557 12665 21591 12699
rect 24225 12665 24259 12699
rect 5733 12597 5767 12631
rect 10885 12597 10919 12631
rect 11621 12597 11655 12631
rect 14105 12597 14139 12631
rect 15853 12597 15887 12631
rect 16313 12597 16347 12631
rect 17601 12597 17635 12631
rect 18797 12597 18831 12631
rect 20361 12597 20395 12631
rect 20637 12597 20671 12631
rect 22201 12597 22235 12631
rect 22937 12597 22971 12631
rect 24593 12597 24627 12631
rect 8677 12393 8711 12427
rect 9413 12393 9447 12427
rect 10057 12393 10091 12427
rect 10609 12393 10643 12427
rect 12541 12393 12575 12427
rect 13645 12393 13679 12427
rect 15577 12393 15611 12427
rect 17049 12393 17083 12427
rect 19579 12393 19613 12427
rect 22201 12393 22235 12427
rect 22661 12393 22695 12427
rect 22845 12393 22879 12427
rect 6285 12325 6319 12359
rect 7849 12325 7883 12359
rect 11621 12325 11655 12359
rect 16450 12325 16484 12359
rect 18061 12325 18095 12359
rect 18889 12325 18923 12359
rect 19257 12325 19291 12359
rect 21373 12325 21407 12359
rect 22017 12325 22051 12359
rect 1444 12257 1478 12291
rect 16129 12257 16163 12291
rect 19441 12257 19475 12291
rect 6193 12189 6227 12223
rect 6837 12189 6871 12223
rect 7113 12189 7147 12223
rect 7757 12189 7791 12223
rect 9689 12189 9723 12223
rect 11529 12189 11563 12223
rect 13277 12189 13311 12223
rect 17969 12189 18003 12223
rect 18245 12189 18279 12223
rect 21281 12189 21315 12223
rect 21925 12189 21959 12223
rect 22753 12257 22787 12291
rect 23213 12257 23247 12291
rect 24384 12257 24418 12291
rect 8309 12121 8343 12155
rect 12081 12121 12115 12155
rect 16037 12121 16071 12155
rect 22017 12121 22051 12155
rect 24455 12121 24489 12155
rect 1547 12053 1581 12087
rect 12909 12053 12943 12087
rect 14197 12053 14231 12087
rect 14473 12053 14507 12087
rect 19993 12053 20027 12087
rect 23765 12053 23799 12087
rect 1593 11849 1627 11883
rect 7849 11849 7883 11883
rect 8217 11849 8251 11883
rect 8953 11849 8987 11883
rect 10977 11849 11011 11883
rect 11437 11849 11471 11883
rect 11805 11849 11839 11883
rect 14197 11849 14231 11883
rect 17785 11849 17819 11883
rect 23811 11849 23845 11883
rect 15485 11781 15519 11815
rect 19533 11781 19567 11815
rect 24409 11781 24443 11815
rect 25237 11781 25271 11815
rect 7205 11713 7239 11747
rect 9781 11713 9815 11747
rect 13277 11713 13311 11747
rect 14473 11713 14507 11747
rect 17141 11713 17175 11747
rect 21833 11713 21867 11747
rect 22201 11713 22235 11747
rect 22753 11713 22787 11747
rect 23121 11713 23155 11747
rect 5089 11645 5123 11679
rect 5825 11645 5859 11679
rect 8468 11645 8502 11679
rect 12817 11645 12851 11679
rect 15301 11645 15335 11679
rect 15853 11645 15887 11679
rect 18337 11645 18371 11679
rect 18429 11645 18463 11679
rect 18889 11645 18923 11679
rect 19993 11645 20027 11679
rect 20913 11645 20947 11679
rect 21557 11645 21591 11679
rect 23581 11645 23615 11679
rect 24752 11645 24786 11679
rect 5917 11577 5951 11611
rect 6193 11577 6227 11611
rect 6929 11577 6963 11611
rect 7021 11577 7055 11611
rect 10102 11577 10136 11611
rect 13185 11577 13219 11611
rect 13639 11577 13673 11611
rect 16497 11577 16531 11611
rect 16589 11577 16623 11611
rect 19165 11577 19199 11611
rect 20314 11577 20348 11611
rect 21925 11577 21959 11611
rect 6561 11509 6595 11543
rect 8539 11509 8573 11543
rect 9321 11509 9355 11543
rect 9597 11509 9631 11543
rect 10701 11509 10735 11543
rect 16313 11509 16347 11543
rect 17417 11509 17451 11543
rect 19809 11509 19843 11543
rect 21189 11509 21223 11543
rect 24823 11509 24857 11543
rect 6285 11305 6319 11339
rect 8539 11305 8573 11339
rect 10103 11305 10137 11339
rect 13277 11305 13311 11339
rect 16313 11305 16347 11339
rect 16773 11305 16807 11339
rect 19993 11305 20027 11339
rect 5457 11237 5491 11271
rect 6009 11237 6043 11271
rect 7021 11237 7055 11271
rect 10425 11237 10459 11271
rect 11161 11237 11195 11271
rect 11713 11237 11747 11271
rect 13553 11237 13587 11271
rect 13645 11237 13679 11271
rect 14197 11237 14231 11271
rect 15485 11237 15519 11271
rect 17049 11237 17083 11271
rect 19394 11237 19428 11271
rect 22017 11237 22051 11271
rect 23581 11237 23615 11271
rect 4169 11169 4203 11203
rect 8401 11169 8435 11203
rect 10032 11169 10066 11203
rect 17509 11169 17543 11203
rect 18061 11169 18095 11203
rect 4399 11101 4433 11135
rect 5365 11101 5399 11135
rect 6929 11101 6963 11135
rect 7205 11101 7239 11135
rect 11069 11101 11103 11135
rect 15393 11101 15427 11135
rect 15669 11101 15703 11135
rect 18245 11101 18279 11135
rect 19073 11101 19107 11135
rect 21925 11101 21959 11135
rect 22201 11101 22235 11135
rect 23478 11101 23512 11135
rect 23765 11101 23799 11135
rect 13001 10965 13035 10999
rect 18521 10965 18555 10999
rect 21281 10965 21315 10999
rect 21649 10965 21683 10999
rect 4261 10761 4295 10795
rect 4721 10761 4755 10795
rect 5089 10761 5123 10795
rect 6561 10761 6595 10795
rect 7941 10761 7975 10795
rect 11299 10761 11333 10795
rect 12173 10761 12207 10795
rect 12587 10761 12621 10795
rect 16405 10761 16439 10795
rect 16727 10761 16761 10795
rect 17509 10761 17543 10795
rect 20821 10761 20855 10795
rect 21189 10761 21223 10795
rect 22845 10761 22879 10795
rect 23489 10761 23523 10795
rect 24593 10761 24627 10795
rect 7481 10693 7515 10727
rect 13277 10693 13311 10727
rect 16037 10693 16071 10727
rect 5917 10625 5951 10659
rect 6929 10625 6963 10659
rect 8493 10625 8527 10659
rect 13553 10625 13587 10659
rect 15577 10625 15611 10659
rect 18797 10625 18831 10659
rect 19901 10625 19935 10659
rect 5825 10557 5859 10591
rect 11228 10557 11262 10591
rect 11713 10557 11747 10591
rect 12516 10557 12550 10591
rect 15025 10557 15059 10591
rect 15485 10557 15519 10591
rect 16656 10557 16690 10591
rect 21649 10557 21683 10591
rect 23724 10557 23758 10591
rect 7021 10489 7055 10523
rect 9689 10489 9723 10523
rect 9781 10489 9815 10523
rect 10333 10489 10367 10523
rect 13645 10489 13679 10523
rect 14197 10489 14231 10523
rect 14933 10489 14967 10523
rect 18153 10489 18187 10523
rect 18245 10489 18279 10523
rect 20263 10489 20297 10523
rect 21970 10489 22004 10523
rect 23811 10489 23845 10523
rect 24225 10489 24259 10523
rect 6285 10421 6319 10455
rect 9045 10421 9079 10455
rect 9505 10421 9539 10455
rect 10701 10421 10735 10455
rect 11069 10421 11103 10455
rect 13001 10421 13035 10455
rect 14473 10421 14507 10455
rect 17141 10421 17175 10455
rect 17877 10421 17911 10455
rect 19165 10421 19199 10455
rect 19717 10421 19751 10455
rect 21465 10421 21499 10455
rect 22569 10421 22603 10455
rect 5273 10217 5307 10251
rect 6837 10217 6871 10251
rect 7665 10217 7699 10251
rect 8585 10217 8619 10251
rect 11069 10217 11103 10251
rect 12449 10217 12483 10251
rect 13829 10217 13863 10251
rect 15117 10217 15151 10251
rect 19809 10217 19843 10251
rect 20177 10217 20211 10251
rect 9873 10149 9907 10183
rect 11345 10149 11379 10183
rect 11437 10149 11471 10183
rect 13271 10149 13305 10183
rect 16037 10149 16071 10183
rect 17049 10149 17083 10183
rect 19533 10149 19567 10183
rect 21649 10149 21683 10183
rect 7389 10081 7423 10115
rect 14289 10081 14323 10115
rect 15301 10081 15335 10115
rect 15577 10081 15611 10115
rect 19073 10081 19107 10115
rect 19257 10081 19291 10115
rect 22201 10081 22235 10115
rect 23121 10081 23155 10115
rect 6469 10013 6503 10047
rect 9781 10013 9815 10047
rect 10057 10013 10091 10047
rect 11621 10013 11655 10047
rect 12909 10013 12943 10047
rect 16957 10013 16991 10047
rect 17601 10013 17635 10047
rect 21557 10013 21591 10047
rect 23029 10013 23063 10047
rect 15393 9945 15427 9979
rect 18245 9945 18279 9979
rect 14565 9877 14599 9911
rect 17969 9877 18003 9911
rect 7757 9673 7791 9707
rect 9045 9673 9079 9707
rect 10425 9673 10459 9707
rect 11161 9673 11195 9707
rect 11805 9673 11839 9707
rect 12173 9673 12207 9707
rect 13461 9673 13495 9707
rect 16313 9673 16347 9707
rect 16635 9673 16669 9707
rect 21649 9673 21683 9707
rect 22247 9673 22281 9707
rect 22661 9673 22695 9707
rect 23121 9673 23155 9707
rect 9229 9605 9263 9639
rect 9321 9605 9355 9639
rect 10701 9605 10735 9639
rect 24731 9605 24765 9639
rect 6837 9469 6871 9503
rect 8677 9469 8711 9503
rect 11345 9537 11379 9571
rect 18153 9537 18187 9571
rect 18797 9537 18831 9571
rect 9505 9469 9539 9503
rect 12449 9469 12483 9503
rect 13001 9469 13035 9503
rect 14473 9469 14507 9503
rect 14933 9469 14967 9503
rect 15209 9469 15243 9503
rect 15393 9469 15427 9503
rect 16564 9469 16598 9503
rect 22176 9469 22210 9503
rect 24660 9469 24694 9503
rect 6285 9401 6319 9435
rect 6653 9401 6687 9435
rect 7199 9401 7233 9435
rect 9229 9401 9263 9435
rect 9826 9401 9860 9435
rect 14105 9401 14139 9435
rect 15669 9401 15703 9435
rect 17877 9401 17911 9435
rect 18245 9401 18279 9435
rect 20637 9401 20671 9435
rect 20729 9401 20763 9435
rect 21281 9401 21315 9435
rect 5917 9333 5951 9367
rect 8125 9333 8159 9367
rect 12541 9333 12575 9367
rect 15945 9333 15979 9367
rect 17049 9333 17083 9367
rect 17325 9333 17359 9367
rect 19073 9333 19107 9367
rect 19441 9333 19475 9367
rect 20453 9333 20487 9367
rect 22017 9333 22051 9367
rect 25145 9333 25179 9367
rect 6745 9129 6779 9163
rect 11161 9129 11195 9163
rect 12909 9129 12943 9163
rect 13277 9129 13311 9163
rect 14289 9129 14323 9163
rect 15485 9129 15519 9163
rect 16589 9129 16623 9163
rect 21281 9129 21315 9163
rect 5825 9061 5859 9095
rect 14933 9061 14967 9095
rect 16031 9061 16065 9095
rect 17601 9061 17635 9095
rect 22845 9061 22879 9095
rect 24409 9061 24443 9095
rect 5089 8993 5123 9027
rect 5365 8993 5399 9027
rect 6193 8993 6227 9027
rect 6837 8993 6871 9027
rect 7389 8993 7423 9027
rect 7665 8993 7699 9027
rect 8033 8993 8067 9027
rect 9908 8993 9942 9027
rect 11161 8993 11195 9027
rect 11621 8993 11655 9027
rect 11897 8993 11931 9027
rect 12265 8993 12299 9027
rect 13369 8993 13403 9027
rect 13645 8993 13679 9027
rect 15669 8993 15703 9027
rect 19073 8993 19107 9027
rect 19441 8993 19475 9027
rect 21833 8993 21867 9027
rect 6561 8925 6595 8959
rect 10011 8925 10045 8959
rect 16865 8925 16899 8959
rect 17509 8925 17543 8959
rect 17785 8925 17819 8959
rect 18429 8925 18463 8959
rect 19717 8925 19751 8959
rect 19993 8925 20027 8959
rect 20913 8925 20947 8959
rect 22753 8925 22787 8959
rect 23029 8925 23063 8959
rect 24317 8925 24351 8959
rect 24593 8925 24627 8959
rect 5181 8857 5215 8891
rect 8493 8857 8527 8891
rect 10425 8857 10459 8891
rect 17325 8857 17359 8891
rect 9413 8789 9447 8823
rect 10701 8789 10735 8823
rect 14657 8789 14691 8823
rect 20545 8789 20579 8823
rect 5825 8585 5859 8619
rect 9229 8585 9263 8619
rect 13553 8585 13587 8619
rect 16313 8585 16347 8619
rect 16957 8585 16991 8619
rect 23029 8585 23063 8619
rect 23397 8585 23431 8619
rect 5181 8517 5215 8551
rect 8309 8517 8343 8551
rect 9505 8517 9539 8551
rect 10977 8517 11011 8551
rect 16635 8517 16669 8551
rect 17785 8517 17819 8551
rect 20637 8517 20671 8551
rect 9873 8449 9907 8483
rect 14105 8449 14139 8483
rect 18889 8449 18923 8483
rect 19717 8449 19751 8483
rect 21833 8449 21867 8483
rect 22753 8449 22787 8483
rect 6929 8381 6963 8415
rect 7389 8381 7423 8415
rect 7941 8381 7975 8415
rect 8125 8381 8159 8415
rect 9413 8381 9447 8415
rect 9689 8381 9723 8415
rect 12265 8381 12299 8415
rect 12633 8381 12667 8415
rect 14381 8381 14415 8415
rect 14657 8381 14691 8415
rect 15117 8381 15151 8415
rect 15393 8381 15427 8415
rect 16564 8381 16598 8415
rect 18153 8381 18187 8415
rect 18705 8381 18739 8415
rect 23673 8381 23707 8415
rect 24317 8381 24351 8415
rect 24844 8381 24878 8415
rect 25237 8381 25271 8415
rect 11345 8313 11379 8347
rect 13277 8313 13311 8347
rect 17417 8313 17451 8347
rect 19533 8313 19567 8347
rect 20038 8313 20072 8347
rect 20913 8313 20947 8347
rect 21557 8313 21591 8347
rect 21649 8313 21683 8347
rect 24593 8313 24627 8347
rect 5549 8245 5583 8279
rect 6285 8245 6319 8279
rect 6653 8245 6687 8279
rect 8677 8245 8711 8279
rect 10609 8245 10643 8279
rect 11897 8245 11931 8279
rect 15393 8245 15427 8279
rect 16037 8245 16071 8279
rect 19257 8245 19291 8279
rect 21281 8245 21315 8279
rect 23857 8245 23891 8279
rect 24915 8245 24949 8279
rect 1593 8041 1627 8075
rect 6929 8041 6963 8075
rect 12449 8041 12483 8075
rect 15117 8041 15151 8075
rect 21557 8041 21591 8075
rect 24455 8041 24489 8075
rect 6745 7973 6779 8007
rect 10425 7973 10459 8007
rect 13185 7973 13219 8007
rect 14381 7973 14415 8007
rect 15939 7973 15973 8007
rect 19901 7973 19935 8007
rect 21097 7973 21131 8007
rect 21925 7973 21959 8007
rect 5892 7905 5926 7939
rect 6837 7905 6871 7939
rect 7389 7905 7423 7939
rect 7665 7905 7699 7939
rect 8217 7905 8251 7939
rect 9689 7905 9723 7939
rect 9935 7905 9969 7939
rect 11529 7905 11563 7939
rect 11897 7905 11931 7939
rect 12081 7905 12115 7939
rect 12633 7905 12667 7939
rect 13921 7905 13955 7939
rect 15577 7905 15611 7939
rect 17325 7905 17359 7939
rect 17785 7905 17819 7939
rect 19165 7905 19199 7939
rect 19625 7905 19659 7939
rect 23340 7905 23374 7939
rect 24384 7905 24418 7939
rect 6377 7837 6411 7871
rect 17877 7837 17911 7871
rect 21833 7837 21867 7871
rect 22109 7837 22143 7871
rect 9137 7769 9171 7803
rect 9781 7769 9815 7803
rect 14657 7769 14691 7803
rect 18337 7769 18371 7803
rect 18981 7769 19015 7803
rect 24133 7769 24167 7803
rect 5963 7701 5997 7735
rect 9413 7701 9447 7735
rect 10885 7701 10919 7735
rect 16497 7701 16531 7735
rect 20269 7701 20303 7735
rect 22845 7701 22879 7735
rect 23443 7701 23477 7735
rect 23857 7701 23891 7735
rect 5917 7497 5951 7531
rect 8125 7497 8159 7531
rect 11621 7497 11655 7531
rect 13369 7497 13403 7531
rect 13921 7497 13955 7531
rect 14657 7497 14691 7531
rect 16313 7497 16347 7531
rect 19349 7497 19383 7531
rect 21465 7497 21499 7531
rect 22569 7497 22603 7531
rect 23029 7497 23063 7531
rect 25789 7497 25823 7531
rect 6929 7361 6963 7395
rect 10333 7361 10367 7395
rect 11897 7361 11931 7395
rect 12541 7361 12575 7395
rect 12817 7361 12851 7395
rect 4972 7293 5006 7327
rect 5365 7293 5399 7327
rect 6653 7293 6687 7327
rect 8677 7293 8711 7327
rect 9413 7293 9447 7327
rect 9505 7293 9539 7327
rect 10149 7225 10183 7259
rect 10654 7225 10688 7259
rect 12633 7225 12667 7259
rect 15301 7429 15335 7463
rect 17785 7429 17819 7463
rect 22201 7429 22235 7463
rect 16589 7361 16623 7395
rect 18705 7361 18739 7395
rect 21649 7361 21683 7395
rect 23489 7361 23523 7395
rect 23765 7361 23799 7395
rect 24133 7361 24167 7395
rect 14248 7293 14282 7327
rect 15209 7293 15243 7327
rect 15485 7293 15519 7327
rect 15945 7293 15979 7327
rect 16900 7293 16934 7327
rect 17325 7293 17359 7327
rect 19993 7293 20027 7327
rect 20361 7293 20395 7327
rect 20637 7293 20671 7327
rect 23673 7293 23707 7327
rect 23949 7293 23983 7327
rect 25304 7293 25338 7327
rect 13461 7225 13495 7259
rect 14335 7225 14369 7259
rect 18429 7225 18463 7259
rect 18521 7225 18555 7259
rect 20913 7225 20947 7259
rect 21741 7225 21775 7259
rect 5043 7157 5077 7191
rect 6285 7157 6319 7191
rect 7297 7157 7331 7191
rect 7849 7157 7883 7191
rect 9873 7157 9907 7191
rect 11253 7157 11287 7191
rect 13369 7157 13403 7191
rect 15117 7157 15151 7191
rect 17003 7157 17037 7191
rect 19809 7157 19843 7191
rect 24685 7157 24719 7191
rect 25375 7157 25409 7191
rect 1593 6953 1627 6987
rect 6101 6953 6135 6987
rect 9137 6953 9171 6987
rect 10885 6953 10919 6987
rect 11897 6953 11931 6987
rect 13461 6953 13495 6987
rect 16865 6953 16899 6987
rect 17417 6953 17451 6987
rect 18153 6953 18187 6987
rect 19533 6953 19567 6987
rect 20729 6953 20763 6987
rect 21005 6953 21039 6987
rect 25283 6953 25317 6987
rect 5089 6885 5123 6919
rect 5181 6885 5215 6919
rect 6745 6885 6779 6919
rect 9413 6885 9447 6919
rect 12173 6885 12207 6919
rect 13001 6885 13035 6919
rect 14381 6885 14415 6919
rect 16129 6885 16163 6919
rect 19165 6885 19199 6919
rect 22201 6885 22235 6919
rect 23765 6885 23799 6919
rect 1409 6817 1443 6851
rect 8125 6817 8159 6851
rect 9689 6817 9723 6851
rect 10425 6817 10459 6851
rect 10701 6817 10735 6851
rect 10977 6817 11011 6851
rect 13645 6817 13679 6851
rect 13921 6817 13955 6851
rect 15393 6817 15427 6851
rect 15669 6817 15703 6851
rect 17785 6817 17819 6851
rect 19844 6817 19878 6851
rect 25145 6817 25179 6851
rect 5733 6749 5767 6783
rect 6653 6749 6687 6783
rect 12081 6749 12115 6783
rect 12725 6749 12759 6783
rect 15117 6749 15151 6783
rect 15485 6749 15519 6783
rect 22109 6749 22143 6783
rect 22385 6749 22419 6783
rect 23673 6749 23707 6783
rect 23949 6749 23983 6783
rect 7205 6681 7239 6715
rect 7941 6681 7975 6715
rect 13737 6681 13771 6715
rect 16497 6681 16531 6715
rect 4905 6613 4939 6647
rect 6469 6613 6503 6647
rect 7573 6613 7607 6647
rect 8263 6613 8297 6647
rect 11529 6613 11563 6647
rect 18705 6613 18739 6647
rect 19947 6613 19981 6647
rect 21649 6613 21683 6647
rect 1823 6409 1857 6443
rect 4077 6409 4111 6443
rect 5089 6409 5123 6443
rect 6653 6409 6687 6443
rect 16129 6409 16163 6443
rect 24777 6409 24811 6443
rect 25237 6409 25271 6443
rect 4721 6341 4755 6375
rect 9229 6341 9263 6375
rect 15761 6341 15795 6375
rect 20729 6341 20763 6375
rect 22569 6341 22603 6375
rect 4307 6273 4341 6307
rect 5273 6273 5307 6307
rect 7481 6273 7515 6307
rect 12817 6273 12851 6307
rect 14381 6273 14415 6307
rect 16497 6273 16531 6307
rect 21649 6273 21683 6307
rect 1752 6205 1786 6239
rect 4220 6205 4254 6239
rect 9965 6205 9999 6239
rect 10333 6205 10367 6239
rect 10609 6205 10643 6239
rect 11069 6205 11103 6239
rect 18061 6205 18095 6239
rect 19809 6205 19843 6239
rect 5365 6137 5399 6171
rect 5917 6137 5951 6171
rect 7205 6137 7239 6171
rect 7297 6137 7331 6171
rect 8677 6137 8711 6171
rect 9597 6137 9631 6171
rect 11897 6137 11931 6171
rect 12541 6137 12575 6171
rect 12633 6137 12667 6171
rect 14094 6137 14128 6171
rect 14197 6137 14231 6171
rect 15025 6137 15059 6171
rect 16589 6137 16623 6171
rect 17141 6137 17175 6171
rect 18382 6137 18416 6171
rect 19257 6137 19291 6171
rect 20130 6137 20164 6171
rect 21741 6137 21775 6171
rect 22293 6137 22327 6171
rect 23765 6137 23799 6171
rect 23857 6137 23891 6171
rect 24409 6137 24443 6171
rect 2237 6069 2271 6103
rect 6193 6069 6227 6103
rect 8217 6069 8251 6103
rect 8585 6069 8619 6103
rect 9965 6069 9999 6103
rect 11437 6069 11471 6103
rect 12173 6069 12207 6103
rect 13737 6069 13771 6103
rect 15393 6069 15427 6103
rect 17417 6069 17451 6103
rect 17785 6069 17819 6103
rect 18981 6069 19015 6103
rect 19625 6069 19659 6103
rect 21465 6069 21499 6103
rect 23121 6069 23155 6103
rect 23397 6069 23431 6103
rect 1961 5865 1995 5899
rect 6653 5865 6687 5899
rect 8125 5865 8159 5899
rect 9137 5865 9171 5899
rect 9965 5865 9999 5899
rect 11529 5865 11563 5899
rect 13001 5865 13035 5899
rect 17049 5865 17083 5899
rect 21833 5865 21867 5899
rect 22109 5865 22143 5899
rect 24041 5865 24075 5899
rect 6193 5797 6227 5831
rect 7205 5797 7239 5831
rect 9505 5797 9539 5831
rect 10562 5797 10596 5831
rect 12173 5797 12207 5831
rect 13553 5797 13587 5831
rect 16681 5797 16715 5831
rect 17871 5797 17905 5831
rect 19441 5797 19475 5831
rect 21234 5797 21268 5831
rect 22753 5797 22787 5831
rect 22845 5797 22879 5831
rect 24409 5797 24443 5831
rect 1409 5729 1443 5763
rect 4445 5729 4479 5763
rect 5273 5729 5307 5763
rect 6101 5729 6135 5763
rect 8620 5729 8654 5763
rect 10241 5729 10275 5763
rect 13645 5729 13679 5763
rect 16129 5729 16163 5763
rect 16497 5729 16531 5763
rect 18705 5729 18739 5763
rect 20913 5729 20947 5763
rect 7113 5661 7147 5695
rect 7389 5661 7423 5695
rect 11897 5661 11931 5695
rect 12081 5661 12115 5695
rect 17509 5661 17543 5695
rect 19349 5661 19383 5695
rect 19993 5661 20027 5695
rect 23029 5661 23063 5695
rect 24317 5661 24351 5695
rect 1593 5593 1627 5627
rect 8723 5593 8757 5627
rect 12633 5593 12667 5627
rect 17417 5593 17451 5627
rect 24869 5593 24903 5627
rect 4583 5525 4617 5559
rect 11161 5525 11195 5559
rect 13461 5525 13495 5559
rect 14565 5525 14599 5559
rect 14933 5525 14967 5559
rect 18429 5525 18463 5559
rect 20269 5525 20303 5559
rect 23765 5525 23799 5559
rect 1823 5321 1857 5355
rect 8585 5321 8619 5355
rect 9137 5321 9171 5355
rect 9689 5321 9723 5355
rect 11805 5321 11839 5355
rect 13553 5321 13587 5355
rect 16037 5321 16071 5355
rect 19441 5321 19475 5355
rect 20269 5321 20303 5355
rect 21649 5321 21683 5355
rect 23029 5321 23063 5355
rect 24685 5321 24719 5355
rect 25053 5321 25087 5355
rect 25375 5321 25409 5355
rect 2237 5253 2271 5287
rect 7941 5253 7975 5287
rect 10701 5253 10735 5287
rect 12265 5253 12299 5287
rect 23765 5253 23799 5287
rect 5917 5185 5951 5219
rect 6285 5185 6319 5219
rect 7389 5185 7423 5219
rect 11529 5185 11563 5219
rect 13185 5185 13219 5219
rect 15669 5185 15703 5219
rect 17141 5185 17175 5219
rect 18429 5185 18463 5219
rect 19809 5185 19843 5219
rect 22201 5185 22235 5219
rect 24133 5185 24167 5219
rect 1752 5117 1786 5151
rect 4537 5117 4571 5151
rect 5089 5117 5123 5151
rect 5825 5117 5859 5151
rect 9321 5117 9355 5151
rect 11437 5117 11471 5151
rect 14289 5117 14323 5151
rect 14473 5117 14507 5151
rect 16681 5117 16715 5151
rect 16957 5117 16991 5151
rect 20453 5117 20487 5151
rect 22661 5117 22695 5151
rect 23489 5117 23523 5151
rect 23673 5117 23707 5151
rect 23949 5117 23983 5151
rect 25304 5117 25338 5151
rect 25789 5117 25823 5151
rect 7205 5049 7239 5083
rect 7481 5049 7515 5083
rect 12541 5049 12575 5083
rect 12633 5049 12667 5083
rect 15117 5049 15151 5083
rect 18153 5049 18187 5083
rect 18245 5049 18279 5083
rect 19073 5049 19107 5083
rect 6653 4981 6687 5015
rect 10241 4981 10275 5015
rect 17509 4981 17543 5015
rect 20821 4981 20855 5015
rect 21373 4981 21407 5015
rect 1593 4777 1627 4811
rect 7849 4777 7883 4811
rect 8125 4777 8159 4811
rect 9505 4777 9539 4811
rect 14841 4777 14875 4811
rect 15439 4777 15473 4811
rect 17509 4777 17543 4811
rect 18613 4777 18647 4811
rect 21373 4777 21407 4811
rect 23765 4777 23799 4811
rect 7205 4709 7239 4743
rect 8769 4709 8803 4743
rect 10977 4709 11011 4743
rect 11529 4709 11563 4743
rect 13829 4709 13863 4743
rect 18429 4709 18463 4743
rect 19993 4709 20027 4743
rect 20453 4709 20487 4743
rect 22385 4709 22419 4743
rect 5984 4641 6018 4675
rect 10609 4641 10643 4675
rect 12265 4641 12299 4675
rect 13001 4641 13035 4675
rect 13921 4641 13955 4675
rect 15368 4641 15402 4675
rect 16773 4641 16807 4675
rect 18220 4641 18254 4675
rect 6469 4573 6503 4607
rect 6929 4573 6963 4607
rect 9781 4573 9815 4607
rect 10885 4573 10919 4607
rect 12357 4573 12391 4607
rect 16313 4573 16347 4607
rect 19257 4641 19291 4675
rect 19809 4641 19843 4675
rect 20980 4641 21014 4675
rect 21741 4573 21775 4607
rect 22293 4573 22327 4607
rect 6055 4505 6089 4539
rect 13369 4505 13403 4539
rect 14105 4505 14139 4539
rect 18291 4505 18325 4539
rect 18429 4505 18463 4539
rect 21051 4505 21085 4539
rect 22845 4505 22879 4539
rect 6837 4437 6871 4471
rect 9045 4437 9079 4471
rect 10333 4437 10367 4471
rect 11805 4437 11839 4471
rect 14473 4437 14507 4471
rect 16037 4437 16071 4471
rect 18061 4437 18095 4471
rect 6193 4233 6227 4267
rect 13737 4233 13771 4267
rect 15853 4233 15887 4267
rect 17509 4233 17543 4267
rect 19257 4233 19291 4267
rect 21465 4233 21499 4267
rect 22661 4233 22695 4267
rect 23029 4233 23063 4267
rect 24731 4233 24765 4267
rect 13093 4165 13127 4199
rect 20637 4165 20671 4199
rect 22293 4165 22327 4199
rect 8493 4097 8527 4131
rect 11713 4097 11747 4131
rect 13737 4097 13771 4131
rect 14013 4097 14047 4131
rect 18153 4097 18187 4131
rect 18521 4097 18555 4131
rect 20269 4097 20303 4131
rect 21189 4097 21223 4131
rect 21741 4097 21775 4131
rect 5089 4029 5123 4063
rect 5825 4029 5859 4063
rect 6929 4029 6963 4063
rect 7389 4029 7423 4063
rect 7757 4029 7791 4063
rect 8125 4029 8159 4063
rect 8677 4029 8711 4063
rect 9873 4029 9907 4063
rect 10517 4029 10551 4063
rect 10701 4029 10735 4063
rect 11253 4029 11287 4063
rect 13553 4029 13587 4063
rect 14105 4029 14139 4063
rect 14565 4029 14599 4063
rect 14933 4029 14967 4063
rect 15485 4029 15519 4063
rect 19901 4029 19935 4063
rect 20085 4029 20119 4063
rect 24660 4029 24694 4063
rect 5917 3961 5951 3995
rect 8493 3961 8527 3995
rect 9781 3961 9815 3995
rect 11345 3961 11379 3995
rect 12541 3961 12575 3995
rect 12633 3961 12667 3995
rect 15577 3961 15611 3995
rect 16497 3961 16531 3995
rect 16589 3961 16623 3995
rect 17141 3961 17175 3995
rect 18245 3961 18279 3995
rect 21833 3961 21867 3995
rect 6561 3893 6595 3927
rect 7021 3893 7055 3927
rect 9321 3893 9355 3927
rect 12265 3893 12299 3927
rect 16313 3893 16347 3927
rect 17785 3893 17819 3927
rect 25145 3893 25179 3927
rect 9505 3689 9539 3723
rect 9965 3689 9999 3723
rect 11437 3689 11471 3723
rect 13001 3689 13035 3723
rect 14565 3689 14599 3723
rect 18429 3689 18463 3723
rect 20085 3689 20119 3723
rect 21373 3689 21407 3723
rect 5273 3621 5307 3655
rect 7481 3621 7515 3655
rect 8401 3621 8435 3655
rect 12081 3621 12115 3655
rect 12173 3621 12207 3655
rect 13553 3621 13587 3655
rect 15663 3621 15697 3655
rect 16589 3621 16623 3655
rect 17233 3621 17267 3655
rect 4525 3553 4559 3587
rect 4813 3553 4847 3587
rect 6193 3553 6227 3587
rect 7113 3553 7147 3587
rect 7665 3553 7699 3587
rect 7941 3553 7975 3587
rect 9689 3553 9723 3587
rect 10425 3553 10459 3587
rect 10517 3553 10551 3587
rect 11069 3553 11103 3587
rect 13645 3553 13679 3587
rect 16221 3553 16255 3587
rect 18705 3553 18739 3587
rect 20913 3553 20947 3587
rect 21005 3553 21039 3587
rect 21189 3553 21223 3587
rect 22477 3553 22511 3587
rect 23540 3553 23574 3587
rect 8677 3485 8711 3519
rect 15301 3485 15335 3519
rect 17141 3485 17175 3519
rect 17417 3485 17451 3519
rect 18613 3485 18647 3519
rect 23627 3485 23661 3519
rect 4629 3417 4663 3451
rect 7757 3417 7791 3451
rect 12633 3417 12667 3451
rect 16957 3417 16991 3451
rect 21925 3417 21959 3451
rect 5549 3349 5583 3383
rect 6561 3349 6595 3383
rect 9137 3349 9171 3383
rect 11897 3349 11931 3383
rect 13461 3349 13495 3383
rect 15117 3349 15151 3383
rect 18153 3349 18187 3383
rect 19717 3349 19751 3383
rect 22615 3349 22649 3383
rect 1547 3145 1581 3179
rect 3709 3145 3743 3179
rect 6561 3145 6595 3179
rect 12081 3145 12115 3179
rect 16313 3145 16347 3179
rect 17417 3145 17451 3179
rect 20913 3145 20947 3179
rect 24731 3145 24765 3179
rect 4307 3077 4341 3111
rect 10149 3077 10183 3111
rect 10517 3077 10551 3111
rect 13553 3077 13587 3111
rect 15485 3077 15519 3111
rect 19717 3077 19751 3111
rect 21281 3077 21315 3111
rect 5917 3009 5951 3043
rect 8217 3009 8251 3043
rect 9137 3009 9171 3043
rect 10609 3009 10643 3043
rect 12541 3009 12575 3043
rect 12817 3009 12851 3043
rect 16497 3009 16531 3043
rect 17141 3009 17175 3043
rect 18153 3009 18187 3043
rect 18429 3009 18463 3043
rect 20085 3009 20119 3043
rect 21649 3009 21683 3043
rect 1476 2941 1510 2975
rect 1869 2941 1903 2975
rect 4077 2941 4111 2975
rect 4204 2941 4238 2975
rect 5089 2941 5123 2975
rect 5825 2941 5859 2975
rect 6009 2941 6043 2975
rect 7481 2941 7515 2975
rect 7573 2941 7607 2975
rect 7757 2941 7791 2975
rect 8493 2941 8527 2975
rect 9781 2941 9815 2975
rect 14013 2941 14047 2975
rect 14105 2941 14139 2975
rect 14565 2941 14599 2975
rect 14933 2941 14967 2975
rect 15485 2941 15519 2975
rect 19165 2941 19199 2975
rect 19625 2941 19659 2975
rect 19901 2941 19935 2975
rect 21189 2941 21223 2975
rect 21465 2941 21499 2975
rect 22201 2941 22235 2975
rect 24660 2941 24694 2975
rect 6193 2873 6227 2907
rect 7297 2873 7331 2907
rect 9229 2873 9263 2907
rect 12633 2873 12667 2907
rect 16589 2873 16623 2907
rect 17877 2873 17911 2907
rect 18245 2873 18279 2907
rect 22937 2873 22971 2907
rect 4629 2805 4663 2839
rect 6009 2805 6043 2839
rect 8861 2805 8895 2839
rect 10977 2805 11011 2839
rect 11529 2805 11563 2839
rect 15853 2805 15887 2839
rect 19441 2805 19475 2839
rect 22661 2805 22695 2839
rect 23857 2805 23891 2839
rect 25145 2805 25179 2839
rect 3893 2601 3927 2635
rect 4537 2601 4571 2635
rect 7113 2601 7147 2635
rect 13645 2601 13679 2635
rect 14473 2601 14507 2635
rect 14933 2601 14967 2635
rect 16405 2601 16439 2635
rect 17233 2601 17267 2635
rect 19717 2601 19751 2635
rect 20545 2601 20579 2635
rect 21373 2601 21407 2635
rect 3525 2533 3559 2567
rect 4813 2533 4847 2567
rect 7481 2533 7515 2567
rect 7941 2533 7975 2567
rect 8769 2533 8803 2567
rect 10194 2533 10228 2567
rect 11069 2533 11103 2567
rect 12725 2533 12759 2567
rect 12817 2533 12851 2567
rect 14197 2533 14231 2567
rect 15806 2533 15840 2567
rect 18061 2533 18095 2567
rect 18521 2533 18555 2567
rect 3040 2465 3074 2499
rect 4328 2465 4362 2499
rect 5181 2465 5215 2499
rect 5365 2465 5399 2499
rect 6929 2465 6963 2499
rect 8033 2465 8067 2499
rect 8309 2465 8343 2499
rect 9873 2465 9907 2499
rect 11437 2465 11471 2499
rect 12449 2465 12483 2499
rect 14289 2465 14323 2499
rect 15485 2465 15519 2499
rect 16681 2465 16715 2499
rect 17785 2465 17819 2499
rect 19901 2465 19935 2499
rect 20913 2465 20947 2499
rect 21649 2465 21683 2499
rect 22201 2465 22235 2499
rect 22788 2465 22822 2499
rect 23213 2465 23247 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 5273 2397 5307 2431
rect 6285 2397 6319 2431
rect 6653 2397 6687 2431
rect 8125 2397 8159 2431
rect 11989 2397 12023 2431
rect 17141 2397 17175 2431
rect 17877 2397 17911 2431
rect 18429 2397 18463 2431
rect 3111 2329 3145 2363
rect 9045 2329 9079 2363
rect 10793 2329 10827 2363
rect 13277 2329 13311 2363
rect 15209 2329 15243 2363
rect 18981 2329 19015 2363
rect 20085 2329 20119 2363
rect 21833 2329 21867 2363
rect 24777 2329 24811 2363
rect 9505 2261 9539 2295
rect 17877 2261 17911 2295
rect 22891 2261 22925 2295
<< metal1 >>
rect 8294 27480 8300 27532
rect 8352 27520 8358 27532
rect 9582 27520 9588 27532
rect 8352 27492 9588 27520
rect 8352 27480 8358 27492
rect 9582 27480 9588 27492
rect 9640 27480 9646 27532
rect 11054 27480 11060 27532
rect 11112 27520 11118 27532
rect 11698 27520 11704 27532
rect 11112 27492 11704 27520
rect 11112 27480 11118 27492
rect 11698 27480 11704 27492
rect 11756 27480 11762 27532
rect 15746 27480 15752 27532
rect 15804 27520 15810 27532
rect 18230 27520 18236 27532
rect 15804 27492 18236 27520
rect 15804 27480 15810 27492
rect 18230 27480 18236 27492
rect 18288 27480 18294 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 22830 24265 22836 24268
rect 22808 24259 22836 24265
rect 22808 24256 22820 24259
rect 22743 24228 22820 24256
rect 22808 24225 22820 24228
rect 22888 24256 22894 24268
rect 24670 24256 24676 24268
rect 22888 24228 24676 24256
rect 22808 24219 22836 24225
rect 22830 24216 22836 24219
rect 22888 24216 22894 24228
rect 24670 24216 24676 24228
rect 24728 24216 24734 24268
rect 21082 24012 21088 24064
rect 21140 24052 21146 24064
rect 22879 24055 22937 24061
rect 22879 24052 22891 24055
rect 21140 24024 22891 24052
rect 21140 24012 21146 24024
rect 22879 24021 22891 24024
rect 22925 24021 22937 24055
rect 22879 24015 22937 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 7009 23851 7067 23857
rect 7009 23817 7021 23851
rect 7055 23848 7067 23851
rect 7466 23848 7472 23860
rect 7055 23820 7472 23848
rect 7055 23817 7067 23820
rect 7009 23811 7067 23817
rect 7466 23808 7472 23820
rect 7524 23808 7530 23860
rect 21913 23851 21971 23857
rect 21913 23817 21925 23851
rect 21959 23848 21971 23851
rect 22462 23848 22468 23860
rect 21959 23820 22468 23848
rect 21959 23817 21971 23820
rect 21913 23811 21971 23817
rect 22462 23808 22468 23820
rect 22520 23808 22526 23860
rect 22830 23848 22836 23860
rect 22791 23820 22836 23848
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 24210 23848 24216 23860
rect 24171 23820 24216 23848
rect 24210 23808 24216 23820
rect 24268 23808 24274 23860
rect 25225 23851 25283 23857
rect 25225 23817 25237 23851
rect 25271 23848 25283 23851
rect 26786 23848 26792 23860
rect 25271 23820 26792 23848
rect 25271 23817 25283 23820
rect 25225 23811 25283 23817
rect 22738 23740 22744 23792
rect 22796 23780 22802 23792
rect 24811 23783 24869 23789
rect 24811 23780 24823 23783
rect 22796 23752 24823 23780
rect 22796 23740 22802 23752
rect 24811 23749 24823 23752
rect 24857 23749 24869 23783
rect 24811 23743 24869 23749
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 6914 23644 6920 23656
rect 6871 23616 6920 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 6914 23604 6920 23616
rect 6972 23644 6978 23656
rect 7377 23647 7435 23653
rect 7377 23644 7389 23647
rect 6972 23616 7389 23644
rect 6972 23604 6978 23616
rect 7377 23613 7389 23616
rect 7423 23613 7435 23647
rect 7377 23607 7435 23613
rect 9192 23647 9250 23653
rect 9192 23613 9204 23647
rect 9238 23644 9250 23647
rect 9582 23644 9588 23656
rect 9238 23616 9588 23644
rect 9238 23613 9250 23616
rect 9192 23607 9250 23613
rect 9582 23604 9588 23616
rect 9640 23604 9646 23656
rect 10321 23647 10379 23653
rect 10321 23613 10333 23647
rect 10367 23644 10379 23647
rect 10870 23644 10876 23656
rect 10367 23616 10876 23644
rect 10367 23613 10379 23616
rect 10321 23607 10379 23613
rect 10870 23604 10876 23616
rect 10928 23604 10934 23656
rect 21542 23604 21548 23656
rect 21600 23644 21606 23656
rect 21729 23647 21787 23653
rect 21729 23644 21741 23647
rect 21600 23616 21741 23644
rect 21600 23604 21606 23616
rect 21729 23613 21741 23616
rect 21775 23644 21787 23647
rect 22281 23647 22339 23653
rect 22281 23644 22293 23647
rect 21775 23616 22293 23644
rect 21775 23613 21787 23616
rect 21729 23607 21787 23613
rect 22281 23613 22293 23616
rect 22327 23613 22339 23647
rect 22281 23607 22339 23613
rect 23712 23647 23770 23653
rect 23712 23613 23724 23647
rect 23758 23644 23770 23647
rect 24210 23644 24216 23656
rect 23758 23616 24216 23644
rect 23758 23613 23770 23616
rect 23712 23607 23770 23613
rect 24210 23604 24216 23616
rect 24268 23604 24274 23656
rect 24740 23647 24798 23653
rect 24740 23613 24752 23647
rect 24786 23644 24798 23647
rect 25240 23644 25268 23811
rect 26786 23808 26792 23820
rect 26844 23808 26850 23860
rect 24786 23616 25268 23644
rect 24786 23613 24798 23616
rect 24740 23607 24798 23613
rect 22462 23536 22468 23588
rect 22520 23576 22526 23588
rect 23799 23579 23857 23585
rect 23799 23576 23811 23579
rect 22520 23548 23811 23576
rect 22520 23536 22526 23548
rect 23799 23545 23811 23548
rect 23845 23545 23857 23579
rect 23799 23539 23857 23545
rect 9263 23511 9321 23517
rect 9263 23477 9275 23511
rect 9309 23508 9321 23511
rect 9398 23508 9404 23520
rect 9309 23480 9404 23508
rect 9309 23477 9321 23480
rect 9263 23471 9321 23477
rect 9398 23468 9404 23480
rect 9456 23468 9462 23520
rect 10042 23468 10048 23520
rect 10100 23508 10106 23520
rect 10505 23511 10563 23517
rect 10505 23508 10517 23511
rect 10100 23480 10517 23508
rect 10100 23468 10106 23480
rect 10505 23477 10517 23480
rect 10551 23477 10563 23511
rect 10505 23471 10563 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 5258 23264 5264 23316
rect 5316 23304 5322 23316
rect 10042 23304 10048 23316
rect 5316 23276 10048 23304
rect 5316 23264 5322 23276
rect 10042 23264 10048 23276
rect 10100 23264 10106 23316
rect 10870 23264 10876 23316
rect 10928 23304 10934 23316
rect 11011 23307 11069 23313
rect 11011 23304 11023 23307
rect 10928 23276 11023 23304
rect 10928 23264 10934 23276
rect 11011 23273 11023 23276
rect 11057 23273 11069 23307
rect 11011 23267 11069 23273
rect 22830 23177 22836 23180
rect 22808 23171 22836 23177
rect 22808 23168 22820 23171
rect 22743 23140 22820 23168
rect 22808 23137 22820 23140
rect 22888 23168 22894 23180
rect 23198 23168 23204 23180
rect 22888 23140 23204 23168
rect 22808 23131 22836 23137
rect 22830 23128 22836 23131
rect 22888 23128 22894 23140
rect 23198 23128 23204 23140
rect 23256 23128 23262 23180
rect 10778 22964 10784 22976
rect 10739 22936 10784 22964
rect 10778 22924 10784 22936
rect 10836 22924 10842 22976
rect 22094 22924 22100 22976
rect 22152 22964 22158 22976
rect 22879 22967 22937 22973
rect 22879 22964 22891 22967
rect 22152 22936 22891 22964
rect 22152 22924 22158 22936
rect 22879 22933 22891 22936
rect 22925 22933 22937 22967
rect 22879 22927 22937 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 22830 22760 22836 22772
rect 22791 22732 22836 22760
rect 22830 22720 22836 22732
rect 22888 22720 22894 22772
rect 25130 22760 25136 22772
rect 25091 22732 25136 22760
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 1394 22556 1400 22568
rect 1355 22528 1400 22556
rect 1394 22516 1400 22528
rect 1452 22556 1458 22568
rect 1949 22559 2007 22565
rect 1949 22556 1961 22559
rect 1452 22528 1961 22556
rect 1452 22516 1458 22528
rect 1949 22525 1961 22528
rect 1995 22525 2007 22559
rect 1949 22519 2007 22525
rect 24632 22559 24690 22565
rect 24632 22525 24644 22559
rect 24678 22556 24690 22559
rect 25130 22556 25136 22568
rect 24678 22528 25136 22556
rect 24678 22525 24690 22528
rect 24632 22519 24690 22525
rect 25130 22516 25136 22528
rect 25188 22516 25194 22568
rect 18874 22448 18880 22500
rect 18932 22488 18938 22500
rect 24719 22491 24777 22497
rect 24719 22488 24731 22491
rect 18932 22460 24731 22488
rect 18932 22448 18938 22460
rect 24719 22457 24731 22460
rect 24765 22457 24777 22491
rect 24719 22451 24777 22457
rect 14 22380 20 22432
rect 72 22420 78 22432
rect 1581 22423 1639 22429
rect 1581 22420 1593 22423
rect 72 22392 1593 22420
rect 72 22380 78 22392
rect 1581 22389 1593 22392
rect 1627 22389 1639 22423
rect 1581 22383 1639 22389
rect 10778 22380 10784 22432
rect 10836 22420 10842 22432
rect 10965 22423 11023 22429
rect 10965 22420 10977 22423
rect 10836 22392 10977 22420
rect 10836 22380 10842 22392
rect 10965 22389 10977 22392
rect 11011 22420 11023 22423
rect 11606 22420 11612 22432
rect 11011 22392 11612 22420
rect 11011 22389 11023 22392
rect 10965 22383 11023 22389
rect 11606 22380 11612 22392
rect 11664 22380 11670 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 1443 21440 2084 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 2056 21341 2084 21440
rect 2041 21335 2099 21341
rect 2041 21301 2053 21335
rect 2087 21332 2099 21335
rect 2130 21332 2136 21344
rect 2087 21304 2136 21332
rect 2087 21301 2099 21304
rect 2041 21295 2099 21301
rect 2130 21292 2136 21304
rect 2188 21292 2194 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 19797 21131 19855 21137
rect 19797 21097 19809 21131
rect 19843 21128 19855 21131
rect 19978 21128 19984 21140
rect 19843 21100 19984 21128
rect 19843 21097 19855 21100
rect 19797 21091 19855 21097
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 19610 20992 19616 21004
rect 19571 20964 19616 20992
rect 19610 20952 19616 20964
rect 19668 20952 19674 21004
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 18739 20519 18797 20525
rect 18739 20485 18751 20519
rect 18785 20516 18797 20519
rect 19610 20516 19616 20528
rect 18785 20488 19616 20516
rect 18785 20485 18797 20488
rect 18739 20479 18797 20485
rect 19610 20476 19616 20488
rect 19668 20476 19674 20528
rect 18414 20340 18420 20392
rect 18472 20380 18478 20392
rect 18668 20383 18726 20389
rect 18668 20380 18680 20383
rect 18472 20352 18680 20380
rect 18472 20340 18478 20352
rect 18668 20349 18680 20352
rect 18714 20380 18726 20383
rect 19061 20383 19119 20389
rect 19061 20380 19073 20383
rect 18714 20352 19073 20380
rect 18714 20349 18726 20352
rect 18668 20343 18726 20349
rect 19061 20349 19073 20352
rect 19107 20349 19119 20383
rect 19061 20343 19119 20349
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 12250 19864 12256 19916
rect 12308 19904 12314 19916
rect 12596 19907 12654 19913
rect 12596 19904 12608 19907
rect 12308 19876 12608 19904
rect 12308 19864 12314 19876
rect 12596 19873 12608 19876
rect 12642 19904 12654 19907
rect 13906 19904 13912 19916
rect 12642 19876 13912 19904
rect 12642 19873 12654 19876
rect 12596 19867 12654 19873
rect 13906 19864 13912 19876
rect 13964 19864 13970 19916
rect 14550 19864 14556 19916
rect 14608 19904 14614 19916
rect 15324 19907 15382 19913
rect 15324 19904 15336 19907
rect 14608 19876 15336 19904
rect 14608 19864 14614 19876
rect 15324 19873 15336 19876
rect 15370 19873 15382 19907
rect 15324 19867 15382 19873
rect 13722 19796 13728 19848
rect 13780 19836 13786 19848
rect 14001 19839 14059 19845
rect 14001 19836 14013 19839
rect 13780 19808 14013 19836
rect 13780 19796 13786 19808
rect 14001 19805 14013 19808
rect 14047 19805 14059 19839
rect 14001 19799 14059 19805
rect 12667 19703 12725 19709
rect 12667 19669 12679 19703
rect 12713 19700 12725 19703
rect 13630 19700 13636 19712
rect 12713 19672 13636 19700
rect 12713 19669 12725 19672
rect 12667 19663 12725 19669
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 15427 19703 15485 19709
rect 15427 19669 15439 19703
rect 15473 19700 15485 19703
rect 15562 19700 15568 19712
rect 15473 19672 15568 19700
rect 15473 19669 15485 19672
rect 15427 19663 15485 19669
rect 15562 19660 15568 19672
rect 15620 19660 15626 19712
rect 16025 19703 16083 19709
rect 16025 19669 16037 19703
rect 16071 19700 16083 19703
rect 16482 19700 16488 19712
rect 16071 19672 16488 19700
rect 16071 19669 16083 19672
rect 16025 19663 16083 19669
rect 16482 19660 16488 19672
rect 16540 19660 16546 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 12250 19496 12256 19508
rect 12211 19468 12256 19496
rect 12250 19456 12256 19468
rect 12308 19456 12314 19508
rect 13630 19456 13636 19508
rect 13688 19496 13694 19508
rect 13725 19499 13783 19505
rect 13725 19496 13737 19499
rect 13688 19468 13737 19496
rect 13688 19456 13694 19468
rect 13725 19465 13737 19468
rect 13771 19465 13783 19499
rect 13725 19459 13783 19465
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 12802 19292 12808 19304
rect 1443 19264 2084 19292
rect 12763 19264 12808 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 2056 19165 2084 19264
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 12894 19252 12900 19304
rect 12952 19292 12958 19304
rect 14956 19295 15014 19301
rect 14956 19292 14968 19295
rect 12952 19264 14968 19292
rect 12952 19252 12958 19264
rect 14956 19261 14968 19264
rect 15002 19292 15014 19295
rect 15381 19295 15439 19301
rect 15381 19292 15393 19295
rect 15002 19264 15393 19292
rect 15002 19261 15014 19264
rect 14956 19255 15014 19261
rect 15381 19261 15393 19264
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 15933 19295 15991 19301
rect 15933 19261 15945 19295
rect 15979 19261 15991 19295
rect 16482 19292 16488 19304
rect 16395 19264 16488 19292
rect 15933 19255 15991 19261
rect 13446 19224 13452 19236
rect 13407 19196 13452 19224
rect 13446 19184 13452 19196
rect 13504 19184 13510 19236
rect 15470 19184 15476 19236
rect 15528 19224 15534 19236
rect 15749 19227 15807 19233
rect 15749 19224 15761 19227
rect 15528 19196 15761 19224
rect 15528 19184 15534 19196
rect 15749 19193 15761 19196
rect 15795 19224 15807 19227
rect 15948 19224 15976 19255
rect 16482 19252 16488 19264
rect 16540 19292 16546 19304
rect 19058 19292 19064 19304
rect 16540 19264 19064 19292
rect 16540 19252 16546 19264
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 16666 19224 16672 19236
rect 15795 19196 15976 19224
rect 16627 19196 16672 19224
rect 15795 19193 15807 19196
rect 15749 19187 15807 19193
rect 16666 19184 16672 19196
rect 16724 19184 16730 19236
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19156 2099 19159
rect 2406 19156 2412 19168
rect 2087 19128 2412 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 2406 19116 2412 19128
rect 2464 19116 2470 19168
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 14737 19159 14795 19165
rect 14737 19156 14749 19159
rect 14608 19128 14749 19156
rect 14608 19116 14614 19128
rect 14737 19125 14749 19128
rect 14783 19125 14795 19159
rect 14737 19119 14795 19125
rect 15059 19159 15117 19165
rect 15059 19125 15071 19159
rect 15105 19156 15117 19159
rect 15654 19156 15660 19168
rect 15105 19128 15660 19156
rect 15105 19125 15117 19128
rect 15059 19119 15117 19125
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 9950 18952 9956 18964
rect 9911 18924 9956 18952
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 12802 18952 12808 18964
rect 12763 18924 12808 18952
rect 12802 18912 12808 18924
rect 12860 18912 12866 18964
rect 13630 18952 13636 18964
rect 13280 18924 13636 18952
rect 10870 18844 10876 18896
rect 10928 18884 10934 18896
rect 13280 18893 13308 18924
rect 13630 18912 13636 18924
rect 13688 18912 13694 18964
rect 13722 18912 13728 18964
rect 13780 18952 13786 18964
rect 14185 18955 14243 18961
rect 14185 18952 14197 18955
rect 13780 18924 14197 18952
rect 13780 18912 13786 18924
rect 14185 18921 14197 18924
rect 14231 18952 14243 18955
rect 14274 18952 14280 18964
rect 14231 18924 14280 18952
rect 14231 18921 14243 18924
rect 14185 18915 14243 18921
rect 14274 18912 14280 18924
rect 14332 18912 14338 18964
rect 17218 18952 17224 18964
rect 17052 18924 17224 18952
rect 11793 18887 11851 18893
rect 11793 18884 11805 18887
rect 10928 18856 11805 18884
rect 10928 18844 10934 18856
rect 11793 18853 11805 18856
rect 11839 18853 11851 18887
rect 11793 18847 11851 18853
rect 13265 18887 13323 18893
rect 13265 18853 13277 18887
rect 13311 18853 13323 18887
rect 13265 18847 13323 18853
rect 13357 18887 13415 18893
rect 13357 18853 13369 18887
rect 13403 18884 13415 18887
rect 13446 18884 13452 18896
rect 13403 18856 13452 18884
rect 13403 18853 13415 18856
rect 13357 18847 13415 18853
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 17052 18893 17080 18924
rect 17218 18912 17224 18924
rect 17276 18952 17282 18964
rect 21082 18952 21088 18964
rect 17276 18924 21088 18952
rect 17276 18912 17282 18924
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 21542 18912 21548 18964
rect 21600 18952 21606 18964
rect 21637 18955 21695 18961
rect 21637 18952 21649 18955
rect 21600 18924 21649 18952
rect 21600 18912 21606 18924
rect 21637 18921 21649 18924
rect 21683 18921 21695 18955
rect 24762 18952 24768 18964
rect 24723 18924 24768 18952
rect 21637 18915 21695 18921
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 17037 18887 17095 18893
rect 17037 18853 17049 18887
rect 17083 18853 17095 18887
rect 17037 18847 17095 18853
rect 17126 18844 17132 18896
rect 17184 18884 17190 18896
rect 17184 18856 17229 18884
rect 17184 18844 17190 18856
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 1486 18816 1492 18828
rect 1443 18788 1492 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 1486 18776 1492 18788
rect 1544 18776 1550 18828
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18816 7895 18819
rect 7926 18816 7932 18828
rect 7883 18788 7932 18816
rect 7883 18785 7895 18788
rect 7837 18779 7895 18785
rect 7926 18776 7932 18788
rect 7984 18816 7990 18828
rect 8294 18816 8300 18828
rect 7984 18788 8300 18816
rect 7984 18776 7990 18788
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 9769 18819 9827 18825
rect 9769 18785 9781 18819
rect 9815 18816 9827 18819
rect 9858 18816 9864 18828
rect 9815 18788 9864 18816
rect 9815 18785 9827 18788
rect 9769 18779 9827 18785
rect 9858 18776 9864 18788
rect 9916 18776 9922 18828
rect 15378 18816 15384 18828
rect 15339 18788 15384 18816
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 15838 18816 15844 18828
rect 15799 18788 15844 18816
rect 15838 18776 15844 18788
rect 15896 18776 15902 18828
rect 21428 18819 21486 18825
rect 21428 18785 21440 18819
rect 21474 18816 21486 18819
rect 21726 18816 21732 18828
rect 21474 18788 21732 18816
rect 21474 18785 21486 18788
rect 21428 18779 21486 18785
rect 21726 18776 21732 18788
rect 21784 18776 21790 18828
rect 24581 18819 24639 18825
rect 24581 18785 24593 18819
rect 24627 18816 24639 18819
rect 24670 18816 24676 18828
rect 24627 18788 24676 18816
rect 24627 18785 24639 18788
rect 24581 18779 24639 18785
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 11698 18748 11704 18760
rect 11659 18720 11704 18748
rect 11698 18708 11704 18720
rect 11756 18708 11762 18760
rect 11974 18748 11980 18760
rect 11935 18720 11980 18748
rect 11974 18708 11980 18720
rect 12032 18708 12038 18760
rect 13722 18748 13728 18760
rect 13683 18720 13728 18748
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18748 16175 18751
rect 17402 18748 17408 18760
rect 16163 18720 17408 18748
rect 16163 18717 16175 18720
rect 16117 18711 16175 18717
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 17681 18751 17739 18757
rect 17681 18717 17693 18751
rect 17727 18748 17739 18751
rect 17770 18748 17776 18760
rect 17727 18720 17776 18748
rect 17727 18717 17739 18720
rect 17681 18711 17739 18717
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 8018 18680 8024 18692
rect 7979 18652 8024 18680
rect 8018 18640 8024 18652
rect 8076 18640 8082 18692
rect 16206 18640 16212 18692
rect 16264 18680 16270 18692
rect 16761 18683 16819 18689
rect 16761 18680 16773 18683
rect 16264 18652 16773 18680
rect 16264 18640 16270 18652
rect 16761 18649 16773 18652
rect 16807 18649 16819 18683
rect 16761 18643 16819 18649
rect 1535 18615 1593 18621
rect 1535 18581 1547 18615
rect 1581 18612 1593 18615
rect 8294 18612 8300 18624
rect 1581 18584 8300 18612
rect 1581 18581 1593 18584
rect 1535 18575 1593 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 16390 18612 16396 18624
rect 16351 18584 16396 18612
rect 16390 18572 16396 18584
rect 16448 18572 16454 18624
rect 18046 18612 18052 18624
rect 18007 18584 18052 18612
rect 18046 18572 18052 18584
rect 18104 18572 18110 18624
rect 21910 18612 21916 18624
rect 21871 18584 21916 18612
rect 21910 18572 21916 18584
rect 21968 18572 21974 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1486 18368 1492 18420
rect 1544 18408 1550 18420
rect 1857 18411 1915 18417
rect 1857 18408 1869 18411
rect 1544 18380 1869 18408
rect 1544 18368 1550 18380
rect 1857 18377 1869 18380
rect 1903 18377 1915 18411
rect 7926 18408 7932 18420
rect 7887 18380 7932 18408
rect 1857 18371 1915 18377
rect 7926 18368 7932 18380
rect 7984 18408 7990 18420
rect 11793 18411 11851 18417
rect 11793 18408 11805 18411
rect 7984 18380 11805 18408
rect 7984 18368 7990 18380
rect 1854 18272 1860 18284
rect 1479 18244 1860 18272
rect 1479 18213 1507 18244
rect 1854 18232 1860 18244
rect 1912 18272 1918 18284
rect 2225 18275 2283 18281
rect 2225 18272 2237 18275
rect 1912 18244 2237 18272
rect 1912 18232 1918 18244
rect 2225 18241 2237 18244
rect 2271 18241 2283 18275
rect 8938 18272 8944 18284
rect 2225 18235 2283 18241
rect 4126 18244 8944 18272
rect 1448 18207 1507 18213
rect 1448 18173 1460 18207
rect 1494 18176 1507 18207
rect 1535 18207 1593 18213
rect 1494 18173 1506 18176
rect 1448 18167 1506 18173
rect 1535 18173 1547 18207
rect 1581 18204 1593 18207
rect 4126 18204 4154 18244
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 11399 18213 11427 18380
rect 11793 18377 11805 18380
rect 11839 18408 11851 18411
rect 12894 18408 12900 18420
rect 11839 18380 12900 18408
rect 11839 18377 11851 18380
rect 11793 18371 11851 18377
rect 12894 18368 12900 18380
rect 12952 18368 12958 18420
rect 13446 18368 13452 18420
rect 13504 18408 13510 18420
rect 13633 18411 13691 18417
rect 13633 18408 13645 18411
rect 13504 18380 13645 18408
rect 13504 18368 13510 18380
rect 13633 18377 13645 18380
rect 13679 18377 13691 18411
rect 13633 18371 13691 18377
rect 14274 18272 14280 18284
rect 14235 18244 14280 18272
rect 14274 18232 14280 18244
rect 14332 18232 14338 18284
rect 14550 18272 14556 18284
rect 14511 18244 14556 18272
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 16206 18272 16212 18284
rect 16167 18244 16212 18272
rect 16206 18232 16212 18244
rect 16264 18232 16270 18284
rect 20806 18232 20812 18284
rect 20864 18272 20870 18284
rect 24581 18275 24639 18281
rect 24581 18272 24593 18275
rect 20864 18244 24593 18272
rect 20864 18232 20870 18244
rect 24581 18241 24593 18244
rect 24627 18272 24639 18275
rect 24670 18272 24676 18284
rect 24627 18244 24676 18272
rect 24627 18241 24639 18244
rect 24581 18235 24639 18241
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 1581 18176 4154 18204
rect 9636 18207 9694 18213
rect 1581 18173 1593 18176
rect 1535 18167 1593 18173
rect 9636 18173 9648 18207
rect 9682 18204 9694 18207
rect 11384 18207 11442 18213
rect 9682 18176 10548 18204
rect 9682 18173 9694 18176
rect 9636 18167 9694 18173
rect 9723 18139 9781 18145
rect 9723 18136 9735 18139
rect 4126 18108 9735 18136
rect 2406 18028 2412 18080
rect 2464 18068 2470 18080
rect 4126 18068 4154 18108
rect 9723 18105 9735 18108
rect 9769 18105 9781 18139
rect 9723 18099 9781 18105
rect 2464 18040 4154 18068
rect 2464 18028 2470 18040
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 10520 18077 10548 18176
rect 11384 18173 11396 18207
rect 11430 18173 11442 18207
rect 11384 18167 11442 18173
rect 17865 18207 17923 18213
rect 17865 18173 17877 18207
rect 17911 18204 17923 18207
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17911 18176 18061 18204
rect 17911 18173 17923 18176
rect 17865 18167 17923 18173
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 11471 18139 11529 18145
rect 11471 18105 11483 18139
rect 11517 18136 11529 18139
rect 12710 18136 12716 18148
rect 11517 18108 12716 18136
rect 11517 18105 11529 18108
rect 11471 18099 11529 18105
rect 12710 18096 12716 18108
rect 12768 18096 12774 18148
rect 12802 18096 12808 18148
rect 12860 18136 12866 18148
rect 13357 18139 13415 18145
rect 12860 18108 12905 18136
rect 12860 18096 12866 18108
rect 13357 18105 13369 18139
rect 13403 18136 13415 18139
rect 13722 18136 13728 18148
rect 13403 18108 13728 18136
rect 13403 18105 13415 18108
rect 13357 18099 13415 18105
rect 13722 18096 13728 18108
rect 13780 18096 13786 18148
rect 14093 18139 14151 18145
rect 14093 18105 14105 18139
rect 14139 18136 14151 18139
rect 14366 18136 14372 18148
rect 14139 18108 14372 18136
rect 14139 18105 14151 18108
rect 14093 18099 14151 18105
rect 14366 18096 14372 18108
rect 14424 18096 14430 18148
rect 16301 18139 16359 18145
rect 16301 18105 16313 18139
rect 16347 18136 16359 18139
rect 16390 18136 16396 18148
rect 16347 18108 16396 18136
rect 16347 18105 16359 18108
rect 16301 18099 16359 18105
rect 16390 18096 16396 18108
rect 16448 18096 16454 18148
rect 16850 18136 16856 18148
rect 16811 18108 16856 18136
rect 16850 18096 16856 18108
rect 16908 18096 16914 18148
rect 18064 18136 18092 18167
rect 18138 18164 18144 18216
rect 18196 18204 18202 18216
rect 18509 18207 18567 18213
rect 18509 18204 18521 18207
rect 18196 18176 18521 18204
rect 18196 18164 18202 18176
rect 18509 18173 18521 18176
rect 18555 18173 18567 18207
rect 18509 18167 18567 18173
rect 18782 18136 18788 18148
rect 18064 18108 18788 18136
rect 18782 18096 18788 18108
rect 18840 18096 18846 18148
rect 21361 18139 21419 18145
rect 21361 18105 21373 18139
rect 21407 18136 21419 18139
rect 21726 18136 21732 18148
rect 21407 18108 21732 18136
rect 21407 18105 21419 18108
rect 21361 18099 21419 18105
rect 21726 18096 21732 18108
rect 21784 18096 21790 18148
rect 21910 18136 21916 18148
rect 21871 18108 21916 18136
rect 21910 18096 21916 18108
rect 21968 18096 21974 18148
rect 22005 18139 22063 18145
rect 22005 18105 22017 18139
rect 22051 18105 22063 18139
rect 22005 18099 22063 18105
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9916 18040 10057 18068
rect 9916 18028 9922 18040
rect 10045 18037 10057 18040
rect 10091 18037 10103 18071
rect 10045 18031 10103 18037
rect 10505 18071 10563 18077
rect 10505 18037 10517 18071
rect 10551 18068 10563 18071
rect 10778 18068 10784 18080
rect 10551 18040 10784 18068
rect 10551 18037 10563 18040
rect 10505 18031 10563 18037
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 10870 18028 10876 18080
rect 10928 18068 10934 18080
rect 11149 18071 11207 18077
rect 11149 18068 11161 18071
rect 10928 18040 11161 18068
rect 10928 18028 10934 18040
rect 11149 18037 11161 18040
rect 11195 18037 11207 18071
rect 11149 18031 11207 18037
rect 12253 18071 12311 18077
rect 12253 18037 12265 18071
rect 12299 18068 12311 18071
rect 12820 18068 12848 18096
rect 15378 18068 15384 18080
rect 12299 18040 12848 18068
rect 15339 18040 15384 18068
rect 12299 18037 12311 18040
rect 12253 18031 12311 18037
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 15838 18068 15844 18080
rect 15799 18040 15844 18068
rect 15838 18028 15844 18040
rect 15896 18028 15902 18080
rect 17034 18028 17040 18080
rect 17092 18068 17098 18080
rect 17129 18071 17187 18077
rect 17129 18068 17141 18071
rect 17092 18040 17141 18068
rect 17092 18028 17098 18040
rect 17129 18037 17141 18040
rect 17175 18037 17187 18071
rect 17129 18031 17187 18037
rect 17954 18028 17960 18080
rect 18012 18068 18018 18080
rect 18141 18071 18199 18077
rect 18141 18068 18153 18071
rect 18012 18040 18153 18068
rect 18012 18028 18018 18040
rect 18141 18037 18153 18040
rect 18187 18037 18199 18071
rect 18141 18031 18199 18037
rect 21637 18071 21695 18077
rect 21637 18037 21649 18071
rect 21683 18068 21695 18071
rect 22020 18068 22048 18099
rect 22186 18096 22192 18148
rect 22244 18136 22250 18148
rect 22557 18139 22615 18145
rect 22557 18136 22569 18139
rect 22244 18108 22569 18136
rect 22244 18096 22250 18108
rect 22557 18105 22569 18108
rect 22603 18136 22615 18139
rect 24946 18136 24952 18148
rect 22603 18108 24952 18136
rect 22603 18105 22615 18108
rect 22557 18099 22615 18105
rect 24946 18096 24952 18108
rect 25004 18096 25010 18148
rect 22922 18068 22928 18080
rect 21683 18040 22928 18068
rect 21683 18037 21695 18040
rect 21637 18031 21695 18037
rect 22922 18028 22928 18040
rect 22980 18028 22986 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 12158 17864 12164 17876
rect 12119 17836 12164 17864
rect 12158 17824 12164 17836
rect 12216 17824 12222 17876
rect 12713 17867 12771 17873
rect 12713 17833 12725 17867
rect 12759 17864 12771 17867
rect 12802 17864 12808 17876
rect 12759 17836 12808 17864
rect 12759 17833 12771 17836
rect 12713 17827 12771 17833
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 15654 17824 15660 17876
rect 15712 17864 15718 17876
rect 15933 17867 15991 17873
rect 15933 17864 15945 17867
rect 15712 17836 15945 17864
rect 15712 17824 15718 17836
rect 15933 17833 15945 17836
rect 15979 17833 15991 17867
rect 17218 17864 17224 17876
rect 17179 17836 17224 17864
rect 15933 17827 15991 17833
rect 17218 17824 17224 17836
rect 17276 17824 17282 17876
rect 22094 17864 22100 17876
rect 22055 17836 22100 17864
rect 22094 17824 22100 17836
rect 22152 17824 22158 17876
rect 22462 17824 22468 17876
rect 22520 17864 22526 17876
rect 24762 17864 24768 17876
rect 22520 17836 22600 17864
rect 24723 17836 24768 17864
rect 22520 17824 22526 17836
rect 9398 17756 9404 17808
rect 9456 17796 9462 17808
rect 10321 17799 10379 17805
rect 10321 17796 10333 17799
rect 9456 17768 10333 17796
rect 9456 17756 9462 17768
rect 10321 17765 10333 17768
rect 10367 17765 10379 17799
rect 10321 17759 10379 17765
rect 10413 17799 10471 17805
rect 10413 17765 10425 17799
rect 10459 17796 10471 17799
rect 10686 17796 10692 17808
rect 10459 17768 10692 17796
rect 10459 17765 10471 17768
rect 10413 17759 10471 17765
rect 10686 17756 10692 17768
rect 10744 17756 10750 17808
rect 10965 17799 11023 17805
rect 10965 17765 10977 17799
rect 11011 17796 11023 17799
rect 11974 17796 11980 17808
rect 11011 17768 11980 17796
rect 11011 17765 11023 17768
rect 10965 17759 11023 17765
rect 11974 17756 11980 17768
rect 12032 17756 12038 17808
rect 13814 17756 13820 17808
rect 13872 17796 13878 17808
rect 14369 17799 14427 17805
rect 13872 17768 13917 17796
rect 13872 17756 13878 17768
rect 14369 17765 14381 17799
rect 14415 17796 14427 17799
rect 14550 17796 14556 17808
rect 14415 17768 14556 17796
rect 14415 17765 14427 17768
rect 14369 17759 14427 17765
rect 14550 17756 14556 17768
rect 14608 17756 14614 17808
rect 16298 17796 16304 17808
rect 16259 17768 16304 17796
rect 16298 17756 16304 17768
rect 16356 17756 16362 17808
rect 17862 17796 17868 17808
rect 17823 17768 17868 17796
rect 17862 17756 17868 17768
rect 17920 17756 17926 17808
rect 18414 17796 18420 17808
rect 18375 17768 18420 17796
rect 18414 17756 18420 17768
rect 18472 17756 18478 17808
rect 22572 17805 22600 17836
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 22557 17799 22615 17805
rect 22557 17765 22569 17799
rect 22603 17765 22615 17799
rect 22557 17759 22615 17765
rect 22649 17799 22707 17805
rect 22649 17765 22661 17799
rect 22695 17796 22707 17799
rect 23014 17796 23020 17808
rect 22695 17768 23020 17796
rect 22695 17765 22707 17768
rect 22649 17759 22707 17765
rect 23014 17756 23020 17768
rect 23072 17756 23078 17808
rect 11698 17728 11704 17740
rect 11659 17700 11704 17728
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 11790 17660 11796 17672
rect 11751 17632 11796 17660
rect 11790 17620 11796 17632
rect 11848 17620 11854 17672
rect 11992 17660 12020 17756
rect 12710 17688 12716 17740
rect 12768 17728 12774 17740
rect 13357 17731 13415 17737
rect 13357 17728 13369 17731
rect 12768 17700 13369 17728
rect 12768 17688 12774 17700
rect 13357 17697 13369 17700
rect 13403 17697 13415 17731
rect 13357 17691 13415 17697
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 25038 17728 25044 17740
rect 24627 17700 25044 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 25038 17688 25044 17700
rect 25096 17688 25102 17740
rect 13538 17660 13544 17672
rect 11992 17632 13544 17660
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 13722 17660 13728 17672
rect 13683 17632 13728 17660
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 16209 17663 16267 17669
rect 16209 17629 16221 17663
rect 16255 17629 16267 17663
rect 16850 17660 16856 17672
rect 16763 17632 16856 17660
rect 16209 17623 16267 17629
rect 16114 17552 16120 17604
rect 16172 17592 16178 17604
rect 16224 17592 16252 17623
rect 16850 17620 16856 17632
rect 16908 17660 16914 17672
rect 17770 17660 17776 17672
rect 16908 17632 17776 17660
rect 16908 17620 16914 17632
rect 17770 17620 17776 17632
rect 17828 17620 17834 17672
rect 20990 17660 20996 17672
rect 20951 17632 20996 17660
rect 20990 17620 20996 17632
rect 21048 17620 21054 17672
rect 22830 17660 22836 17672
rect 22791 17632 22836 17660
rect 22830 17620 22836 17632
rect 22888 17620 22894 17672
rect 16172 17564 16252 17592
rect 16172 17552 16178 17564
rect 11238 17524 11244 17536
rect 11199 17496 11244 17524
rect 11238 17484 11244 17496
rect 11296 17484 11302 17536
rect 12802 17484 12808 17536
rect 12860 17524 12866 17536
rect 12989 17527 13047 17533
rect 12989 17524 13001 17527
rect 12860 17496 13001 17524
rect 12860 17484 12866 17496
rect 12989 17493 13001 17496
rect 13035 17493 13047 17527
rect 12989 17487 13047 17493
rect 20530 17484 20536 17536
rect 20588 17524 20594 17536
rect 21223 17527 21281 17533
rect 21223 17524 21235 17527
rect 20588 17496 21235 17524
rect 20588 17484 20594 17496
rect 21223 17493 21235 17496
rect 21269 17493 21281 17527
rect 21223 17487 21281 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 9398 17280 9404 17332
rect 9456 17320 9462 17332
rect 9585 17323 9643 17329
rect 9585 17320 9597 17323
rect 9456 17292 9597 17320
rect 9456 17280 9462 17292
rect 9585 17289 9597 17292
rect 9631 17289 9643 17323
rect 9585 17283 9643 17289
rect 17770 17280 17776 17332
rect 17828 17320 17834 17332
rect 19061 17323 19119 17329
rect 19061 17320 19073 17323
rect 17828 17292 19073 17320
rect 17828 17280 17834 17292
rect 19061 17289 19073 17292
rect 19107 17289 19119 17323
rect 21450 17320 21456 17332
rect 19061 17283 19119 17289
rect 21100 17292 21456 17320
rect 21100 17261 21128 17292
rect 21450 17280 21456 17292
rect 21508 17320 21514 17332
rect 22186 17320 22192 17332
rect 21508 17292 22192 17320
rect 21508 17280 21514 17292
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 22278 17280 22284 17332
rect 22336 17320 22342 17332
rect 23014 17320 23020 17332
rect 22336 17292 23020 17320
rect 22336 17280 22342 17292
rect 23014 17280 23020 17292
rect 23072 17280 23078 17332
rect 21085 17255 21143 17261
rect 21085 17221 21097 17255
rect 21131 17221 21143 17255
rect 21085 17215 21143 17221
rect 21174 17212 21180 17264
rect 21232 17252 21238 17264
rect 22830 17252 22836 17264
rect 21232 17224 22836 17252
rect 21232 17212 21238 17224
rect 9907 17187 9965 17193
rect 9907 17153 9919 17187
rect 9953 17184 9965 17187
rect 10873 17187 10931 17193
rect 10873 17184 10885 17187
rect 9953 17156 10885 17184
rect 9953 17153 9965 17156
rect 9907 17147 9965 17153
rect 10873 17153 10885 17156
rect 10919 17184 10931 17187
rect 11238 17184 11244 17196
rect 10919 17156 11244 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 14366 17184 14372 17196
rect 14327 17156 14372 17184
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 15654 17144 15660 17196
rect 15712 17184 15718 17196
rect 16301 17187 16359 17193
rect 16301 17184 16313 17187
rect 15712 17156 16313 17184
rect 15712 17144 15718 17156
rect 16301 17153 16313 17156
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 16945 17187 17003 17193
rect 16945 17153 16957 17187
rect 16991 17184 17003 17187
rect 18230 17184 18236 17196
rect 16991 17156 18236 17184
rect 16991 17153 17003 17156
rect 16945 17147 17003 17153
rect 18230 17144 18236 17156
rect 18288 17184 18294 17196
rect 18417 17187 18475 17193
rect 18417 17184 18429 17187
rect 18288 17156 18429 17184
rect 18288 17144 18294 17156
rect 18417 17153 18429 17156
rect 18463 17153 18475 17187
rect 20530 17184 20536 17196
rect 20491 17156 20536 17184
rect 18417 17147 18475 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 20990 17144 20996 17196
rect 21048 17184 21054 17196
rect 21453 17187 21511 17193
rect 21453 17184 21465 17187
rect 21048 17156 21465 17184
rect 21048 17144 21054 17156
rect 21453 17153 21465 17156
rect 21499 17184 21511 17187
rect 21542 17184 21548 17196
rect 21499 17156 21548 17184
rect 21499 17153 21511 17156
rect 21453 17147 21511 17153
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 22094 17184 22100 17196
rect 22055 17156 22100 17184
rect 22094 17144 22100 17156
rect 22152 17144 22158 17196
rect 22388 17193 22416 17224
rect 22830 17212 22836 17224
rect 22888 17212 22894 17264
rect 22373 17187 22431 17193
rect 22373 17153 22385 17187
rect 22419 17153 22431 17187
rect 22373 17147 22431 17153
rect 24210 17144 24216 17196
rect 24268 17184 24274 17196
rect 24719 17187 24777 17193
rect 24719 17184 24731 17187
rect 24268 17156 24731 17184
rect 24268 17144 24274 17156
rect 24719 17153 24731 17156
rect 24765 17153 24777 17187
rect 24719 17147 24777 17153
rect 9820 17119 9878 17125
rect 9820 17085 9832 17119
rect 9866 17116 9878 17119
rect 9866 17085 9904 17116
rect 9820 17079 9904 17085
rect 9876 16992 9904 17079
rect 12066 17076 12072 17128
rect 12124 17116 12130 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 12124 17088 12633 17116
rect 12124 17076 12130 17088
rect 12621 17085 12633 17088
rect 12667 17116 12679 17119
rect 12802 17116 12808 17128
rect 12667 17088 12808 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 12802 17076 12808 17088
rect 12860 17076 12866 17128
rect 13541 17119 13599 17125
rect 13541 17085 13553 17119
rect 13587 17116 13599 17119
rect 13814 17116 13820 17128
rect 13587 17088 13820 17116
rect 13587 17085 13599 17088
rect 13541 17079 13599 17085
rect 13814 17076 13820 17088
rect 13872 17116 13878 17128
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13872 17088 13921 17116
rect 13872 17076 13878 17088
rect 13909 17085 13921 17088
rect 13955 17116 13967 17119
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 13955 17088 14289 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 14277 17085 14289 17088
rect 14323 17116 14335 17119
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 14323 17088 14473 17116
rect 14323 17085 14335 17088
rect 14277 17079 14335 17085
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 24632 17119 24690 17125
rect 24632 17085 24644 17119
rect 24678 17116 24690 17119
rect 24854 17116 24860 17128
rect 24678 17088 24860 17116
rect 24678 17085 24690 17088
rect 24632 17079 24690 17085
rect 24854 17076 24860 17088
rect 24912 17116 24918 17128
rect 25409 17119 25467 17125
rect 25409 17116 25421 17119
rect 24912 17088 25421 17116
rect 24912 17076 24918 17088
rect 25409 17085 25421 17088
rect 25455 17085 25467 17119
rect 25409 17079 25467 17085
rect 10965 17051 11023 17057
rect 10965 17017 10977 17051
rect 11011 17017 11023 17051
rect 11514 17048 11520 17060
rect 11475 17020 11520 17048
rect 10965 17011 11023 17017
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 9916 16952 10241 16980
rect 9916 16940 9922 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 10229 16943 10287 16949
rect 10689 16983 10747 16989
rect 10689 16949 10701 16983
rect 10735 16980 10747 16983
rect 10870 16980 10876 16992
rect 10735 16952 10876 16980
rect 10735 16949 10747 16952
rect 10689 16943 10747 16949
rect 10870 16940 10876 16952
rect 10928 16980 10934 16992
rect 10980 16980 11008 17011
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 11885 17051 11943 17057
rect 11885 17017 11897 17051
rect 11931 17048 11943 17051
rect 12158 17048 12164 17060
rect 11931 17020 12164 17048
rect 11931 17017 11943 17020
rect 11885 17011 11943 17017
rect 12158 17008 12164 17020
rect 12216 17048 12222 17060
rect 12253 17051 12311 17057
rect 12253 17048 12265 17051
rect 12216 17020 12265 17048
rect 12216 17008 12222 17020
rect 12253 17017 12265 17020
rect 12299 17048 12311 17051
rect 12983 17051 13041 17057
rect 12983 17048 12995 17051
rect 12299 17020 12995 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12983 17017 12995 17020
rect 13029 17048 13041 17051
rect 13354 17048 13360 17060
rect 13029 17020 13360 17048
rect 13029 17017 13041 17020
rect 12983 17011 13041 17017
rect 13354 17008 13360 17020
rect 13412 17008 13418 17060
rect 16117 17051 16175 17057
rect 16117 17017 16129 17051
rect 16163 17048 16175 17051
rect 16393 17051 16451 17057
rect 16393 17048 16405 17051
rect 16163 17020 16405 17048
rect 16163 17017 16175 17020
rect 16117 17011 16175 17017
rect 16393 17017 16405 17020
rect 16439 17048 16451 17051
rect 17034 17048 17040 17060
rect 16439 17020 17040 17048
rect 16439 17017 16451 17020
rect 16393 17011 16451 17017
rect 17034 17008 17040 17020
rect 17092 17008 17098 17060
rect 18141 17051 18199 17057
rect 18141 17017 18153 17051
rect 18187 17017 18199 17051
rect 18141 17011 18199 17017
rect 18233 17051 18291 17057
rect 18233 17017 18245 17051
rect 18279 17048 18291 17051
rect 18322 17048 18328 17060
rect 18279 17020 18328 17048
rect 18279 17017 18291 17020
rect 18233 17011 18291 17017
rect 10928 16952 11008 16980
rect 15749 16983 15807 16989
rect 10928 16940 10934 16952
rect 15749 16949 15761 16983
rect 15795 16980 15807 16983
rect 16298 16980 16304 16992
rect 15795 16952 16304 16980
rect 15795 16949 15807 16952
rect 15749 16943 15807 16949
rect 16298 16940 16304 16952
rect 16356 16980 16362 16992
rect 17310 16980 17316 16992
rect 16356 16952 17316 16980
rect 16356 16940 16362 16952
rect 17310 16940 17316 16952
rect 17368 16980 17374 16992
rect 17405 16983 17463 16989
rect 17405 16980 17417 16983
rect 17368 16952 17417 16980
rect 17368 16940 17374 16952
rect 17405 16949 17417 16952
rect 17451 16949 17463 16983
rect 17770 16980 17776 16992
rect 17731 16952 17776 16980
rect 17405 16943 17463 16949
rect 17770 16940 17776 16952
rect 17828 16980 17834 16992
rect 18156 16980 18184 17011
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 20349 17051 20407 17057
rect 20349 17017 20361 17051
rect 20395 17048 20407 17051
rect 20625 17051 20683 17057
rect 20625 17048 20637 17051
rect 20395 17020 20637 17048
rect 20395 17017 20407 17020
rect 20349 17011 20407 17017
rect 20625 17017 20637 17020
rect 20671 17048 20683 17051
rect 20990 17048 20996 17060
rect 20671 17020 20996 17048
rect 20671 17017 20683 17020
rect 20625 17011 20683 17017
rect 20990 17008 20996 17020
rect 21048 17048 21054 17060
rect 22094 17048 22100 17060
rect 21048 17020 22100 17048
rect 21048 17008 21054 17020
rect 22094 17008 22100 17020
rect 22152 17008 22158 17060
rect 22189 17051 22247 17057
rect 22189 17017 22201 17051
rect 22235 17017 22247 17051
rect 22189 17011 22247 17017
rect 17828 16952 18184 16980
rect 21913 16983 21971 16989
rect 17828 16940 17834 16952
rect 21913 16949 21925 16983
rect 21959 16980 21971 16983
rect 22204 16980 22232 17011
rect 22278 16980 22284 16992
rect 21959 16952 22284 16980
rect 21959 16949 21971 16952
rect 21913 16943 21971 16949
rect 22278 16940 22284 16952
rect 22336 16940 22342 16992
rect 25038 16980 25044 16992
rect 24999 16952 25044 16980
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 13722 16776 13728 16788
rect 13683 16748 13728 16776
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 15654 16776 15660 16788
rect 15615 16748 15660 16776
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 16114 16776 16120 16788
rect 16075 16748 16120 16776
rect 16114 16736 16120 16748
rect 16172 16736 16178 16788
rect 16942 16776 16948 16788
rect 16903 16748 16948 16776
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 17497 16779 17555 16785
rect 17497 16745 17509 16779
rect 17543 16776 17555 16779
rect 17862 16776 17868 16788
rect 17543 16748 17868 16776
rect 17543 16745 17555 16748
rect 17497 16739 17555 16745
rect 17862 16736 17868 16748
rect 17920 16776 17926 16788
rect 18417 16779 18475 16785
rect 18417 16776 18429 16779
rect 17920 16748 18429 16776
rect 17920 16736 17926 16748
rect 18417 16745 18429 16748
rect 18463 16745 18475 16779
rect 20530 16776 20536 16788
rect 20491 16748 20536 16776
rect 18417 16739 18475 16745
rect 20530 16736 20536 16748
rect 20588 16736 20594 16788
rect 22462 16776 22468 16788
rect 22423 16748 22468 16776
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 10226 16668 10232 16720
rect 10284 16708 10290 16720
rect 10597 16711 10655 16717
rect 10597 16708 10609 16711
rect 10284 16680 10609 16708
rect 10284 16668 10290 16680
rect 10597 16677 10609 16680
rect 10643 16708 10655 16711
rect 10686 16708 10692 16720
rect 10643 16680 10692 16708
rect 10643 16677 10655 16680
rect 10597 16671 10655 16677
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 12894 16708 12900 16720
rect 12855 16680 12900 16708
rect 12894 16668 12900 16680
rect 12952 16668 12958 16720
rect 17310 16668 17316 16720
rect 17368 16708 17374 16720
rect 18322 16708 18328 16720
rect 17368 16680 18328 16708
rect 17368 16668 17374 16680
rect 18322 16668 18328 16680
rect 18380 16668 18386 16720
rect 21266 16708 21272 16720
rect 21227 16680 21272 16708
rect 21266 16668 21272 16680
rect 21324 16668 21330 16720
rect 22738 16708 22744 16720
rect 22699 16680 22744 16708
rect 22738 16668 22744 16680
rect 22796 16668 22802 16720
rect 22833 16711 22891 16717
rect 22833 16677 22845 16711
rect 22879 16708 22891 16711
rect 22922 16708 22928 16720
rect 22879 16680 22928 16708
rect 22879 16677 22891 16680
rect 22833 16671 22891 16677
rect 22922 16668 22928 16680
rect 22980 16668 22986 16720
rect 24397 16711 24455 16717
rect 24397 16708 24409 16711
rect 23446 16680 24409 16708
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16640 15531 16643
rect 15562 16640 15568 16652
rect 15519 16612 15568 16640
rect 15519 16609 15531 16612
rect 15473 16603 15531 16609
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16640 16635 16643
rect 16666 16640 16672 16652
rect 16623 16612 16672 16640
rect 16623 16609 16635 16612
rect 16577 16603 16635 16609
rect 16666 16600 16672 16612
rect 16724 16600 16730 16652
rect 19058 16640 19064 16652
rect 19019 16612 19064 16640
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 19242 16640 19248 16652
rect 19203 16612 19248 16640
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 10134 16572 10140 16584
rect 8619 16544 10140 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 10134 16532 10140 16544
rect 10192 16572 10198 16584
rect 10505 16575 10563 16581
rect 10505 16572 10517 16575
rect 10192 16544 10517 16572
rect 10192 16532 10198 16544
rect 10505 16541 10517 16544
rect 10551 16541 10563 16575
rect 11146 16572 11152 16584
rect 11059 16544 11152 16572
rect 10505 16535 10563 16541
rect 11146 16532 11152 16544
rect 11204 16572 11210 16584
rect 11514 16572 11520 16584
rect 11204 16544 11520 16572
rect 11204 16532 11210 16544
rect 11514 16532 11520 16544
rect 11572 16572 11578 16584
rect 12802 16572 12808 16584
rect 11572 16544 12808 16572
rect 11572 16532 11578 16544
rect 12802 16532 12808 16544
rect 12860 16532 12866 16584
rect 13446 16572 13452 16584
rect 13407 16544 13452 16572
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 19518 16572 19524 16584
rect 19479 16544 19524 16572
rect 19518 16532 19524 16544
rect 19576 16532 19582 16584
rect 21174 16572 21180 16584
rect 21135 16544 21180 16572
rect 21174 16532 21180 16544
rect 21232 16572 21238 16584
rect 23017 16575 23075 16581
rect 23017 16572 23029 16575
rect 21232 16544 23029 16572
rect 21232 16532 21238 16544
rect 23017 16541 23029 16544
rect 23063 16541 23075 16575
rect 23017 16535 23075 16541
rect 21726 16504 21732 16516
rect 21687 16476 21732 16504
rect 21726 16464 21732 16476
rect 21784 16464 21790 16516
rect 22278 16464 22284 16516
rect 22336 16504 22342 16516
rect 23446 16504 23474 16680
rect 24397 16677 24409 16680
rect 24443 16708 24455 16711
rect 24670 16708 24676 16720
rect 24443 16680 24676 16708
rect 24443 16677 24455 16680
rect 24397 16671 24455 16677
rect 24670 16668 24676 16680
rect 24728 16668 24734 16720
rect 24946 16708 24952 16720
rect 24907 16680 24952 16708
rect 24946 16668 24952 16680
rect 25004 16668 25010 16720
rect 24305 16575 24363 16581
rect 24305 16541 24317 16575
rect 24351 16541 24363 16575
rect 24305 16535 24363 16541
rect 22336 16476 23474 16504
rect 22336 16464 22342 16476
rect 24210 16464 24216 16516
rect 24268 16504 24274 16516
rect 24320 16504 24348 16535
rect 24268 16476 24348 16504
rect 24268 16464 24274 16476
rect 10226 16436 10232 16448
rect 10187 16408 10232 16436
rect 10226 16396 10232 16408
rect 10284 16396 10290 16448
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 11790 16436 11796 16448
rect 11296 16408 11796 16436
rect 11296 16396 11302 16408
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 18138 16436 18144 16448
rect 18099 16408 18144 16436
rect 18138 16396 18144 16408
rect 18196 16396 18202 16448
rect 22094 16436 22100 16448
rect 22055 16408 22100 16436
rect 22094 16396 22100 16408
rect 22152 16396 22158 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 10134 16232 10140 16244
rect 10095 16204 10140 16232
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 12802 16192 12808 16244
rect 12860 16232 12866 16244
rect 13909 16235 13967 16241
rect 13909 16232 13921 16235
rect 12860 16204 13921 16232
rect 12860 16192 12866 16204
rect 13909 16201 13921 16204
rect 13955 16201 13967 16235
rect 13909 16195 13967 16201
rect 14185 16235 14243 16241
rect 14185 16201 14197 16235
rect 14231 16232 14243 16235
rect 15562 16232 15568 16244
rect 14231 16204 15332 16232
rect 15523 16204 15568 16232
rect 14231 16201 14243 16204
rect 14185 16195 14243 16201
rect 10226 16124 10232 16176
rect 10284 16164 10290 16176
rect 11701 16167 11759 16173
rect 11701 16164 11713 16167
rect 10284 16136 11713 16164
rect 10284 16124 10290 16136
rect 11701 16133 11713 16136
rect 11747 16133 11759 16167
rect 11701 16127 11759 16133
rect 13446 16124 13452 16176
rect 13504 16164 13510 16176
rect 15105 16167 15163 16173
rect 15105 16164 15117 16167
rect 13504 16136 15117 16164
rect 13504 16124 13510 16136
rect 15105 16133 15117 16136
rect 15151 16133 15163 16167
rect 15304 16164 15332 16204
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 16666 16192 16672 16244
rect 16724 16232 16730 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 16724 16204 17417 16232
rect 16724 16192 16730 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 20717 16235 20775 16241
rect 20717 16201 20729 16235
rect 20763 16232 20775 16235
rect 21085 16235 21143 16241
rect 21085 16232 21097 16235
rect 20763 16204 21097 16232
rect 20763 16201 20775 16204
rect 20717 16195 20775 16201
rect 21085 16201 21097 16204
rect 21131 16232 21143 16235
rect 21266 16232 21272 16244
rect 21131 16204 21272 16232
rect 21131 16201 21143 16204
rect 21085 16195 21143 16201
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 22738 16192 22744 16244
rect 22796 16232 22802 16244
rect 23109 16235 23167 16241
rect 23109 16232 23121 16235
rect 22796 16204 23121 16232
rect 22796 16192 22802 16204
rect 23109 16201 23121 16204
rect 23155 16201 23167 16235
rect 24670 16232 24676 16244
rect 24631 16204 24676 16232
rect 23109 16195 23167 16201
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 15841 16167 15899 16173
rect 15841 16164 15853 16167
rect 15304 16136 15853 16164
rect 15105 16127 15163 16133
rect 15841 16133 15853 16136
rect 15887 16164 15899 16167
rect 16206 16164 16212 16176
rect 15887 16136 16212 16164
rect 15887 16133 15899 16136
rect 15841 16127 15899 16133
rect 16206 16124 16212 16136
rect 16264 16124 16270 16176
rect 22833 16167 22891 16173
rect 22833 16133 22845 16167
rect 22879 16164 22891 16167
rect 22922 16164 22928 16176
rect 22879 16136 22928 16164
rect 22879 16133 22891 16136
rect 22833 16127 22891 16133
rect 22922 16124 22928 16136
rect 22980 16124 22986 16176
rect 11057 16099 11115 16105
rect 11057 16065 11069 16099
rect 11103 16096 11115 16099
rect 11146 16096 11152 16108
rect 11103 16068 11152 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 12158 16056 12164 16108
rect 12216 16096 12222 16108
rect 12216 16068 13400 16096
rect 12216 16056 12222 16068
rect 7650 15988 7656 16040
rect 7708 16028 7714 16040
rect 9344 16031 9402 16037
rect 9344 16028 9356 16031
rect 7708 16000 9356 16028
rect 7708 15988 7714 16000
rect 9344 15997 9356 16000
rect 9390 16028 9402 16031
rect 9769 16031 9827 16037
rect 9769 16028 9781 16031
rect 9390 16000 9781 16028
rect 9390 15997 9402 16000
rect 9344 15991 9402 15997
rect 9769 15997 9781 16000
rect 9815 15997 9827 16031
rect 9769 15991 9827 15997
rect 12805 16031 12863 16037
rect 12805 15997 12817 16031
rect 12851 16028 12863 16031
rect 13170 16028 13176 16040
rect 12851 16000 13176 16028
rect 12851 15997 12863 16000
rect 12805 15991 12863 15997
rect 13170 15988 13176 16000
rect 13228 15988 13234 16040
rect 13372 16037 13400 16068
rect 13538 16056 13544 16108
rect 13596 16096 13602 16108
rect 14550 16096 14556 16108
rect 13596 16068 14556 16096
rect 13596 16056 13602 16068
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 14918 16056 14924 16108
rect 14976 16096 14982 16108
rect 16393 16099 16451 16105
rect 16393 16096 16405 16099
rect 14976 16068 16405 16096
rect 14976 16056 14982 16068
rect 16393 16065 16405 16068
rect 16439 16065 16451 16099
rect 16393 16059 16451 16065
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 19797 16099 19855 16105
rect 19797 16096 19809 16099
rect 19576 16068 19809 16096
rect 19576 16056 19582 16068
rect 19797 16065 19809 16068
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 13357 16031 13415 16037
rect 13357 15997 13369 16031
rect 13403 15997 13415 16031
rect 18046 16028 18052 16040
rect 13357 15991 13415 15997
rect 17880 16000 18052 16028
rect 9447 15963 9505 15969
rect 9447 15929 9459 15963
rect 9493 15960 9505 15963
rect 10042 15960 10048 15972
rect 9493 15932 10048 15960
rect 9493 15929 9505 15932
rect 9447 15923 9505 15929
rect 10042 15920 10048 15932
rect 10100 15960 10106 15972
rect 10413 15963 10471 15969
rect 10413 15960 10425 15963
rect 10100 15932 10425 15960
rect 10100 15920 10106 15932
rect 10413 15929 10425 15932
rect 10459 15929 10471 15963
rect 10413 15923 10471 15929
rect 10505 15963 10563 15969
rect 10505 15929 10517 15963
rect 10551 15960 10563 15963
rect 11425 15963 11483 15969
rect 11425 15960 11437 15963
rect 10551 15932 11437 15960
rect 10551 15929 10563 15932
rect 10505 15923 10563 15929
rect 11425 15929 11437 15932
rect 11471 15960 11483 15963
rect 13906 15960 13912 15972
rect 11471 15932 13912 15960
rect 11471 15929 11483 15932
rect 11425 15923 11483 15929
rect 8202 15852 8208 15904
rect 8260 15892 8266 15904
rect 10520 15892 10548 15923
rect 13906 15920 13912 15932
rect 13964 15960 13970 15972
rect 14185 15963 14243 15969
rect 14185 15960 14197 15963
rect 13964 15932 14197 15960
rect 13964 15920 13970 15932
rect 14185 15929 14197 15932
rect 14231 15929 14243 15963
rect 14185 15923 14243 15929
rect 14645 15963 14703 15969
rect 14645 15929 14657 15963
rect 14691 15929 14703 15963
rect 16114 15960 16120 15972
rect 16075 15932 16120 15960
rect 14645 15923 14703 15929
rect 12158 15892 12164 15904
rect 8260 15864 10548 15892
rect 12119 15864 12164 15892
rect 8260 15852 8266 15864
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 13170 15892 13176 15904
rect 13131 15864 13176 15892
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 14274 15892 14280 15904
rect 14235 15864 14280 15892
rect 14274 15852 14280 15864
rect 14332 15892 14338 15904
rect 14660 15892 14688 15923
rect 16114 15920 16120 15932
rect 16172 15920 16178 15972
rect 16206 15920 16212 15972
rect 16264 15960 16270 15972
rect 16264 15932 16309 15960
rect 16264 15920 16270 15932
rect 17880 15904 17908 16000
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 18138 15988 18144 16040
rect 18196 16028 18202 16040
rect 18601 16031 18659 16037
rect 18601 16028 18613 16031
rect 18196 16000 18613 16028
rect 18196 15988 18202 16000
rect 18601 15997 18613 16000
rect 18647 16028 18659 16031
rect 18966 16028 18972 16040
rect 18647 16000 18972 16028
rect 18647 15997 18659 16000
rect 18601 15991 18659 15997
rect 18966 15988 18972 16000
rect 19024 15988 19030 16040
rect 21082 15988 21088 16040
rect 21140 16028 21146 16040
rect 21545 16031 21603 16037
rect 21545 16028 21557 16031
rect 21140 16000 21557 16028
rect 21140 15988 21146 16000
rect 21545 15997 21557 16000
rect 21591 16028 21603 16031
rect 22094 16028 22100 16040
rect 21591 16000 22100 16028
rect 21591 15997 21603 16000
rect 21545 15991 21603 15997
rect 22094 15988 22100 16000
rect 22152 15988 22158 16040
rect 20159 15963 20217 15969
rect 20159 15929 20171 15963
rect 20205 15929 20217 15963
rect 21866 15963 21924 15969
rect 21866 15960 21878 15963
rect 20159 15923 20217 15929
rect 21376 15932 21878 15960
rect 14332 15864 14688 15892
rect 14332 15852 14338 15864
rect 16942 15852 16948 15904
rect 17000 15892 17006 15904
rect 17037 15895 17095 15901
rect 17037 15892 17049 15895
rect 17000 15864 17049 15892
rect 17000 15852 17006 15864
rect 17037 15861 17049 15864
rect 17083 15861 17095 15895
rect 17862 15892 17868 15904
rect 17823 15864 17868 15892
rect 17037 15855 17095 15861
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 18138 15892 18144 15904
rect 18099 15864 18144 15892
rect 18138 15852 18144 15864
rect 18196 15852 18202 15904
rect 19058 15892 19064 15904
rect 19019 15864 19064 15892
rect 19058 15852 19064 15864
rect 19116 15852 19122 15904
rect 19705 15895 19763 15901
rect 19705 15861 19717 15895
rect 19751 15892 19763 15895
rect 20174 15892 20202 15923
rect 20254 15892 20260 15904
rect 19751 15864 20260 15892
rect 19751 15861 19763 15864
rect 19705 15855 19763 15861
rect 20254 15852 20260 15864
rect 20312 15892 20318 15904
rect 21376 15901 21404 15932
rect 21866 15929 21878 15932
rect 21912 15929 21924 15963
rect 21866 15923 21924 15929
rect 21361 15895 21419 15901
rect 21361 15892 21373 15895
rect 20312 15864 21373 15892
rect 20312 15852 20318 15864
rect 21361 15861 21373 15864
rect 21407 15861 21419 15895
rect 22462 15892 22468 15904
rect 22423 15864 22468 15892
rect 21361 15855 21419 15861
rect 22462 15852 22468 15864
rect 22520 15852 22526 15904
rect 24210 15892 24216 15904
rect 24171 15864 24216 15892
rect 24210 15852 24216 15864
rect 24268 15852 24274 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 10042 15688 10048 15700
rect 10003 15660 10048 15688
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 12805 15691 12863 15697
rect 12805 15657 12817 15691
rect 12851 15688 12863 15691
rect 12894 15688 12900 15700
rect 12851 15660 12900 15688
rect 12851 15657 12863 15660
rect 12805 15651 12863 15657
rect 12894 15648 12900 15660
rect 12952 15688 12958 15700
rect 13817 15691 13875 15697
rect 13817 15688 13829 15691
rect 12952 15660 13829 15688
rect 12952 15648 12958 15660
rect 13817 15657 13829 15660
rect 13863 15657 13875 15691
rect 14550 15688 14556 15700
rect 14511 15660 14556 15688
rect 13817 15651 13875 15657
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 15381 15691 15439 15697
rect 15381 15657 15393 15691
rect 15427 15688 15439 15691
rect 17770 15688 17776 15700
rect 15427 15660 17776 15688
rect 15427 15657 15439 15660
rect 15381 15651 15439 15657
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 19242 15688 19248 15700
rect 19203 15660 19248 15688
rect 19242 15648 19248 15660
rect 19300 15648 19306 15700
rect 19518 15648 19524 15700
rect 19576 15688 19582 15700
rect 19797 15691 19855 15697
rect 19797 15688 19809 15691
rect 19576 15660 19809 15688
rect 19576 15648 19582 15660
rect 19797 15657 19809 15660
rect 19843 15657 19855 15691
rect 21174 15688 21180 15700
rect 21135 15660 21180 15688
rect 19797 15651 19855 15657
rect 21174 15648 21180 15660
rect 21232 15648 21238 15700
rect 23109 15691 23167 15697
rect 23109 15657 23121 15691
rect 23155 15688 23167 15691
rect 24210 15688 24216 15700
rect 23155 15660 24216 15688
rect 23155 15657 23167 15660
rect 23109 15651 23167 15657
rect 24210 15648 24216 15660
rect 24268 15648 24274 15700
rect 8202 15620 8208 15632
rect 8163 15592 8208 15620
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 10410 15620 10416 15632
rect 10371 15592 10416 15620
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 13259 15623 13317 15629
rect 13259 15589 13271 15623
rect 13305 15620 13317 15623
rect 13354 15620 13360 15632
rect 13305 15592 13360 15620
rect 13305 15589 13317 15592
rect 13259 15583 13317 15589
rect 13354 15580 13360 15592
rect 13412 15580 13418 15632
rect 15930 15580 15936 15632
rect 15988 15620 15994 15632
rect 16714 15623 16772 15629
rect 16714 15620 16726 15623
rect 15988 15592 16726 15620
rect 15988 15580 15994 15592
rect 16714 15589 16726 15592
rect 16760 15620 16772 15623
rect 16942 15620 16948 15632
rect 16760 15592 16948 15620
rect 16760 15589 16772 15592
rect 16714 15583 16772 15589
rect 16942 15580 16948 15592
rect 17000 15580 17006 15632
rect 17494 15620 17500 15632
rect 17328 15592 17500 15620
rect 11952 15555 12010 15561
rect 11952 15521 11964 15555
rect 11998 15552 12010 15555
rect 12250 15552 12256 15564
rect 11998 15524 12256 15552
rect 11998 15521 12010 15524
rect 11952 15515 12010 15521
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 17328 15561 17356 15592
rect 17494 15580 17500 15592
rect 17552 15620 17558 15632
rect 18325 15623 18383 15629
rect 18325 15620 18337 15623
rect 17552 15592 18337 15620
rect 17552 15580 17558 15592
rect 18325 15589 18337 15592
rect 18371 15589 18383 15623
rect 18325 15583 18383 15589
rect 21634 15580 21640 15632
rect 21692 15620 21698 15632
rect 21729 15623 21787 15629
rect 21729 15620 21741 15623
rect 21692 15592 21741 15620
rect 21692 15580 21698 15592
rect 21729 15589 21741 15592
rect 21775 15620 21787 15623
rect 22462 15620 22468 15632
rect 21775 15592 22468 15620
rect 21775 15589 21787 15592
rect 21729 15583 21787 15589
rect 22462 15580 22468 15592
rect 22520 15580 22526 15632
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15484 8171 15487
rect 8202 15484 8208 15496
rect 8159 15456 8208 15484
rect 8159 15453 8171 15456
rect 8113 15447 8171 15453
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 8389 15487 8447 15493
rect 8389 15484 8401 15487
rect 8352 15456 8401 15484
rect 8352 15444 8358 15456
rect 8389 15453 8401 15456
rect 8435 15484 8447 15487
rect 10321 15487 10379 15493
rect 10321 15484 10333 15487
rect 8435 15456 10333 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 10321 15453 10333 15456
rect 10367 15484 10379 15487
rect 11054 15484 11060 15496
rect 10367 15456 11060 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 11054 15444 11060 15456
rect 11112 15444 11118 15496
rect 12894 15484 12900 15496
rect 12855 15456 12900 15484
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15484 16451 15487
rect 17218 15484 17224 15496
rect 16439 15456 17224 15484
rect 16439 15453 16451 15456
rect 16393 15447 16451 15453
rect 17218 15444 17224 15456
rect 17276 15484 17282 15496
rect 17954 15484 17960 15496
rect 17276 15456 17960 15484
rect 17276 15444 17282 15456
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 18230 15484 18236 15496
rect 18191 15456 18236 15484
rect 18230 15444 18236 15456
rect 18288 15444 18294 15496
rect 18414 15444 18420 15496
rect 18472 15484 18478 15496
rect 18509 15487 18567 15493
rect 18509 15484 18521 15487
rect 18472 15456 18521 15484
rect 18472 15444 18478 15456
rect 18509 15453 18521 15456
rect 18555 15453 18567 15487
rect 18509 15447 18567 15453
rect 21450 15444 21456 15496
rect 21508 15484 21514 15496
rect 21637 15487 21695 15493
rect 21637 15484 21649 15487
rect 21508 15456 21649 15484
rect 21508 15444 21514 15456
rect 21637 15453 21649 15456
rect 21683 15453 21695 15487
rect 21637 15447 21695 15453
rect 21726 15444 21732 15496
rect 21784 15484 21790 15496
rect 22281 15487 22339 15493
rect 22281 15484 22293 15487
rect 21784 15456 22293 15484
rect 21784 15444 21790 15456
rect 22281 15453 22293 15456
rect 22327 15484 22339 15487
rect 22830 15484 22836 15496
rect 22327 15456 22836 15484
rect 22327 15453 22339 15456
rect 22281 15447 22339 15453
rect 22830 15444 22836 15456
rect 22888 15444 22894 15496
rect 10778 15376 10784 15428
rect 10836 15416 10842 15428
rect 10873 15419 10931 15425
rect 10873 15416 10885 15419
rect 10836 15388 10885 15416
rect 10836 15376 10842 15388
rect 10873 15385 10885 15388
rect 10919 15416 10931 15419
rect 13446 15416 13452 15428
rect 10919 15388 13452 15416
rect 10919 15385 10931 15388
rect 10873 15379 10931 15385
rect 13446 15376 13452 15388
rect 13504 15376 13510 15428
rect 15933 15419 15991 15425
rect 15933 15385 15945 15419
rect 15979 15416 15991 15419
rect 16114 15416 16120 15428
rect 15979 15388 16120 15416
rect 15979 15385 15991 15388
rect 15933 15379 15991 15385
rect 16114 15376 16120 15388
rect 16172 15416 16178 15428
rect 20070 15416 20076 15428
rect 16172 15388 20076 15416
rect 16172 15376 16178 15388
rect 20070 15376 20076 15388
rect 20128 15376 20134 15428
rect 12023 15351 12081 15357
rect 12023 15317 12035 15351
rect 12069 15348 12081 15351
rect 12526 15348 12532 15360
rect 12069 15320 12532 15348
rect 12069 15317 12081 15320
rect 12023 15311 12081 15317
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 16206 15348 16212 15360
rect 16167 15320 16212 15348
rect 16206 15308 16212 15320
rect 16264 15308 16270 15360
rect 20438 15348 20444 15360
rect 20399 15320 20444 15348
rect 20438 15308 20444 15320
rect 20496 15308 20502 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 7837 15147 7895 15153
rect 7837 15113 7849 15147
rect 7883 15144 7895 15147
rect 8110 15144 8116 15156
rect 7883 15116 8116 15144
rect 7883 15113 7895 15116
rect 7837 15107 7895 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 10410 15104 10416 15156
rect 10468 15144 10474 15156
rect 10686 15144 10692 15156
rect 10468 15116 10692 15144
rect 10468 15104 10474 15116
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 11054 15144 11060 15156
rect 11015 15116 11060 15144
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 14093 15147 14151 15153
rect 14093 15113 14105 15147
rect 14139 15144 14151 15147
rect 14274 15144 14280 15156
rect 14139 15116 14280 15144
rect 14139 15113 14151 15116
rect 14093 15107 14151 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 15470 15144 15476 15156
rect 15431 15116 15476 15144
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 15841 15147 15899 15153
rect 15841 15144 15853 15147
rect 15804 15116 15853 15144
rect 15804 15104 15810 15116
rect 15841 15113 15853 15116
rect 15887 15113 15899 15147
rect 17494 15144 17500 15156
rect 17455 15116 17500 15144
rect 15841 15107 15899 15113
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 18230 15144 18236 15156
rect 17788 15116 18236 15144
rect 17037 15079 17095 15085
rect 17037 15045 17049 15079
rect 17083 15076 17095 15079
rect 17788 15076 17816 15116
rect 18230 15104 18236 15116
rect 18288 15104 18294 15156
rect 21634 15144 21640 15156
rect 21595 15116 21640 15144
rect 21634 15104 21640 15116
rect 21692 15104 21698 15156
rect 21910 15104 21916 15156
rect 21968 15144 21974 15156
rect 22235 15147 22293 15153
rect 22235 15144 22247 15147
rect 21968 15116 22247 15144
rect 21968 15104 21974 15116
rect 22235 15113 22247 15116
rect 22281 15113 22293 15147
rect 22646 15144 22652 15156
rect 22607 15116 22652 15144
rect 22235 15107 22293 15113
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 19061 15079 19119 15085
rect 19061 15076 19073 15079
rect 17083 15048 17816 15076
rect 18156 15048 19073 15076
rect 17083 15045 17095 15048
rect 17037 15039 17095 15045
rect 8294 15008 8300 15020
rect 8255 14980 8300 15008
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 10134 15008 10140 15020
rect 8864 14980 10140 15008
rect 7101 14875 7159 14881
rect 7101 14841 7113 14875
rect 7147 14872 7159 14875
rect 8018 14872 8024 14884
rect 7147 14844 8024 14872
rect 7147 14841 7159 14844
rect 7101 14835 7159 14841
rect 8018 14832 8024 14844
rect 8076 14832 8082 14884
rect 8113 14875 8171 14881
rect 8113 14841 8125 14875
rect 8159 14872 8171 14875
rect 8864 14872 8892 14980
rect 10134 14968 10140 14980
rect 10192 15008 10198 15020
rect 13170 15008 13176 15020
rect 10192 14980 10456 15008
rect 13131 14980 13176 15008
rect 10192 14968 10198 14980
rect 10428 14949 10456 14980
rect 13170 14968 13176 14980
rect 13228 15008 13234 15020
rect 14737 15011 14795 15017
rect 14737 15008 14749 15011
rect 13228 14980 14749 15008
rect 13228 14968 13234 14980
rect 14737 14977 14749 14980
rect 14783 14977 14795 15011
rect 14737 14971 14795 14977
rect 16206 14968 16212 15020
rect 16264 15008 16270 15020
rect 16485 15011 16543 15017
rect 16485 15008 16497 15011
rect 16264 14980 16497 15008
rect 16264 14968 16270 14980
rect 16485 14977 16497 14980
rect 16531 14977 16543 15011
rect 16485 14971 16543 14977
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18156 15017 18184 15048
rect 19061 15045 19073 15048
rect 19107 15045 19119 15079
rect 19061 15039 19119 15045
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 18012 14980 18153 15008
rect 18012 14968 18018 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18414 15008 18420 15020
rect 18375 14980 18420 15008
rect 18141 14971 18199 14977
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 21450 14968 21456 15020
rect 21508 15008 21514 15020
rect 21913 15011 21971 15017
rect 21913 15008 21925 15011
rect 21508 14980 21925 15008
rect 21508 14968 21514 14980
rect 21913 14977 21925 14980
rect 21959 14977 21971 15011
rect 21913 14971 21971 14977
rect 9493 14943 9551 14949
rect 9493 14940 9505 14943
rect 8159 14844 8892 14872
rect 8956 14912 9505 14940
rect 8159 14841 8171 14844
rect 8113 14835 8171 14841
rect 7469 14807 7527 14813
rect 7469 14773 7481 14807
rect 7515 14804 7527 14807
rect 8128 14804 8156 14835
rect 8956 14816 8984 14912
rect 9493 14909 9505 14912
rect 9539 14909 9551 14943
rect 10413 14943 10471 14949
rect 9493 14903 9551 14909
rect 9692 14912 9858 14940
rect 9692 14816 9720 14912
rect 9830 14881 9858 14912
rect 10413 14909 10425 14943
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 11384 14943 11442 14949
rect 11384 14909 11396 14943
rect 11430 14940 11442 14943
rect 11885 14943 11943 14949
rect 11885 14940 11897 14943
rect 11430 14912 11897 14940
rect 11430 14909 11442 14912
rect 11384 14903 11442 14909
rect 11885 14909 11897 14912
rect 11931 14940 11943 14943
rect 12250 14940 12256 14952
rect 11931 14912 12256 14940
rect 11931 14909 11943 14912
rect 11885 14903 11943 14909
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 14642 14900 14648 14952
rect 14700 14940 14706 14952
rect 15289 14943 15347 14949
rect 15289 14940 15301 14943
rect 14700 14912 15301 14940
rect 14700 14900 14706 14912
rect 15289 14909 15301 14912
rect 15335 14940 15347 14943
rect 15746 14940 15752 14952
rect 15335 14912 15752 14940
rect 15335 14909 15347 14912
rect 15289 14903 15347 14909
rect 15746 14900 15752 14912
rect 15804 14900 15810 14952
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 20349 14943 20407 14949
rect 20349 14940 20361 14943
rect 19392 14912 20361 14940
rect 19392 14900 19398 14912
rect 20349 14909 20361 14912
rect 20395 14940 20407 14943
rect 20438 14940 20444 14952
rect 20395 14912 20444 14940
rect 20395 14909 20407 14912
rect 20349 14903 20407 14909
rect 20438 14900 20444 14912
rect 20496 14900 20502 14952
rect 22164 14943 22222 14949
rect 22164 14909 22176 14943
rect 22210 14940 22222 14943
rect 22646 14940 22652 14952
rect 22210 14912 22652 14940
rect 22210 14909 22222 14912
rect 22164 14903 22222 14909
rect 22646 14900 22652 14912
rect 22704 14940 22710 14952
rect 23290 14940 23296 14952
rect 22704 14912 23296 14940
rect 22704 14900 22710 14912
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 9815 14875 9873 14881
rect 9815 14841 9827 14875
rect 9861 14841 9873 14875
rect 9815 14835 9873 14841
rect 13494 14875 13552 14881
rect 13494 14841 13506 14875
rect 13540 14841 13552 14875
rect 13494 14835 13552 14841
rect 8938 14804 8944 14816
rect 7515 14776 8156 14804
rect 8899 14776 8944 14804
rect 7515 14773 7527 14776
rect 7469 14767 7527 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 9401 14807 9459 14813
rect 9401 14773 9413 14807
rect 9447 14804 9459 14807
rect 9674 14804 9680 14816
rect 9447 14776 9680 14804
rect 9447 14773 9459 14776
rect 9401 14767 9459 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 10042 14764 10048 14816
rect 10100 14804 10106 14816
rect 11471 14807 11529 14813
rect 11471 14804 11483 14807
rect 10100 14776 11483 14804
rect 10100 14764 10106 14776
rect 11471 14773 11483 14776
rect 11517 14773 11529 14807
rect 11471 14767 11529 14773
rect 12989 14807 13047 14813
rect 12989 14773 13001 14807
rect 13035 14804 13047 14807
rect 13354 14804 13360 14816
rect 13035 14776 13360 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 13354 14764 13360 14776
rect 13412 14804 13418 14816
rect 13509 14804 13537 14835
rect 16482 14832 16488 14884
rect 16540 14872 16546 14884
rect 16577 14875 16635 14881
rect 16577 14872 16589 14875
rect 16540 14844 16589 14872
rect 16540 14832 16546 14844
rect 16577 14841 16589 14844
rect 16623 14841 16635 14875
rect 16577 14835 16635 14841
rect 18233 14875 18291 14881
rect 18233 14841 18245 14875
rect 18279 14841 18291 14875
rect 20670 14875 20728 14881
rect 20670 14872 20682 14875
rect 18233 14835 18291 14841
rect 20272 14844 20682 14872
rect 13998 14804 14004 14816
rect 13412 14776 14004 14804
rect 13412 14764 13418 14776
rect 13998 14764 14004 14776
rect 14056 14804 14062 14816
rect 14461 14807 14519 14813
rect 14461 14804 14473 14807
rect 14056 14776 14473 14804
rect 14056 14764 14062 14776
rect 14461 14773 14473 14776
rect 14507 14804 14519 14807
rect 15930 14804 15936 14816
rect 14507 14776 15936 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 15930 14764 15936 14776
rect 15988 14804 15994 14816
rect 16209 14807 16267 14813
rect 16209 14804 16221 14807
rect 15988 14776 16221 14804
rect 15988 14764 15994 14776
rect 16209 14773 16221 14776
rect 16255 14773 16267 14807
rect 16209 14767 16267 14773
rect 17865 14807 17923 14813
rect 17865 14773 17877 14807
rect 17911 14804 17923 14807
rect 18248 14804 18276 14835
rect 20272 14816 20300 14844
rect 20670 14841 20682 14844
rect 20716 14841 20728 14875
rect 20670 14835 20728 14841
rect 18322 14804 18328 14816
rect 17911 14776 18328 14804
rect 17911 14773 17923 14776
rect 17865 14767 17923 14773
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 20254 14804 20260 14816
rect 20215 14776 20260 14804
rect 20254 14764 20260 14776
rect 20312 14764 20318 14816
rect 21269 14807 21327 14813
rect 21269 14773 21281 14807
rect 21315 14804 21327 14807
rect 21818 14804 21824 14816
rect 21315 14776 21824 14804
rect 21315 14773 21327 14776
rect 21269 14767 21327 14773
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 10686 14600 10692 14612
rect 10643 14572 10692 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 11514 14600 11520 14612
rect 11475 14572 11520 14600
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 12529 14603 12587 14609
rect 12529 14569 12541 14603
rect 12575 14600 12587 14603
rect 12710 14600 12716 14612
rect 12575 14572 12716 14600
rect 12575 14569 12587 14572
rect 12529 14563 12587 14569
rect 12710 14560 12716 14572
rect 12768 14600 12774 14612
rect 12894 14600 12900 14612
rect 12768 14572 12900 14600
rect 12768 14560 12774 14572
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 13354 14600 13360 14612
rect 13315 14572 13360 14600
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 13906 14600 13912 14612
rect 13867 14572 13912 14600
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 15930 14560 15936 14612
rect 15988 14600 15994 14612
rect 16025 14603 16083 14609
rect 16025 14600 16037 14603
rect 15988 14572 16037 14600
rect 15988 14560 15994 14572
rect 16025 14569 16037 14572
rect 16071 14569 16083 14603
rect 16025 14563 16083 14569
rect 16482 14560 16488 14612
rect 16540 14600 16546 14612
rect 16850 14600 16856 14612
rect 16540 14572 16856 14600
rect 16540 14560 16546 14572
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 17218 14600 17224 14612
rect 17179 14572 17224 14600
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 17770 14600 17776 14612
rect 17731 14572 17776 14600
rect 17770 14560 17776 14572
rect 17828 14560 17834 14612
rect 18322 14600 18328 14612
rect 18283 14572 18328 14600
rect 18322 14560 18328 14572
rect 18380 14560 18386 14612
rect 21266 14600 21272 14612
rect 21227 14572 21272 14600
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 8757 14535 8815 14541
rect 8757 14501 8769 14535
rect 8803 14532 8815 14535
rect 8938 14532 8944 14544
rect 8803 14504 8944 14532
rect 8803 14501 8815 14504
rect 8757 14495 8815 14501
rect 8938 14492 8944 14504
rect 8996 14492 9002 14544
rect 9766 14492 9772 14544
rect 9824 14532 9830 14544
rect 9998 14535 10056 14541
rect 9998 14532 10010 14535
rect 9824 14504 10010 14532
rect 9824 14492 9830 14504
rect 9998 14501 10010 14504
rect 10044 14501 10056 14535
rect 9998 14495 10056 14501
rect 18230 14492 18236 14544
rect 18288 14532 18294 14544
rect 18601 14535 18659 14541
rect 18601 14532 18613 14535
rect 18288 14504 18613 14532
rect 18288 14492 18294 14504
rect 18601 14501 18613 14504
rect 18647 14501 18659 14535
rect 18601 14495 18659 14501
rect 19889 14535 19947 14541
rect 19889 14501 19901 14535
rect 19935 14532 19947 14535
rect 21082 14532 21088 14544
rect 19935 14504 21088 14532
rect 19935 14501 19947 14504
rect 19889 14495 19947 14501
rect 21082 14492 21088 14504
rect 21140 14492 21146 14544
rect 21818 14492 21824 14544
rect 21876 14532 21882 14544
rect 22833 14535 22891 14541
rect 22833 14532 22845 14535
rect 21876 14504 22845 14532
rect 21876 14492 21882 14504
rect 22833 14501 22845 14504
rect 22879 14532 22891 14535
rect 23014 14532 23020 14544
rect 22879 14504 23020 14532
rect 22879 14501 22891 14504
rect 22833 14495 22891 14501
rect 23014 14492 23020 14504
rect 23072 14492 23078 14544
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 1670 14464 1676 14476
rect 1443 14436 1676 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 1670 14424 1676 14436
rect 1728 14424 1734 14476
rect 8110 14464 8116 14476
rect 8071 14436 8116 14464
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 9122 14464 9128 14476
rect 8619 14436 9128 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 9122 14424 9128 14436
rect 9180 14424 9186 14476
rect 11422 14464 11428 14476
rect 11383 14436 11428 14464
rect 11422 14424 11428 14436
rect 11480 14424 11486 14476
rect 11790 14424 11796 14476
rect 11848 14464 11854 14476
rect 11885 14467 11943 14473
rect 11885 14464 11897 14467
rect 11848 14436 11897 14464
rect 11848 14424 11854 14436
rect 11885 14433 11897 14436
rect 11931 14464 11943 14467
rect 12158 14464 12164 14476
rect 11931 14436 12164 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 12158 14424 12164 14436
rect 12216 14464 12222 14476
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12216 14436 12817 14464
rect 12216 14424 12222 14436
rect 12805 14433 12817 14436
rect 12851 14464 12863 14467
rect 13262 14464 13268 14476
rect 12851 14436 13268 14464
rect 12851 14433 12863 14436
rect 12805 14427 12863 14433
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 15565 14467 15623 14473
rect 15565 14433 15577 14467
rect 15611 14464 15623 14467
rect 15657 14467 15715 14473
rect 15657 14464 15669 14467
rect 15611 14436 15669 14464
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 15657 14433 15669 14436
rect 15703 14464 15715 14467
rect 18138 14464 18144 14476
rect 15703 14436 18144 14464
rect 15703 14433 15715 14436
rect 15657 14427 15715 14433
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 18782 14424 18788 14476
rect 18840 14464 18846 14476
rect 19153 14467 19211 14473
rect 19153 14464 19165 14467
rect 18840 14436 19165 14464
rect 18840 14424 18846 14436
rect 19153 14433 19165 14436
rect 19199 14433 19211 14467
rect 19153 14427 19211 14433
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 19613 14467 19671 14473
rect 19613 14464 19625 14467
rect 19300 14436 19625 14464
rect 19300 14424 19306 14436
rect 19613 14433 19625 14436
rect 19659 14433 19671 14467
rect 19613 14427 19671 14433
rect 9674 14396 9680 14408
rect 9635 14368 9680 14396
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 12250 14356 12256 14408
rect 12308 14396 12314 14408
rect 12989 14399 13047 14405
rect 12989 14396 13001 14399
rect 12308 14368 13001 14396
rect 12308 14356 12314 14368
rect 12989 14365 13001 14368
rect 13035 14396 13047 14399
rect 14458 14396 14464 14408
rect 13035 14368 14464 14396
rect 13035 14365 13047 14368
rect 12989 14359 13047 14365
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 17402 14396 17408 14408
rect 17363 14368 17408 14396
rect 17402 14356 17408 14368
rect 17460 14356 17466 14408
rect 20622 14356 20628 14408
rect 20680 14396 20686 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20680 14368 20913 14396
rect 20680 14356 20686 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 22738 14396 22744 14408
rect 22699 14368 22744 14396
rect 20901 14359 20959 14365
rect 22738 14356 22744 14368
rect 22796 14356 22802 14408
rect 22830 14356 22836 14408
rect 22888 14396 22894 14408
rect 23017 14399 23075 14405
rect 23017 14396 23029 14399
rect 22888 14368 23029 14396
rect 22888 14356 22894 14368
rect 23017 14365 23029 14368
rect 23063 14365 23075 14399
rect 23017 14359 23075 14365
rect 7193 14263 7251 14269
rect 7193 14229 7205 14263
rect 7239 14260 7251 14263
rect 7282 14260 7288 14272
rect 7239 14232 7288 14260
rect 7239 14229 7251 14232
rect 7193 14223 7251 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 7929 14263 7987 14269
rect 7929 14229 7941 14263
rect 7975 14260 7987 14263
rect 8202 14260 8208 14272
rect 7975 14232 8208 14260
rect 7975 14229 7987 14232
rect 7929 14223 7987 14229
rect 8202 14220 8208 14232
rect 8260 14260 8266 14272
rect 9214 14260 9220 14272
rect 8260 14232 9220 14260
rect 8260 14220 8266 14232
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 16577 14263 16635 14269
rect 16577 14229 16589 14263
rect 16623 14260 16635 14263
rect 17218 14260 17224 14272
rect 16623 14232 17224 14260
rect 16623 14229 16635 14232
rect 16577 14223 16635 14229
rect 17218 14220 17224 14232
rect 17276 14220 17282 14272
rect 20162 14260 20168 14272
rect 20123 14232 20168 14260
rect 20162 14220 20168 14232
rect 20220 14220 20226 14272
rect 21821 14263 21879 14269
rect 21821 14229 21833 14263
rect 21867 14260 21879 14263
rect 22278 14260 22284 14272
rect 21867 14232 22284 14260
rect 21867 14229 21879 14232
rect 21821 14223 21879 14229
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 7282 14016 7288 14068
rect 7340 14056 7346 14068
rect 9585 14059 9643 14065
rect 9585 14056 9597 14059
rect 7340 14028 9597 14056
rect 7340 14016 7346 14028
rect 9585 14025 9597 14028
rect 9631 14025 9643 14059
rect 9585 14019 9643 14025
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 9950 14056 9956 14068
rect 9824 14028 9956 14056
rect 9824 14016 9830 14028
rect 9950 14016 9956 14028
rect 10008 14056 10014 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 10008 14028 10057 14056
rect 10008 14016 10014 14028
rect 10045 14025 10057 14028
rect 10091 14056 10103 14059
rect 10410 14056 10416 14068
rect 10091 14028 10416 14056
rect 10091 14025 10103 14028
rect 10045 14019 10103 14025
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 12250 14056 12256 14068
rect 12211 14028 12256 14056
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 17402 14016 17408 14068
rect 17460 14056 17466 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17460 14028 17785 14056
rect 17460 14016 17466 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 20990 14016 20996 14068
rect 21048 14056 21054 14068
rect 21085 14059 21143 14065
rect 21085 14056 21097 14059
rect 21048 14028 21097 14056
rect 21048 14016 21054 14028
rect 21085 14025 21097 14028
rect 21131 14056 21143 14059
rect 21821 14059 21879 14065
rect 21821 14056 21833 14059
rect 21131 14028 21833 14056
rect 21131 14025 21143 14028
rect 21085 14019 21143 14025
rect 21821 14025 21833 14028
rect 21867 14056 21879 14059
rect 22186 14056 22192 14068
rect 21867 14028 22192 14056
rect 21867 14025 21879 14028
rect 21821 14019 21879 14025
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 23014 14056 23020 14068
rect 22975 14028 23020 14056
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 25406 14056 25412 14068
rect 25367 14028 25412 14056
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 11422 13988 11428 14000
rect 10192 13960 11428 13988
rect 10192 13948 10198 13960
rect 11422 13948 11428 13960
rect 11480 13948 11486 14000
rect 14277 13991 14335 13997
rect 14277 13988 14289 13991
rect 14108 13960 14289 13988
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 8294 13920 8300 13932
rect 7883 13892 8300 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 8846 13920 8852 13932
rect 8772 13892 8852 13920
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 8772 13861 8800 13892
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9398 13920 9404 13932
rect 9311 13892 9404 13920
rect 9398 13880 9404 13892
rect 9456 13920 9462 13932
rect 9674 13920 9680 13932
rect 9456 13892 9680 13920
rect 9456 13880 9462 13892
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10686 13920 10692 13932
rect 10275 13892 10692 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10686 13880 10692 13892
rect 10744 13920 10750 13932
rect 11514 13920 11520 13932
rect 10744 13892 11520 13920
rect 10744 13880 10750 13892
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13920 13967 13923
rect 13998 13920 14004 13932
rect 13955 13892 14004 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8260 13824 8585 13852
rect 8260 13812 8266 13824
rect 8573 13821 8585 13824
rect 8619 13852 8631 13855
rect 8757 13855 8815 13861
rect 8757 13852 8769 13855
rect 8619 13824 8769 13852
rect 8619 13821 8631 13824
rect 8573 13815 8631 13821
rect 8757 13821 8769 13824
rect 8803 13821 8815 13855
rect 9122 13852 9128 13864
rect 9083 13824 9128 13852
rect 8757 13815 8815 13821
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13852 9643 13855
rect 10870 13852 10876 13864
rect 9631 13824 10876 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 10870 13812 10876 13824
rect 10928 13852 10934 13864
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 10928 13824 11161 13852
rect 10928 13812 10934 13824
rect 11149 13821 11161 13824
rect 11195 13821 11207 13855
rect 11149 13815 11207 13821
rect 12713 13855 12771 13861
rect 12713 13821 12725 13855
rect 12759 13852 12771 13855
rect 13078 13852 13084 13864
rect 12759 13824 13084 13852
rect 12759 13821 12771 13824
rect 12713 13815 12771 13821
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 13262 13852 13268 13864
rect 13223 13824 13268 13852
rect 13262 13812 13268 13824
rect 13320 13852 13326 13864
rect 13814 13852 13820 13864
rect 13320 13824 13820 13852
rect 13320 13812 13326 13824
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 6641 13787 6699 13793
rect 6641 13753 6653 13787
rect 6687 13784 6699 13787
rect 7190 13784 7196 13796
rect 6687 13756 7196 13784
rect 6687 13753 6699 13756
rect 6641 13747 6699 13753
rect 7190 13744 7196 13756
rect 7248 13744 7254 13796
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 7340 13756 7385 13784
rect 7340 13744 7346 13756
rect 8018 13744 8024 13796
rect 8076 13784 8082 13796
rect 10042 13784 10048 13796
rect 8076 13756 10048 13784
rect 8076 13744 8082 13756
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 10410 13744 10416 13796
rect 10468 13784 10474 13796
rect 10591 13787 10649 13793
rect 10591 13784 10603 13787
rect 10468 13756 10603 13784
rect 10468 13744 10474 13756
rect 10591 13753 10603 13756
rect 10637 13784 10649 13787
rect 13924 13784 13952 13883
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 10637 13756 13952 13784
rect 10637 13753 10649 13756
rect 10591 13747 10649 13753
rect 1670 13716 1676 13728
rect 1631 13688 1676 13716
rect 1670 13676 1676 13688
rect 1728 13676 1734 13728
rect 8110 13716 8116 13728
rect 8071 13688 8116 13716
rect 8110 13676 8116 13688
rect 8168 13676 8174 13728
rect 11790 13716 11796 13728
rect 11751 13688 11796 13716
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 12897 13719 12955 13725
rect 12897 13716 12909 13719
rect 12768 13688 12909 13716
rect 12768 13676 12774 13688
rect 12897 13685 12909 13688
rect 12943 13685 12955 13719
rect 12897 13679 12955 13685
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 14108 13716 14136 13960
rect 14277 13957 14289 13960
rect 14323 13988 14335 13991
rect 20254 13988 20260 14000
rect 14323 13960 14688 13988
rect 20167 13960 20260 13988
rect 14323 13957 14335 13960
rect 14277 13951 14335 13957
rect 14660 13861 14688 13960
rect 20254 13948 20260 13960
rect 20312 13988 20318 14000
rect 21266 13988 21272 14000
rect 20312 13960 21272 13988
rect 20312 13948 20318 13960
rect 21266 13948 21272 13960
rect 21324 13948 21330 14000
rect 22922 13948 22928 14000
rect 22980 13988 22986 14000
rect 23477 13991 23535 13997
rect 23477 13988 23489 13991
rect 22980 13960 23489 13988
rect 22980 13948 22986 13960
rect 23477 13957 23489 13960
rect 23523 13988 23535 13991
rect 23842 13988 23848 14000
rect 23523 13960 23848 13988
rect 23523 13957 23535 13960
rect 23477 13951 23535 13957
rect 23842 13948 23848 13960
rect 23900 13948 23906 14000
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 20162 13920 20168 13932
rect 19300 13892 20168 13920
rect 19300 13880 19306 13892
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 22738 13920 22744 13932
rect 22699 13892 22744 13920
rect 22738 13880 22744 13892
rect 22796 13920 22802 13932
rect 23382 13920 23388 13932
rect 22796 13892 23388 13920
rect 22796 13880 22802 13892
rect 23382 13880 23388 13892
rect 23440 13920 23446 13932
rect 24029 13923 24087 13929
rect 24029 13920 24041 13923
rect 23440 13892 24041 13920
rect 23440 13880 23446 13892
rect 24029 13889 24041 13892
rect 24075 13889 24087 13923
rect 24029 13883 24087 13889
rect 14645 13855 14703 13861
rect 14645 13821 14657 13855
rect 14691 13821 14703 13855
rect 14826 13852 14832 13864
rect 14787 13824 14832 13852
rect 14645 13815 14703 13821
rect 14660 13784 14688 13815
rect 14826 13812 14832 13824
rect 14884 13812 14890 13864
rect 16301 13855 16359 13861
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16347 13824 16681 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 16669 13821 16681 13824
rect 16715 13852 16727 13855
rect 16758 13852 16764 13864
rect 16715 13824 16764 13852
rect 16715 13821 16727 13824
rect 16669 13815 16727 13821
rect 16316 13784 16344 13815
rect 16758 13812 16764 13824
rect 16816 13812 16822 13864
rect 16853 13855 16911 13861
rect 16853 13821 16865 13855
rect 16899 13852 16911 13855
rect 16899 13824 16933 13852
rect 16899 13821 16911 13824
rect 16853 13815 16911 13821
rect 14660 13756 16344 13784
rect 16482 13744 16488 13796
rect 16540 13784 16546 13796
rect 16868 13784 16896 13815
rect 18322 13812 18328 13864
rect 18380 13852 18386 13864
rect 18417 13855 18475 13861
rect 18417 13852 18429 13855
rect 18380 13824 18429 13852
rect 18380 13812 18386 13824
rect 18417 13821 18429 13824
rect 18463 13852 18475 13855
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18463 13824 18613 13852
rect 18463 13821 18475 13824
rect 18417 13815 18475 13821
rect 18601 13821 18613 13824
rect 18647 13821 18659 13855
rect 18601 13815 18659 13821
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 19150 13852 19156 13864
rect 18840 13824 19156 13852
rect 18840 13812 18846 13824
rect 19150 13812 19156 13824
rect 19208 13812 19214 13864
rect 19334 13852 19340 13864
rect 19295 13824 19340 13852
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 24946 13812 24952 13864
rect 25004 13852 25010 13864
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 25004 13824 25237 13852
rect 25004 13812 25010 13824
rect 25225 13821 25237 13824
rect 25271 13852 25283 13855
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 25271 13824 25789 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 25777 13821 25789 13824
rect 25823 13821 25835 13855
rect 25777 13815 25835 13821
rect 16540 13756 16896 13784
rect 17129 13787 17187 13793
rect 16540 13744 16546 13756
rect 17129 13753 17141 13787
rect 17175 13784 17187 13787
rect 20254 13784 20260 13796
rect 17175 13756 20260 13784
rect 17175 13753 17187 13756
rect 17129 13747 17187 13753
rect 20254 13744 20260 13756
rect 20312 13744 20318 13796
rect 20527 13787 20585 13793
rect 20527 13753 20539 13787
rect 20573 13753 20585 13787
rect 22094 13784 22100 13796
rect 22055 13756 22100 13784
rect 20527 13747 20585 13753
rect 14458 13716 14464 13728
rect 13412 13688 14136 13716
rect 14419 13688 14464 13716
rect 13412 13676 13418 13688
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 15749 13719 15807 13725
rect 15749 13685 15761 13719
rect 15795 13716 15807 13719
rect 15838 13716 15844 13728
rect 15795 13688 15844 13716
rect 15795 13685 15807 13688
rect 15749 13679 15807 13685
rect 15838 13676 15844 13688
rect 15896 13716 15902 13728
rect 17405 13719 17463 13725
rect 17405 13716 17417 13719
rect 15896 13688 17417 13716
rect 15896 13676 15902 13688
rect 17405 13685 17417 13688
rect 17451 13716 17463 13719
rect 17770 13716 17776 13728
rect 17451 13688 17776 13716
rect 17451 13685 17463 13688
rect 17405 13679 17463 13685
rect 17770 13676 17776 13688
rect 17828 13676 17834 13728
rect 18690 13676 18696 13728
rect 18748 13716 18754 13728
rect 19613 13719 19671 13725
rect 19613 13716 19625 13719
rect 18748 13688 19625 13716
rect 18748 13676 18754 13688
rect 19613 13685 19625 13688
rect 19659 13685 19671 13719
rect 19613 13679 19671 13685
rect 20073 13719 20131 13725
rect 20073 13685 20085 13719
rect 20119 13716 20131 13719
rect 20542 13716 20570 13747
rect 22094 13744 22100 13756
rect 22152 13744 22158 13796
rect 22186 13744 22192 13796
rect 22244 13784 22250 13796
rect 23753 13787 23811 13793
rect 22244 13756 22289 13784
rect 22244 13744 22250 13756
rect 23753 13753 23765 13787
rect 23799 13753 23811 13787
rect 23753 13747 23811 13753
rect 20714 13716 20720 13728
rect 20119 13688 20720 13716
rect 20119 13685 20131 13688
rect 20073 13679 20131 13685
rect 20714 13676 20720 13688
rect 20772 13716 20778 13728
rect 21266 13716 21272 13728
rect 20772 13688 21272 13716
rect 20772 13676 20778 13688
rect 21266 13676 21272 13688
rect 21324 13716 21330 13728
rect 21361 13719 21419 13725
rect 21361 13716 21373 13719
rect 21324 13688 21373 13716
rect 21324 13676 21330 13688
rect 21361 13685 21373 13688
rect 21407 13685 21419 13719
rect 21361 13679 21419 13685
rect 23658 13676 23664 13728
rect 23716 13716 23722 13728
rect 23768 13716 23796 13747
rect 23842 13744 23848 13796
rect 23900 13784 23906 13796
rect 23900 13756 23945 13784
rect 23900 13744 23906 13756
rect 23716 13688 23796 13716
rect 23716 13676 23722 13688
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 5583 13515 5641 13521
rect 5583 13512 5595 13515
rect 1728 13484 5595 13512
rect 1728 13472 1734 13484
rect 5583 13481 5595 13484
rect 5629 13481 5641 13515
rect 9398 13512 9404 13524
rect 9359 13484 9404 13512
rect 5583 13475 5641 13481
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 10597 13515 10655 13521
rect 10597 13481 10609 13515
rect 10643 13512 10655 13515
rect 10686 13512 10692 13524
rect 10643 13484 10692 13512
rect 10643 13481 10655 13484
rect 10597 13475 10655 13481
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 11422 13472 11428 13524
rect 11480 13512 11486 13524
rect 11480 13484 13537 13512
rect 11480 13472 11486 13484
rect 2774 13404 2780 13456
rect 2832 13444 2838 13456
rect 2832 13416 7087 13444
rect 2832 13404 2838 13416
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1670 13376 1676 13388
rect 1443 13348 1676 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 5445 13379 5503 13385
rect 5445 13345 5457 13379
rect 5491 13376 5503 13379
rect 5534 13376 5540 13388
rect 5491 13348 5540 13376
rect 5491 13345 5503 13348
rect 5445 13339 5503 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 7059 13385 7087 13416
rect 9214 13404 9220 13456
rect 9272 13444 9278 13456
rect 9815 13447 9873 13453
rect 9815 13444 9827 13447
rect 9272 13416 9827 13444
rect 9272 13404 9278 13416
rect 9815 13413 9827 13416
rect 9861 13413 9873 13447
rect 11333 13447 11391 13453
rect 11333 13444 11345 13447
rect 9815 13407 9873 13413
rect 10606 13416 11345 13444
rect 7044 13379 7102 13385
rect 7044 13345 7056 13379
rect 7090 13376 7102 13379
rect 7374 13376 7380 13388
rect 7090 13348 7380 13376
rect 7090 13345 7102 13348
rect 7044 13339 7102 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 8294 13376 8300 13388
rect 8255 13348 8300 13376
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8386 13336 8392 13388
rect 8444 13376 8450 13388
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 8444 13348 8493 13376
rect 8444 13336 8450 13348
rect 8481 13345 8493 13348
rect 8527 13345 8539 13379
rect 9712 13379 9770 13385
rect 9712 13376 9724 13379
rect 8481 13339 8539 13345
rect 8588 13348 9724 13376
rect 7392 13308 7420 13336
rect 8588 13308 8616 13348
rect 9712 13345 9724 13348
rect 9758 13376 9770 13379
rect 10502 13376 10508 13388
rect 9758 13348 10508 13376
rect 9758 13345 9770 13348
rect 9712 13339 9770 13345
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 7392 13280 8616 13308
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13308 8815 13311
rect 9490 13308 9496 13320
rect 8803 13280 9496 13308
rect 8803 13277 8815 13280
rect 8757 13271 8815 13277
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 10606 13308 10634 13416
rect 11333 13413 11345 13416
rect 11379 13444 11391 13447
rect 11882 13444 11888 13456
rect 11379 13416 11888 13444
rect 11379 13413 11391 13416
rect 11333 13407 11391 13413
rect 11882 13404 11888 13416
rect 11940 13404 11946 13456
rect 13509 13444 13537 13484
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14369 13515 14427 13521
rect 14369 13512 14381 13515
rect 13872 13484 14381 13512
rect 13872 13472 13878 13484
rect 14369 13481 14381 13484
rect 14415 13512 14427 13515
rect 14826 13512 14832 13524
rect 14415 13484 14832 13512
rect 14415 13481 14427 13484
rect 14369 13475 14427 13481
rect 14826 13472 14832 13484
rect 14884 13472 14890 13524
rect 19153 13515 19211 13521
rect 19153 13481 19165 13515
rect 19199 13512 19211 13515
rect 19242 13512 19248 13524
rect 19199 13484 19248 13512
rect 19199 13481 19211 13484
rect 19153 13475 19211 13481
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 22557 13515 22615 13521
rect 22557 13481 22569 13515
rect 22603 13512 22615 13515
rect 22603 13484 23428 13512
rect 22603 13481 22615 13484
rect 22557 13475 22615 13481
rect 23400 13456 23428 13484
rect 15562 13444 15568 13456
rect 13509 13416 15568 13444
rect 15562 13404 15568 13416
rect 15620 13444 15626 13456
rect 17218 13444 17224 13456
rect 15620 13416 15976 13444
rect 17179 13416 17224 13444
rect 15620 13404 15626 13416
rect 13078 13376 13084 13388
rect 13039 13348 13084 13376
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 13262 13336 13268 13388
rect 13320 13376 13326 13388
rect 13357 13379 13415 13385
rect 13357 13376 13369 13379
rect 13320 13348 13369 13376
rect 13320 13336 13326 13348
rect 13357 13345 13369 13348
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15746 13376 15752 13388
rect 15436 13348 15752 13376
rect 15436 13336 15442 13348
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 15948 13385 15976 13416
rect 17218 13404 17224 13416
rect 17276 13404 17282 13456
rect 18782 13404 18788 13456
rect 18840 13444 18846 13456
rect 18840 13416 19380 13444
rect 18840 13404 18846 13416
rect 15933 13379 15991 13385
rect 15933 13345 15945 13379
rect 15979 13345 15991 13379
rect 15933 13339 15991 13345
rect 18414 13336 18420 13388
rect 18472 13376 18478 13388
rect 19352 13385 19380 13416
rect 20714 13404 20720 13456
rect 20772 13444 20778 13456
rect 21222 13447 21280 13453
rect 21222 13444 21234 13447
rect 20772 13416 21234 13444
rect 20772 13404 20778 13416
rect 21222 13413 21234 13416
rect 21268 13413 21280 13447
rect 21222 13407 21280 13413
rect 22278 13404 22284 13456
rect 22336 13444 22342 13456
rect 22833 13447 22891 13453
rect 22833 13444 22845 13447
rect 22336 13416 22845 13444
rect 22336 13404 22342 13416
rect 22833 13413 22845 13416
rect 22879 13444 22891 13447
rect 23198 13444 23204 13456
rect 22879 13416 23204 13444
rect 22879 13413 22891 13416
rect 22833 13407 22891 13413
rect 23198 13404 23204 13416
rect 23256 13404 23262 13456
rect 23382 13444 23388 13456
rect 23343 13416 23388 13444
rect 23382 13404 23388 13416
rect 23440 13404 23446 13456
rect 18877 13379 18935 13385
rect 18877 13376 18889 13379
rect 18472 13348 18889 13376
rect 18472 13336 18478 13348
rect 18877 13345 18889 13348
rect 18923 13345 18935 13379
rect 18877 13339 18935 13345
rect 19337 13379 19395 13385
rect 19337 13345 19349 13379
rect 19383 13376 19395 13379
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 19383 13348 19901 13376
rect 19383 13345 19395 13348
rect 19337 13339 19395 13345
rect 19889 13345 19901 13348
rect 19935 13345 19947 13379
rect 19889 13339 19947 13345
rect 20254 13336 20260 13388
rect 20312 13376 20318 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20312 13348 20913 13376
rect 20312 13336 20318 13348
rect 20901 13345 20913 13348
rect 20947 13376 20959 13379
rect 21818 13376 21824 13388
rect 20947 13348 21824 13376
rect 20947 13345 20959 13348
rect 20901 13339 20959 13345
rect 21818 13336 21824 13348
rect 21876 13336 21882 13388
rect 24264 13379 24322 13385
rect 24264 13345 24276 13379
rect 24310 13376 24322 13379
rect 24762 13376 24768 13388
rect 24310 13348 24768 13376
rect 24310 13345 24322 13348
rect 24264 13339 24322 13345
rect 24762 13336 24768 13348
rect 24820 13336 24826 13388
rect 10152 13280 10634 13308
rect 7147 13175 7205 13181
rect 7147 13141 7159 13175
rect 7193 13172 7205 13175
rect 7742 13172 7748 13184
rect 7193 13144 7748 13172
rect 7193 13141 7205 13144
rect 7147 13135 7205 13141
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 7929 13175 7987 13181
rect 7929 13141 7941 13175
rect 7975 13172 7987 13175
rect 9122 13172 9128 13184
rect 7975 13144 9128 13172
rect 7975 13141 7987 13144
rect 7929 13135 7987 13141
rect 9122 13132 9128 13144
rect 9180 13172 9186 13184
rect 9674 13172 9680 13184
rect 9180 13144 9680 13172
rect 9180 13132 9186 13144
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 10152 13181 10180 13280
rect 10870 13268 10876 13320
rect 10928 13308 10934 13320
rect 11241 13311 11299 13317
rect 11241 13308 11253 13311
rect 10928 13280 11253 13308
rect 10928 13268 10934 13280
rect 11241 13277 11253 13280
rect 11287 13277 11299 13311
rect 13446 13308 13452 13320
rect 13407 13280 13452 13308
rect 11241 13271 11299 13277
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 16114 13308 16120 13320
rect 16075 13280 16120 13308
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 17126 13308 17132 13320
rect 17087 13280 17132 13308
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13308 17831 13311
rect 17954 13308 17960 13320
rect 17819 13280 17960 13308
rect 17819 13277 17831 13280
rect 17773 13271 17831 13277
rect 17954 13268 17960 13280
rect 18012 13308 18018 13320
rect 18230 13308 18236 13320
rect 18012 13280 18236 13308
rect 18012 13268 18018 13280
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 22738 13308 22744 13320
rect 22699 13280 22744 13308
rect 22738 13268 22744 13280
rect 22796 13308 22802 13320
rect 24351 13311 24409 13317
rect 24351 13308 24363 13311
rect 22796 13280 24363 13308
rect 22796 13268 22802 13280
rect 24351 13277 24363 13280
rect 24397 13277 24409 13311
rect 24351 13271 24409 13277
rect 11790 13240 11796 13252
rect 11751 13212 11796 13240
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 16666 13200 16672 13252
rect 16724 13240 16730 13252
rect 17678 13240 17684 13252
rect 16724 13212 17684 13240
rect 16724 13200 16730 13212
rect 17678 13200 17684 13212
rect 17736 13240 17742 13252
rect 18690 13240 18696 13252
rect 17736 13212 18696 13240
rect 17736 13200 17742 13212
rect 18690 13200 18696 13212
rect 18748 13200 18754 13252
rect 21821 13243 21879 13249
rect 21821 13209 21833 13243
rect 21867 13240 21879 13243
rect 22922 13240 22928 13252
rect 21867 13212 22928 13240
rect 21867 13209 21879 13212
rect 21821 13203 21879 13209
rect 22922 13200 22928 13212
rect 22980 13200 22986 13252
rect 10137 13175 10195 13181
rect 10137 13172 10149 13175
rect 9824 13144 10149 13172
rect 9824 13132 9830 13144
rect 10137 13141 10149 13144
rect 10183 13141 10195 13175
rect 12710 13172 12716 13184
rect 12671 13144 12716 13172
rect 10137 13135 10195 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 16022 13132 16028 13184
rect 16080 13172 16086 13184
rect 16482 13172 16488 13184
rect 16080 13144 16488 13172
rect 16080 13132 16086 13144
rect 16482 13132 16488 13144
rect 16540 13172 16546 13184
rect 18601 13175 18659 13181
rect 18601 13172 18613 13175
rect 16540 13144 18613 13172
rect 16540 13132 16546 13144
rect 18601 13141 18613 13144
rect 18647 13172 18659 13175
rect 18782 13172 18788 13184
rect 18647 13144 18788 13172
rect 18647 13141 18659 13144
rect 18601 13135 18659 13141
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 20622 13172 20628 13184
rect 20583 13144 20628 13172
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 22186 13172 22192 13184
rect 22147 13144 22192 13172
rect 22186 13132 22192 13144
rect 22244 13132 22250 13184
rect 23658 13172 23664 13184
rect 23619 13144 23664 13172
rect 23658 13132 23664 13144
rect 23716 13132 23722 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7055 12971 7113 12977
rect 7055 12968 7067 12971
rect 6972 12940 7067 12968
rect 6972 12928 6978 12940
rect 7055 12937 7067 12940
rect 7101 12937 7113 12971
rect 7374 12968 7380 12980
rect 7335 12940 7380 12968
rect 7055 12931 7113 12937
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 9033 12971 9091 12977
rect 9033 12968 9045 12971
rect 8352 12940 9045 12968
rect 8352 12928 8358 12940
rect 9033 12937 9045 12940
rect 9079 12968 9091 12971
rect 10134 12968 10140 12980
rect 9079 12940 10140 12968
rect 9079 12937 9091 12940
rect 9033 12931 9091 12937
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 10502 12968 10508 12980
rect 10463 12940 10508 12968
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 11882 12968 11888 12980
rect 11843 12940 11888 12968
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 13078 12928 13084 12980
rect 13136 12968 13142 12980
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 13136 12940 13645 12968
rect 13136 12928 13142 12940
rect 13633 12937 13645 12940
rect 13679 12968 13691 12971
rect 16666 12968 16672 12980
rect 13679 12940 16672 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 16666 12928 16672 12940
rect 16724 12928 16730 12980
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17218 12968 17224 12980
rect 17179 12940 17224 12968
rect 17218 12928 17224 12940
rect 17276 12928 17282 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 18966 12968 18972 12980
rect 18748 12940 18972 12968
rect 18748 12928 18754 12940
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 21818 12968 21824 12980
rect 21779 12940 21824 12968
rect 21818 12928 21824 12940
rect 21876 12928 21882 12980
rect 22186 12928 22192 12980
rect 22244 12968 22250 12980
rect 22511 12971 22569 12977
rect 22511 12968 22523 12971
rect 22244 12940 22523 12968
rect 22244 12928 22250 12940
rect 22511 12937 22523 12940
rect 22557 12937 22569 12971
rect 23198 12968 23204 12980
rect 23159 12940 23204 12968
rect 22511 12931 22569 12937
rect 23198 12928 23204 12940
rect 23256 12928 23262 12980
rect 23658 12928 23664 12980
rect 23716 12968 23722 12980
rect 23799 12971 23857 12977
rect 23799 12968 23811 12971
rect 23716 12940 23811 12968
rect 23716 12928 23722 12940
rect 23799 12937 23811 12940
rect 23845 12937 23857 12971
rect 23799 12931 23857 12937
rect 7190 12860 7196 12912
rect 7248 12900 7254 12912
rect 11195 12903 11253 12909
rect 11195 12900 11207 12903
rect 7248 12872 11207 12900
rect 7248 12860 7254 12872
rect 11195 12869 11207 12872
rect 11241 12869 11253 12903
rect 11195 12863 11253 12869
rect 11514 12860 11520 12912
rect 11572 12900 11578 12912
rect 15470 12900 15476 12912
rect 11572 12872 13032 12900
rect 15383 12872 15476 12900
rect 11572 12860 11578 12872
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 9398 12832 9404 12844
rect 7800 12804 9404 12832
rect 7800 12792 7806 12804
rect 9398 12792 9404 12804
rect 9456 12832 9462 12844
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 9456 12804 9597 12832
rect 9456 12792 9462 12804
rect 9585 12801 9597 12804
rect 9631 12801 9643 12835
rect 10042 12832 10048 12844
rect 10003 12804 10048 12832
rect 9585 12795 9643 12801
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 12526 12792 12532 12844
rect 12584 12832 12590 12844
rect 13004 12841 13032 12872
rect 15470 12860 15476 12872
rect 15528 12900 15534 12912
rect 15746 12900 15752 12912
rect 15528 12872 15752 12900
rect 15528 12860 15534 12872
rect 15746 12860 15752 12872
rect 15804 12900 15810 12912
rect 17862 12900 17868 12912
rect 15804 12872 17868 12900
rect 15804 12860 15810 12872
rect 17862 12860 17868 12872
rect 17920 12900 17926 12912
rect 22646 12900 22652 12912
rect 17920 12872 22652 12900
rect 17920 12860 17926 12872
rect 22646 12860 22652 12872
rect 22704 12860 22710 12912
rect 12713 12835 12771 12841
rect 12713 12832 12725 12835
rect 12584 12804 12725 12832
rect 12584 12792 12590 12804
rect 12713 12801 12725 12804
rect 12759 12801 12771 12835
rect 12713 12795 12771 12801
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 14550 12832 14556 12844
rect 14511 12804 14556 12832
rect 12989 12795 13047 12801
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 17494 12832 17500 12844
rect 15620 12804 17500 12832
rect 15620 12792 15626 12804
rect 17494 12792 17500 12804
rect 17552 12832 17558 12844
rect 18414 12832 18420 12844
rect 17552 12804 18420 12832
rect 17552 12792 17558 12804
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 18598 12792 18604 12844
rect 18656 12832 18662 12844
rect 24811 12835 24869 12841
rect 24811 12832 24823 12835
rect 18656 12804 24823 12832
rect 18656 12792 18662 12804
rect 24811 12801 24823 12804
rect 24857 12801 24869 12835
rect 24811 12795 24869 12801
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 6952 12767 7010 12773
rect 6952 12764 6964 12767
rect 6687 12736 6964 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 6952 12733 6964 12736
rect 6998 12764 7010 12767
rect 7190 12764 7196 12776
rect 6998 12736 7196 12764
rect 6998 12733 7010 12736
rect 6952 12727 7010 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 8202 12764 8208 12776
rect 7883 12736 8208 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 8386 12764 8392 12776
rect 8347 12736 8392 12764
rect 8386 12724 8392 12736
rect 8444 12764 8450 12776
rect 9214 12764 9220 12776
rect 8444 12736 9220 12764
rect 8444 12724 8450 12736
rect 9214 12724 9220 12736
rect 9272 12764 9278 12776
rect 9309 12767 9367 12773
rect 9309 12764 9321 12767
rect 9272 12736 9321 12764
rect 9272 12724 9278 12736
rect 9309 12733 9321 12736
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 11124 12767 11182 12773
rect 11124 12733 11136 12767
rect 11170 12764 11182 12767
rect 15930 12764 15936 12776
rect 11170 12736 11652 12764
rect 15891 12736 15936 12764
rect 11170 12733 11182 12736
rect 11124 12727 11182 12733
rect 5534 12696 5540 12708
rect 5447 12668 5540 12696
rect 5534 12656 5540 12668
rect 5592 12696 5598 12708
rect 8478 12696 8484 12708
rect 5592 12668 8484 12696
rect 5592 12656 5598 12668
rect 8478 12656 8484 12668
rect 8536 12656 8542 12708
rect 8665 12699 8723 12705
rect 8665 12665 8677 12699
rect 8711 12696 8723 12699
rect 9582 12696 9588 12708
rect 8711 12668 9588 12696
rect 8711 12665 8723 12668
rect 8665 12659 8723 12665
rect 9582 12656 9588 12668
rect 9640 12656 9646 12708
rect 9677 12699 9735 12705
rect 9677 12665 9689 12699
rect 9723 12696 9735 12699
rect 9766 12696 9772 12708
rect 9723 12668 9772 12696
rect 9723 12665 9735 12668
rect 9677 12659 9735 12665
rect 9766 12656 9772 12668
rect 9824 12656 9830 12708
rect 11624 12640 11652 12736
rect 15930 12724 15936 12736
rect 15988 12724 15994 12776
rect 18969 12767 19027 12773
rect 18969 12764 18981 12767
rect 18800 12736 18981 12764
rect 12710 12656 12716 12708
rect 12768 12696 12774 12708
rect 12805 12699 12863 12705
rect 12805 12696 12817 12699
rect 12768 12668 12817 12696
rect 12768 12656 12774 12668
rect 12805 12665 12817 12668
rect 12851 12665 12863 12699
rect 14274 12696 14280 12708
rect 14235 12668 14280 12696
rect 12805 12659 12863 12665
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 14369 12699 14427 12705
rect 14369 12665 14381 12699
rect 14415 12665 14427 12699
rect 14369 12659 14427 12665
rect 5721 12631 5779 12637
rect 5721 12597 5733 12631
rect 5767 12628 5779 12631
rect 6270 12628 6276 12640
rect 5767 12600 6276 12628
rect 5767 12597 5779 12600
rect 5721 12591 5779 12597
rect 6270 12588 6276 12600
rect 6328 12588 6334 12640
rect 10870 12628 10876 12640
rect 10831 12600 10876 12628
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 11606 12628 11612 12640
rect 11567 12600 11612 12628
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 14093 12631 14151 12637
rect 14093 12597 14105 12631
rect 14139 12628 14151 12631
rect 14182 12628 14188 12640
rect 14139 12600 14188 12628
rect 14139 12597 14151 12600
rect 14093 12591 14151 12597
rect 14182 12588 14188 12600
rect 14240 12628 14246 12640
rect 14384 12628 14412 12659
rect 15838 12628 15844 12640
rect 14240 12600 14412 12628
rect 15751 12600 15844 12628
rect 14240 12588 14246 12600
rect 15838 12588 15844 12600
rect 15896 12628 15902 12640
rect 16298 12628 16304 12640
rect 15896 12600 16304 12628
rect 15896 12588 15902 12600
rect 16298 12588 16304 12600
rect 16356 12588 16362 12640
rect 17126 12588 17132 12640
rect 17184 12628 17190 12640
rect 17589 12631 17647 12637
rect 17589 12628 17601 12631
rect 17184 12600 17601 12628
rect 17184 12588 17190 12600
rect 17589 12597 17601 12600
rect 17635 12628 17647 12631
rect 18138 12628 18144 12640
rect 17635 12600 18144 12628
rect 17635 12597 17647 12600
rect 17589 12591 17647 12597
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 18690 12588 18696 12640
rect 18748 12628 18754 12640
rect 18800 12637 18828 12736
rect 18969 12733 18981 12736
rect 19015 12733 19027 12767
rect 18969 12727 19027 12733
rect 19242 12724 19248 12776
rect 19300 12764 19306 12776
rect 19429 12767 19487 12773
rect 19429 12764 19441 12767
rect 19300 12736 19441 12764
rect 19300 12724 19306 12736
rect 19429 12733 19441 12736
rect 19475 12733 19487 12767
rect 19429 12727 19487 12733
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12764 19763 12767
rect 20622 12764 20628 12776
rect 19751 12736 20628 12764
rect 19751 12733 19763 12736
rect 19705 12727 19763 12733
rect 20622 12724 20628 12736
rect 20680 12724 20686 12776
rect 22440 12767 22498 12773
rect 22440 12733 22452 12767
rect 22486 12764 22498 12767
rect 23728 12767 23786 12773
rect 22486 12736 22968 12764
rect 22486 12733 22498 12736
rect 22440 12727 22498 12733
rect 20898 12696 20904 12708
rect 20859 12668 20904 12696
rect 20898 12656 20904 12668
rect 20956 12656 20962 12708
rect 20993 12699 21051 12705
rect 20993 12665 21005 12699
rect 21039 12696 21051 12699
rect 21174 12696 21180 12708
rect 21039 12668 21180 12696
rect 21039 12665 21051 12668
rect 20993 12659 21051 12665
rect 21174 12656 21180 12668
rect 21232 12656 21238 12708
rect 21542 12696 21548 12708
rect 21503 12668 21548 12696
rect 21542 12656 21548 12668
rect 21600 12656 21606 12708
rect 18785 12631 18843 12637
rect 18785 12628 18797 12631
rect 18748 12600 18797 12628
rect 18748 12588 18754 12600
rect 18785 12597 18797 12600
rect 18831 12597 18843 12631
rect 20346 12628 20352 12640
rect 20307 12600 20352 12628
rect 18785 12591 18843 12597
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 20622 12628 20628 12640
rect 20583 12600 20628 12628
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 20916 12628 20944 12656
rect 22940 12640 22968 12736
rect 23728 12733 23740 12767
rect 23774 12764 23786 12767
rect 24724 12767 24782 12773
rect 23774 12736 24256 12764
rect 23774 12733 23786 12736
rect 23728 12727 23786 12733
rect 24228 12705 24256 12736
rect 24724 12733 24736 12767
rect 24770 12764 24782 12767
rect 25130 12764 25136 12776
rect 24770 12736 25136 12764
rect 24770 12733 24782 12736
rect 24724 12727 24782 12733
rect 25130 12724 25136 12736
rect 25188 12724 25194 12776
rect 24213 12699 24271 12705
rect 24213 12665 24225 12699
rect 24259 12696 24271 12699
rect 25222 12696 25228 12708
rect 24259 12668 25228 12696
rect 24259 12665 24271 12668
rect 24213 12659 24271 12665
rect 25222 12656 25228 12668
rect 25280 12656 25286 12708
rect 22189 12631 22247 12637
rect 22189 12628 22201 12631
rect 20916 12600 22201 12628
rect 22189 12597 22201 12600
rect 22235 12597 22247 12631
rect 22922 12628 22928 12640
rect 22883 12600 22928 12628
rect 22189 12591 22247 12597
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 24581 12631 24639 12637
rect 24581 12597 24593 12631
rect 24627 12628 24639 12631
rect 24762 12628 24768 12640
rect 24627 12600 24768 12628
rect 24627 12597 24639 12600
rect 24581 12591 24639 12597
rect 24762 12588 24768 12600
rect 24820 12588 24826 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 8665 12427 8723 12433
rect 8665 12424 8677 12427
rect 8444 12396 8677 12424
rect 8444 12384 8450 12396
rect 8665 12393 8677 12396
rect 8711 12393 8723 12427
rect 9398 12424 9404 12436
rect 9359 12396 9404 12424
rect 8665 12387 8723 12393
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 9950 12384 9956 12436
rect 10008 12424 10014 12436
rect 10045 12427 10103 12433
rect 10045 12424 10057 12427
rect 10008 12396 10057 12424
rect 10008 12384 10014 12396
rect 10045 12393 10057 12396
rect 10091 12393 10103 12427
rect 10045 12387 10103 12393
rect 10597 12427 10655 12433
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 11422 12424 11428 12436
rect 10643 12396 11428 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 11422 12384 11428 12396
rect 11480 12424 11486 12436
rect 12526 12424 12532 12436
rect 11480 12396 11652 12424
rect 12487 12396 12532 12424
rect 11480 12384 11486 12396
rect 6178 12316 6184 12368
rect 6236 12356 6242 12368
rect 6273 12359 6331 12365
rect 6273 12356 6285 12359
rect 6236 12328 6285 12356
rect 6236 12316 6242 12328
rect 6273 12325 6285 12328
rect 6319 12325 6331 12359
rect 7834 12356 7840 12368
rect 7795 12328 7840 12356
rect 6273 12319 6331 12325
rect 7834 12316 7840 12328
rect 7892 12316 7898 12368
rect 11624 12365 11652 12396
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 13630 12424 13636 12436
rect 13591 12396 13636 12424
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 15562 12424 15568 12436
rect 15523 12396 15568 12424
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 17034 12424 17040 12436
rect 16995 12396 17040 12424
rect 17034 12384 17040 12396
rect 17092 12424 17098 12436
rect 17770 12424 17776 12436
rect 17092 12396 17776 12424
rect 17092 12384 17098 12396
rect 17770 12384 17776 12396
rect 17828 12424 17834 12436
rect 17828 12396 18092 12424
rect 17828 12384 17834 12396
rect 11609 12359 11667 12365
rect 11609 12325 11621 12359
rect 11655 12325 11667 12359
rect 11609 12319 11667 12325
rect 16298 12316 16304 12368
rect 16356 12356 16362 12368
rect 18064 12365 18092 12396
rect 18138 12384 18144 12436
rect 18196 12424 18202 12436
rect 19567 12427 19625 12433
rect 19567 12424 19579 12427
rect 18196 12396 19579 12424
rect 18196 12384 18202 12396
rect 19567 12393 19579 12396
rect 19613 12393 19625 12427
rect 19567 12387 19625 12393
rect 21542 12384 21548 12436
rect 21600 12424 21606 12436
rect 21818 12424 21824 12436
rect 21600 12396 21824 12424
rect 21600 12384 21606 12396
rect 21818 12384 21824 12396
rect 21876 12424 21882 12436
rect 22189 12427 22247 12433
rect 22189 12424 22201 12427
rect 21876 12396 22201 12424
rect 21876 12384 21882 12396
rect 22189 12393 22201 12396
rect 22235 12393 22247 12427
rect 22189 12387 22247 12393
rect 22649 12427 22707 12433
rect 22649 12393 22661 12427
rect 22695 12424 22707 12427
rect 22738 12424 22744 12436
rect 22695 12396 22744 12424
rect 22695 12393 22707 12396
rect 22649 12387 22707 12393
rect 22738 12384 22744 12396
rect 22796 12384 22802 12436
rect 22833 12427 22891 12433
rect 22833 12393 22845 12427
rect 22879 12393 22891 12427
rect 22833 12387 22891 12393
rect 16438 12359 16496 12365
rect 16438 12356 16450 12359
rect 16356 12328 16450 12356
rect 16356 12316 16362 12328
rect 16438 12325 16450 12328
rect 16484 12325 16496 12359
rect 16438 12319 16496 12325
rect 18049 12359 18107 12365
rect 18049 12325 18061 12359
rect 18095 12325 18107 12359
rect 18049 12319 18107 12325
rect 18782 12316 18788 12368
rect 18840 12356 18846 12368
rect 18877 12359 18935 12365
rect 18877 12356 18889 12359
rect 18840 12328 18889 12356
rect 18840 12316 18846 12328
rect 18877 12325 18889 12328
rect 18923 12356 18935 12359
rect 19242 12356 19248 12368
rect 18923 12328 19248 12356
rect 18923 12325 18935 12328
rect 18877 12319 18935 12325
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 21358 12356 21364 12368
rect 21319 12328 21364 12356
rect 21358 12316 21364 12328
rect 21416 12316 21422 12368
rect 22005 12359 22063 12365
rect 22005 12325 22017 12359
rect 22051 12356 22063 12359
rect 22848 12356 22876 12387
rect 22051 12328 22876 12356
rect 22051 12325 22063 12328
rect 22005 12319 22063 12325
rect 23106 12316 23112 12368
rect 23164 12356 23170 12368
rect 23164 12328 23244 12356
rect 23164 12316 23170 12328
rect 1210 12248 1216 12300
rect 1268 12288 1274 12300
rect 1432 12291 1490 12297
rect 1432 12288 1444 12291
rect 1268 12260 1444 12288
rect 1268 12248 1274 12260
rect 1432 12257 1444 12260
rect 1478 12257 1490 12291
rect 16114 12288 16120 12300
rect 16075 12260 16120 12288
rect 1432 12251 1490 12257
rect 16114 12248 16120 12260
rect 16172 12248 16178 12300
rect 19429 12291 19487 12297
rect 19429 12257 19441 12291
rect 19475 12288 19487 12291
rect 19518 12288 19524 12300
rect 19475 12260 19524 12288
rect 19475 12257 19487 12260
rect 19429 12251 19487 12257
rect 19518 12248 19524 12260
rect 19576 12248 19582 12300
rect 22738 12288 22744 12300
rect 22699 12260 22744 12288
rect 22738 12248 22744 12260
rect 22796 12248 22802 12300
rect 23216 12297 23244 12328
rect 23201 12291 23259 12297
rect 23201 12257 23213 12291
rect 23247 12257 23259 12291
rect 23201 12251 23259 12257
rect 24372 12291 24430 12297
rect 24372 12257 24384 12291
rect 24418 12288 24430 12291
rect 24670 12288 24676 12300
rect 24418 12260 24676 12288
rect 24418 12257 24430 12260
rect 24372 12251 24430 12257
rect 24670 12248 24676 12260
rect 24728 12248 24734 12300
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6270 12220 6276 12232
rect 6227 12192 6276 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 6914 12220 6920 12232
rect 6871 12192 6920 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 6914 12180 6920 12192
rect 6972 12220 6978 12232
rect 7101 12223 7159 12229
rect 7101 12220 7113 12223
rect 6972 12192 7113 12220
rect 6972 12180 6978 12192
rect 7101 12189 7113 12192
rect 7147 12189 7159 12223
rect 7101 12183 7159 12189
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 8202 12220 8208 12232
rect 7791 12192 8208 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 9674 12220 9680 12232
rect 9635 12192 9680 12220
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 11514 12220 11520 12232
rect 10100 12192 11520 12220
rect 10100 12180 10106 12192
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12220 13323 12223
rect 13722 12220 13728 12232
rect 13311 12192 13728 12220
rect 13311 12189 13323 12192
rect 13265 12183 13323 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 17957 12223 18015 12229
rect 17957 12220 17969 12223
rect 17460 12192 17969 12220
rect 17460 12180 17466 12192
rect 17957 12189 17969 12192
rect 18003 12189 18015 12223
rect 18230 12220 18236 12232
rect 18191 12192 18236 12220
rect 17957 12183 18015 12189
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 21266 12220 21272 12232
rect 21227 12192 21272 12220
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12220 21971 12223
rect 22186 12220 22192 12232
rect 21959 12192 22192 12220
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 22186 12180 22192 12192
rect 22244 12180 22250 12232
rect 25130 12220 25136 12232
rect 23308 12192 25136 12220
rect 7466 12112 7472 12164
rect 7524 12152 7530 12164
rect 8297 12155 8355 12161
rect 8297 12152 8309 12155
rect 7524 12124 8309 12152
rect 7524 12112 7530 12124
rect 8297 12121 8309 12124
rect 8343 12121 8355 12155
rect 8297 12115 8355 12121
rect 8478 12112 8484 12164
rect 8536 12152 8542 12164
rect 12069 12155 12127 12161
rect 12069 12152 12081 12155
rect 8536 12124 12081 12152
rect 8536 12112 8542 12124
rect 12069 12121 12081 12124
rect 12115 12152 12127 12155
rect 14550 12152 14556 12164
rect 12115 12124 14556 12152
rect 12115 12121 12127 12124
rect 12069 12115 12127 12121
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 15930 12112 15936 12164
rect 15988 12152 15994 12164
rect 16025 12155 16083 12161
rect 16025 12152 16037 12155
rect 15988 12124 16037 12152
rect 15988 12112 15994 12124
rect 16025 12121 16037 12124
rect 16071 12152 16083 12155
rect 22005 12155 22063 12161
rect 22005 12152 22017 12155
rect 16071 12124 22017 12152
rect 16071 12121 16083 12124
rect 16025 12115 16083 12121
rect 22005 12121 22017 12124
rect 22051 12121 22063 12155
rect 22204 12152 22232 12180
rect 23308 12152 23336 12192
rect 25130 12180 25136 12192
rect 25188 12180 25194 12232
rect 24443 12155 24501 12161
rect 24443 12152 24455 12155
rect 22204 12124 23336 12152
rect 23446 12124 24455 12152
rect 22005 12115 22063 12121
rect 1535 12087 1593 12093
rect 1535 12053 1547 12087
rect 1581 12084 1593 12087
rect 8570 12084 8576 12096
rect 1581 12056 8576 12084
rect 1581 12053 1593 12056
rect 1535 12047 1593 12053
rect 8570 12044 8576 12056
rect 8628 12044 8634 12096
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 12434 12084 12440 12096
rect 9272 12056 12440 12084
rect 9272 12044 9278 12056
rect 12434 12044 12440 12056
rect 12492 12084 12498 12096
rect 12897 12087 12955 12093
rect 12897 12084 12909 12087
rect 12492 12056 12909 12084
rect 12492 12044 12498 12056
rect 12897 12053 12909 12056
rect 12943 12084 12955 12087
rect 13262 12084 13268 12096
rect 12943 12056 13268 12084
rect 12943 12053 12955 12056
rect 12897 12047 12955 12053
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 14185 12087 14243 12093
rect 14185 12084 14197 12087
rect 14056 12056 14197 12084
rect 14056 12044 14062 12056
rect 14185 12053 14197 12056
rect 14231 12053 14243 12087
rect 14185 12047 14243 12053
rect 14274 12044 14280 12096
rect 14332 12084 14338 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 14332 12056 14473 12084
rect 14332 12044 14338 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 19978 12084 19984 12096
rect 19939 12056 19984 12084
rect 14461 12047 14519 12053
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 22094 12044 22100 12096
rect 22152 12084 22158 12096
rect 23446 12084 23474 12124
rect 24443 12121 24455 12124
rect 24489 12121 24501 12155
rect 24443 12115 24501 12121
rect 23750 12084 23756 12096
rect 22152 12056 23474 12084
rect 23711 12056 23756 12084
rect 22152 12044 22158 12056
rect 23750 12044 23756 12056
rect 23808 12044 23814 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1210 11840 1216 11892
rect 1268 11880 1274 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 1268 11852 1593 11880
rect 1268 11840 1274 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 7834 11880 7840 11892
rect 7795 11852 7840 11880
rect 1581 11843 1639 11849
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 8202 11880 8208 11892
rect 8163 11852 8208 11880
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8941 11883 8999 11889
rect 8941 11849 8953 11883
rect 8987 11880 8999 11883
rect 9306 11880 9312 11892
rect 8987 11852 9312 11880
rect 8987 11849 8999 11852
rect 8941 11843 8999 11849
rect 7852 11812 7880 11840
rect 6288 11784 7880 11812
rect 5074 11676 5080 11688
rect 4987 11648 5080 11676
rect 5074 11636 5080 11648
rect 5132 11676 5138 11688
rect 5813 11679 5871 11685
rect 5813 11676 5825 11679
rect 5132 11648 5825 11676
rect 5132 11636 5138 11648
rect 5813 11645 5825 11648
rect 5859 11676 5871 11679
rect 6288 11676 6316 11784
rect 7190 11744 7196 11756
rect 7151 11716 7196 11744
rect 7190 11704 7196 11716
rect 7248 11704 7254 11756
rect 5859 11648 6316 11676
rect 8456 11679 8514 11685
rect 5859 11645 5871 11648
rect 5813 11639 5871 11645
rect 8456 11645 8468 11679
rect 8502 11676 8514 11679
rect 8956 11676 8984 11843
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 9732 11852 10977 11880
rect 9732 11840 9738 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 11422 11880 11428 11892
rect 11383 11852 11428 11880
rect 10965 11843 11023 11849
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11572 11852 11805 11880
rect 11572 11840 11578 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 14182 11880 14188 11892
rect 14143 11852 14188 11880
rect 11793 11843 11851 11849
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 17770 11880 17776 11892
rect 17731 11852 17776 11880
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 20070 11840 20076 11892
rect 20128 11880 20134 11892
rect 23198 11880 23204 11892
rect 20128 11852 23204 11880
rect 20128 11840 20134 11852
rect 23198 11840 23204 11852
rect 23256 11840 23262 11892
rect 23799 11883 23857 11889
rect 23799 11849 23811 11883
rect 23845 11880 23857 11883
rect 24946 11880 24952 11892
rect 23845 11852 24952 11880
rect 23845 11849 23857 11852
rect 23799 11843 23857 11849
rect 24946 11840 24952 11852
rect 25004 11840 25010 11892
rect 9030 11772 9036 11824
rect 9088 11812 9094 11824
rect 15473 11815 15531 11821
rect 15473 11812 15485 11815
rect 9088 11784 15485 11812
rect 9088 11772 9094 11784
rect 15473 11781 15485 11784
rect 15519 11781 15531 11815
rect 19518 11812 19524 11824
rect 19431 11784 19524 11812
rect 15473 11775 15531 11781
rect 19518 11772 19524 11784
rect 19576 11812 19582 11824
rect 24397 11815 24455 11821
rect 24397 11812 24409 11815
rect 19576 11784 24409 11812
rect 19576 11772 19582 11784
rect 24397 11781 24409 11784
rect 24443 11812 24455 11815
rect 24670 11812 24676 11824
rect 24443 11784 24676 11812
rect 24443 11781 24455 11784
rect 24397 11775 24455 11781
rect 24670 11772 24676 11784
rect 24728 11772 24734 11824
rect 25222 11812 25228 11824
rect 25183 11784 25228 11812
rect 25222 11772 25228 11784
rect 25280 11772 25286 11824
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9548 11716 9781 11744
rect 9548 11704 9554 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11744 13323 11747
rect 13446 11744 13452 11756
rect 13311 11716 13452 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 13446 11704 13452 11716
rect 13504 11744 13510 11756
rect 14461 11747 14519 11753
rect 14461 11744 14473 11747
rect 13504 11716 14473 11744
rect 13504 11704 13510 11716
rect 14461 11713 14473 11716
rect 14507 11713 14519 11747
rect 14461 11707 14519 11713
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11744 17187 11747
rect 18230 11744 18236 11756
rect 17175 11716 18236 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 18230 11704 18236 11716
rect 18288 11704 18294 11756
rect 19886 11744 19892 11756
rect 18432 11716 19892 11744
rect 8502 11648 8984 11676
rect 12805 11679 12863 11685
rect 8502 11645 8514 11648
rect 8456 11639 8514 11645
rect 12805 11645 12817 11679
rect 12851 11676 12863 11679
rect 13722 11676 13728 11688
rect 12851 11648 13728 11676
rect 12851 11645 12863 11648
rect 12805 11639 12863 11645
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 15289 11679 15347 11685
rect 15289 11645 15301 11679
rect 15335 11676 15347 11679
rect 15746 11676 15752 11688
rect 15335 11648 15752 11676
rect 15335 11645 15347 11648
rect 15289 11639 15347 11645
rect 15746 11636 15752 11648
rect 15804 11676 15810 11688
rect 15841 11679 15899 11685
rect 15841 11676 15853 11679
rect 15804 11648 15853 11676
rect 15804 11636 15810 11648
rect 15841 11645 15853 11648
rect 15887 11645 15899 11679
rect 18322 11676 18328 11688
rect 18235 11648 18328 11676
rect 15841 11639 15899 11645
rect 18322 11636 18328 11648
rect 18380 11676 18386 11688
rect 18432 11685 18460 11716
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 21818 11744 21824 11756
rect 21779 11716 21824 11744
rect 21818 11704 21824 11716
rect 21876 11704 21882 11756
rect 22186 11744 22192 11756
rect 22147 11716 22192 11744
rect 22186 11704 22192 11716
rect 22244 11704 22250 11756
rect 22738 11744 22744 11756
rect 22699 11716 22744 11744
rect 22738 11704 22744 11716
rect 22796 11704 22802 11756
rect 23106 11744 23112 11756
rect 23067 11716 23112 11744
rect 23106 11704 23112 11716
rect 23164 11704 23170 11756
rect 18417 11679 18475 11685
rect 18417 11676 18429 11679
rect 18380 11648 18429 11676
rect 18380 11636 18386 11648
rect 18417 11645 18429 11648
rect 18463 11645 18475 11679
rect 18417 11639 18475 11645
rect 18506 11636 18512 11688
rect 18564 11676 18570 11688
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 18564 11648 18889 11676
rect 18564 11636 18570 11648
rect 18877 11645 18889 11648
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 19518 11636 19524 11688
rect 19576 11676 19582 11688
rect 19978 11676 19984 11688
rect 19576 11648 19984 11676
rect 19576 11636 19582 11648
rect 19978 11636 19984 11648
rect 20036 11636 20042 11688
rect 20901 11679 20959 11685
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 21545 11679 21603 11685
rect 21545 11676 21557 11679
rect 20947 11648 21557 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 21545 11645 21557 11648
rect 21591 11645 21603 11679
rect 21545 11639 21603 11645
rect 23569 11679 23627 11685
rect 23569 11645 23581 11679
rect 23615 11676 23627 11679
rect 23750 11676 23756 11688
rect 23615 11648 23756 11676
rect 23615 11645 23627 11648
rect 23569 11639 23627 11645
rect 5905 11611 5963 11617
rect 5905 11577 5917 11611
rect 5951 11608 5963 11611
rect 6178 11608 6184 11620
rect 5951 11580 6184 11608
rect 5951 11577 5963 11580
rect 5905 11571 5963 11577
rect 6178 11568 6184 11580
rect 6236 11568 6242 11620
rect 6914 11608 6920 11620
rect 6875 11580 6920 11608
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 7009 11611 7067 11617
rect 7009 11577 7021 11611
rect 7055 11577 7067 11611
rect 9950 11608 9956 11620
rect 7009 11571 7067 11577
rect 9600 11580 9956 11608
rect 6546 11540 6552 11552
rect 6507 11512 6552 11540
rect 6546 11500 6552 11512
rect 6604 11540 6610 11552
rect 7024 11540 7052 11571
rect 6604 11512 7052 11540
rect 6604 11500 6610 11512
rect 7926 11500 7932 11552
rect 7984 11540 7990 11552
rect 8527 11543 8585 11549
rect 8527 11540 8539 11543
rect 7984 11512 8539 11540
rect 7984 11500 7990 11512
rect 8527 11509 8539 11512
rect 8573 11509 8585 11543
rect 9306 11540 9312 11552
rect 9267 11512 9312 11540
rect 8527 11503 8585 11509
rect 9306 11500 9312 11512
rect 9364 11540 9370 11552
rect 9600 11549 9628 11580
rect 9950 11568 9956 11580
rect 10008 11608 10014 11620
rect 10090 11611 10148 11617
rect 10090 11608 10102 11611
rect 10008 11580 10102 11608
rect 10008 11568 10014 11580
rect 10090 11577 10102 11580
rect 10136 11577 10148 11611
rect 10090 11571 10148 11577
rect 13173 11611 13231 11617
rect 13173 11577 13185 11611
rect 13219 11608 13231 11611
rect 13262 11608 13268 11620
rect 13219 11580 13268 11608
rect 13219 11577 13231 11580
rect 13173 11571 13231 11577
rect 13262 11568 13268 11580
rect 13320 11608 13326 11620
rect 13630 11617 13636 11620
rect 13627 11608 13636 11617
rect 13320 11580 13636 11608
rect 13320 11568 13326 11580
rect 13627 11571 13636 11580
rect 13688 11608 13694 11620
rect 16482 11608 16488 11620
rect 13688 11580 16344 11608
rect 16443 11580 16488 11608
rect 13630 11568 13636 11571
rect 13688 11568 13694 11580
rect 16316 11552 16344 11580
rect 16482 11568 16488 11580
rect 16540 11568 16546 11620
rect 16577 11611 16635 11617
rect 16577 11577 16589 11611
rect 16623 11608 16635 11611
rect 16850 11608 16856 11620
rect 16623 11580 16856 11608
rect 16623 11577 16635 11580
rect 16577 11571 16635 11577
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 19150 11608 19156 11620
rect 19111 11580 19156 11608
rect 19150 11568 19156 11580
rect 19208 11568 19214 11620
rect 20302 11611 20360 11617
rect 20302 11577 20314 11611
rect 20348 11608 20360 11611
rect 20622 11608 20628 11620
rect 20348 11580 20628 11608
rect 20348 11577 20360 11580
rect 20302 11571 20360 11577
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9364 11512 9597 11540
rect 9364 11500 9370 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 9824 11512 10701 11540
rect 9824 11500 9830 11512
rect 10689 11509 10701 11512
rect 10735 11509 10747 11543
rect 16298 11540 16304 11552
rect 16259 11512 16304 11540
rect 10689 11503 10747 11509
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 17402 11540 17408 11552
rect 17363 11512 17408 11540
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 19242 11500 19248 11552
rect 19300 11540 19306 11552
rect 19797 11543 19855 11549
rect 19797 11540 19809 11543
rect 19300 11512 19809 11540
rect 19300 11500 19306 11512
rect 19797 11509 19809 11512
rect 19843 11540 19855 11543
rect 20317 11540 20345 11571
rect 20622 11568 20628 11580
rect 20680 11568 20686 11620
rect 19843 11512 20345 11540
rect 19843 11509 19855 11512
rect 19797 11503 19855 11509
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 21177 11543 21235 11549
rect 21177 11540 21189 11543
rect 20864 11512 21189 11540
rect 20864 11500 20870 11512
rect 21177 11509 21189 11512
rect 21223 11540 21235 11543
rect 21358 11540 21364 11552
rect 21223 11512 21364 11540
rect 21223 11509 21235 11512
rect 21177 11503 21235 11509
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 21560 11540 21588 11639
rect 23750 11636 23756 11648
rect 23808 11636 23814 11688
rect 24740 11679 24798 11685
rect 24740 11645 24752 11679
rect 24786 11676 24798 11679
rect 25240 11676 25268 11772
rect 24786 11648 25268 11676
rect 24786 11645 24798 11648
rect 24740 11639 24798 11645
rect 21913 11611 21971 11617
rect 21913 11577 21925 11611
rect 21959 11577 21971 11611
rect 21913 11571 21971 11577
rect 21928 11540 21956 11571
rect 21560 11512 21956 11540
rect 24670 11500 24676 11552
rect 24728 11540 24734 11552
rect 24811 11543 24869 11549
rect 24811 11540 24823 11543
rect 24728 11512 24823 11540
rect 24728 11500 24734 11512
rect 24811 11509 24823 11512
rect 24857 11509 24869 11543
rect 24811 11503 24869 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 6270 11336 6276 11348
rect 6231 11308 6276 11336
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 8527 11339 8585 11345
rect 8527 11336 8539 11339
rect 8260 11308 8539 11336
rect 8260 11296 8266 11308
rect 8527 11305 8539 11308
rect 8573 11305 8585 11339
rect 8527 11299 8585 11305
rect 10091 11339 10149 11345
rect 10091 11305 10103 11339
rect 10137 11336 10149 11339
rect 10870 11336 10876 11348
rect 10137 11308 10876 11336
rect 10137 11305 10149 11308
rect 10091 11299 10149 11305
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 11330 11336 11336 11348
rect 11072 11308 11336 11336
rect 5074 11228 5080 11280
rect 5132 11268 5138 11280
rect 5445 11271 5503 11277
rect 5445 11268 5457 11271
rect 5132 11240 5457 11268
rect 5132 11228 5138 11240
rect 5445 11237 5457 11240
rect 5491 11237 5503 11271
rect 5445 11231 5503 11237
rect 5997 11271 6055 11277
rect 5997 11237 6009 11271
rect 6043 11268 6055 11271
rect 6914 11268 6920 11280
rect 6043 11240 6920 11268
rect 6043 11237 6055 11240
rect 5997 11231 6055 11237
rect 6914 11228 6920 11240
rect 6972 11228 6978 11280
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 7064 11240 7109 11268
rect 7064 11228 7070 11240
rect 9490 11228 9496 11280
rect 9548 11268 9554 11280
rect 10413 11271 10471 11277
rect 10413 11268 10425 11271
rect 9548 11240 10425 11268
rect 9548 11228 9554 11240
rect 10413 11237 10425 11240
rect 10459 11237 10471 11271
rect 11072 11268 11100 11308
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 13262 11336 13268 11348
rect 13223 11308 13268 11336
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 16114 11296 16120 11348
rect 16172 11336 16178 11348
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 16172 11308 16313 11336
rect 16172 11296 16178 11308
rect 16301 11305 16313 11308
rect 16347 11305 16359 11339
rect 16301 11299 16359 11305
rect 16761 11339 16819 11345
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16850 11336 16856 11348
rect 16807 11308 16856 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 19981 11339 20039 11345
rect 19981 11305 19993 11339
rect 20027 11336 20039 11339
rect 20346 11336 20352 11348
rect 20027 11308 20352 11336
rect 20027 11305 20039 11308
rect 19981 11299 20039 11305
rect 20346 11296 20352 11308
rect 20404 11336 20410 11348
rect 20404 11308 21220 11336
rect 20404 11296 20410 11308
rect 21192 11280 21220 11308
rect 10413 11231 10471 11237
rect 10704 11240 11100 11268
rect 11149 11271 11207 11277
rect 10704 11212 10732 11240
rect 11149 11237 11161 11271
rect 11195 11268 11207 11271
rect 11422 11268 11428 11280
rect 11195 11240 11428 11268
rect 11195 11237 11207 11240
rect 11149 11231 11207 11237
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 11701 11271 11759 11277
rect 11701 11237 11713 11271
rect 11747 11268 11759 11271
rect 11790 11268 11796 11280
rect 11747 11240 11796 11268
rect 11747 11237 11759 11240
rect 11701 11231 11759 11237
rect 11790 11228 11796 11240
rect 11848 11268 11854 11280
rect 13541 11271 13599 11277
rect 13541 11268 13553 11271
rect 11848 11240 13553 11268
rect 11848 11228 11854 11240
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11200 4215 11203
rect 4246 11200 4252 11212
rect 4203 11172 4252 11200
rect 4203 11169 4215 11172
rect 4157 11163 4215 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 8478 11200 8484 11212
rect 8435 11172 8484 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 10020 11203 10078 11209
rect 10020 11169 10032 11203
rect 10066 11200 10078 11203
rect 10686 11200 10692 11212
rect 10066 11172 10692 11200
rect 10066 11169 10078 11172
rect 10020 11163 10078 11169
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 4387 11135 4445 11141
rect 4387 11101 4399 11135
rect 4433 11132 4445 11135
rect 4706 11132 4712 11144
rect 4433 11104 4712 11132
rect 4433 11101 4445 11104
rect 4387 11095 4445 11101
rect 4706 11092 4712 11104
rect 4764 11132 4770 11144
rect 5353 11135 5411 11141
rect 5353 11132 5365 11135
rect 4764 11104 5365 11132
rect 4764 11092 4770 11104
rect 5353 11101 5365 11104
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11101 6975 11135
rect 7190 11132 7196 11144
rect 7151 11104 7196 11132
rect 6917 11095 6975 11101
rect 6932 11064 6960 11095
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 11054 11132 11060 11144
rect 11015 11104 11060 11132
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 7466 11064 7472 11076
rect 6932 11036 7472 11064
rect 7466 11024 7472 11036
rect 7524 11024 7530 11076
rect 13372 11064 13400 11240
rect 13541 11237 13553 11240
rect 13587 11237 13599 11271
rect 13541 11231 13599 11237
rect 13633 11271 13691 11277
rect 13633 11237 13645 11271
rect 13679 11268 13691 11271
rect 13998 11268 14004 11280
rect 13679 11240 14004 11268
rect 13679 11237 13691 11240
rect 13633 11231 13691 11237
rect 13998 11228 14004 11240
rect 14056 11228 14062 11280
rect 14185 11271 14243 11277
rect 14185 11237 14197 11271
rect 14231 11268 14243 11271
rect 14550 11268 14556 11280
rect 14231 11240 14556 11268
rect 14231 11237 14243 11240
rect 14185 11231 14243 11237
rect 14550 11228 14556 11240
rect 14608 11228 14614 11280
rect 15470 11268 15476 11280
rect 15431 11240 15476 11268
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 16482 11228 16488 11280
rect 16540 11268 16546 11280
rect 17037 11271 17095 11277
rect 17037 11268 17049 11271
rect 16540 11240 17049 11268
rect 16540 11228 16546 11240
rect 17037 11237 17049 11240
rect 17083 11237 17095 11271
rect 17037 11231 17095 11237
rect 19242 11228 19248 11280
rect 19300 11268 19306 11280
rect 19382 11271 19440 11277
rect 19382 11268 19394 11271
rect 19300 11240 19394 11268
rect 19300 11228 19306 11240
rect 19382 11237 19394 11240
rect 19428 11237 19440 11271
rect 19382 11231 19440 11237
rect 21174 11228 21180 11280
rect 21232 11268 21238 11280
rect 22005 11271 22063 11277
rect 22005 11268 22017 11271
rect 21232 11240 22017 11268
rect 21232 11228 21238 11240
rect 22005 11237 22017 11240
rect 22051 11268 22063 11271
rect 23566 11268 23572 11280
rect 22051 11240 23572 11268
rect 22051 11237 22063 11240
rect 22005 11231 22063 11237
rect 23566 11228 23572 11240
rect 23624 11228 23630 11280
rect 17494 11200 17500 11212
rect 17455 11172 17500 11200
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11200 18107 11203
rect 18506 11200 18512 11212
rect 18095 11172 18512 11200
rect 18095 11169 18107 11172
rect 18049 11163 18107 11169
rect 18506 11160 18512 11172
rect 18564 11160 18570 11212
rect 15378 11132 15384 11144
rect 15339 11104 15384 11132
rect 15378 11092 15384 11104
rect 15436 11092 15442 11144
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11132 18291 11135
rect 19058 11132 19064 11144
rect 18279 11104 19064 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 13372 11036 13814 11064
rect 12986 10996 12992 11008
rect 12947 10968 12992 10996
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 13786 10996 13814 11036
rect 15672 10996 15700 11095
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 21910 11132 21916 11144
rect 21871 11104 21916 11132
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11101 22247 11135
rect 23466 11135 23524 11141
rect 23466 11132 23478 11135
rect 22189 11095 22247 11101
rect 23446 11101 23478 11132
rect 23512 11101 23524 11135
rect 23750 11132 23756 11144
rect 23711 11104 23756 11132
rect 23446 11095 23524 11101
rect 21542 11024 21548 11076
rect 21600 11064 21606 11076
rect 22204 11064 22232 11095
rect 21600 11036 22232 11064
rect 21600 11024 21606 11036
rect 18506 10996 18512 11008
rect 13786 10968 15700 10996
rect 18467 10968 18512 10996
rect 18506 10956 18512 10968
rect 18564 10956 18570 11008
rect 21266 10996 21272 11008
rect 21227 10968 21272 10996
rect 21266 10956 21272 10968
rect 21324 10956 21330 11008
rect 21358 10956 21364 11008
rect 21416 10996 21422 11008
rect 21637 10999 21695 11005
rect 21637 10996 21649 10999
rect 21416 10968 21649 10996
rect 21416 10956 21422 10968
rect 21637 10965 21649 10968
rect 21683 10965 21695 10999
rect 23446 10996 23474 11095
rect 23750 11092 23756 11104
rect 23808 11092 23814 11144
rect 24670 10996 24676 11008
rect 23446 10968 24676 10996
rect 21637 10959 21695 10965
rect 24670 10956 24676 10968
rect 24728 10956 24734 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 4246 10792 4252 10804
rect 4207 10764 4252 10792
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4706 10792 4712 10804
rect 4667 10764 4712 10792
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 5074 10792 5080 10804
rect 5035 10764 5080 10792
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 6178 10752 6184 10804
rect 6236 10792 6242 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 6236 10764 6561 10792
rect 6236 10752 6242 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 7926 10792 7932 10804
rect 7887 10764 7932 10792
rect 6549 10755 6607 10761
rect 6564 10724 6592 10755
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11287 10795 11345 10801
rect 11287 10792 11299 10795
rect 11112 10764 11299 10792
rect 11112 10752 11118 10764
rect 11287 10761 11299 10764
rect 11333 10761 11345 10795
rect 11287 10755 11345 10761
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 11848 10764 12173 10792
rect 11848 10752 11854 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 12161 10755 12219 10761
rect 12575 10795 12633 10801
rect 12575 10761 12587 10795
rect 12621 10792 12633 10795
rect 15378 10792 15384 10804
rect 12621 10764 15384 10792
rect 12621 10761 12633 10764
rect 12575 10755 12633 10761
rect 15378 10752 15384 10764
rect 15436 10792 15442 10804
rect 16393 10795 16451 10801
rect 16393 10792 16405 10795
rect 15436 10764 16405 10792
rect 15436 10752 15442 10764
rect 16393 10761 16405 10764
rect 16439 10761 16451 10795
rect 16393 10755 16451 10761
rect 16482 10752 16488 10804
rect 16540 10792 16546 10804
rect 16715 10795 16773 10801
rect 16715 10792 16727 10795
rect 16540 10764 16727 10792
rect 16540 10752 16546 10764
rect 16715 10761 16727 10764
rect 16761 10761 16773 10795
rect 16715 10755 16773 10761
rect 17218 10752 17224 10804
rect 17276 10792 17282 10804
rect 17494 10792 17500 10804
rect 17276 10764 17500 10792
rect 17276 10752 17282 10764
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 20806 10792 20812 10804
rect 20767 10764 20812 10792
rect 20806 10752 20812 10764
rect 20864 10752 20870 10804
rect 21174 10792 21180 10804
rect 21135 10764 21180 10792
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 21910 10752 21916 10804
rect 21968 10792 21974 10804
rect 22833 10795 22891 10801
rect 22833 10792 22845 10795
rect 21968 10764 22845 10792
rect 21968 10752 21974 10764
rect 22833 10761 22845 10764
rect 22879 10761 22891 10795
rect 22833 10755 22891 10761
rect 23477 10795 23535 10801
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 23566 10792 23572 10804
rect 23523 10764 23572 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 23566 10752 23572 10764
rect 23624 10752 23630 10804
rect 24581 10795 24639 10801
rect 24581 10761 24593 10795
rect 24627 10792 24639 10795
rect 24670 10792 24676 10804
rect 24627 10764 24676 10792
rect 24627 10761 24639 10764
rect 24581 10755 24639 10761
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 7466 10724 7472 10736
rect 6564 10696 6684 10724
rect 7427 10696 7472 10724
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 6546 10656 6552 10668
rect 5951 10628 6552 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10588 5871 10591
rect 5859 10560 6316 10588
rect 5859 10557 5871 10560
rect 5813 10551 5871 10557
rect 6288 10464 6316 10560
rect 6656 10520 6684 10696
rect 7466 10684 7472 10696
rect 7524 10684 7530 10736
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7944 10656 7972 10752
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 13265 10727 13323 10733
rect 13265 10724 13277 10727
rect 12768 10696 13277 10724
rect 12768 10684 12774 10696
rect 13265 10693 13277 10696
rect 13311 10724 13323 10727
rect 13630 10724 13636 10736
rect 13311 10696 13636 10724
rect 13311 10693 13323 10696
rect 13265 10687 13323 10693
rect 13630 10684 13636 10696
rect 13688 10724 13694 10736
rect 15470 10724 15476 10736
rect 13688 10696 15476 10724
rect 13688 10684 13694 10696
rect 15470 10684 15476 10696
rect 15528 10724 15534 10736
rect 16025 10727 16083 10733
rect 16025 10724 16037 10727
rect 15528 10696 16037 10724
rect 15528 10684 15534 10696
rect 16025 10693 16037 10696
rect 16071 10693 16083 10727
rect 16025 10687 16083 10693
rect 8478 10656 8484 10668
rect 6963 10628 7972 10656
rect 8439 10628 8484 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13538 10656 13544 10668
rect 13044 10628 13544 10656
rect 13044 10616 13050 10628
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 13722 10616 13728 10668
rect 13780 10656 13786 10668
rect 15565 10659 15623 10665
rect 15565 10656 15577 10659
rect 13780 10628 15577 10656
rect 13780 10616 13786 10628
rect 15565 10625 15577 10628
rect 15611 10625 15623 10659
rect 18782 10656 18788 10668
rect 18743 10628 18788 10656
rect 15565 10619 15623 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 19150 10616 19156 10668
rect 19208 10656 19214 10668
rect 19889 10659 19947 10665
rect 19889 10656 19901 10659
rect 19208 10628 19901 10656
rect 19208 10616 19214 10628
rect 19889 10625 19901 10628
rect 19935 10656 19947 10659
rect 20162 10656 20168 10668
rect 19935 10628 20168 10656
rect 19935 10625 19947 10628
rect 19889 10619 19947 10625
rect 20162 10616 20168 10628
rect 20220 10616 20226 10668
rect 11216 10591 11274 10597
rect 11216 10557 11228 10591
rect 11262 10588 11274 10591
rect 11606 10588 11612 10600
rect 11262 10560 11612 10588
rect 11262 10557 11274 10560
rect 11216 10551 11274 10557
rect 11606 10548 11612 10560
rect 11664 10588 11670 10600
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 11664 10560 11713 10588
rect 11664 10548 11670 10560
rect 11701 10557 11713 10560
rect 11747 10588 11759 10591
rect 11790 10588 11796 10600
rect 11747 10560 11796 10588
rect 11747 10557 11759 10560
rect 11701 10551 11759 10557
rect 11790 10548 11796 10560
rect 11848 10548 11854 10600
rect 12504 10591 12562 10597
rect 12504 10557 12516 10591
rect 12550 10588 12562 10591
rect 15013 10591 15071 10597
rect 12550 10560 13032 10588
rect 12550 10557 12562 10560
rect 12504 10551 12562 10557
rect 7009 10523 7067 10529
rect 7009 10520 7021 10523
rect 6656 10492 7021 10520
rect 7009 10489 7021 10492
rect 7055 10489 7067 10523
rect 9677 10523 9735 10529
rect 9677 10520 9689 10523
rect 7009 10483 7067 10489
rect 9048 10492 9689 10520
rect 9048 10464 9076 10492
rect 9677 10489 9689 10492
rect 9723 10489 9735 10523
rect 9677 10483 9735 10489
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 10321 10523 10379 10529
rect 9824 10492 9917 10520
rect 9824 10480 9830 10492
rect 10321 10489 10333 10523
rect 10367 10520 10379 10523
rect 11514 10520 11520 10532
rect 10367 10492 11520 10520
rect 10367 10489 10379 10492
rect 10321 10483 10379 10489
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 6270 10452 6276 10464
rect 6231 10424 6276 10452
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 9030 10452 9036 10464
rect 8991 10424 9036 10452
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 9784 10452 9812 10480
rect 10686 10452 10692 10464
rect 9539 10424 9812 10452
rect 10647 10424 10692 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 11057 10455 11115 10461
rect 11057 10421 11069 10455
rect 11103 10452 11115 10455
rect 11422 10452 11428 10464
rect 11103 10424 11428 10452
rect 11103 10421 11115 10424
rect 11057 10415 11115 10421
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 13004 10461 13032 10560
rect 15013 10557 15025 10591
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 13630 10520 13636 10532
rect 13591 10492 13636 10520
rect 13630 10480 13636 10492
rect 13688 10480 13694 10532
rect 14182 10520 14188 10532
rect 14143 10492 14188 10520
rect 14182 10480 14188 10492
rect 14240 10480 14246 10532
rect 14921 10523 14979 10529
rect 14921 10489 14933 10523
rect 14967 10520 14979 10523
rect 15028 10520 15056 10551
rect 15102 10548 15108 10600
rect 15160 10588 15166 10600
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 15160 10560 15485 10588
rect 15160 10548 15166 10560
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 16644 10591 16702 10597
rect 16644 10557 16656 10591
rect 16690 10588 16702 10591
rect 16690 10560 17172 10588
rect 16690 10557 16702 10560
rect 16644 10551 16702 10557
rect 15562 10520 15568 10532
rect 14967 10492 15568 10520
rect 14967 10489 14979 10492
rect 14921 10483 14979 10489
rect 15562 10480 15568 10492
rect 15620 10480 15626 10532
rect 17144 10464 17172 10560
rect 21358 10548 21364 10600
rect 21416 10588 21422 10600
rect 21637 10591 21695 10597
rect 21637 10588 21649 10591
rect 21416 10560 21649 10588
rect 21416 10548 21422 10560
rect 21637 10557 21649 10560
rect 21683 10557 21695 10591
rect 21637 10551 21695 10557
rect 22922 10548 22928 10600
rect 22980 10588 22986 10600
rect 23712 10591 23770 10597
rect 23712 10588 23724 10591
rect 22980 10560 23724 10588
rect 22980 10548 22986 10560
rect 23712 10557 23724 10560
rect 23758 10588 23770 10591
rect 23758 10560 24256 10588
rect 23758 10557 23770 10560
rect 23712 10551 23770 10557
rect 24228 10532 24256 10560
rect 18138 10520 18144 10532
rect 18099 10492 18144 10520
rect 18138 10480 18144 10492
rect 18196 10480 18202 10532
rect 18233 10523 18291 10529
rect 18233 10489 18245 10523
rect 18279 10520 18291 10523
rect 18322 10520 18328 10532
rect 18279 10492 18328 10520
rect 18279 10489 18291 10492
rect 18233 10483 18291 10489
rect 12989 10455 13047 10461
rect 12989 10421 13001 10455
rect 13035 10452 13047 10455
rect 13078 10452 13084 10464
rect 13035 10424 13084 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 13078 10412 13084 10424
rect 13136 10412 13142 10464
rect 13998 10412 14004 10464
rect 14056 10452 14062 10464
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 14056 10424 14473 10452
rect 14056 10412 14062 10424
rect 14461 10421 14473 10424
rect 14507 10421 14519 10455
rect 17126 10452 17132 10464
rect 17087 10424 17132 10452
rect 14461 10415 14519 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17865 10455 17923 10461
rect 17865 10421 17877 10455
rect 17911 10452 17923 10455
rect 18248 10452 18276 10483
rect 18322 10480 18328 10492
rect 18380 10480 18386 10532
rect 20251 10523 20309 10529
rect 20251 10489 20263 10523
rect 20297 10489 20309 10523
rect 21958 10523 22016 10529
rect 21958 10520 21970 10523
rect 20251 10483 20309 10489
rect 21468 10492 21970 10520
rect 17911 10424 18276 10452
rect 19153 10455 19211 10461
rect 17911 10421 17923 10424
rect 17865 10415 17923 10421
rect 19153 10421 19165 10455
rect 19199 10452 19211 10455
rect 19242 10452 19248 10464
rect 19199 10424 19248 10452
rect 19199 10421 19211 10424
rect 19153 10415 19211 10421
rect 19242 10412 19248 10424
rect 19300 10452 19306 10464
rect 19705 10455 19763 10461
rect 19705 10452 19717 10455
rect 19300 10424 19717 10452
rect 19300 10412 19306 10424
rect 19705 10421 19717 10424
rect 19751 10452 19763 10455
rect 20266 10452 20294 10483
rect 21468 10461 21496 10492
rect 21958 10489 21970 10492
rect 22004 10489 22016 10523
rect 21958 10483 22016 10489
rect 23382 10480 23388 10532
rect 23440 10520 23446 10532
rect 23799 10523 23857 10529
rect 23799 10520 23811 10523
rect 23440 10492 23811 10520
rect 23440 10480 23446 10492
rect 23799 10489 23811 10492
rect 23845 10489 23857 10523
rect 24210 10520 24216 10532
rect 24171 10492 24216 10520
rect 23799 10483 23857 10489
rect 24210 10480 24216 10492
rect 24268 10480 24274 10532
rect 21453 10455 21511 10461
rect 21453 10452 21465 10455
rect 19751 10424 21465 10452
rect 19751 10421 19763 10424
rect 19705 10415 19763 10421
rect 21453 10421 21465 10424
rect 21499 10421 21511 10455
rect 22554 10452 22560 10464
rect 22515 10424 22560 10452
rect 21453 10415 21511 10421
rect 22554 10412 22560 10424
rect 22612 10412 22618 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10248 5319 10251
rect 6270 10248 6276 10260
rect 5307 10220 6276 10248
rect 5307 10217 5319 10220
rect 5261 10211 5319 10217
rect 6270 10208 6276 10220
rect 6328 10208 6334 10260
rect 6825 10251 6883 10257
rect 6825 10217 6837 10251
rect 6871 10248 6883 10251
rect 7282 10248 7288 10260
rect 6871 10220 7288 10248
rect 6871 10217 6883 10220
rect 6825 10211 6883 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 7524 10220 7665 10248
rect 7524 10208 7530 10220
rect 7653 10217 7665 10220
rect 7699 10217 7711 10251
rect 7653 10211 7711 10217
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 11054 10248 11060 10260
rect 8619 10220 10685 10248
rect 11015 10220 11060 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 9858 10180 9864 10192
rect 9819 10152 9864 10180
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 10657 10180 10685 10220
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 12434 10248 12440 10260
rect 12395 10220 12440 10248
rect 12434 10208 12440 10220
rect 12492 10248 12498 10260
rect 12986 10248 12992 10260
rect 12492 10220 12992 10248
rect 12492 10208 12498 10220
rect 12986 10208 12992 10220
rect 13044 10248 13050 10260
rect 13044 10220 13400 10248
rect 13044 10208 13050 10220
rect 11330 10180 11336 10192
rect 10657 10152 11336 10180
rect 11330 10140 11336 10152
rect 11388 10140 11394 10192
rect 11422 10140 11428 10192
rect 11480 10180 11486 10192
rect 13262 10189 13268 10192
rect 13259 10180 13268 10189
rect 11480 10152 11525 10180
rect 13223 10152 13268 10180
rect 11480 10140 11486 10152
rect 13259 10143 13268 10152
rect 13262 10140 13268 10143
rect 13320 10140 13326 10192
rect 13372 10180 13400 10220
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13817 10251 13875 10257
rect 13817 10248 13829 10251
rect 13688 10220 13829 10248
rect 13688 10208 13694 10220
rect 13817 10217 13829 10220
rect 13863 10217 13875 10251
rect 15102 10248 15108 10260
rect 15063 10220 15108 10248
rect 13817 10211 13875 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 16114 10248 16120 10260
rect 15620 10220 16120 10248
rect 15620 10208 15626 10220
rect 16114 10208 16120 10220
rect 16172 10248 16178 10260
rect 16172 10220 17540 10248
rect 16172 10208 16178 10220
rect 15120 10180 15148 10208
rect 16022 10180 16028 10192
rect 13372 10152 15148 10180
rect 15983 10152 16028 10180
rect 16022 10140 16028 10152
rect 16080 10140 16086 10192
rect 17037 10183 17095 10189
rect 17037 10149 17049 10183
rect 17083 10180 17095 10183
rect 17310 10180 17316 10192
rect 17083 10152 17316 10180
rect 17083 10149 17095 10152
rect 17037 10143 17095 10149
rect 17310 10140 17316 10152
rect 17368 10140 17374 10192
rect 17512 10180 17540 10220
rect 19058 10208 19064 10260
rect 19116 10248 19122 10260
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 19116 10220 19809 10248
rect 19116 10208 19122 10220
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 20162 10248 20168 10260
rect 20123 10220 20168 10248
rect 19797 10211 19855 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 23014 10208 23020 10260
rect 23072 10248 23078 10260
rect 23750 10248 23756 10260
rect 23072 10220 23756 10248
rect 23072 10208 23078 10220
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 19334 10180 19340 10192
rect 17512 10152 19340 10180
rect 19076 10124 19104 10152
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 19521 10183 19579 10189
rect 19521 10149 19533 10183
rect 19567 10180 19579 10183
rect 21358 10180 21364 10192
rect 19567 10152 21364 10180
rect 19567 10149 19579 10152
rect 19521 10143 19579 10149
rect 21358 10140 21364 10152
rect 21416 10140 21422 10192
rect 21634 10180 21640 10192
rect 21547 10152 21640 10180
rect 21634 10140 21640 10152
rect 21692 10180 21698 10192
rect 22554 10180 22560 10192
rect 21692 10152 22560 10180
rect 21692 10140 21698 10152
rect 22554 10140 22560 10152
rect 22612 10140 22618 10192
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 7834 10112 7840 10124
rect 7423 10084 7840 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 14182 10112 14188 10124
rect 11992 10084 14188 10112
rect 6454 10044 6460 10056
rect 6415 10016 6460 10044
rect 6454 10004 6460 10016
rect 6512 10004 6518 10056
rect 9769 10047 9827 10053
rect 9769 10013 9781 10047
rect 9815 10013 9827 10047
rect 10042 10044 10048 10056
rect 10003 10016 10048 10044
rect 9769 10007 9827 10013
rect 4430 9936 4436 9988
rect 4488 9976 4494 9988
rect 9784 9976 9812 10007
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 11514 10004 11520 10056
rect 11572 10044 11578 10056
rect 11609 10047 11667 10053
rect 11609 10044 11621 10047
rect 11572 10016 11621 10044
rect 11572 10004 11578 10016
rect 11609 10013 11621 10016
rect 11655 10044 11667 10047
rect 11992 10044 12020 10084
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 14277 10115 14335 10121
rect 14277 10081 14289 10115
rect 14323 10112 14335 10115
rect 15286 10112 15292 10124
rect 14323 10084 15292 10112
rect 14323 10081 14335 10084
rect 14277 10075 14335 10081
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 15562 10112 15568 10124
rect 15523 10084 15568 10112
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 19058 10112 19064 10124
rect 19019 10084 19064 10112
rect 19058 10072 19064 10084
rect 19116 10072 19122 10124
rect 19150 10072 19156 10124
rect 19208 10112 19214 10124
rect 19245 10115 19303 10121
rect 19245 10112 19257 10115
rect 19208 10084 19257 10112
rect 19208 10072 19214 10084
rect 19245 10081 19257 10084
rect 19291 10081 19303 10115
rect 19245 10075 19303 10081
rect 22186 10072 22192 10124
rect 22244 10112 22250 10124
rect 23106 10112 23112 10124
rect 22244 10084 22289 10112
rect 23067 10084 23112 10112
rect 22244 10072 22250 10084
rect 23106 10072 23112 10084
rect 23164 10072 23170 10124
rect 12894 10044 12900 10056
rect 11655 10016 12020 10044
rect 12855 10016 12900 10044
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 16942 10044 16948 10056
rect 13786 10016 15700 10044
rect 16903 10016 16948 10044
rect 10686 9976 10692 9988
rect 4488 9948 10692 9976
rect 4488 9936 4494 9948
rect 10686 9936 10692 9948
rect 10744 9936 10750 9988
rect 11974 9936 11980 9988
rect 12032 9976 12038 9988
rect 13786 9976 13814 10016
rect 15378 9976 15384 9988
rect 12032 9948 13814 9976
rect 15339 9948 15384 9976
rect 12032 9936 12038 9948
rect 15378 9936 15384 9948
rect 15436 9936 15442 9988
rect 15672 9976 15700 10016
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17586 10044 17592 10056
rect 17547 10016 17592 10044
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 21542 10044 21548 10056
rect 21503 10016 21548 10044
rect 21542 10004 21548 10016
rect 21600 10004 21606 10056
rect 23017 10047 23075 10053
rect 23017 10044 23029 10047
rect 21652 10016 23029 10044
rect 18138 9976 18144 9988
rect 15672 9948 18144 9976
rect 18138 9936 18144 9948
rect 18196 9976 18202 9988
rect 18233 9979 18291 9985
rect 18233 9976 18245 9979
rect 18196 9948 18245 9976
rect 18196 9936 18202 9948
rect 18233 9945 18245 9948
rect 18279 9945 18291 9979
rect 18233 9939 18291 9945
rect 18322 9936 18328 9988
rect 18380 9976 18386 9988
rect 21652 9976 21680 10016
rect 23017 10013 23029 10016
rect 23063 10013 23075 10047
rect 23017 10007 23075 10013
rect 18380 9948 21680 9976
rect 18380 9936 18386 9948
rect 8110 9868 8116 9920
rect 8168 9908 8174 9920
rect 12158 9908 12164 9920
rect 8168 9880 12164 9908
rect 8168 9868 8174 9880
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 14550 9908 14556 9920
rect 14511 9880 14556 9908
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 17957 9911 18015 9917
rect 17957 9877 17969 9911
rect 18003 9908 18015 9911
rect 18506 9908 18512 9920
rect 18003 9880 18512 9908
rect 18003 9877 18015 9880
rect 17957 9871 18015 9877
rect 18506 9868 18512 9880
rect 18564 9908 18570 9920
rect 19150 9908 19156 9920
rect 18564 9880 19156 9908
rect 18564 9868 18570 9880
rect 19150 9868 19156 9880
rect 19208 9868 19214 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 6270 9664 6276 9716
rect 6328 9704 6334 9716
rect 7006 9704 7012 9716
rect 6328 9676 7012 9704
rect 6328 9664 6334 9676
rect 7006 9664 7012 9676
rect 7064 9704 7070 9716
rect 7745 9707 7803 9713
rect 7745 9704 7757 9707
rect 7064 9676 7757 9704
rect 7064 9664 7070 9676
rect 7745 9673 7757 9676
rect 7791 9673 7803 9707
rect 7745 9667 7803 9673
rect 9033 9707 9091 9713
rect 9033 9673 9045 9707
rect 9079 9704 9091 9707
rect 9858 9704 9864 9716
rect 9079 9676 9864 9704
rect 9079 9673 9091 9676
rect 9033 9667 9091 9673
rect 9858 9664 9864 9676
rect 9916 9704 9922 9716
rect 10413 9707 10471 9713
rect 10413 9704 10425 9707
rect 9916 9676 10425 9704
rect 9916 9664 9922 9676
rect 10413 9673 10425 9676
rect 10459 9704 10471 9707
rect 11149 9707 11207 9713
rect 11149 9704 11161 9707
rect 10459 9676 11161 9704
rect 10459 9673 10471 9676
rect 10413 9667 10471 9673
rect 11149 9673 11161 9676
rect 11195 9673 11207 9707
rect 11149 9667 11207 9673
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 9217 9639 9275 9645
rect 9217 9636 9229 9639
rect 7340 9608 9229 9636
rect 7340 9596 7346 9608
rect 9217 9605 9229 9608
rect 9263 9636 9275 9639
rect 9306 9636 9312 9648
rect 9263 9608 9312 9636
rect 9263 9605 9275 9608
rect 9217 9599 9275 9605
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 10686 9636 10692 9648
rect 10647 9608 10692 9636
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 11164 9636 11192 9667
rect 11330 9664 11336 9716
rect 11388 9704 11394 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11388 9676 11805 9704
rect 11388 9664 11394 9676
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 12158 9704 12164 9716
rect 12119 9676 12164 9704
rect 11793 9667 11851 9673
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 13320 9676 13461 9704
rect 13320 9664 13326 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 13449 9667 13507 9673
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 16301 9707 16359 9713
rect 16301 9704 16313 9707
rect 15344 9676 16313 9704
rect 15344 9664 15350 9676
rect 16301 9673 16313 9676
rect 16347 9673 16359 9707
rect 16301 9667 16359 9673
rect 16623 9707 16681 9713
rect 16623 9673 16635 9707
rect 16669 9704 16681 9707
rect 17402 9704 17408 9716
rect 16669 9676 17408 9704
rect 16669 9673 16681 9676
rect 16623 9667 16681 9673
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 18690 9704 18696 9716
rect 17512 9676 18696 9704
rect 11422 9636 11428 9648
rect 11164 9608 11428 9636
rect 11422 9596 11428 9608
rect 11480 9596 11486 9648
rect 1670 9528 1676 9580
rect 1728 9568 1734 9580
rect 9030 9568 9036 9580
rect 1728 9540 9036 9568
rect 1728 9528 1734 9540
rect 9030 9528 9036 9540
rect 9088 9528 9094 9580
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11974 9568 11980 9580
rect 11379 9540 11980 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12176 9568 12204 9664
rect 17512 9636 17540 9676
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 21634 9704 21640 9716
rect 21595 9676 21640 9704
rect 21634 9664 21640 9676
rect 21692 9664 21698 9716
rect 21910 9664 21916 9716
rect 21968 9704 21974 9716
rect 22235 9707 22293 9713
rect 22235 9704 22247 9707
rect 21968 9676 22247 9704
rect 21968 9664 21974 9676
rect 22235 9673 22247 9676
rect 22281 9673 22293 9707
rect 22646 9704 22652 9716
rect 22607 9676 22652 9704
rect 22235 9667 22293 9673
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 23106 9704 23112 9716
rect 23067 9676 23112 9704
rect 23106 9664 23112 9676
rect 23164 9664 23170 9716
rect 13786 9608 17540 9636
rect 12176 9540 12480 9568
rect 12452 9509 12480 9540
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 8665 9503 8723 9509
rect 6871 9472 8156 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 6273 9435 6331 9441
rect 6273 9401 6285 9435
rect 6319 9432 6331 9435
rect 6641 9435 6699 9441
rect 6641 9432 6653 9435
rect 6319 9404 6653 9432
rect 6319 9401 6331 9404
rect 6273 9395 6331 9401
rect 6641 9401 6653 9404
rect 6687 9432 6699 9435
rect 7187 9435 7245 9441
rect 7187 9432 7199 9435
rect 6687 9404 7199 9432
rect 6687 9401 6699 9404
rect 6641 9395 6699 9401
rect 7187 9401 7199 9404
rect 7233 9432 7245 9435
rect 7282 9432 7288 9444
rect 7233 9404 7288 9432
rect 7233 9401 7245 9404
rect 7187 9395 7245 9401
rect 7282 9392 7288 9404
rect 7340 9392 7346 9444
rect 8128 9376 8156 9472
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 9493 9503 9551 9509
rect 9493 9500 9505 9503
rect 8711 9472 9505 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 9493 9469 9505 9472
rect 9539 9500 9551 9503
rect 12437 9503 12495 9509
rect 9539 9472 12296 9500
rect 9539 9469 9551 9472
rect 9493 9463 9551 9469
rect 9217 9435 9275 9441
rect 9217 9401 9229 9435
rect 9263 9432 9275 9435
rect 9814 9435 9872 9441
rect 9814 9432 9826 9435
rect 9263 9404 9826 9432
rect 9263 9401 9275 9404
rect 9217 9395 9275 9401
rect 9814 9401 9826 9404
rect 9860 9401 9872 9435
rect 9814 9395 9872 9401
rect 5902 9364 5908 9376
rect 5863 9336 5908 9364
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 8110 9364 8116 9376
rect 8071 9336 8116 9364
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 12268 9364 12296 9472
rect 12437 9469 12449 9503
rect 12483 9469 12495 9503
rect 12986 9500 12992 9512
rect 12947 9472 12992 9500
rect 12437 9463 12495 9469
rect 12452 9432 12480 9463
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 13786 9432 13814 9608
rect 18598 9596 18604 9648
rect 18656 9636 18662 9648
rect 24719 9639 24777 9645
rect 24719 9636 24731 9639
rect 18656 9608 24731 9636
rect 18656 9596 18662 9608
rect 24719 9605 24731 9608
rect 24765 9605 24777 9639
rect 24719 9599 24777 9605
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 17644 9540 18153 9568
rect 17644 9528 17650 9540
rect 18141 9537 18153 9540
rect 18187 9537 18199 9571
rect 18782 9568 18788 9580
rect 18743 9540 18788 9568
rect 18141 9531 18199 9537
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 23106 9568 23112 9580
rect 19720 9540 23112 9568
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 14550 9500 14556 9512
rect 14507 9472 14556 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 14550 9460 14556 9472
rect 14608 9460 14614 9512
rect 14921 9503 14979 9509
rect 14921 9469 14933 9503
rect 14967 9469 14979 9503
rect 15194 9500 15200 9512
rect 15155 9472 15200 9500
rect 14921 9463 14979 9469
rect 12452 9404 13814 9432
rect 14093 9435 14151 9441
rect 14093 9401 14105 9435
rect 14139 9432 14151 9435
rect 14936 9432 14964 9463
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 15381 9503 15439 9509
rect 15381 9469 15393 9503
rect 15427 9469 15439 9503
rect 15381 9463 15439 9469
rect 16552 9503 16610 9509
rect 16552 9469 16564 9503
rect 16598 9469 16610 9503
rect 16552 9463 16610 9469
rect 15286 9432 15292 9444
rect 14139 9404 15292 9432
rect 14139 9401 14151 9404
rect 14093 9395 14151 9401
rect 15286 9392 15292 9404
rect 15344 9392 15350 9444
rect 12529 9367 12587 9373
rect 12529 9364 12541 9367
rect 12268 9336 12541 9364
rect 12529 9333 12541 9336
rect 12575 9333 12587 9367
rect 12529 9327 12587 9333
rect 13538 9324 13544 9376
rect 13596 9364 13602 9376
rect 14642 9364 14648 9376
rect 13596 9336 14648 9364
rect 13596 9324 13602 9336
rect 14642 9324 14648 9336
rect 14700 9364 14706 9376
rect 15396 9364 15424 9463
rect 15654 9432 15660 9444
rect 15615 9404 15660 9432
rect 15654 9392 15660 9404
rect 15712 9392 15718 9444
rect 14700 9336 15424 9364
rect 14700 9324 14706 9336
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 15933 9367 15991 9373
rect 15933 9364 15945 9367
rect 15620 9336 15945 9364
rect 15620 9324 15626 9336
rect 15933 9333 15945 9336
rect 15979 9333 15991 9367
rect 16567 9364 16595 9463
rect 16666 9392 16672 9444
rect 16724 9432 16730 9444
rect 17865 9435 17923 9441
rect 17865 9432 17877 9435
rect 16724 9404 17877 9432
rect 16724 9392 16730 9404
rect 17865 9401 17877 9404
rect 17911 9432 17923 9435
rect 18233 9435 18291 9441
rect 18233 9432 18245 9435
rect 17911 9404 18245 9432
rect 17911 9401 17923 9404
rect 17865 9395 17923 9401
rect 18233 9401 18245 9404
rect 18279 9432 18291 9435
rect 19720 9432 19748 9540
rect 23106 9528 23112 9540
rect 23164 9528 23170 9580
rect 23198 9528 23204 9580
rect 23256 9568 23262 9580
rect 23934 9568 23940 9580
rect 23256 9540 23940 9568
rect 23256 9528 23262 9540
rect 23934 9528 23940 9540
rect 23992 9528 23998 9580
rect 22002 9460 22008 9512
rect 22060 9500 22066 9512
rect 22164 9503 22222 9509
rect 22164 9500 22176 9503
rect 22060 9472 22176 9500
rect 22060 9460 22066 9472
rect 22164 9469 22176 9472
rect 22210 9500 22222 9503
rect 22646 9500 22652 9512
rect 22210 9472 22652 9500
rect 22210 9469 22222 9472
rect 22164 9463 22222 9469
rect 22646 9460 22652 9472
rect 22704 9460 22710 9512
rect 24648 9503 24706 9509
rect 24648 9469 24660 9503
rect 24694 9500 24706 9503
rect 24694 9472 25176 9500
rect 24694 9469 24706 9472
rect 24648 9463 24706 9469
rect 20622 9432 20628 9444
rect 18279 9404 19748 9432
rect 20583 9404 20628 9432
rect 18279 9401 18291 9404
rect 18233 9395 18291 9401
rect 20622 9392 20628 9404
rect 20680 9392 20686 9444
rect 20714 9392 20720 9444
rect 20772 9432 20778 9444
rect 21266 9432 21272 9444
rect 20772 9404 20817 9432
rect 21179 9404 21272 9432
rect 20772 9392 20778 9404
rect 21266 9392 21272 9404
rect 21324 9432 21330 9444
rect 23014 9432 23020 9444
rect 21324 9404 23020 9432
rect 21324 9392 21330 9404
rect 23014 9392 23020 9404
rect 23072 9392 23078 9444
rect 17034 9364 17040 9376
rect 16567 9336 17040 9364
rect 15933 9327 15991 9333
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 17310 9364 17316 9376
rect 17271 9336 17316 9364
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 19058 9364 19064 9376
rect 19019 9336 19064 9364
rect 19058 9324 19064 9336
rect 19116 9324 19122 9376
rect 19150 9324 19156 9376
rect 19208 9364 19214 9376
rect 19429 9367 19487 9373
rect 19429 9364 19441 9367
rect 19208 9336 19441 9364
rect 19208 9324 19214 9336
rect 19429 9333 19441 9336
rect 19475 9333 19487 9367
rect 19429 9327 19487 9333
rect 20441 9367 20499 9373
rect 20441 9333 20453 9367
rect 20487 9364 20499 9367
rect 20732 9364 20760 9392
rect 25148 9376 25176 9472
rect 20487 9336 20760 9364
rect 20487 9333 20499 9336
rect 20441 9327 20499 9333
rect 21542 9324 21548 9376
rect 21600 9364 21606 9376
rect 22005 9367 22063 9373
rect 22005 9364 22017 9367
rect 21600 9336 22017 9364
rect 21600 9324 21606 9336
rect 22005 9333 22017 9336
rect 22051 9364 22063 9367
rect 22186 9364 22192 9376
rect 22051 9336 22192 9364
rect 22051 9333 22063 9336
rect 22005 9327 22063 9333
rect 22186 9324 22192 9336
rect 22244 9324 22250 9376
rect 25130 9364 25136 9376
rect 25091 9336 25136 9364
rect 25130 9324 25136 9336
rect 25188 9324 25194 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 5902 9120 5908 9172
rect 5960 9160 5966 9172
rect 6454 9160 6460 9172
rect 5960 9132 6460 9160
rect 5960 9120 5966 9132
rect 6454 9120 6460 9132
rect 6512 9160 6518 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6512 9132 6745 9160
rect 6512 9120 6518 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 11149 9163 11207 9169
rect 11149 9129 11161 9163
rect 11195 9160 11207 9163
rect 11238 9160 11244 9172
rect 11195 9132 11244 9160
rect 11195 9129 11207 9132
rect 11149 9123 11207 9129
rect 11238 9120 11244 9132
rect 11296 9120 11302 9172
rect 12894 9160 12900 9172
rect 12855 9132 12900 9160
rect 12894 9120 12900 9132
rect 12952 9160 12958 9172
rect 13265 9163 13323 9169
rect 13265 9160 13277 9163
rect 12952 9132 13277 9160
rect 12952 9120 12958 9132
rect 13265 9129 13277 9132
rect 13311 9129 13323 9163
rect 13265 9123 13323 9129
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9160 14335 9163
rect 14642 9160 14648 9172
rect 14323 9132 14648 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 14642 9120 14648 9132
rect 14700 9160 14706 9172
rect 15378 9160 15384 9172
rect 14700 9132 15384 9160
rect 14700 9120 14706 9132
rect 15378 9120 15384 9132
rect 15436 9160 15442 9172
rect 15473 9163 15531 9169
rect 15473 9160 15485 9163
rect 15436 9132 15485 9160
rect 15436 9120 15442 9132
rect 15473 9129 15485 9132
rect 15519 9129 15531 9163
rect 15473 9123 15531 9129
rect 16577 9163 16635 9169
rect 16577 9129 16589 9163
rect 16623 9160 16635 9163
rect 16666 9160 16672 9172
rect 16623 9132 16672 9160
rect 16623 9129 16635 9132
rect 16577 9123 16635 9129
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 21174 9120 21180 9172
rect 21232 9160 21238 9172
rect 21269 9163 21327 9169
rect 21269 9160 21281 9163
rect 21232 9132 21281 9160
rect 21232 9120 21238 9132
rect 21269 9129 21281 9132
rect 21315 9129 21327 9163
rect 21269 9123 21327 9129
rect 5813 9095 5871 9101
rect 5813 9061 5825 9095
rect 5859 9092 5871 9095
rect 6086 9092 6092 9104
rect 5859 9064 6092 9092
rect 5859 9061 5871 9064
rect 5813 9055 5871 9061
rect 6086 9052 6092 9064
rect 6144 9052 6150 9104
rect 12986 9052 12992 9104
rect 13044 9092 13050 9104
rect 13044 9064 13676 9092
rect 13044 9052 13050 9064
rect 5074 9024 5080 9036
rect 5035 8996 5080 9024
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5166 8984 5172 9036
rect 5224 9024 5230 9036
rect 5353 9027 5411 9033
rect 5353 9024 5365 9027
rect 5224 8996 5365 9024
rect 5224 8984 5230 8996
rect 5353 8993 5365 8996
rect 5399 8993 5411 9027
rect 5353 8987 5411 8993
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 6822 9024 6828 9036
rect 6227 8996 6828 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7374 9024 7380 9036
rect 7335 8996 7380 9024
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 7650 9024 7656 9036
rect 7611 8996 7656 9024
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 8018 9024 8024 9036
rect 7979 8996 8024 9024
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 9896 9027 9954 9033
rect 9896 8993 9908 9027
rect 9942 8993 9954 9027
rect 11146 9024 11152 9036
rect 11107 8996 11152 9024
rect 9896 8987 9954 8993
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8956 6607 8959
rect 7668 8956 7696 8984
rect 6595 8928 7696 8956
rect 6595 8925 6607 8928
rect 6549 8919 6607 8925
rect 5169 8891 5227 8897
rect 5169 8857 5181 8891
rect 5215 8888 5227 8891
rect 5534 8888 5540 8900
rect 5215 8860 5540 8888
rect 5215 8857 5227 8860
rect 5169 8851 5227 8857
rect 5534 8848 5540 8860
rect 5592 8848 5598 8900
rect 8481 8891 8539 8897
rect 8481 8857 8493 8891
rect 8527 8888 8539 8891
rect 9911 8888 9939 8987
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 11609 9027 11667 9033
rect 11609 8993 11621 9027
rect 11655 9024 11667 9027
rect 11790 9024 11796 9036
rect 11655 8996 11796 9024
rect 11655 8993 11667 8996
rect 11609 8987 11667 8993
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 11885 9027 11943 9033
rect 11885 8993 11897 9027
rect 11931 9024 11943 9027
rect 11974 9024 11980 9036
rect 11931 8996 11980 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 12250 9024 12256 9036
rect 12211 8996 12256 9024
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 13354 9024 13360 9036
rect 13315 8996 13360 9024
rect 13354 8984 13360 8996
rect 13412 8984 13418 9036
rect 13648 9033 13676 9064
rect 14366 9052 14372 9104
rect 14424 9092 14430 9104
rect 14550 9092 14556 9104
rect 14424 9064 14556 9092
rect 14424 9052 14430 9064
rect 14550 9052 14556 9064
rect 14608 9092 14614 9104
rect 14921 9095 14979 9101
rect 14921 9092 14933 9095
rect 14608 9064 14933 9092
rect 14608 9052 14614 9064
rect 14921 9061 14933 9064
rect 14967 9061 14979 9095
rect 14921 9055 14979 9061
rect 16019 9095 16077 9101
rect 16019 9061 16031 9095
rect 16065 9092 16077 9095
rect 16298 9092 16304 9104
rect 16065 9064 16304 9092
rect 16065 9061 16077 9064
rect 16019 9055 16077 9061
rect 16298 9052 16304 9064
rect 16356 9052 16362 9104
rect 17494 9052 17500 9104
rect 17552 9092 17558 9104
rect 17589 9095 17647 9101
rect 17589 9092 17601 9095
rect 17552 9064 17601 9092
rect 17552 9052 17558 9064
rect 17589 9061 17601 9064
rect 17635 9061 17647 9095
rect 22830 9092 22836 9104
rect 17589 9055 17647 9061
rect 21836 9064 22836 9092
rect 13633 9027 13691 9033
rect 13633 8993 13645 9027
rect 13679 8993 13691 9027
rect 15654 9024 15660 9036
rect 15615 8996 15660 9024
rect 13633 8987 13691 8993
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 18690 8984 18696 9036
rect 18748 9024 18754 9036
rect 19061 9027 19119 9033
rect 19061 9024 19073 9027
rect 18748 8996 19073 9024
rect 18748 8984 18754 8996
rect 19061 8993 19073 8996
rect 19107 8993 19119 9027
rect 19061 8987 19119 8993
rect 9999 8959 10057 8965
rect 9999 8925 10011 8959
rect 10045 8956 10057 8959
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 10045 8928 16865 8956
rect 10045 8925 10057 8928
rect 9999 8919 10057 8925
rect 16853 8925 16865 8928
rect 16899 8956 16911 8959
rect 16942 8956 16948 8968
rect 16899 8928 16948 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 17497 8959 17555 8965
rect 17497 8925 17509 8959
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 10413 8891 10471 8897
rect 10413 8888 10425 8891
rect 8527 8860 9536 8888
rect 9911 8860 10425 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 9398 8820 9404 8832
rect 9359 8792 9404 8820
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 9508 8820 9536 8860
rect 10413 8857 10425 8860
rect 10459 8888 10471 8891
rect 17313 8891 17371 8897
rect 10459 8860 11376 8888
rect 10459 8857 10471 8860
rect 10413 8851 10471 8857
rect 9858 8820 9864 8832
rect 9508 8792 9864 8820
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 10686 8820 10692 8832
rect 10647 8792 10692 8820
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 11348 8820 11376 8860
rect 17313 8857 17325 8891
rect 17359 8888 17371 8891
rect 17512 8888 17540 8919
rect 17586 8916 17592 8968
rect 17644 8956 17650 8968
rect 17773 8959 17831 8965
rect 17773 8956 17785 8959
rect 17644 8928 17785 8956
rect 17644 8916 17650 8928
rect 17773 8925 17785 8928
rect 17819 8956 17831 8959
rect 18417 8959 18475 8965
rect 18417 8956 18429 8959
rect 17819 8928 18429 8956
rect 17819 8925 17831 8928
rect 17773 8919 17831 8925
rect 18417 8925 18429 8928
rect 18463 8925 18475 8959
rect 19076 8956 19104 8987
rect 19150 8984 19156 9036
rect 19208 9024 19214 9036
rect 21836 9033 21864 9064
rect 22830 9052 22836 9064
rect 22888 9052 22894 9104
rect 24118 9052 24124 9104
rect 24176 9092 24182 9104
rect 24397 9095 24455 9101
rect 24397 9092 24409 9095
rect 24176 9064 24409 9092
rect 24176 9052 24182 9064
rect 24397 9061 24409 9064
rect 24443 9061 24455 9095
rect 24397 9055 24455 9061
rect 19429 9027 19487 9033
rect 19429 9024 19441 9027
rect 19208 8996 19441 9024
rect 19208 8984 19214 8996
rect 19429 8993 19441 8996
rect 19475 8993 19487 9027
rect 19429 8987 19487 8993
rect 21821 9027 21879 9033
rect 21821 8993 21833 9027
rect 21867 8993 21879 9027
rect 21821 8987 21879 8993
rect 19334 8956 19340 8968
rect 19076 8928 19340 8956
rect 18417 8919 18475 8925
rect 19334 8916 19340 8928
rect 19392 8916 19398 8968
rect 19702 8956 19708 8968
rect 19615 8928 19708 8956
rect 19702 8916 19708 8928
rect 19760 8956 19766 8968
rect 19981 8959 20039 8965
rect 19981 8956 19993 8959
rect 19760 8928 19993 8956
rect 19760 8916 19766 8928
rect 19981 8925 19993 8928
rect 20027 8925 20039 8959
rect 20898 8956 20904 8968
rect 20859 8928 20904 8956
rect 19981 8919 20039 8925
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 22738 8956 22744 8968
rect 22699 8928 22744 8956
rect 22738 8916 22744 8928
rect 22796 8916 22802 8968
rect 23014 8956 23020 8968
rect 22975 8928 23020 8956
rect 23014 8916 23020 8928
rect 23072 8916 23078 8968
rect 23382 8916 23388 8968
rect 23440 8956 23446 8968
rect 24305 8959 24363 8965
rect 24305 8956 24317 8959
rect 23440 8928 24317 8956
rect 23440 8916 23446 8928
rect 24305 8925 24317 8928
rect 24351 8925 24363 8959
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 24305 8919 24363 8925
rect 24412 8928 24593 8956
rect 18230 8888 18236 8900
rect 17359 8860 18236 8888
rect 17359 8857 17371 8860
rect 17313 8851 17371 8857
rect 18230 8848 18236 8860
rect 18288 8848 18294 8900
rect 14458 8820 14464 8832
rect 11348 8792 14464 8820
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 14645 8823 14703 8829
rect 14645 8789 14657 8823
rect 14691 8820 14703 8823
rect 15286 8820 15292 8832
rect 14691 8792 15292 8820
rect 14691 8789 14703 8792
rect 14645 8783 14703 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15838 8780 15844 8832
rect 15896 8820 15902 8832
rect 20533 8823 20591 8829
rect 20533 8820 20545 8823
rect 15896 8792 20545 8820
rect 15896 8780 15902 8792
rect 20533 8789 20545 8792
rect 20579 8820 20591 8823
rect 20622 8820 20628 8832
rect 20579 8792 20628 8820
rect 20579 8789 20591 8792
rect 20533 8783 20591 8789
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 22186 8780 22192 8832
rect 22244 8820 22250 8832
rect 24412 8820 24440 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 22244 8792 24440 8820
rect 22244 8780 22250 8792
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 5132 8588 5825 8616
rect 5132 8576 5138 8588
rect 5813 8585 5825 8588
rect 5859 8616 5871 8619
rect 7558 8616 7564 8628
rect 5859 8588 7564 8616
rect 5859 8585 5871 8588
rect 5813 8579 5871 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 8036 8588 9229 8616
rect 5166 8548 5172 8560
rect 5127 8520 5172 8548
rect 5166 8508 5172 8520
rect 5224 8548 5230 8560
rect 8036 8548 8064 8588
rect 9217 8585 9229 8588
rect 9263 8616 9275 8619
rect 9674 8616 9680 8628
rect 9263 8588 9680 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 11606 8616 11612 8628
rect 10008 8588 11612 8616
rect 10008 8576 10014 8588
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 13412 8588 13553 8616
rect 13412 8576 13418 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 13541 8579 13599 8585
rect 15654 8576 15660 8628
rect 15712 8616 15718 8628
rect 16301 8619 16359 8625
rect 16301 8616 16313 8619
rect 15712 8588 16313 8616
rect 15712 8576 15718 8588
rect 16301 8585 16313 8588
rect 16347 8585 16359 8619
rect 16301 8579 16359 8585
rect 16482 8576 16488 8628
rect 16540 8616 16546 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 16540 8588 16957 8616
rect 16540 8576 16546 8588
rect 5224 8520 8064 8548
rect 5224 8508 5230 8520
rect 8110 8508 8116 8560
rect 8168 8548 8174 8560
rect 8297 8551 8355 8557
rect 8297 8548 8309 8551
rect 8168 8520 8309 8548
rect 8168 8508 8174 8520
rect 8297 8517 8309 8520
rect 8343 8517 8355 8551
rect 8297 8511 8355 8517
rect 8662 8508 8668 8560
rect 8720 8548 8726 8560
rect 9493 8551 9551 8557
rect 9493 8548 9505 8551
rect 8720 8520 9505 8548
rect 8720 8508 8726 8520
rect 9493 8517 9505 8520
rect 9539 8548 9551 8551
rect 10962 8548 10968 8560
rect 9539 8520 9996 8548
rect 10875 8520 10968 8548
rect 9539 8517 9551 8520
rect 9493 8511 9551 8517
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9180 8452 9873 8480
rect 9180 8440 9186 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9968 8480 9996 8520
rect 10962 8508 10968 8520
rect 11020 8548 11026 8560
rect 12250 8548 12256 8560
rect 11020 8520 12256 8548
rect 11020 8508 11026 8520
rect 12250 8508 12256 8520
rect 12308 8548 12314 8560
rect 12308 8520 14136 8548
rect 12308 8508 12314 8520
rect 14108 8489 14136 8520
rect 16206 8508 16212 8560
rect 16264 8548 16270 8560
rect 16623 8551 16681 8557
rect 16623 8548 16635 8551
rect 16264 8520 16635 8548
rect 16264 8508 16270 8520
rect 16623 8517 16635 8520
rect 16669 8517 16681 8551
rect 16623 8511 16681 8517
rect 14093 8483 14151 8489
rect 9968 8452 11008 8480
rect 9861 8443 9919 8449
rect 6822 8372 6828 8424
rect 6880 8412 6886 8424
rect 6917 8415 6975 8421
rect 6917 8412 6929 8415
rect 6880 8384 6929 8412
rect 6880 8372 6886 8384
rect 6917 8381 6929 8384
rect 6963 8381 6975 8415
rect 7374 8412 7380 8424
rect 7335 8384 7380 8412
rect 6917 8375 6975 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7708 8384 7941 8412
rect 7708 8372 7714 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 8110 8412 8116 8424
rect 8071 8384 8116 8412
rect 7929 8375 7987 8381
rect 7944 8344 7972 8375
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 9398 8412 9404 8424
rect 9311 8384 9404 8412
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 10042 8412 10048 8424
rect 9732 8384 10048 8412
rect 9732 8372 9738 8384
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10980 8412 11008 8452
rect 14093 8449 14105 8483
rect 14139 8480 14151 8483
rect 14139 8452 15240 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 10980 8384 12265 8412
rect 12253 8381 12265 8384
rect 12299 8412 12311 8415
rect 12618 8412 12624 8424
rect 12299 8384 12624 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12618 8372 12624 8384
rect 12676 8412 12682 8424
rect 14366 8412 14372 8424
rect 12676 8384 13814 8412
rect 14327 8384 14372 8412
rect 12676 8372 12682 8384
rect 8478 8344 8484 8356
rect 7944 8316 8484 8344
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 9416 8344 9444 8372
rect 10778 8344 10784 8356
rect 9416 8316 10784 8344
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 11333 8347 11391 8353
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 12526 8344 12532 8356
rect 11379 8316 12532 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 13262 8344 13268 8356
rect 13223 8316 13268 8344
rect 13262 8304 13268 8316
rect 13320 8304 13326 8356
rect 13786 8344 13814 8384
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 14642 8412 14648 8424
rect 14603 8384 14648 8412
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 15105 8415 15163 8421
rect 15105 8381 15117 8415
rect 15151 8381 15163 8415
rect 15212 8412 15240 8452
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 15212 8384 15393 8412
rect 15105 8375 15163 8381
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 16552 8415 16610 8421
rect 16552 8381 16564 8415
rect 16598 8412 16610 8415
rect 16776 8412 16804 8588
rect 16945 8585 16957 8588
rect 16991 8616 17003 8619
rect 16991 8588 21772 8616
rect 16991 8585 17003 8588
rect 16945 8579 17003 8585
rect 17678 8508 17684 8560
rect 17736 8548 17742 8560
rect 17773 8551 17831 8557
rect 17773 8548 17785 8551
rect 17736 8520 17785 8548
rect 17736 8508 17742 8520
rect 17773 8517 17785 8520
rect 17819 8517 17831 8551
rect 17773 8511 17831 8517
rect 20625 8551 20683 8557
rect 20625 8517 20637 8551
rect 20671 8548 20683 8551
rect 20714 8548 20720 8560
rect 20671 8520 20720 8548
rect 20671 8517 20683 8520
rect 20625 8511 20683 8517
rect 16598 8384 16804 8412
rect 17788 8412 17816 8511
rect 20714 8508 20720 8520
rect 20772 8548 20778 8560
rect 21634 8548 21640 8560
rect 20772 8520 21640 8548
rect 20772 8508 20778 8520
rect 21634 8508 21640 8520
rect 21692 8508 21698 8560
rect 21744 8548 21772 8588
rect 22738 8576 22744 8628
rect 22796 8616 22802 8628
rect 23017 8619 23075 8625
rect 23017 8616 23029 8619
rect 22796 8588 23029 8616
rect 22796 8576 22802 8588
rect 23017 8585 23029 8588
rect 23063 8585 23075 8619
rect 23382 8616 23388 8628
rect 23343 8588 23388 8616
rect 23017 8579 23075 8585
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 21744 8520 23474 8548
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 19518 8480 19524 8492
rect 18923 8452 19524 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 19518 8440 19524 8452
rect 19576 8440 19582 8492
rect 19702 8480 19708 8492
rect 19663 8452 19708 8480
rect 19702 8440 19708 8452
rect 19760 8440 19766 8492
rect 21818 8480 21824 8492
rect 21779 8452 21824 8480
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 22741 8483 22799 8489
rect 22741 8449 22753 8483
rect 22787 8480 22799 8483
rect 22830 8480 22836 8492
rect 22787 8452 22836 8480
rect 22787 8449 22799 8452
rect 22741 8443 22799 8449
rect 22830 8440 22836 8452
rect 22888 8440 22894 8492
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 17788 8384 18153 8412
rect 16598 8381 16610 8384
rect 16552 8375 16610 8381
rect 18141 8381 18153 8384
rect 18187 8412 18199 8415
rect 18598 8412 18604 8424
rect 18187 8384 18604 8412
rect 18187 8381 18199 8384
rect 18141 8375 18199 8381
rect 14660 8344 14688 8372
rect 13786 8316 14688 8344
rect 15120 8344 15148 8375
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 18693 8415 18751 8421
rect 18693 8381 18705 8415
rect 18739 8412 18751 8415
rect 19150 8412 19156 8424
rect 18739 8384 19156 8412
rect 18739 8381 18751 8384
rect 18693 8375 18751 8381
rect 19150 8372 19156 8384
rect 19208 8372 19214 8424
rect 19242 8372 19248 8424
rect 19300 8372 19306 8424
rect 23446 8412 23474 8520
rect 23661 8415 23719 8421
rect 23661 8412 23673 8415
rect 23446 8384 23673 8412
rect 23661 8381 23673 8384
rect 23707 8412 23719 8415
rect 24305 8415 24363 8421
rect 24305 8412 24317 8415
rect 23707 8384 24317 8412
rect 23707 8381 23719 8384
rect 23661 8375 23719 8381
rect 24305 8381 24317 8384
rect 24351 8412 24363 8415
rect 24832 8415 24890 8421
rect 24832 8412 24844 8415
rect 24351 8384 24844 8412
rect 24351 8381 24363 8384
rect 24305 8375 24363 8381
rect 24832 8381 24844 8384
rect 24878 8412 24890 8415
rect 25225 8415 25283 8421
rect 25225 8412 25237 8415
rect 24878 8384 25237 8412
rect 24878 8381 24890 8384
rect 24832 8375 24890 8381
rect 25225 8381 25237 8384
rect 25271 8381 25283 8415
rect 25225 8375 25283 8381
rect 15286 8344 15292 8356
rect 15120 8316 15292 8344
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 15470 8304 15476 8356
rect 15528 8344 15534 8356
rect 17405 8347 17463 8353
rect 17405 8344 17417 8347
rect 15528 8316 17417 8344
rect 15528 8304 15534 8316
rect 17405 8313 17417 8316
rect 17451 8344 17463 8347
rect 17494 8344 17500 8356
rect 17451 8316 17500 8344
rect 17451 8313 17463 8316
rect 17405 8307 17463 8313
rect 17494 8304 17500 8316
rect 17552 8304 17558 8356
rect 19260 8344 19288 8372
rect 19521 8347 19579 8353
rect 19521 8344 19533 8347
rect 18385 8316 19533 8344
rect 5534 8276 5540 8288
rect 5447 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8276 5598 8288
rect 6273 8279 6331 8285
rect 6273 8276 6285 8279
rect 5592 8248 6285 8276
rect 5592 8236 5598 8248
rect 6273 8245 6285 8248
rect 6319 8276 6331 8279
rect 6454 8276 6460 8288
rect 6319 8248 6460 8276
rect 6319 8245 6331 8248
rect 6273 8239 6331 8245
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 6638 8276 6644 8288
rect 6599 8248 6644 8276
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 8662 8276 8668 8288
rect 8623 8248 8668 8276
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 10042 8236 10048 8288
rect 10100 8276 10106 8288
rect 10597 8279 10655 8285
rect 10597 8276 10609 8279
rect 10100 8248 10609 8276
rect 10100 8236 10106 8248
rect 10597 8245 10609 8248
rect 10643 8276 10655 8279
rect 11146 8276 11152 8288
rect 10643 8248 11152 8276
rect 10643 8245 10655 8248
rect 10597 8239 10655 8245
rect 11146 8236 11152 8248
rect 11204 8276 11210 8288
rect 11514 8276 11520 8288
rect 11204 8248 11520 8276
rect 11204 8236 11210 8248
rect 11514 8236 11520 8248
rect 11572 8236 11578 8288
rect 11882 8276 11888 8288
rect 11795 8248 11888 8276
rect 11882 8236 11888 8248
rect 11940 8276 11946 8288
rect 13280 8276 13308 8304
rect 11940 8248 13308 8276
rect 11940 8236 11946 8248
rect 15102 8236 15108 8288
rect 15160 8276 15166 8288
rect 15381 8279 15439 8285
rect 15381 8276 15393 8279
rect 15160 8248 15393 8276
rect 15160 8236 15166 8248
rect 15381 8245 15393 8248
rect 15427 8245 15439 8279
rect 15381 8239 15439 8245
rect 16025 8279 16083 8285
rect 16025 8245 16037 8279
rect 16071 8276 16083 8279
rect 16298 8276 16304 8288
rect 16071 8248 16304 8276
rect 16071 8245 16083 8248
rect 16025 8239 16083 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 18138 8236 18144 8288
rect 18196 8276 18202 8288
rect 18385 8276 18413 8316
rect 19521 8313 19533 8316
rect 19567 8344 19579 8347
rect 20026 8347 20084 8353
rect 20026 8344 20038 8347
rect 19567 8316 20038 8344
rect 19567 8313 19579 8316
rect 19521 8307 19579 8313
rect 20026 8313 20038 8316
rect 20072 8344 20084 8347
rect 20901 8347 20959 8353
rect 20901 8344 20913 8347
rect 20072 8316 20913 8344
rect 20072 8313 20084 8316
rect 20026 8307 20084 8313
rect 20901 8313 20913 8316
rect 20947 8344 20959 8347
rect 21174 8344 21180 8356
rect 20947 8316 21180 8344
rect 20947 8313 20959 8316
rect 20901 8307 20959 8313
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 21545 8347 21603 8353
rect 21545 8344 21557 8347
rect 21284 8316 21557 8344
rect 18196 8248 18413 8276
rect 19245 8279 19303 8285
rect 18196 8236 18202 8248
rect 19245 8245 19257 8279
rect 19291 8276 19303 8279
rect 19334 8276 19340 8288
rect 19291 8248 19340 8276
rect 19291 8245 19303 8248
rect 19245 8239 19303 8245
rect 19334 8236 19340 8248
rect 19392 8236 19398 8288
rect 20990 8236 20996 8288
rect 21048 8276 21054 8288
rect 21284 8285 21312 8316
rect 21545 8313 21557 8316
rect 21591 8313 21603 8347
rect 21545 8307 21603 8313
rect 21634 8304 21640 8356
rect 21692 8344 21698 8356
rect 24118 8344 24124 8356
rect 21692 8316 24124 8344
rect 21692 8304 21698 8316
rect 24118 8304 24124 8316
rect 24176 8344 24182 8356
rect 24581 8347 24639 8353
rect 24581 8344 24593 8347
rect 24176 8316 24593 8344
rect 24176 8304 24182 8316
rect 24581 8313 24593 8316
rect 24627 8313 24639 8347
rect 24581 8307 24639 8313
rect 21269 8279 21327 8285
rect 21269 8276 21281 8279
rect 21048 8248 21281 8276
rect 21048 8236 21054 8248
rect 21269 8245 21281 8248
rect 21315 8245 21327 8279
rect 21269 8239 21327 8245
rect 23845 8279 23903 8285
rect 23845 8245 23857 8279
rect 23891 8276 23903 8279
rect 24210 8276 24216 8288
rect 23891 8248 24216 8276
rect 23891 8245 23903 8248
rect 23845 8239 23903 8245
rect 24210 8236 24216 8248
rect 24268 8236 24274 8288
rect 24670 8236 24676 8288
rect 24728 8276 24734 8288
rect 24903 8279 24961 8285
rect 24903 8276 24915 8279
rect 24728 8248 24915 8276
rect 24728 8236 24734 8248
rect 24903 8245 24915 8248
rect 24949 8245 24961 8279
rect 24903 8239 24961 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 6914 8072 6920 8084
rect 6875 8044 6920 8072
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 7650 8072 7656 8084
rect 7162 8044 7656 8072
rect 6733 8007 6791 8013
rect 6733 7973 6745 8007
rect 6779 8004 6791 8007
rect 7162 8004 7190 8044
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 10962 8072 10968 8084
rect 9830 8044 10968 8072
rect 6779 7976 7190 8004
rect 6779 7973 6791 7976
rect 6733 7967 6791 7973
rect 8018 7964 8024 8016
rect 8076 8004 8082 8016
rect 9830 8004 9858 8044
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12437 8075 12495 8081
rect 12437 8072 12449 8075
rect 12124 8044 12449 8072
rect 12124 8032 12130 8044
rect 12437 8041 12449 8044
rect 12483 8041 12495 8075
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 12437 8035 12495 8041
rect 15102 8032 15108 8044
rect 15160 8072 15166 8084
rect 21545 8075 21603 8081
rect 15160 8044 15608 8072
rect 15160 8032 15166 8044
rect 8076 7976 9858 8004
rect 10413 8007 10471 8013
rect 8076 7964 8082 7976
rect 5880 7939 5938 7945
rect 5880 7905 5892 7939
rect 5926 7936 5938 7939
rect 5994 7936 6000 7948
rect 5926 7908 6000 7936
rect 5926 7905 5938 7908
rect 5880 7899 5938 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6822 7936 6828 7948
rect 6783 7908 6828 7936
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 7374 7936 7380 7948
rect 7335 7908 7380 7936
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 7558 7896 7564 7948
rect 7616 7936 7622 7948
rect 8220 7945 8248 7976
rect 10413 7973 10425 8007
rect 10459 8004 10471 8007
rect 12986 8004 12992 8016
rect 10459 7976 12992 8004
rect 10459 7973 10471 7976
rect 10413 7967 10471 7973
rect 12986 7964 12992 7976
rect 13044 8004 13050 8016
rect 13173 8007 13231 8013
rect 13173 8004 13185 8007
rect 13044 7976 13185 8004
rect 13044 7964 13050 7976
rect 13173 7973 13185 7976
rect 13219 7973 13231 8007
rect 13173 7967 13231 7973
rect 14369 8007 14427 8013
rect 14369 7973 14381 8007
rect 14415 8004 14427 8007
rect 15470 8004 15476 8016
rect 14415 7976 15476 8004
rect 14415 7973 14427 7976
rect 14369 7967 14427 7973
rect 15470 7964 15476 7976
rect 15528 7964 15534 8016
rect 7653 7939 7711 7945
rect 7653 7936 7665 7939
rect 7616 7908 7665 7936
rect 7616 7896 7622 7908
rect 7653 7905 7665 7908
rect 7699 7905 7711 7939
rect 7653 7899 7711 7905
rect 8205 7939 8263 7945
rect 8205 7905 8217 7939
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 9923 7939 9981 7945
rect 9923 7936 9935 7939
rect 9732 7908 9777 7936
rect 9732 7896 9738 7908
rect 9911 7905 9935 7936
rect 9969 7905 9981 7939
rect 11514 7936 11520 7948
rect 11475 7908 11520 7936
rect 9911 7899 9981 7905
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 8110 7868 8116 7880
rect 6411 7840 8116 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 9911 7812 9939 7899
rect 11514 7896 11520 7908
rect 11572 7896 11578 7948
rect 11882 7936 11888 7948
rect 11843 7908 11888 7936
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 12066 7936 12072 7948
rect 12027 7908 12072 7936
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7936 12679 7939
rect 13538 7936 13544 7948
rect 12667 7908 13544 7936
rect 12667 7905 12679 7908
rect 12621 7899 12679 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 13906 7936 13912 7948
rect 13867 7908 13912 7936
rect 13906 7896 13912 7908
rect 13964 7896 13970 7948
rect 15580 7945 15608 8044
rect 21545 8041 21557 8075
rect 21591 8072 21603 8075
rect 21634 8072 21640 8084
rect 21591 8044 21640 8072
rect 21591 8041 21603 8044
rect 21545 8035 21603 8041
rect 21634 8032 21640 8044
rect 21692 8032 21698 8084
rect 22738 8032 22744 8084
rect 22796 8072 22802 8084
rect 24443 8075 24501 8081
rect 24443 8072 24455 8075
rect 22796 8044 24455 8072
rect 22796 8032 22802 8044
rect 24443 8041 24455 8044
rect 24489 8041 24501 8075
rect 24443 8035 24501 8041
rect 15927 8007 15985 8013
rect 15927 7973 15939 8007
rect 15973 8004 15985 8007
rect 16298 8004 16304 8016
rect 15973 7976 16304 8004
rect 15973 7973 15985 7976
rect 15927 7967 15985 7973
rect 16298 7964 16304 7976
rect 16356 7964 16362 8016
rect 17494 8004 17500 8016
rect 17328 7976 17500 8004
rect 17328 7945 17356 7976
rect 17494 7964 17500 7976
rect 17552 7964 17558 8016
rect 19889 8007 19947 8013
rect 19889 7973 19901 8007
rect 19935 8004 19947 8007
rect 20898 8004 20904 8016
rect 19935 7976 20904 8004
rect 19935 7973 19947 7976
rect 19889 7967 19947 7973
rect 20898 7964 20904 7976
rect 20956 8004 20962 8016
rect 21085 8007 21143 8013
rect 21085 8004 21097 8007
rect 20956 7976 21097 8004
rect 20956 7964 20962 7976
rect 21085 7973 21097 7976
rect 21131 7973 21143 8007
rect 21085 7967 21143 7973
rect 21913 8007 21971 8013
rect 21913 7973 21925 8007
rect 21959 8004 21971 8007
rect 22554 8004 22560 8016
rect 21959 7976 22560 8004
rect 21959 7973 21971 7976
rect 21913 7967 21971 7973
rect 22554 7964 22560 7976
rect 22612 8004 22618 8016
rect 22830 8004 22836 8016
rect 22612 7976 22836 8004
rect 22612 7964 22618 7976
rect 22830 7964 22836 7976
rect 22888 7964 22894 8016
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7905 15623 7939
rect 15565 7899 15623 7905
rect 17313 7939 17371 7945
rect 17313 7905 17325 7939
rect 17359 7905 17371 7939
rect 17313 7899 17371 7905
rect 17402 7896 17408 7948
rect 17460 7936 17466 7948
rect 17773 7939 17831 7945
rect 17773 7936 17785 7939
rect 17460 7908 17785 7936
rect 17460 7896 17466 7908
rect 17773 7905 17785 7908
rect 17819 7936 17831 7939
rect 17819 7908 18368 7936
rect 17819 7905 17831 7908
rect 17773 7899 17831 7905
rect 14550 7828 14556 7880
rect 14608 7868 14614 7880
rect 17678 7868 17684 7880
rect 14608 7840 17684 7868
rect 14608 7828 14614 7840
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 17862 7868 17868 7880
rect 17823 7840 17868 7868
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 18340 7868 18368 7908
rect 18966 7896 18972 7948
rect 19024 7936 19030 7948
rect 19153 7939 19211 7945
rect 19153 7936 19165 7939
rect 19024 7908 19165 7936
rect 19024 7896 19030 7908
rect 19153 7905 19165 7908
rect 19199 7905 19211 7939
rect 19153 7899 19211 7905
rect 19242 7896 19248 7948
rect 19300 7936 19306 7948
rect 19613 7939 19671 7945
rect 19613 7936 19625 7939
rect 19300 7908 19625 7936
rect 19300 7896 19306 7908
rect 19613 7905 19625 7908
rect 19659 7905 19671 7939
rect 19613 7899 19671 7905
rect 22462 7896 22468 7948
rect 22520 7936 22526 7948
rect 23014 7936 23020 7948
rect 22520 7908 23020 7936
rect 22520 7896 22526 7908
rect 23014 7896 23020 7908
rect 23072 7936 23078 7948
rect 23328 7939 23386 7945
rect 23328 7936 23340 7939
rect 23072 7908 23340 7936
rect 23072 7896 23078 7908
rect 23328 7905 23340 7908
rect 23374 7905 23386 7939
rect 23328 7899 23386 7905
rect 24372 7939 24430 7945
rect 24372 7905 24384 7939
rect 24418 7905 24430 7939
rect 24372 7899 24430 7905
rect 21821 7871 21879 7877
rect 18340 7840 20300 7868
rect 9125 7803 9183 7809
rect 9125 7769 9137 7803
rect 9171 7800 9183 7803
rect 9766 7800 9772 7812
rect 9171 7772 9772 7800
rect 9171 7769 9183 7772
rect 9125 7763 9183 7769
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 9858 7760 9864 7812
rect 9916 7800 9939 7812
rect 14366 7800 14372 7812
rect 9916 7772 14372 7800
rect 9916 7760 9922 7772
rect 14366 7760 14372 7772
rect 14424 7800 14430 7812
rect 14645 7803 14703 7809
rect 14645 7800 14657 7803
rect 14424 7772 14657 7800
rect 14424 7760 14430 7772
rect 14645 7769 14657 7772
rect 14691 7769 14703 7803
rect 14645 7763 14703 7769
rect 15930 7760 15936 7812
rect 15988 7800 15994 7812
rect 18325 7803 18383 7809
rect 18325 7800 18337 7803
rect 15988 7772 18337 7800
rect 15988 7760 15994 7772
rect 18325 7769 18337 7772
rect 18371 7800 18383 7803
rect 18969 7803 19027 7809
rect 18969 7800 18981 7803
rect 18371 7772 18981 7800
rect 18371 7769 18383 7772
rect 18325 7763 18383 7769
rect 18969 7769 18981 7772
rect 19015 7800 19027 7803
rect 19150 7800 19156 7812
rect 19015 7772 19156 7800
rect 19015 7769 19027 7772
rect 18969 7763 19027 7769
rect 19150 7760 19156 7772
rect 19208 7760 19214 7812
rect 20272 7744 20300 7840
rect 21821 7837 21833 7871
rect 21867 7837 21879 7871
rect 21821 7831 21879 7837
rect 5951 7735 6009 7741
rect 5951 7701 5963 7735
rect 5997 7732 6009 7735
rect 6178 7732 6184 7744
rect 5997 7704 6184 7732
rect 5997 7701 6009 7704
rect 5951 7695 6009 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 6454 7692 6460 7744
rect 6512 7732 6518 7744
rect 7374 7732 7380 7744
rect 6512 7704 7380 7732
rect 6512 7692 6518 7704
rect 7374 7692 7380 7704
rect 7432 7732 7438 7744
rect 8662 7732 8668 7744
rect 7432 7704 8668 7732
rect 7432 7692 7438 7704
rect 8662 7692 8668 7704
rect 8720 7732 8726 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 8720 7704 9413 7732
rect 8720 7692 8726 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 9401 7695 9459 7701
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 10873 7735 10931 7741
rect 10873 7732 10885 7735
rect 10836 7704 10885 7732
rect 10836 7692 10842 7704
rect 10873 7701 10885 7704
rect 10919 7701 10931 7735
rect 10873 7695 10931 7701
rect 13906 7692 13912 7744
rect 13964 7732 13970 7744
rect 16485 7735 16543 7741
rect 16485 7732 16497 7735
rect 13964 7704 16497 7732
rect 13964 7692 13970 7704
rect 16485 7701 16497 7704
rect 16531 7732 16543 7735
rect 17310 7732 17316 7744
rect 16531 7704 17316 7732
rect 16531 7701 16543 7704
rect 16485 7695 16543 7701
rect 17310 7692 17316 7704
rect 17368 7692 17374 7744
rect 20254 7732 20260 7744
rect 20215 7704 20260 7732
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 21836 7732 21864 7831
rect 21910 7828 21916 7880
rect 21968 7868 21974 7880
rect 22097 7871 22155 7877
rect 22097 7868 22109 7871
rect 21968 7840 22109 7868
rect 21968 7828 21974 7840
rect 22097 7837 22109 7840
rect 22143 7837 22155 7871
rect 24387 7868 24415 7899
rect 24670 7868 24676 7880
rect 24387 7840 24676 7868
rect 22097 7831 22155 7837
rect 24670 7828 24676 7840
rect 24728 7828 24734 7880
rect 23658 7760 23664 7812
rect 23716 7800 23722 7812
rect 24121 7803 24179 7809
rect 24121 7800 24133 7803
rect 23716 7772 24133 7800
rect 23716 7760 23722 7772
rect 24121 7769 24133 7772
rect 24167 7769 24179 7803
rect 24121 7763 24179 7769
rect 22830 7732 22836 7744
rect 21836 7704 22836 7732
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 22922 7692 22928 7744
rect 22980 7732 22986 7744
rect 23431 7735 23489 7741
rect 23431 7732 23443 7735
rect 22980 7704 23443 7732
rect 22980 7692 22986 7704
rect 23431 7701 23443 7704
rect 23477 7701 23489 7735
rect 23842 7732 23848 7744
rect 23803 7704 23848 7732
rect 23431 7695 23489 7701
rect 23842 7692 23848 7704
rect 23900 7692 23906 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 5994 7528 6000 7540
rect 5951 7500 6000 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 7742 7528 7748 7540
rect 7616 7500 7748 7528
rect 7616 7488 7622 7500
rect 7742 7488 7748 7500
rect 7800 7528 7806 7540
rect 8113 7531 8171 7537
rect 8113 7528 8125 7531
rect 7800 7500 8125 7528
rect 7800 7488 7806 7500
rect 8113 7497 8125 7500
rect 8159 7528 8171 7531
rect 9674 7528 9680 7540
rect 8159 7500 9680 7528
rect 8159 7497 8171 7500
rect 8113 7491 8171 7497
rect 9674 7488 9680 7500
rect 9732 7528 9738 7540
rect 9858 7528 9864 7540
rect 9732 7500 9864 7528
rect 9732 7488 9738 7500
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 11514 7488 11520 7540
rect 11572 7528 11578 7540
rect 11609 7531 11667 7537
rect 11609 7528 11621 7531
rect 11572 7500 11621 7528
rect 11572 7488 11578 7500
rect 11609 7497 11621 7500
rect 11655 7528 11667 7531
rect 13357 7531 13415 7537
rect 13357 7528 13369 7531
rect 11655 7500 13369 7528
rect 11655 7497 11667 7500
rect 11609 7491 11667 7497
rect 13357 7497 13369 7500
rect 13403 7497 13415 7531
rect 13906 7528 13912 7540
rect 13867 7500 13912 7528
rect 13357 7491 13415 7497
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 14645 7531 14703 7537
rect 14645 7528 14657 7531
rect 14516 7500 14657 7528
rect 14516 7488 14522 7500
rect 14645 7497 14657 7500
rect 14691 7497 14703 7531
rect 16298 7528 16304 7540
rect 16211 7500 16304 7528
rect 14645 7491 14703 7497
rect 16298 7488 16304 7500
rect 16356 7528 16362 7540
rect 18138 7528 18144 7540
rect 16356 7500 18144 7528
rect 16356 7488 16362 7500
rect 18138 7488 18144 7500
rect 18196 7488 18202 7540
rect 18966 7488 18972 7540
rect 19024 7528 19030 7540
rect 19337 7531 19395 7537
rect 19337 7528 19349 7531
rect 19024 7500 19349 7528
rect 19024 7488 19030 7500
rect 19337 7497 19349 7500
rect 19383 7528 19395 7531
rect 20070 7528 20076 7540
rect 19383 7500 20076 7528
rect 19383 7497 19395 7500
rect 19337 7491 19395 7497
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 21453 7531 21511 7537
rect 21453 7497 21465 7531
rect 21499 7528 21511 7531
rect 21818 7528 21824 7540
rect 21499 7500 21824 7528
rect 21499 7497 21511 7500
rect 21453 7491 21511 7497
rect 21818 7488 21824 7500
rect 21876 7528 21882 7540
rect 22554 7528 22560 7540
rect 21876 7500 22560 7528
rect 21876 7488 21882 7500
rect 22554 7488 22560 7500
rect 22612 7488 22618 7540
rect 23014 7528 23020 7540
rect 22975 7500 23020 7528
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 25774 7528 25780 7540
rect 25735 7500 25780 7528
rect 25774 7488 25780 7500
rect 25832 7488 25838 7540
rect 6178 7420 6184 7472
rect 6236 7460 6242 7472
rect 12986 7460 12992 7472
rect 6236 7432 12992 7460
rect 6236 7420 6242 7432
rect 6914 7392 6920 7404
rect 6875 7364 6920 7392
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7392 10379 7395
rect 10686 7392 10692 7404
rect 10367 7364 10692 7392
rect 10367 7361 10379 7364
rect 10321 7355 10379 7361
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 10778 7352 10784 7404
rect 10836 7392 10842 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 10836 7364 11897 7392
rect 10836 7352 10842 7364
rect 11885 7361 11897 7364
rect 11931 7392 11943 7395
rect 12066 7392 12072 7404
rect 11931 7364 12072 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12544 7401 12572 7432
rect 12986 7420 12992 7432
rect 13044 7420 13050 7472
rect 13262 7420 13268 7472
rect 13320 7460 13326 7472
rect 15289 7463 15347 7469
rect 15289 7460 15301 7463
rect 13320 7432 15301 7460
rect 13320 7420 13326 7432
rect 15289 7429 15301 7432
rect 15335 7460 15347 7463
rect 15470 7460 15476 7472
rect 15335 7432 15476 7460
rect 15335 7429 15347 7432
rect 15289 7423 15347 7429
rect 15470 7420 15476 7432
rect 15528 7420 15534 7472
rect 17494 7420 17500 7472
rect 17552 7460 17558 7472
rect 17773 7463 17831 7469
rect 17773 7460 17785 7463
rect 17552 7432 17785 7460
rect 17552 7420 17558 7432
rect 17773 7429 17785 7432
rect 17819 7460 17831 7463
rect 19242 7460 19248 7472
rect 17819 7432 19248 7460
rect 17819 7429 17831 7432
rect 17773 7423 17831 7429
rect 19242 7420 19248 7432
rect 19300 7420 19306 7472
rect 22186 7460 22192 7472
rect 22147 7432 22192 7460
rect 22186 7420 22192 7432
rect 22244 7420 22250 7472
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7361 12587 7395
rect 12802 7392 12808 7404
rect 12763 7364 12808 7392
rect 12529 7355 12587 7361
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 16577 7395 16635 7401
rect 16577 7392 16589 7395
rect 15212 7364 16589 7392
rect 3418 7284 3424 7336
rect 3476 7324 3482 7336
rect 4960 7327 5018 7333
rect 4960 7324 4972 7327
rect 3476 7296 4972 7324
rect 3476 7284 3482 7296
rect 4960 7293 4972 7296
rect 5006 7324 5018 7327
rect 5353 7327 5411 7333
rect 5353 7324 5365 7327
rect 5006 7296 5365 7324
rect 5006 7293 5018 7296
rect 4960 7287 5018 7293
rect 5353 7293 5365 7296
rect 5399 7293 5411 7327
rect 6638 7324 6644 7336
rect 6551 7296 6644 7324
rect 5353 7287 5411 7293
rect 6638 7284 6644 7296
rect 6696 7324 6702 7336
rect 8018 7324 8024 7336
rect 6696 7296 8024 7324
rect 6696 7284 6702 7296
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7324 8723 7327
rect 9398 7324 9404 7336
rect 8711 7296 9404 7324
rect 8711 7293 8723 7296
rect 8665 7287 8723 7293
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 9493 7327 9551 7333
rect 9493 7293 9505 7327
rect 9539 7324 9551 7327
rect 12342 7324 12348 7336
rect 9539 7296 12348 7324
rect 9539 7293 9551 7296
rect 9493 7287 9551 7293
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 14236 7327 14294 7333
rect 14236 7293 14248 7327
rect 14282 7324 14294 7327
rect 14458 7324 14464 7336
rect 14282 7296 14464 7324
rect 14282 7293 14294 7296
rect 14236 7287 14294 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 15212 7333 15240 7364
rect 16577 7361 16589 7364
rect 16623 7361 16635 7395
rect 16577 7355 16635 7361
rect 18230 7352 18236 7404
rect 18288 7392 18294 7404
rect 18693 7395 18751 7401
rect 18693 7392 18705 7395
rect 18288 7364 18705 7392
rect 18288 7352 18294 7364
rect 18693 7361 18705 7364
rect 18739 7361 18751 7395
rect 18693 7355 18751 7361
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 21637 7395 21695 7401
rect 21637 7392 21649 7395
rect 20772 7364 21649 7392
rect 20772 7352 20778 7364
rect 21637 7361 21649 7364
rect 21683 7392 21695 7395
rect 22922 7392 22928 7404
rect 21683 7364 22928 7392
rect 21683 7361 21695 7364
rect 21637 7355 21695 7361
rect 22922 7352 22928 7364
rect 22980 7352 22986 7404
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 23750 7392 23756 7404
rect 23523 7364 23756 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 23750 7352 23756 7364
rect 23808 7352 23814 7404
rect 24118 7392 24124 7404
rect 24079 7364 24124 7392
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 14884 7296 15209 7324
rect 14884 7284 14890 7296
rect 15197 7293 15209 7296
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 15473 7327 15531 7333
rect 15473 7293 15485 7327
rect 15519 7324 15531 7327
rect 15654 7324 15660 7336
rect 15519 7296 15660 7324
rect 15519 7293 15531 7296
rect 15473 7287 15531 7293
rect 15654 7284 15660 7296
rect 15712 7284 15718 7336
rect 15930 7324 15936 7336
rect 15891 7296 15936 7324
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16666 7284 16672 7336
rect 16724 7324 16730 7336
rect 16888 7327 16946 7333
rect 16888 7324 16900 7327
rect 16724 7296 16900 7324
rect 16724 7284 16730 7296
rect 16888 7293 16900 7296
rect 16934 7324 16946 7327
rect 17034 7324 17040 7336
rect 16934 7296 17040 7324
rect 16934 7293 16946 7296
rect 16888 7287 16946 7293
rect 17034 7284 17040 7296
rect 17092 7324 17098 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 17092 7296 17325 7324
rect 17092 7284 17098 7296
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 19978 7324 19984 7336
rect 19939 7296 19984 7324
rect 17313 7287 17371 7293
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 20254 7284 20260 7336
rect 20312 7324 20318 7336
rect 20349 7327 20407 7333
rect 20349 7324 20361 7327
rect 20312 7296 20361 7324
rect 20312 7284 20318 7296
rect 20349 7293 20361 7296
rect 20395 7293 20407 7327
rect 20622 7324 20628 7336
rect 20583 7296 20628 7324
rect 20349 7287 20407 7293
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 22554 7284 22560 7336
rect 22612 7324 22618 7336
rect 23290 7324 23296 7336
rect 22612 7296 23296 7324
rect 22612 7284 22618 7296
rect 23290 7284 23296 7296
rect 23348 7284 23354 7336
rect 23658 7324 23664 7336
rect 23619 7296 23664 7324
rect 23658 7284 23664 7296
rect 23716 7284 23722 7336
rect 23842 7284 23848 7336
rect 23900 7324 23906 7336
rect 23937 7327 23995 7333
rect 23937 7324 23949 7327
rect 23900 7296 23949 7324
rect 23900 7284 23906 7296
rect 23937 7293 23949 7296
rect 23983 7293 23995 7327
rect 23937 7287 23995 7293
rect 25292 7327 25350 7333
rect 25292 7293 25304 7327
rect 25338 7324 25350 7327
rect 25774 7324 25780 7336
rect 25338 7296 25780 7324
rect 25338 7293 25350 7296
rect 25292 7287 25350 7293
rect 25774 7284 25780 7296
rect 25832 7284 25838 7336
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 7300 7228 10149 7256
rect 7300 7200 7328 7228
rect 10137 7225 10149 7228
rect 10183 7256 10195 7259
rect 10642 7259 10700 7265
rect 10642 7256 10654 7259
rect 10183 7228 10654 7256
rect 10183 7225 10195 7228
rect 10137 7219 10195 7225
rect 10642 7225 10654 7228
rect 10688 7225 10700 7259
rect 12621 7259 12679 7265
rect 10642 7219 10700 7225
rect 11256 7228 12020 7256
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 5031 7191 5089 7197
rect 5031 7188 5043 7191
rect 4948 7160 5043 7188
rect 4948 7148 4954 7160
rect 5031 7157 5043 7160
rect 5077 7157 5089 7191
rect 5031 7151 5089 7157
rect 6273 7191 6331 7197
rect 6273 7157 6285 7191
rect 6319 7188 6331 7191
rect 6454 7188 6460 7200
rect 6319 7160 6460 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 7282 7188 7288 7200
rect 7243 7160 7288 7188
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 7834 7188 7840 7200
rect 7795 7160 7840 7188
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 9858 7188 9864 7200
rect 9819 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 11256 7197 11284 7228
rect 11241 7191 11299 7197
rect 11241 7157 11253 7191
rect 11287 7157 11299 7191
rect 11992 7188 12020 7228
rect 12621 7225 12633 7259
rect 12667 7256 12679 7259
rect 13449 7259 13507 7265
rect 13449 7256 13461 7259
rect 12667 7228 13461 7256
rect 12667 7225 12679 7228
rect 12621 7219 12679 7225
rect 13449 7225 13461 7228
rect 13495 7225 13507 7259
rect 13449 7219 13507 7225
rect 14323 7259 14381 7265
rect 14323 7225 14335 7259
rect 14369 7256 14381 7259
rect 18417 7259 18475 7265
rect 18417 7256 18429 7259
rect 14369 7228 18429 7256
rect 14369 7225 14381 7228
rect 14323 7219 14381 7225
rect 18417 7225 18429 7228
rect 18463 7225 18475 7259
rect 18417 7219 18475 7225
rect 12434 7188 12440 7200
rect 11992 7160 12440 7188
rect 11241 7151 11299 7157
rect 12434 7148 12440 7160
rect 12492 7188 12498 7200
rect 12636 7188 12664 7219
rect 12492 7160 12664 7188
rect 13357 7191 13415 7197
rect 12492 7148 12498 7160
rect 13357 7157 13369 7191
rect 13403 7188 13415 7191
rect 15105 7191 15163 7197
rect 15105 7188 15117 7191
rect 13403 7160 15117 7188
rect 13403 7157 13415 7160
rect 13357 7151 13415 7157
rect 15105 7157 15117 7160
rect 15151 7188 15163 7191
rect 15654 7188 15660 7200
rect 15151 7160 15660 7188
rect 15151 7157 15163 7160
rect 15105 7151 15163 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 16850 7148 16856 7200
rect 16908 7188 16914 7200
rect 16991 7191 17049 7197
rect 16991 7188 17003 7191
rect 16908 7160 17003 7188
rect 16908 7148 16914 7160
rect 16991 7157 17003 7160
rect 17037 7157 17049 7191
rect 18432 7188 18460 7219
rect 18506 7216 18512 7268
rect 18564 7256 18570 7268
rect 20901 7259 20959 7265
rect 20901 7256 20913 7259
rect 18564 7228 18609 7256
rect 19168 7228 20913 7256
rect 18564 7216 18570 7228
rect 19168 7188 19196 7228
rect 20901 7225 20913 7228
rect 20947 7225 20959 7259
rect 20901 7219 20959 7225
rect 21729 7259 21787 7265
rect 21729 7225 21741 7259
rect 21775 7256 21787 7259
rect 21818 7256 21824 7268
rect 21775 7228 21824 7256
rect 21775 7225 21787 7228
rect 21729 7219 21787 7225
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 18432 7160 19196 7188
rect 19797 7191 19855 7197
rect 16991 7151 17049 7157
rect 19797 7157 19809 7191
rect 19843 7188 19855 7191
rect 19978 7188 19984 7200
rect 19843 7160 19984 7188
rect 19843 7157 19855 7160
rect 19797 7151 19855 7157
rect 19978 7148 19984 7160
rect 20036 7188 20042 7200
rect 21082 7188 21088 7200
rect 20036 7160 21088 7188
rect 20036 7148 20042 7160
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 24670 7188 24676 7200
rect 24631 7160 24676 7188
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 24762 7148 24768 7200
rect 24820 7188 24826 7200
rect 25363 7191 25421 7197
rect 25363 7188 25375 7191
rect 24820 7160 25375 7188
rect 24820 7148 24826 7160
rect 25363 7157 25375 7160
rect 25409 7157 25421 7191
rect 25363 7151 25421 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 6089 6987 6147 6993
rect 6089 6953 6101 6987
rect 6135 6984 6147 6987
rect 6914 6984 6920 6996
rect 6135 6956 6920 6984
rect 6135 6953 6147 6956
rect 6089 6947 6147 6953
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 8110 6944 8116 6996
rect 8168 6984 8174 6996
rect 9125 6987 9183 6993
rect 8168 6956 8651 6984
rect 8168 6944 8174 6956
rect 4890 6916 4896 6928
rect 4126 6888 4896 6916
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 4126 6792 4154 6888
rect 4890 6876 4896 6888
rect 4948 6916 4954 6928
rect 5077 6919 5135 6925
rect 5077 6916 5089 6919
rect 4948 6888 5089 6916
rect 4948 6876 4954 6888
rect 5077 6885 5089 6888
rect 5123 6885 5135 6919
rect 5077 6879 5135 6885
rect 5166 6876 5172 6928
rect 5224 6916 5230 6928
rect 6730 6916 6736 6928
rect 5224 6888 6736 6916
rect 5224 6876 5230 6888
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 8623 6916 8651 6956
rect 9125 6953 9137 6987
rect 9171 6984 9183 6987
rect 9674 6984 9680 6996
rect 9171 6956 9680 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9674 6944 9680 6956
rect 9732 6984 9738 6996
rect 9950 6984 9956 6996
rect 9732 6956 9956 6984
rect 9732 6944 9738 6956
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 10686 6944 10692 6996
rect 10744 6984 10750 6996
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 10744 6956 10885 6984
rect 10744 6944 10750 6956
rect 10873 6953 10885 6956
rect 10919 6953 10931 6987
rect 11882 6984 11888 6996
rect 11843 6956 11888 6984
rect 10873 6947 10931 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 13449 6987 13507 6993
rect 13449 6984 13461 6987
rect 12400 6956 13461 6984
rect 12400 6944 12406 6956
rect 13449 6953 13461 6956
rect 13495 6953 13507 6987
rect 16850 6984 16856 6996
rect 16811 6956 16856 6984
rect 13449 6947 13507 6953
rect 9401 6919 9459 6925
rect 9401 6916 9413 6919
rect 8623 6888 9413 6916
rect 9401 6885 9413 6888
rect 9447 6885 9459 6919
rect 9401 6879 9459 6885
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8202 6848 8208 6860
rect 8159 6820 8208 6848
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 4062 6740 4068 6792
rect 4120 6752 4154 6792
rect 5721 6783 5779 6789
rect 4120 6740 4126 6752
rect 5721 6749 5733 6783
rect 5767 6780 5779 6783
rect 5994 6780 6000 6792
rect 5767 6752 6000 6780
rect 5767 6749 5779 6752
rect 5721 6743 5779 6749
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6638 6780 6644 6792
rect 6599 6752 6644 6780
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 7190 6712 7196 6724
rect 7151 6684 7196 6712
rect 7190 6672 7196 6684
rect 7248 6712 7254 6724
rect 7929 6715 7987 6721
rect 7929 6712 7941 6715
rect 7248 6684 7941 6712
rect 7248 6672 7254 6684
rect 7929 6681 7941 6684
rect 7975 6681 7987 6715
rect 9416 6712 9444 6879
rect 9858 6876 9864 6928
rect 9916 6916 9922 6928
rect 12161 6919 12219 6925
rect 9916 6888 10732 6916
rect 9916 6876 9922 6888
rect 10704 6860 10732 6888
rect 12161 6885 12173 6919
rect 12207 6916 12219 6919
rect 12250 6916 12256 6928
rect 12207 6888 12256 6916
rect 12207 6885 12219 6888
rect 12161 6879 12219 6885
rect 12250 6876 12256 6888
rect 12308 6876 12314 6928
rect 12986 6916 12992 6928
rect 12947 6888 12992 6916
rect 12986 6876 12992 6888
rect 13044 6876 13050 6928
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 9692 6780 9720 6811
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 10410 6848 10416 6860
rect 9824 6820 10416 6848
rect 9824 6808 9830 6820
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 10686 6848 10692 6860
rect 10647 6820 10692 6848
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 10962 6848 10968 6860
rect 10923 6820 10968 6848
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 10042 6780 10048 6792
rect 9692 6752 10048 6780
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 11514 6740 11520 6792
rect 11572 6780 11578 6792
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 11572 6752 12081 6780
rect 11572 6740 11578 6752
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12710 6780 12716 6792
rect 12671 6752 12716 6780
rect 12069 6743 12127 6749
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 13464 6712 13492 6947
rect 16850 6944 16856 6956
rect 16908 6944 16914 6996
rect 17402 6984 17408 6996
rect 17363 6956 17408 6984
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 18138 6984 18144 6996
rect 18099 6956 18144 6984
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 19518 6984 19524 6996
rect 18564 6956 19524 6984
rect 18564 6944 18570 6956
rect 19518 6944 19524 6956
rect 19576 6944 19582 6996
rect 20714 6984 20720 6996
rect 20675 6956 20720 6984
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 20990 6984 20996 6996
rect 20951 6956 20996 6984
rect 20990 6944 20996 6956
rect 21048 6944 21054 6996
rect 22830 6944 22836 6996
rect 22888 6984 22894 6996
rect 25271 6987 25329 6993
rect 25271 6984 25283 6987
rect 22888 6956 25283 6984
rect 22888 6944 22894 6956
rect 25271 6953 25283 6956
rect 25317 6953 25329 6987
rect 25271 6947 25329 6953
rect 14369 6919 14427 6925
rect 14369 6885 14381 6919
rect 14415 6916 14427 6919
rect 14550 6916 14556 6928
rect 14415 6888 14556 6916
rect 14415 6885 14427 6888
rect 14369 6879 14427 6885
rect 14550 6876 14556 6888
rect 14608 6876 14614 6928
rect 16117 6919 16175 6925
rect 16117 6885 16129 6919
rect 16163 6916 16175 6919
rect 17034 6916 17040 6928
rect 16163 6888 17040 6916
rect 16163 6885 16175 6888
rect 16117 6879 16175 6885
rect 17034 6876 17040 6888
rect 17092 6916 17098 6928
rect 17420 6916 17448 6944
rect 19150 6916 19156 6928
rect 17092 6888 17448 6916
rect 19111 6888 19156 6916
rect 17092 6876 17098 6888
rect 19150 6876 19156 6888
rect 19208 6876 19214 6928
rect 22186 6916 22192 6928
rect 22147 6888 22192 6916
rect 22186 6876 22192 6888
rect 22244 6876 22250 6928
rect 23753 6919 23811 6925
rect 23753 6885 23765 6919
rect 23799 6916 23811 6919
rect 24026 6916 24032 6928
rect 23799 6888 24032 6916
rect 23799 6885 23811 6888
rect 23753 6879 23811 6885
rect 24026 6876 24032 6888
rect 24084 6876 24090 6928
rect 13538 6808 13544 6860
rect 13596 6848 13602 6860
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 13596 6820 13645 6848
rect 13596 6808 13602 6820
rect 13633 6817 13645 6820
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 13909 6851 13967 6857
rect 13909 6848 13921 6851
rect 13780 6820 13921 6848
rect 13780 6808 13786 6820
rect 13909 6817 13921 6820
rect 13955 6817 13967 6851
rect 15378 6848 15384 6860
rect 15339 6820 15384 6848
rect 13909 6811 13967 6817
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 15654 6848 15660 6860
rect 15615 6820 15660 6848
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 17773 6851 17831 6857
rect 17773 6817 17785 6851
rect 17819 6848 17831 6851
rect 17862 6848 17868 6860
rect 17819 6820 17868 6848
rect 17819 6817 17831 6820
rect 17773 6811 17831 6817
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 19610 6808 19616 6860
rect 19668 6848 19674 6860
rect 19832 6851 19890 6857
rect 19832 6848 19844 6851
rect 19668 6820 19844 6848
rect 19668 6808 19674 6820
rect 19832 6817 19844 6820
rect 19878 6817 19890 6851
rect 19832 6811 19890 6817
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6848 25191 6851
rect 25222 6848 25228 6860
rect 25179 6820 25228 6848
rect 25179 6817 25191 6820
rect 25133 6811 25191 6817
rect 25222 6808 25228 6820
rect 25280 6808 25286 6860
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6780 15163 6783
rect 15470 6780 15476 6792
rect 15151 6752 15476 6780
rect 15151 6749 15163 6752
rect 15105 6743 15163 6749
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 21266 6780 21272 6792
rect 15580 6752 21272 6780
rect 13725 6715 13783 6721
rect 13725 6712 13737 6715
rect 9416 6684 11284 6712
rect 13464 6684 13737 6712
rect 7929 6675 7987 6681
rect 11256 6656 11284 6684
rect 13725 6681 13737 6684
rect 13771 6712 13783 6715
rect 15580 6712 15608 6752
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 22094 6780 22100 6792
rect 22055 6752 22100 6780
rect 22094 6740 22100 6752
rect 22152 6740 22158 6792
rect 22373 6783 22431 6789
rect 22373 6749 22385 6783
rect 22419 6749 22431 6783
rect 23658 6780 23664 6792
rect 23619 6752 23664 6780
rect 22373 6743 22431 6749
rect 13771 6684 15608 6712
rect 16485 6715 16543 6721
rect 13771 6681 13783 6684
rect 13725 6675 13783 6681
rect 16485 6681 16497 6715
rect 16531 6712 16543 6715
rect 16574 6712 16580 6724
rect 16531 6684 16580 6712
rect 16531 6681 16543 6684
rect 16485 6675 16543 6681
rect 16574 6672 16580 6684
rect 16632 6712 16638 6724
rect 22388 6712 22416 6743
rect 23658 6740 23664 6752
rect 23716 6740 23722 6792
rect 23937 6783 23995 6789
rect 23937 6780 23949 6783
rect 23768 6752 23949 6780
rect 23014 6712 23020 6724
rect 16632 6684 18736 6712
rect 16632 6672 16638 6684
rect 18708 6656 18736 6684
rect 21652 6684 23020 6712
rect 21652 6656 21680 6684
rect 23014 6672 23020 6684
rect 23072 6712 23078 6724
rect 23768 6712 23796 6752
rect 23937 6749 23949 6752
rect 23983 6749 23995 6783
rect 23937 6743 23995 6749
rect 23072 6684 23796 6712
rect 23072 6672 23078 6684
rect 4890 6644 4896 6656
rect 4851 6616 4896 6644
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 6457 6647 6515 6653
rect 6457 6613 6469 6647
rect 6503 6644 6515 6647
rect 6822 6644 6828 6656
rect 6503 6616 6828 6644
rect 6503 6613 6515 6616
rect 6457 6607 6515 6613
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 7561 6647 7619 6653
rect 7561 6644 7573 6647
rect 7340 6616 7573 6644
rect 7340 6604 7346 6616
rect 7561 6613 7573 6616
rect 7607 6613 7619 6647
rect 7561 6607 7619 6613
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 8251 6647 8309 6653
rect 8251 6644 8263 6647
rect 8168 6616 8263 6644
rect 8168 6604 8174 6616
rect 8251 6613 8263 6616
rect 8297 6613 8309 6647
rect 8251 6607 8309 6613
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11517 6647 11575 6653
rect 11517 6644 11529 6647
rect 11296 6616 11529 6644
rect 11296 6604 11302 6616
rect 11517 6613 11529 6616
rect 11563 6644 11575 6647
rect 13538 6644 13544 6656
rect 11563 6616 13544 6644
rect 11563 6613 11575 6616
rect 11517 6607 11575 6613
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 18690 6644 18696 6656
rect 18651 6616 18696 6644
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 19935 6647 19993 6653
rect 19935 6613 19947 6647
rect 19981 6644 19993 6647
rect 21450 6644 21456 6656
rect 19981 6616 21456 6644
rect 19981 6613 19993 6616
rect 19935 6607 19993 6613
rect 21450 6604 21456 6616
rect 21508 6604 21514 6656
rect 21634 6644 21640 6656
rect 21595 6616 21640 6644
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1811 6443 1869 6449
rect 1811 6440 1823 6443
rect 1452 6412 1823 6440
rect 1452 6400 1458 6412
rect 1811 6409 1823 6412
rect 1857 6440 1869 6443
rect 1946 6440 1952 6452
rect 1857 6412 1952 6440
rect 1857 6409 1869 6412
rect 1811 6403 1869 6409
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 4062 6440 4068 6452
rect 4023 6412 4068 6440
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 5077 6443 5135 6449
rect 5077 6409 5089 6443
rect 5123 6440 5135 6443
rect 5166 6440 5172 6452
rect 5123 6412 5172 6440
rect 5123 6409 5135 6412
rect 5077 6403 5135 6409
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 6730 6440 6736 6452
rect 6687 6412 6736 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 8352 6412 13814 6440
rect 8352 6400 8358 6412
rect 4709 6375 4767 6381
rect 4709 6372 4721 6375
rect 4223 6344 4721 6372
rect 4223 6245 4251 6344
rect 4709 6341 4721 6344
rect 4755 6372 4767 6375
rect 9122 6372 9128 6384
rect 4755 6344 9128 6372
rect 4755 6341 4767 6344
rect 4709 6335 4767 6341
rect 9122 6332 9128 6344
rect 9180 6332 9186 6384
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 10410 6372 10416 6384
rect 9272 6344 9674 6372
rect 10323 6344 10416 6372
rect 9272 6332 9278 6344
rect 4295 6307 4353 6313
rect 4295 6273 4307 6307
rect 4341 6304 4353 6307
rect 4890 6304 4896 6316
rect 4341 6276 4896 6304
rect 4341 6273 4353 6276
rect 4295 6267 4353 6273
rect 4890 6264 4896 6276
rect 4948 6304 4954 6316
rect 5261 6307 5319 6313
rect 5261 6304 5273 6307
rect 4948 6276 5273 6304
rect 4948 6264 4954 6276
rect 5261 6273 5273 6276
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 7432 6276 7481 6304
rect 7432 6264 7438 6276
rect 7469 6273 7481 6276
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 1740 6239 1798 6245
rect 1740 6205 1752 6239
rect 1786 6236 1798 6239
rect 4208 6239 4266 6245
rect 1786 6208 2268 6236
rect 1786 6205 1798 6208
rect 1740 6199 1798 6205
rect 2240 6112 2268 6208
rect 4208 6205 4220 6239
rect 4254 6205 4266 6239
rect 9646 6236 9674 6344
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9646 6208 9965 6236
rect 4208 6199 4266 6205
rect 9953 6205 9965 6208
rect 9999 6236 10011 6239
rect 10042 6236 10048 6248
rect 9999 6208 10048 6236
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 10336 6245 10364 6344
rect 10410 6332 10416 6344
rect 10468 6372 10474 6384
rect 11882 6372 11888 6384
rect 10468 6344 11888 6372
rect 10468 6332 10474 6344
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 13786 6372 13814 6412
rect 15470 6400 15476 6452
rect 15528 6440 15534 6452
rect 16117 6443 16175 6449
rect 16117 6440 16129 6443
rect 15528 6412 16129 6440
rect 15528 6400 15534 6412
rect 16117 6409 16129 6412
rect 16163 6409 16175 6443
rect 16117 6403 16175 6409
rect 18690 6400 18696 6452
rect 18748 6440 18754 6452
rect 23106 6440 23112 6452
rect 18748 6412 23112 6440
rect 18748 6400 18754 6412
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 23658 6400 23664 6452
rect 23716 6440 23722 6452
rect 24762 6440 24768 6452
rect 23716 6412 24768 6440
rect 23716 6400 23722 6412
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 25222 6440 25228 6452
rect 25135 6412 25228 6440
rect 25222 6400 25228 6412
rect 25280 6440 25286 6452
rect 27614 6440 27620 6452
rect 25280 6412 27620 6440
rect 25280 6400 25286 6412
rect 27614 6400 27620 6412
rect 27672 6400 27678 6452
rect 15378 6372 15384 6384
rect 13786 6344 15384 6372
rect 15378 6332 15384 6344
rect 15436 6372 15442 6384
rect 15749 6375 15807 6381
rect 15749 6372 15761 6375
rect 15436 6344 15761 6372
rect 15436 6332 15442 6344
rect 15749 6341 15761 6344
rect 15795 6341 15807 6375
rect 15749 6335 15807 6341
rect 19518 6332 19524 6384
rect 19576 6372 19582 6384
rect 20717 6375 20775 6381
rect 20717 6372 20729 6375
rect 19576 6344 20729 6372
rect 19576 6332 19582 6344
rect 20717 6341 20729 6344
rect 20763 6372 20775 6375
rect 22186 6372 22192 6384
rect 20763 6344 22192 6372
rect 20763 6341 20775 6344
rect 20717 6335 20775 6341
rect 22186 6332 22192 6344
rect 22244 6372 22250 6384
rect 22557 6375 22615 6381
rect 22557 6372 22569 6375
rect 22244 6344 22569 6372
rect 22244 6332 22250 6344
rect 22557 6341 22569 6344
rect 22603 6372 22615 6375
rect 24394 6372 24400 6384
rect 22603 6344 24400 6372
rect 22603 6341 22615 6344
rect 22557 6335 22615 6341
rect 24394 6332 24400 6344
rect 24452 6332 24458 6384
rect 11514 6264 11520 6316
rect 11572 6304 11578 6316
rect 12802 6304 12808 6316
rect 11572 6276 12808 6304
rect 11572 6264 11578 6276
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 14369 6307 14427 6313
rect 14369 6304 14381 6307
rect 13228 6276 14381 6304
rect 13228 6264 13234 6276
rect 14369 6273 14381 6276
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6304 16543 6307
rect 16850 6304 16856 6316
rect 16531 6276 16856 6304
rect 16531 6273 16543 6276
rect 16485 6267 16543 6273
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 21634 6304 21640 6316
rect 21595 6276 21640 6304
rect 21634 6264 21640 6276
rect 21692 6264 21698 6316
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6205 10379 6239
rect 10321 6199 10379 6205
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6236 10655 6239
rect 10686 6236 10692 6248
rect 10643 6208 10692 6236
rect 10643 6205 10655 6208
rect 10597 6199 10655 6205
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 11238 6236 11244 6248
rect 11103 6208 11244 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17736 6208 18061 6236
rect 17736 6196 17742 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 19797 6239 19855 6245
rect 19797 6205 19809 6239
rect 19843 6236 19855 6239
rect 20254 6236 20260 6248
rect 19843 6208 20260 6236
rect 19843 6205 19855 6208
rect 19797 6199 19855 6205
rect 20254 6196 20260 6208
rect 20312 6196 20318 6248
rect 5350 6168 5356 6180
rect 5311 6140 5356 6168
rect 5350 6128 5356 6140
rect 5408 6128 5414 6180
rect 5902 6168 5908 6180
rect 5863 6140 5908 6168
rect 5902 6128 5908 6140
rect 5960 6128 5966 6180
rect 7190 6168 7196 6180
rect 6196 6140 7098 6168
rect 7151 6140 7196 6168
rect 6196 6112 6224 6140
rect 2222 6100 2228 6112
rect 2183 6072 2228 6100
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 6178 6100 6184 6112
rect 6139 6072 6184 6100
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 7070 6100 7098 6140
rect 7190 6128 7196 6140
rect 7248 6128 7254 6180
rect 7285 6171 7343 6177
rect 7285 6137 7297 6171
rect 7331 6137 7343 6171
rect 7285 6131 7343 6137
rect 7300 6100 7328 6131
rect 7926 6128 7932 6180
rect 7984 6168 7990 6180
rect 8665 6171 8723 6177
rect 8665 6168 8677 6171
rect 7984 6140 8677 6168
rect 7984 6128 7990 6140
rect 8665 6137 8677 6140
rect 8711 6137 8723 6171
rect 8665 6131 8723 6137
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 9585 6171 9643 6177
rect 9585 6168 9597 6171
rect 8812 6140 9597 6168
rect 8812 6128 8818 6140
rect 9585 6137 9597 6140
rect 9631 6168 9643 6171
rect 10870 6168 10876 6180
rect 9631 6140 10876 6168
rect 9631 6137 9643 6140
rect 9585 6131 9643 6137
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 11885 6171 11943 6177
rect 11885 6137 11897 6171
rect 11931 6168 11943 6171
rect 12250 6168 12256 6180
rect 11931 6140 12256 6168
rect 11931 6137 11943 6140
rect 11885 6131 11943 6137
rect 12250 6128 12256 6140
rect 12308 6128 12314 6180
rect 12526 6168 12532 6180
rect 12487 6140 12532 6168
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 12621 6171 12679 6177
rect 12621 6137 12633 6171
rect 12667 6168 12679 6171
rect 13906 6168 13912 6180
rect 12667 6140 13912 6168
rect 12667 6137 12679 6140
rect 12621 6131 12679 6137
rect 8202 6100 8208 6112
rect 7070 6072 7328 6100
rect 8163 6072 8208 6100
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8570 6100 8576 6112
rect 8531 6072 8576 6100
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 9950 6100 9956 6112
rect 9911 6072 9956 6100
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 10686 6060 10692 6112
rect 10744 6100 10750 6112
rect 11425 6103 11483 6109
rect 11425 6100 11437 6103
rect 10744 6072 11437 6100
rect 10744 6060 10750 6072
rect 11425 6069 11437 6072
rect 11471 6069 11483 6103
rect 11425 6063 11483 6069
rect 12066 6060 12072 6112
rect 12124 6100 12130 6112
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 12124 6072 12173 6100
rect 12124 6060 12130 6072
rect 12161 6069 12173 6072
rect 12207 6100 12219 6103
rect 12636 6100 12664 6131
rect 13906 6128 13912 6140
rect 13964 6128 13970 6180
rect 14082 6171 14140 6177
rect 14082 6137 14094 6171
rect 14128 6137 14140 6171
rect 14082 6131 14140 6137
rect 13722 6100 13728 6112
rect 12207 6072 12664 6100
rect 13683 6072 13728 6100
rect 12207 6069 12219 6072
rect 12161 6063 12219 6069
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 14108 6100 14136 6131
rect 14182 6128 14188 6180
rect 14240 6168 14246 6180
rect 15013 6171 15071 6177
rect 15013 6168 15025 6171
rect 14240 6140 15025 6168
rect 14240 6128 14246 6140
rect 15013 6137 15025 6140
rect 15059 6137 15071 6171
rect 16574 6168 16580 6180
rect 16535 6140 16580 6168
rect 15013 6131 15071 6137
rect 16574 6128 16580 6140
rect 16632 6128 16638 6180
rect 17129 6171 17187 6177
rect 17129 6137 17141 6171
rect 17175 6168 17187 6171
rect 18230 6168 18236 6180
rect 17175 6140 18236 6168
rect 17175 6137 17187 6140
rect 17129 6131 17187 6137
rect 18230 6128 18236 6140
rect 18288 6128 18294 6180
rect 18370 6171 18428 6177
rect 18370 6137 18382 6171
rect 18416 6168 18428 6171
rect 19245 6171 19303 6177
rect 19245 6168 19257 6171
rect 18416 6140 19257 6168
rect 18416 6137 18428 6140
rect 18370 6131 18428 6137
rect 19245 6137 19257 6140
rect 19291 6168 19303 6171
rect 19978 6168 19984 6180
rect 19291 6140 19984 6168
rect 19291 6137 19303 6140
rect 19245 6131 19303 6137
rect 14550 6100 14556 6112
rect 14108 6072 14556 6100
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 15378 6100 15384 6112
rect 15339 6072 15384 6100
rect 15378 6060 15384 6072
rect 15436 6100 15442 6112
rect 15654 6100 15660 6112
rect 15436 6072 15660 6100
rect 15436 6060 15442 6072
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 17402 6100 17408 6112
rect 17363 6072 17408 6100
rect 17402 6060 17408 6072
rect 17460 6100 17466 6112
rect 17773 6103 17831 6109
rect 17773 6100 17785 6103
rect 17460 6072 17785 6100
rect 17460 6060 17466 6072
rect 17773 6069 17785 6072
rect 17819 6100 17831 6103
rect 18138 6100 18144 6112
rect 17819 6072 18144 6100
rect 17819 6069 17831 6072
rect 17773 6063 17831 6069
rect 18138 6060 18144 6072
rect 18196 6100 18202 6112
rect 18385 6100 18413 6131
rect 19978 6128 19984 6140
rect 20036 6168 20042 6180
rect 20118 6171 20176 6177
rect 20118 6168 20130 6171
rect 20036 6140 20130 6168
rect 20036 6128 20042 6140
rect 20118 6137 20130 6140
rect 20164 6137 20176 6171
rect 20118 6131 20176 6137
rect 21729 6171 21787 6177
rect 21729 6137 21741 6171
rect 21775 6137 21787 6171
rect 22278 6168 22284 6180
rect 22239 6140 22284 6168
rect 21729 6131 21787 6137
rect 18966 6100 18972 6112
rect 18196 6072 18413 6100
rect 18927 6072 18972 6100
rect 18196 6060 18202 6072
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 19518 6060 19524 6112
rect 19576 6100 19582 6112
rect 19613 6103 19671 6109
rect 19613 6100 19625 6103
rect 19576 6072 19625 6100
rect 19576 6060 19582 6072
rect 19613 6069 19625 6072
rect 19659 6069 19671 6103
rect 19613 6063 19671 6069
rect 21453 6103 21511 6109
rect 21453 6069 21465 6103
rect 21499 6100 21511 6103
rect 21744 6100 21772 6131
rect 22278 6128 22284 6140
rect 22336 6128 22342 6180
rect 23753 6171 23811 6177
rect 23753 6168 23765 6171
rect 23446 6140 23765 6168
rect 23446 6112 23474 6140
rect 23753 6137 23765 6140
rect 23799 6137 23811 6171
rect 23753 6131 23811 6137
rect 23845 6171 23903 6177
rect 23845 6137 23857 6171
rect 23891 6168 23903 6171
rect 24026 6168 24032 6180
rect 23891 6140 24032 6168
rect 23891 6137 23903 6140
rect 23845 6131 23903 6137
rect 24026 6128 24032 6140
rect 24084 6128 24090 6180
rect 24397 6171 24455 6177
rect 24397 6137 24409 6171
rect 24443 6168 24455 6171
rect 24854 6168 24860 6180
rect 24443 6140 24860 6168
rect 24443 6137 24455 6140
rect 24397 6131 24455 6137
rect 24854 6128 24860 6140
rect 24912 6128 24918 6180
rect 21818 6100 21824 6112
rect 21499 6072 21824 6100
rect 21499 6069 21511 6072
rect 21453 6063 21511 6069
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 23106 6100 23112 6112
rect 23067 6072 23112 6100
rect 23106 6060 23112 6072
rect 23164 6060 23170 6112
rect 23382 6100 23388 6112
rect 23343 6072 23388 6100
rect 23382 6060 23388 6072
rect 23440 6072 23474 6112
rect 23440 6060 23446 6072
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 6638 5896 6644 5908
rect 6551 5868 6644 5896
rect 6638 5856 6644 5868
rect 6696 5896 6702 5908
rect 7926 5896 7932 5908
rect 6696 5868 7932 5896
rect 6696 5856 6702 5868
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 8110 5896 8116 5908
rect 8071 5868 8116 5896
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8628 5868 9137 5896
rect 8628 5856 8634 5868
rect 9125 5865 9137 5868
rect 9171 5896 9183 5899
rect 9766 5896 9772 5908
rect 9171 5868 9772 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 9953 5899 10011 5905
rect 9953 5865 9965 5899
rect 9999 5896 10011 5899
rect 10042 5896 10048 5908
rect 9999 5868 10048 5896
rect 9999 5865 10011 5868
rect 9953 5859 10011 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 11514 5896 11520 5908
rect 11475 5868 11520 5896
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 12526 5856 12532 5908
rect 12584 5896 12590 5908
rect 12989 5899 13047 5905
rect 12989 5896 13001 5899
rect 12584 5868 13001 5896
rect 12584 5856 12590 5868
rect 12989 5865 13001 5868
rect 13035 5865 13047 5899
rect 17034 5896 17040 5908
rect 12989 5859 13047 5865
rect 16500 5868 17040 5896
rect 6181 5831 6239 5837
rect 6181 5797 6193 5831
rect 6227 5828 6239 5831
rect 6730 5828 6736 5840
rect 6227 5800 6736 5828
rect 6227 5797 6239 5800
rect 6181 5791 6239 5797
rect 6730 5788 6736 5800
rect 6788 5788 6794 5840
rect 7098 5788 7104 5840
rect 7156 5828 7162 5840
rect 7193 5831 7251 5837
rect 7193 5828 7205 5831
rect 7156 5800 7205 5828
rect 7156 5788 7162 5800
rect 7193 5797 7205 5800
rect 7239 5797 7251 5831
rect 7193 5791 7251 5797
rect 9493 5831 9551 5837
rect 9493 5797 9505 5831
rect 9539 5828 9551 5831
rect 9858 5828 9864 5840
rect 9539 5800 9864 5828
rect 9539 5797 9551 5800
rect 9493 5791 9551 5797
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 10550 5831 10608 5837
rect 10550 5797 10562 5831
rect 10596 5828 10608 5831
rect 11054 5828 11060 5840
rect 10596 5800 11060 5828
rect 10596 5797 10608 5800
rect 10550 5791 10608 5797
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 12158 5828 12164 5840
rect 12119 5800 12164 5828
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 12250 5788 12256 5840
rect 12308 5828 12314 5840
rect 13541 5831 13599 5837
rect 13541 5828 13553 5831
rect 12308 5800 13553 5828
rect 12308 5788 12314 5800
rect 13541 5797 13553 5800
rect 13587 5797 13599 5831
rect 13541 5791 13599 5797
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 4522 5760 4528 5772
rect 4479 5732 4528 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 5350 5760 5356 5772
rect 5307 5732 5356 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 5350 5720 5356 5732
rect 5408 5760 5414 5772
rect 6089 5763 6147 5769
rect 6089 5760 6101 5763
rect 5408 5732 6101 5760
rect 5408 5720 5414 5732
rect 6089 5729 6101 5732
rect 6135 5760 6147 5763
rect 6270 5760 6276 5772
rect 6135 5732 6276 5760
rect 6135 5729 6147 5732
rect 6089 5723 6147 5729
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 8608 5763 8666 5769
rect 8608 5760 8620 5763
rect 8444 5732 8620 5760
rect 8444 5720 8450 5732
rect 8608 5729 8620 5732
rect 8654 5729 8666 5763
rect 8608 5723 8666 5729
rect 9950 5720 9956 5772
rect 10008 5760 10014 5772
rect 10229 5763 10287 5769
rect 10229 5760 10241 5763
rect 10008 5732 10241 5760
rect 10008 5720 10014 5732
rect 10229 5729 10241 5732
rect 10275 5729 10287 5763
rect 13630 5760 13636 5772
rect 13591 5732 13636 5760
rect 10229 5723 10287 5729
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 16114 5760 16120 5772
rect 16075 5732 16120 5760
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 16500 5769 16528 5868
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 21818 5896 21824 5908
rect 17460 5868 17902 5896
rect 21779 5868 21824 5896
rect 17460 5856 17466 5868
rect 16669 5831 16727 5837
rect 16669 5797 16681 5831
rect 16715 5828 16727 5831
rect 17678 5828 17684 5840
rect 16715 5800 17684 5828
rect 16715 5797 16727 5800
rect 16669 5791 16727 5797
rect 17678 5788 17684 5800
rect 17736 5788 17742 5840
rect 17874 5837 17902 5868
rect 21818 5856 21824 5868
rect 21876 5856 21882 5908
rect 22094 5896 22100 5908
rect 22055 5868 22100 5896
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 23106 5856 23112 5908
rect 23164 5896 23170 5908
rect 24026 5896 24032 5908
rect 23164 5868 24032 5896
rect 23164 5856 23170 5868
rect 24026 5856 24032 5868
rect 24084 5856 24090 5908
rect 17859 5831 17917 5837
rect 17859 5797 17871 5831
rect 17905 5797 17917 5831
rect 17859 5791 17917 5797
rect 18966 5788 18972 5840
rect 19024 5828 19030 5840
rect 19426 5828 19432 5840
rect 19024 5800 19432 5828
rect 19024 5788 19030 5800
rect 19426 5788 19432 5800
rect 19484 5788 19490 5840
rect 19978 5788 19984 5840
rect 20036 5828 20042 5840
rect 21222 5831 21280 5837
rect 21222 5828 21234 5831
rect 20036 5800 21234 5828
rect 20036 5788 20042 5800
rect 21222 5797 21234 5800
rect 21268 5797 21280 5831
rect 21222 5791 21280 5797
rect 21450 5788 21456 5840
rect 21508 5828 21514 5840
rect 22738 5828 22744 5840
rect 21508 5800 22744 5828
rect 21508 5788 21514 5800
rect 22738 5788 22744 5800
rect 22796 5788 22802 5840
rect 22830 5788 22836 5840
rect 22888 5828 22894 5840
rect 24394 5828 24400 5840
rect 22888 5800 22933 5828
rect 24355 5800 24400 5828
rect 22888 5788 22894 5800
rect 24394 5788 24400 5800
rect 24452 5828 24458 5840
rect 24670 5828 24676 5840
rect 24452 5800 24676 5828
rect 24452 5788 24458 5800
rect 24670 5788 24676 5800
rect 24728 5788 24734 5840
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5729 16543 5763
rect 17696 5760 17724 5788
rect 18693 5763 18751 5769
rect 18693 5760 18705 5763
rect 17696 5732 18705 5760
rect 16485 5723 16543 5729
rect 18693 5729 18705 5732
rect 18739 5729 18751 5763
rect 18693 5723 18751 5729
rect 20622 5720 20628 5772
rect 20680 5760 20686 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20680 5732 20913 5760
rect 20680 5720 20686 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 5902 5652 5908 5704
rect 5960 5692 5966 5704
rect 7101 5695 7159 5701
rect 7101 5692 7113 5695
rect 5960 5664 7113 5692
rect 5960 5652 5966 5664
rect 7101 5661 7113 5664
rect 7147 5661 7159 5695
rect 7374 5692 7380 5704
rect 7335 5664 7380 5692
rect 7101 5655 7159 5661
rect 1578 5624 1584 5636
rect 1539 5596 1584 5624
rect 1578 5584 1584 5596
rect 1636 5584 1642 5636
rect 7116 5624 7144 5655
rect 7374 5652 7380 5664
rect 7432 5652 7438 5704
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5692 11943 5695
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11931 5664 12081 5692
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 12069 5661 12081 5664
rect 12115 5692 12127 5695
rect 13170 5692 13176 5704
rect 12115 5664 13176 5692
rect 12115 5661 12127 5664
rect 12069 5655 12127 5661
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 18230 5652 18236 5704
rect 18288 5692 18294 5704
rect 19337 5695 19395 5701
rect 19337 5692 19349 5695
rect 18288 5664 19349 5692
rect 18288 5652 18294 5664
rect 19337 5661 19349 5664
rect 19383 5661 19395 5695
rect 19337 5655 19395 5661
rect 19981 5695 20039 5701
rect 19981 5661 19993 5695
rect 20027 5692 20039 5695
rect 22278 5692 22284 5704
rect 20027 5664 22284 5692
rect 20027 5661 20039 5664
rect 19981 5655 20039 5661
rect 7926 5624 7932 5636
rect 7116 5596 7932 5624
rect 7926 5584 7932 5596
rect 7984 5584 7990 5636
rect 8711 5627 8769 5633
rect 8711 5593 8723 5627
rect 8757 5624 8769 5627
rect 11330 5624 11336 5636
rect 8757 5596 11336 5624
rect 8757 5593 8769 5596
rect 8711 5587 8769 5593
rect 11330 5584 11336 5596
rect 11388 5584 11394 5636
rect 12621 5627 12679 5633
rect 12621 5593 12633 5627
rect 12667 5624 12679 5627
rect 12710 5624 12716 5636
rect 12667 5596 12716 5624
rect 12667 5593 12679 5596
rect 12621 5587 12679 5593
rect 4571 5559 4629 5565
rect 4571 5525 4583 5559
rect 4617 5556 4629 5559
rect 5074 5556 5080 5568
rect 4617 5528 5080 5556
rect 4617 5525 4629 5528
rect 4571 5519 4629 5525
rect 5074 5516 5080 5528
rect 5132 5516 5138 5568
rect 11146 5556 11152 5568
rect 11107 5528 11152 5556
rect 11146 5516 11152 5528
rect 11204 5516 11210 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 12636 5556 12664 5587
rect 12710 5584 12716 5596
rect 12768 5584 12774 5636
rect 17405 5627 17463 5633
rect 17405 5593 17417 5627
rect 17451 5624 17463 5627
rect 17862 5624 17868 5636
rect 17451 5596 17868 5624
rect 17451 5593 17463 5596
rect 17405 5587 17463 5593
rect 17862 5584 17868 5596
rect 17920 5584 17926 5636
rect 18322 5584 18328 5636
rect 18380 5624 18386 5636
rect 19996 5624 20024 5655
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 23014 5692 23020 5704
rect 22975 5664 23020 5692
rect 23014 5652 23020 5664
rect 23072 5652 23078 5704
rect 24305 5695 24363 5701
rect 24305 5661 24317 5695
rect 24351 5692 24363 5695
rect 25038 5692 25044 5704
rect 24351 5664 25044 5692
rect 24351 5661 24363 5664
rect 24305 5655 24363 5661
rect 25038 5652 25044 5664
rect 25096 5652 25102 5704
rect 18380 5596 20024 5624
rect 18380 5584 18386 5596
rect 20714 5584 20720 5636
rect 20772 5624 20778 5636
rect 22462 5624 22468 5636
rect 20772 5596 22468 5624
rect 20772 5584 20778 5596
rect 22462 5584 22468 5596
rect 22520 5584 22526 5636
rect 24854 5624 24860 5636
rect 24815 5596 24860 5624
rect 24854 5584 24860 5596
rect 24912 5584 24918 5636
rect 12584 5528 12664 5556
rect 13449 5559 13507 5565
rect 12584 5516 12590 5528
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 13538 5556 13544 5568
rect 13495 5528 13544 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 13538 5516 13544 5528
rect 13596 5556 13602 5568
rect 13906 5556 13912 5568
rect 13596 5528 13912 5556
rect 13596 5516 13602 5528
rect 13906 5516 13912 5528
rect 13964 5516 13970 5568
rect 14550 5556 14556 5568
rect 14511 5528 14556 5556
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 14734 5516 14740 5568
rect 14792 5556 14798 5568
rect 14921 5559 14979 5565
rect 14921 5556 14933 5559
rect 14792 5528 14933 5556
rect 14792 5516 14798 5528
rect 14921 5525 14933 5528
rect 14967 5525 14979 5559
rect 18414 5556 18420 5568
rect 18375 5528 18420 5556
rect 14921 5519 14979 5525
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 20254 5556 20260 5568
rect 20215 5528 20260 5556
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 23753 5559 23811 5565
rect 23753 5525 23765 5559
rect 23799 5556 23811 5559
rect 23842 5556 23848 5568
rect 23799 5528 23848 5556
rect 23799 5525 23811 5528
rect 23753 5519 23811 5525
rect 23842 5516 23848 5528
rect 23900 5516 23906 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1811 5355 1869 5361
rect 1811 5352 1823 5355
rect 1452 5324 1823 5352
rect 1452 5312 1458 5324
rect 1811 5321 1823 5324
rect 1857 5321 1869 5355
rect 7374 5352 7380 5364
rect 1811 5315 1869 5321
rect 4126 5324 7380 5352
rect 2225 5287 2283 5293
rect 2225 5253 2237 5287
rect 2271 5284 2283 5287
rect 4126 5284 4154 5324
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 8386 5312 8392 5364
rect 8444 5352 8450 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 8444 5324 8585 5352
rect 8444 5312 8450 5324
rect 8573 5321 8585 5324
rect 8619 5321 8631 5355
rect 8573 5315 8631 5321
rect 9125 5355 9183 5361
rect 9125 5321 9137 5355
rect 9171 5352 9183 5355
rect 9214 5352 9220 5364
rect 9171 5324 9220 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 9732 5324 9777 5352
rect 9732 5312 9738 5324
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11793 5355 11851 5361
rect 11793 5352 11805 5355
rect 11204 5324 11805 5352
rect 11204 5312 11210 5324
rect 11793 5321 11805 5324
rect 11839 5352 11851 5355
rect 12158 5352 12164 5364
rect 11839 5324 12164 5352
rect 11839 5321 11851 5324
rect 11793 5315 11851 5321
rect 12158 5312 12164 5324
rect 12216 5352 12222 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 12216 5324 13553 5352
rect 12216 5312 12222 5324
rect 13541 5321 13553 5324
rect 13587 5352 13599 5355
rect 13630 5352 13636 5364
rect 13587 5324 13636 5352
rect 13587 5321 13599 5324
rect 13541 5315 13599 5321
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 16025 5355 16083 5361
rect 16025 5321 16037 5355
rect 16071 5352 16083 5355
rect 16114 5352 16120 5364
rect 16071 5324 16120 5352
rect 16071 5321 16083 5324
rect 16025 5315 16083 5321
rect 16114 5312 16120 5324
rect 16172 5312 16178 5364
rect 19426 5352 19432 5364
rect 19387 5324 19432 5352
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 19978 5312 19984 5364
rect 20036 5352 20042 5364
rect 20257 5355 20315 5361
rect 20257 5352 20269 5355
rect 20036 5324 20269 5352
rect 20036 5312 20042 5324
rect 20257 5321 20269 5324
rect 20303 5352 20315 5355
rect 21637 5355 21695 5361
rect 21637 5352 21649 5355
rect 20303 5324 21649 5352
rect 20303 5321 20315 5324
rect 20257 5315 20315 5321
rect 21637 5321 21649 5324
rect 21683 5321 21695 5355
rect 21637 5315 21695 5321
rect 22738 5312 22744 5364
rect 22796 5352 22802 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22796 5324 23029 5352
rect 22796 5312 22802 5324
rect 23017 5321 23029 5324
rect 23063 5321 23075 5355
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 23017 5315 23075 5321
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 25038 5352 25044 5364
rect 24999 5324 25044 5352
rect 25038 5312 25044 5324
rect 25096 5352 25102 5364
rect 25363 5355 25421 5361
rect 25363 5352 25375 5355
rect 25096 5324 25375 5352
rect 25096 5312 25102 5324
rect 25363 5321 25375 5324
rect 25409 5321 25421 5355
rect 25363 5315 25421 5321
rect 2271 5256 4154 5284
rect 2271 5253 2283 5256
rect 2225 5247 2283 5253
rect 1740 5151 1798 5157
rect 1740 5117 1752 5151
rect 1786 5148 1798 5151
rect 2240 5148 2268 5247
rect 7190 5244 7196 5296
rect 7248 5284 7254 5296
rect 7929 5287 7987 5293
rect 7929 5284 7941 5287
rect 7248 5256 7941 5284
rect 7248 5244 7254 5256
rect 7929 5253 7941 5256
rect 7975 5253 7987 5287
rect 7929 5247 7987 5253
rect 10689 5287 10747 5293
rect 10689 5253 10701 5287
rect 10735 5284 10747 5287
rect 12253 5287 12311 5293
rect 12253 5284 12265 5287
rect 10735 5256 12265 5284
rect 10735 5253 10747 5256
rect 10689 5247 10747 5253
rect 5905 5219 5963 5225
rect 5905 5185 5917 5219
rect 5951 5216 5963 5219
rect 6178 5216 6184 5228
rect 5951 5188 6184 5216
rect 5951 5185 5963 5188
rect 5905 5179 5963 5185
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 7377 5219 7435 5225
rect 6328 5188 7236 5216
rect 6328 5176 6334 5188
rect 4522 5148 4528 5160
rect 1786 5120 2268 5148
rect 4483 5120 4528 5148
rect 1786 5117 1798 5120
rect 1740 5111 1798 5117
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5148 5135 5151
rect 5813 5151 5871 5157
rect 5813 5148 5825 5151
rect 5123 5120 5825 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5813 5117 5825 5120
rect 5859 5148 5871 5151
rect 5859 5120 6684 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6656 5024 6684 5120
rect 7208 5089 7236 5188
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 8110 5216 8116 5228
rect 7423 5188 8116 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 9214 5108 9220 5160
rect 9272 5148 9278 5160
rect 11440 5157 11468 5256
rect 12253 5253 12265 5256
rect 12299 5284 12311 5287
rect 12434 5284 12440 5296
rect 12299 5256 12440 5284
rect 12299 5253 12311 5256
rect 12253 5247 12311 5253
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 17218 5284 17224 5296
rect 17052 5256 17224 5284
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5216 11575 5219
rect 12066 5216 12072 5228
rect 11563 5188 12072 5216
rect 11563 5185 11575 5188
rect 11517 5179 11575 5185
rect 12066 5176 12072 5188
rect 12124 5176 12130 5228
rect 13170 5216 13176 5228
rect 13131 5188 13176 5216
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5216 15715 5219
rect 17052 5216 17080 5256
rect 17218 5244 17224 5256
rect 17276 5284 17282 5296
rect 20346 5284 20352 5296
rect 17276 5256 20352 5284
rect 17276 5244 17282 5256
rect 20346 5244 20352 5256
rect 20404 5244 20410 5296
rect 23750 5284 23756 5296
rect 23711 5256 23756 5284
rect 23750 5244 23756 5256
rect 23808 5244 23814 5296
rect 15703 5188 17080 5216
rect 17129 5219 17187 5225
rect 15703 5185 15715 5188
rect 15657 5179 15715 5185
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 9272 5120 9321 5148
rect 9272 5108 9278 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 11425 5151 11483 5157
rect 11425 5117 11437 5151
rect 11471 5117 11483 5151
rect 13998 5148 14004 5160
rect 11425 5111 11483 5117
rect 13786 5120 14004 5148
rect 7193 5083 7251 5089
rect 7193 5049 7205 5083
rect 7239 5080 7251 5083
rect 7469 5083 7527 5089
rect 7469 5080 7481 5083
rect 7239 5052 7481 5080
rect 7239 5049 7251 5052
rect 7193 5043 7251 5049
rect 7469 5049 7481 5052
rect 7515 5080 7527 5083
rect 7834 5080 7840 5092
rect 7515 5052 7840 5080
rect 7515 5049 7527 5052
rect 7469 5043 7527 5049
rect 7834 5040 7840 5052
rect 7892 5040 7898 5092
rect 9398 5040 9404 5092
rect 9456 5080 9462 5092
rect 10962 5080 10968 5092
rect 9456 5052 10968 5080
rect 9456 5040 9462 5052
rect 10962 5040 10968 5052
rect 11020 5040 11026 5092
rect 12526 5080 12532 5092
rect 12487 5052 12532 5080
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 12621 5083 12679 5089
rect 12621 5049 12633 5083
rect 12667 5049 12679 5083
rect 12621 5043 12679 5049
rect 6638 5012 6644 5024
rect 6599 4984 6644 5012
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 7282 4972 7288 5024
rect 7340 5012 7346 5024
rect 10229 5015 10287 5021
rect 10229 5012 10241 5015
rect 7340 4984 10241 5012
rect 7340 4972 7346 4984
rect 10229 4981 10241 4984
rect 10275 4981 10287 5015
rect 10229 4975 10287 4981
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12636 5012 12664 5043
rect 13786 5024 13814 5120
rect 13998 5108 14004 5120
rect 14056 5148 14062 5160
rect 16684 5157 16712 5188
rect 17129 5185 17141 5219
rect 17175 5216 17187 5219
rect 17494 5216 17500 5228
rect 17175 5188 17500 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 17494 5176 17500 5188
rect 17552 5176 17558 5228
rect 18230 5176 18236 5228
rect 18288 5216 18294 5228
rect 18417 5219 18475 5225
rect 18417 5216 18429 5219
rect 18288 5188 18429 5216
rect 18288 5176 18294 5188
rect 18417 5185 18429 5188
rect 18463 5216 18475 5219
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 18463 5188 19809 5216
rect 18463 5185 18475 5188
rect 18417 5179 18475 5185
rect 19797 5185 19809 5188
rect 19843 5185 19855 5219
rect 19797 5179 19855 5185
rect 22189 5219 22247 5225
rect 22189 5185 22201 5219
rect 22235 5216 22247 5219
rect 23382 5216 23388 5228
rect 22235 5188 23388 5216
rect 22235 5185 22247 5188
rect 22189 5179 22247 5185
rect 23382 5176 23388 5188
rect 23440 5176 23446 5228
rect 23842 5176 23848 5228
rect 23900 5216 23906 5228
rect 24118 5216 24124 5228
rect 23900 5188 23980 5216
rect 24079 5188 24124 5216
rect 23900 5176 23906 5188
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 14056 5120 14289 5148
rect 14056 5108 14062 5120
rect 14277 5117 14289 5120
rect 14323 5148 14335 5151
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 14323 5120 14473 5148
rect 14323 5117 14335 5120
rect 14277 5111 14335 5117
rect 14461 5117 14473 5120
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 16945 5151 17003 5157
rect 16945 5117 16957 5151
rect 16991 5148 17003 5151
rect 17034 5148 17040 5160
rect 16991 5120 17040 5148
rect 16991 5117 17003 5120
rect 16945 5111 17003 5117
rect 17034 5108 17040 5120
rect 17092 5108 17098 5160
rect 20438 5148 20444 5160
rect 20399 5120 20444 5148
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 22370 5148 22376 5160
rect 20640 5120 22376 5148
rect 15105 5083 15163 5089
rect 15105 5049 15117 5083
rect 15151 5080 15163 5083
rect 16758 5080 16764 5092
rect 15151 5052 16764 5080
rect 15151 5049 15163 5052
rect 15105 5043 15163 5049
rect 16758 5040 16764 5052
rect 16816 5040 16822 5092
rect 17310 5040 17316 5092
rect 17368 5080 17374 5092
rect 18138 5080 18144 5092
rect 17368 5052 18144 5080
rect 17368 5040 17374 5052
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 18233 5083 18291 5089
rect 18233 5049 18245 5083
rect 18279 5080 18291 5083
rect 18414 5080 18420 5092
rect 18279 5052 18420 5080
rect 18279 5049 18291 5052
rect 18233 5043 18291 5049
rect 18414 5040 18420 5052
rect 18472 5080 18478 5092
rect 19061 5083 19119 5089
rect 19061 5080 19073 5083
rect 18472 5052 19073 5080
rect 18472 5040 18478 5052
rect 19061 5049 19073 5052
rect 19107 5080 19119 5083
rect 20640 5080 20668 5120
rect 22370 5108 22376 5120
rect 22428 5148 22434 5160
rect 22649 5151 22707 5157
rect 22649 5148 22661 5151
rect 22428 5120 22661 5148
rect 22428 5108 22434 5120
rect 22649 5117 22661 5120
rect 22695 5148 22707 5151
rect 22830 5148 22836 5160
rect 22695 5120 22836 5148
rect 22695 5117 22707 5120
rect 22649 5111 22707 5117
rect 22830 5108 22836 5120
rect 22888 5108 22894 5160
rect 23952 5157 23980 5188
rect 24118 5176 24124 5188
rect 24176 5176 24182 5228
rect 23477 5151 23535 5157
rect 23477 5148 23489 5151
rect 22940 5120 23489 5148
rect 19107 5052 20668 5080
rect 19107 5049 19119 5052
rect 19061 5043 19119 5049
rect 20898 5040 20904 5092
rect 20956 5080 20962 5092
rect 22940 5080 22968 5120
rect 23477 5117 23489 5120
rect 23523 5148 23535 5151
rect 23661 5151 23719 5157
rect 23661 5148 23673 5151
rect 23523 5120 23673 5148
rect 23523 5117 23535 5120
rect 23477 5111 23535 5117
rect 23661 5117 23673 5120
rect 23707 5117 23719 5151
rect 23661 5111 23719 5117
rect 23937 5151 23995 5157
rect 23937 5117 23949 5151
rect 23983 5117 23995 5151
rect 23937 5111 23995 5117
rect 25292 5151 25350 5157
rect 25292 5117 25304 5151
rect 25338 5148 25350 5151
rect 25777 5151 25835 5157
rect 25777 5148 25789 5151
rect 25338 5120 25789 5148
rect 25338 5117 25350 5120
rect 25292 5111 25350 5117
rect 25777 5117 25789 5120
rect 25823 5148 25835 5151
rect 27614 5148 27620 5160
rect 25823 5120 27620 5148
rect 25823 5117 25835 5120
rect 25777 5111 25835 5117
rect 27614 5108 27620 5120
rect 27672 5108 27678 5160
rect 20956 5052 22968 5080
rect 20956 5040 20962 5052
rect 12492 4984 12664 5012
rect 12492 4972 12498 4984
rect 13722 4972 13728 5024
rect 13780 4984 13814 5024
rect 13780 4972 13786 4984
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 17402 5012 17408 5024
rect 16172 4984 17408 5012
rect 16172 4972 16178 4984
rect 17402 4972 17408 4984
rect 17460 5012 17466 5024
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 17460 4984 17509 5012
rect 17460 4972 17466 4984
rect 17497 4981 17509 4984
rect 17543 4981 17555 5015
rect 17497 4975 17555 4981
rect 19978 4972 19984 5024
rect 20036 5012 20042 5024
rect 20809 5015 20867 5021
rect 20809 5012 20821 5015
rect 20036 4984 20821 5012
rect 20036 4972 20042 4984
rect 20809 4981 20821 4984
rect 20855 4981 20867 5015
rect 21358 5012 21364 5024
rect 21319 4984 21364 5012
rect 20809 4975 20867 4981
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1394 4768 1400 4820
rect 1452 4808 1458 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1452 4780 1593 4808
rect 1452 4768 1458 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1581 4771 1639 4777
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 7098 4808 7104 4820
rect 6696 4780 7104 4808
rect 6696 4768 6702 4780
rect 7098 4768 7104 4780
rect 7156 4808 7162 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7156 4780 7849 4808
rect 7156 4768 7162 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 7926 4768 7932 4820
rect 7984 4808 7990 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 7984 4780 8125 4808
rect 7984 4768 7990 4780
rect 8113 4777 8125 4780
rect 8159 4777 8171 4811
rect 8113 4771 8171 4777
rect 9493 4811 9551 4817
rect 9493 4777 9505 4811
rect 9539 4808 9551 4811
rect 9950 4808 9956 4820
rect 9539 4780 9956 4808
rect 9539 4777 9551 4780
rect 9493 4771 9551 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 14826 4808 14832 4820
rect 10657 4780 11560 4808
rect 14787 4780 14832 4808
rect 7190 4740 7196 4752
rect 7151 4712 7196 4740
rect 7190 4700 7196 4712
rect 7248 4700 7254 4752
rect 8757 4743 8815 4749
rect 8757 4709 8769 4743
rect 8803 4740 8815 4743
rect 10657 4740 10685 4780
rect 11532 4752 11560 4780
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 15427 4811 15485 4817
rect 15427 4777 15439 4811
rect 15473 4808 15485 4811
rect 17310 4808 17316 4820
rect 15473 4780 17316 4808
rect 15473 4777 15485 4780
rect 15427 4771 15485 4777
rect 17310 4768 17316 4780
rect 17368 4768 17374 4820
rect 17494 4808 17500 4820
rect 17455 4780 17500 4808
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 18138 4768 18144 4820
rect 18196 4808 18202 4820
rect 18601 4811 18659 4817
rect 18601 4808 18613 4811
rect 18196 4780 18613 4808
rect 18196 4768 18202 4780
rect 18601 4777 18613 4780
rect 18647 4777 18659 4811
rect 18601 4771 18659 4777
rect 20622 4768 20628 4820
rect 20680 4808 20686 4820
rect 21361 4811 21419 4817
rect 21361 4808 21373 4811
rect 20680 4780 21373 4808
rect 20680 4768 20686 4780
rect 21361 4777 21373 4780
rect 21407 4777 21419 4811
rect 23750 4808 23756 4820
rect 23711 4780 23756 4808
rect 21361 4771 21419 4777
rect 23750 4768 23756 4780
rect 23808 4768 23814 4820
rect 10962 4740 10968 4752
rect 8803 4712 10685 4740
rect 10923 4712 10968 4740
rect 8803 4709 8815 4712
rect 8757 4703 8815 4709
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 11514 4740 11520 4752
rect 11427 4712 11520 4740
rect 11514 4700 11520 4712
rect 11572 4700 11578 4752
rect 13814 4700 13820 4752
rect 13872 4740 13878 4752
rect 18417 4743 18475 4749
rect 18417 4740 18429 4743
rect 13872 4712 18429 4740
rect 13872 4700 13878 4712
rect 18417 4709 18429 4712
rect 18463 4709 18475 4743
rect 18417 4703 18475 4709
rect 19981 4743 20039 4749
rect 19981 4709 19993 4743
rect 20027 4740 20039 4743
rect 20438 4740 20444 4752
rect 20027 4712 20444 4740
rect 20027 4709 20039 4712
rect 19981 4703 20039 4709
rect 20438 4700 20444 4712
rect 20496 4700 20502 4752
rect 22370 4740 22376 4752
rect 22331 4712 22376 4740
rect 22370 4700 22376 4712
rect 22428 4700 22434 4752
rect 5972 4675 6030 4681
rect 5972 4641 5984 4675
rect 6018 4672 6030 4675
rect 6178 4672 6184 4684
rect 6018 4644 6184 4672
rect 6018 4641 6030 4644
rect 5972 4635 6030 4641
rect 6178 4632 6184 4644
rect 6236 4672 6242 4684
rect 9398 4672 9404 4684
rect 6236 4644 9404 4672
rect 6236 4632 6242 4644
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 9582 4632 9588 4684
rect 9640 4672 9646 4684
rect 9674 4672 9680 4684
rect 9640 4644 9680 4672
rect 9640 4632 9646 4644
rect 9674 4632 9680 4644
rect 9732 4672 9738 4684
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 9732 4644 10609 4672
rect 9732 4632 9738 4644
rect 10597 4641 10609 4644
rect 10643 4641 10655 4675
rect 10597 4635 10655 4641
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4672 12311 4675
rect 12986 4672 12992 4684
rect 12299 4644 12992 4672
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 12986 4632 12992 4644
rect 13044 4632 13050 4684
rect 13909 4675 13967 4681
rect 13909 4641 13921 4675
rect 13955 4672 13967 4675
rect 14550 4672 14556 4684
rect 13955 4644 14556 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 15356 4675 15414 4681
rect 15356 4641 15368 4675
rect 15402 4672 15414 4675
rect 15746 4672 15752 4684
rect 15402 4644 15752 4672
rect 15402 4641 15414 4644
rect 15356 4635 15414 4641
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 16758 4672 16764 4684
rect 16719 4644 16764 4672
rect 16758 4632 16764 4644
rect 16816 4632 16822 4684
rect 18208 4675 18266 4681
rect 18208 4641 18220 4675
rect 18254 4672 18266 4675
rect 18322 4672 18328 4684
rect 18254 4644 18328 4672
rect 18254 4641 18266 4644
rect 18208 4635 18266 4641
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 18598 4632 18604 4684
rect 18656 4672 18662 4684
rect 19242 4672 19248 4684
rect 18656 4644 19248 4672
rect 18656 4632 18662 4644
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 19797 4675 19855 4681
rect 19797 4641 19809 4675
rect 19843 4672 19855 4675
rect 20162 4672 20168 4684
rect 19843 4644 20168 4672
rect 19843 4641 19855 4644
rect 19797 4635 19855 4641
rect 20162 4632 20168 4644
rect 20220 4632 20226 4684
rect 20968 4675 21026 4681
rect 20968 4641 20980 4675
rect 21014 4672 21026 4675
rect 21014 4641 21036 4672
rect 20968 4635 21036 4641
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4604 6515 4607
rect 6917 4607 6975 4613
rect 6917 4604 6929 4607
rect 6503 4576 6929 4604
rect 6503 4573 6515 4576
rect 6457 4567 6515 4573
rect 6917 4573 6929 4576
rect 6963 4604 6975 4607
rect 7006 4604 7012 4616
rect 6963 4576 7012 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 9766 4604 9772 4616
rect 9727 4576 9772 4604
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 12342 4604 12348 4616
rect 12303 4576 12348 4604
rect 10873 4567 10931 4573
rect 6043 4539 6101 4545
rect 6043 4505 6055 4539
rect 6089 4536 6101 4539
rect 10888 4536 10916 4567
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 16298 4604 16304 4616
rect 16259 4576 16304 4604
rect 16298 4564 16304 4576
rect 16356 4564 16362 4616
rect 17770 4564 17776 4616
rect 17828 4604 17834 4616
rect 21008 4604 21036 4635
rect 21729 4607 21787 4613
rect 21729 4604 21741 4607
rect 17828 4576 21741 4604
rect 17828 4564 17834 4576
rect 21729 4573 21741 4576
rect 21775 4573 21787 4607
rect 21729 4567 21787 4573
rect 22281 4607 22339 4613
rect 22281 4573 22293 4607
rect 22327 4604 22339 4607
rect 23014 4604 23020 4616
rect 22327 4576 23020 4604
rect 22327 4573 22339 4576
rect 22281 4567 22339 4573
rect 23014 4564 23020 4576
rect 23072 4564 23078 4616
rect 11330 4536 11336 4548
rect 6089 4508 10732 4536
rect 10888 4508 11336 4536
rect 6089 4505 6101 4508
rect 6043 4499 6101 4505
rect 6822 4468 6828 4480
rect 6783 4440 6828 4468
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 9030 4468 9036 4480
rect 8991 4440 9036 4468
rect 9030 4428 9036 4440
rect 9088 4428 9094 4480
rect 10318 4468 10324 4480
rect 10279 4440 10324 4468
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 10704 4468 10732 4508
rect 11330 4496 11336 4508
rect 11388 4536 11394 4548
rect 13357 4539 13415 4545
rect 13357 4536 13369 4539
rect 11388 4508 13369 4536
rect 11388 4496 11394 4508
rect 13357 4505 13369 4508
rect 13403 4505 13415 4539
rect 13357 4499 13415 4505
rect 14093 4539 14151 4545
rect 14093 4505 14105 4539
rect 14139 4536 14151 4539
rect 14642 4536 14648 4548
rect 14139 4508 14648 4536
rect 14139 4505 14151 4508
rect 14093 4499 14151 4505
rect 14642 4496 14648 4508
rect 14700 4496 14706 4548
rect 15286 4496 15292 4548
rect 15344 4536 15350 4548
rect 18279 4539 18337 4545
rect 18279 4536 18291 4539
rect 15344 4508 18291 4536
rect 15344 4496 15350 4508
rect 18279 4505 18291 4508
rect 18325 4505 18337 4539
rect 18279 4499 18337 4505
rect 18417 4539 18475 4545
rect 18417 4505 18429 4539
rect 18463 4536 18475 4539
rect 21039 4539 21097 4545
rect 21039 4536 21051 4539
rect 18463 4508 21051 4536
rect 18463 4505 18475 4508
rect 18417 4499 18475 4505
rect 21039 4505 21051 4508
rect 21085 4505 21097 4539
rect 21039 4499 21097 4505
rect 22462 4496 22468 4548
rect 22520 4536 22526 4548
rect 22833 4539 22891 4545
rect 22833 4536 22845 4539
rect 22520 4508 22845 4536
rect 22520 4496 22526 4508
rect 22833 4505 22845 4508
rect 22879 4536 22891 4539
rect 24854 4536 24860 4548
rect 22879 4508 24860 4536
rect 22879 4505 22891 4508
rect 22833 4499 22891 4505
rect 24854 4496 24860 4508
rect 24912 4496 24918 4548
rect 11793 4471 11851 4477
rect 11793 4468 11805 4471
rect 10704 4440 11805 4468
rect 11793 4437 11805 4440
rect 11839 4468 11851 4471
rect 12526 4468 12532 4480
rect 11839 4440 12532 4468
rect 11839 4437 11851 4440
rect 11793 4431 11851 4437
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 14274 4428 14280 4480
rect 14332 4468 14338 4480
rect 14461 4471 14519 4477
rect 14461 4468 14473 4471
rect 14332 4440 14473 4468
rect 14332 4428 14338 4440
rect 14461 4437 14473 4440
rect 14507 4437 14519 4471
rect 14461 4431 14519 4437
rect 16025 4471 16083 4477
rect 16025 4437 16037 4471
rect 16071 4468 16083 4471
rect 17034 4468 17040 4480
rect 16071 4440 17040 4468
rect 16071 4437 16083 4440
rect 16025 4431 16083 4437
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 18049 4471 18107 4477
rect 18049 4437 18061 4471
rect 18095 4468 18107 4471
rect 18138 4468 18144 4480
rect 18095 4440 18144 4468
rect 18095 4437 18107 4440
rect 18049 4431 18107 4437
rect 18138 4428 18144 4440
rect 18196 4468 18202 4480
rect 18874 4468 18880 4480
rect 18196 4440 18880 4468
rect 18196 4428 18202 4440
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 22646 4428 22652 4480
rect 22704 4468 22710 4480
rect 23750 4468 23756 4480
rect 22704 4440 23756 4468
rect 22704 4428 22710 4440
rect 23750 4428 23756 4440
rect 23808 4428 23814 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 6178 4264 6184 4276
rect 6139 4236 6184 4264
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 13725 4267 13783 4273
rect 13725 4264 13737 4267
rect 11204 4236 13737 4264
rect 11204 4224 11210 4236
rect 13725 4233 13737 4236
rect 13771 4233 13783 4267
rect 13725 4227 13783 4233
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 15841 4267 15899 4273
rect 15841 4264 15853 4267
rect 15804 4236 15853 4264
rect 15804 4224 15810 4236
rect 15841 4233 15853 4236
rect 15887 4264 15899 4267
rect 16942 4264 16948 4276
rect 15887 4236 16948 4264
rect 15887 4233 15899 4236
rect 15841 4227 15899 4233
rect 16942 4224 16948 4236
rect 17000 4224 17006 4276
rect 17497 4267 17555 4273
rect 17497 4233 17509 4267
rect 17543 4264 17555 4267
rect 18322 4264 18328 4276
rect 17543 4236 18328 4264
rect 17543 4233 17555 4236
rect 17497 4227 17555 4233
rect 18322 4224 18328 4236
rect 18380 4224 18386 4276
rect 19242 4264 19248 4276
rect 19203 4236 19248 4264
rect 19242 4224 19248 4236
rect 19300 4224 19306 4276
rect 21358 4224 21364 4276
rect 21416 4264 21422 4276
rect 21453 4267 21511 4273
rect 21453 4264 21465 4267
rect 21416 4236 21465 4264
rect 21416 4224 21422 4236
rect 21453 4233 21465 4236
rect 21499 4233 21511 4267
rect 21453 4227 21511 4233
rect 22370 4224 22376 4276
rect 22428 4264 22434 4276
rect 22649 4267 22707 4273
rect 22649 4264 22661 4267
rect 22428 4236 22661 4264
rect 22428 4224 22434 4236
rect 22649 4233 22661 4236
rect 22695 4233 22707 4267
rect 23014 4264 23020 4276
rect 22975 4236 23020 4264
rect 22649 4227 22707 4233
rect 23014 4224 23020 4236
rect 23072 4264 23078 4276
rect 24719 4267 24777 4273
rect 24719 4264 24731 4267
rect 23072 4236 24731 4264
rect 23072 4224 23078 4236
rect 24719 4233 24731 4236
rect 24765 4233 24777 4267
rect 24719 4227 24777 4233
rect 12526 4156 12532 4208
rect 12584 4196 12590 4208
rect 13081 4199 13139 4205
rect 13081 4196 13093 4199
rect 12584 4168 13093 4196
rect 12584 4156 12590 4168
rect 13081 4165 13093 4168
rect 13127 4196 13139 4199
rect 14734 4196 14740 4208
rect 13127 4168 14740 4196
rect 13127 4165 13139 4168
rect 13081 4159 13139 4165
rect 14734 4156 14740 4168
rect 14792 4156 14798 4208
rect 20162 4196 20168 4208
rect 20088 4168 20168 4196
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 6512 4100 8493 4128
rect 6512 4088 6518 4100
rect 5077 4063 5135 4069
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5810 4060 5816 4072
rect 5123 4032 5816 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 5092 3924 5120 4023
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 7392 4069 7420 4100
rect 8481 4097 8493 4100
rect 8527 4097 8539 4131
rect 10318 4128 10324 4140
rect 8481 4091 8539 4097
rect 8864 4100 10324 4128
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6880 4032 6929 4060
rect 6880 4020 6886 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 7377 4063 7435 4069
rect 7377 4029 7389 4063
rect 7423 4029 7435 4063
rect 7742 4060 7748 4072
rect 7703 4032 7748 4060
rect 7377 4023 7435 4029
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4060 8171 4063
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8159 4032 8677 4060
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 8665 4029 8677 4032
rect 8711 4060 8723 4063
rect 8864 4060 8892 4100
rect 10318 4088 10324 4100
rect 10376 4128 10382 4140
rect 10376 4100 10824 4128
rect 10376 4088 10382 4100
rect 8711 4032 8892 4060
rect 8711 4029 8723 4032
rect 8665 4023 8723 4029
rect 5905 3995 5963 4001
rect 5905 3961 5917 3995
rect 5951 3992 5963 3995
rect 8128 3992 8156 4023
rect 9582 4020 9588 4072
rect 9640 4060 9646 4072
rect 9861 4063 9919 4069
rect 9861 4060 9873 4063
rect 9640 4032 9873 4060
rect 9640 4020 9646 4032
rect 9861 4029 9873 4032
rect 9907 4029 9919 4063
rect 9861 4023 9919 4029
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4029 10563 4063
rect 10686 4060 10692 4072
rect 10647 4032 10692 4060
rect 10505 4023 10563 4029
rect 5951 3964 8156 3992
rect 8481 3995 8539 4001
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 9769 3995 9827 4001
rect 9769 3992 9781 3995
rect 8527 3964 9781 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 9769 3961 9781 3964
rect 9815 3992 9827 3995
rect 10520 3992 10548 4023
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 10796 4060 10824 4100
rect 10962 4088 10968 4140
rect 11020 4128 11026 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11020 4100 11713 4128
rect 11020 4088 11026 4100
rect 11701 4097 11713 4100
rect 11747 4128 11759 4131
rect 13630 4128 13636 4140
rect 11747 4100 13636 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 13630 4088 13636 4100
rect 13688 4088 13694 4140
rect 13725 4131 13783 4137
rect 13725 4097 13737 4131
rect 13771 4128 13783 4131
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13771 4100 14013 4128
rect 13771 4097 13783 4100
rect 13725 4091 13783 4097
rect 14001 4097 14013 4100
rect 14047 4128 14059 4131
rect 17862 4128 17868 4140
rect 14047 4100 17868 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 11238 4060 11244 4072
rect 10796 4032 11244 4060
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 13541 4063 13599 4069
rect 13541 4029 13553 4063
rect 13587 4060 13599 4063
rect 14090 4060 14096 4072
rect 13587 4032 14096 4060
rect 13587 4029 13599 4032
rect 13541 4023 13599 4029
rect 14090 4020 14096 4032
rect 14148 4020 14154 4072
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 14332 4032 14565 4060
rect 14332 4020 14338 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 14553 4023 14611 4029
rect 14826 4020 14832 4072
rect 14884 4060 14890 4072
rect 15488 4069 15516 4100
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 18138 4128 18144 4140
rect 18099 4100 18144 4128
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 18506 4128 18512 4140
rect 18467 4100 18512 4128
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 14921 4063 14979 4069
rect 14921 4060 14933 4063
rect 14884 4032 14933 4060
rect 14884 4020 14890 4032
rect 14921 4029 14933 4032
rect 14967 4029 14979 4063
rect 14921 4023 14979 4029
rect 15473 4063 15531 4069
rect 15473 4029 15485 4063
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 19889 4063 19947 4069
rect 19889 4029 19901 4063
rect 19935 4060 19947 4063
rect 19978 4060 19984 4072
rect 19935 4032 19984 4060
rect 19935 4029 19947 4032
rect 19889 4023 19947 4029
rect 19978 4020 19984 4032
rect 20036 4020 20042 4072
rect 20088 4069 20116 4168
rect 20162 4156 20168 4168
rect 20220 4196 20226 4208
rect 20625 4199 20683 4205
rect 20625 4196 20637 4199
rect 20220 4168 20637 4196
rect 20220 4156 20226 4168
rect 20625 4165 20637 4168
rect 20671 4165 20683 4199
rect 22278 4196 22284 4208
rect 22239 4168 22284 4196
rect 20625 4159 20683 4165
rect 22278 4156 22284 4168
rect 22336 4156 22342 4208
rect 20254 4128 20260 4140
rect 20215 4100 20260 4128
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 21177 4131 21235 4137
rect 21177 4097 21189 4131
rect 21223 4128 21235 4131
rect 21729 4131 21787 4137
rect 21729 4128 21741 4131
rect 21223 4100 21741 4128
rect 21223 4097 21235 4100
rect 21177 4091 21235 4097
rect 21729 4097 21741 4100
rect 21775 4128 21787 4131
rect 22462 4128 22468 4140
rect 21775 4100 22468 4128
rect 21775 4097 21787 4100
rect 21729 4091 21787 4097
rect 22462 4088 22468 4100
rect 22520 4088 22526 4140
rect 20073 4063 20131 4069
rect 20073 4029 20085 4063
rect 20119 4029 20131 4063
rect 20073 4023 20131 4029
rect 24648 4063 24706 4069
rect 24648 4029 24660 4063
rect 24694 4060 24706 4063
rect 24694 4032 25176 4060
rect 24694 4029 24706 4032
rect 24648 4023 24706 4029
rect 10778 3992 10784 4004
rect 9815 3964 10784 3992
rect 9815 3961 9827 3964
rect 9769 3955 9827 3961
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 11330 3992 11336 4004
rect 11291 3964 11336 3992
rect 11330 3952 11336 3964
rect 11388 3952 11394 4004
rect 12158 3952 12164 4004
rect 12216 3992 12222 4004
rect 12529 3995 12587 4001
rect 12529 3992 12541 3995
rect 12216 3964 12541 3992
rect 12216 3952 12222 3964
rect 12529 3961 12541 3964
rect 12575 3961 12587 3995
rect 12529 3955 12587 3961
rect 12621 3995 12679 4001
rect 12621 3961 12633 3995
rect 12667 3961 12679 3995
rect 15562 3992 15568 4004
rect 15523 3964 15568 3992
rect 12621 3955 12679 3961
rect 3384 3896 5120 3924
rect 3384 3884 3390 3896
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 6512 3896 6561 3924
rect 6512 3884 6518 3896
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 7006 3924 7012 3936
rect 6967 3896 7012 3924
rect 6549 3887 6607 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 9306 3924 9312 3936
rect 8812 3896 9312 3924
rect 8812 3884 8818 3896
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 12253 3927 12311 3933
rect 12253 3893 12265 3927
rect 12299 3924 12311 3927
rect 12434 3924 12440 3936
rect 12299 3896 12440 3924
rect 12299 3893 12311 3896
rect 12253 3887 12311 3893
rect 12434 3884 12440 3896
rect 12492 3924 12498 3936
rect 12636 3924 12664 3955
rect 15562 3952 15568 3964
rect 15620 3952 15626 4004
rect 16482 3992 16488 4004
rect 16443 3964 16488 3992
rect 16482 3952 16488 3964
rect 16540 3952 16546 4004
rect 16577 3995 16635 4001
rect 16577 3961 16589 3995
rect 16623 3961 16635 3995
rect 17126 3992 17132 4004
rect 17087 3964 17132 3992
rect 16577 3955 16635 3961
rect 13538 3924 13544 3936
rect 12492 3896 13544 3924
rect 12492 3884 12498 3896
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 16301 3927 16359 3933
rect 16301 3893 16313 3927
rect 16347 3924 16359 3927
rect 16390 3924 16396 3936
rect 16347 3896 16396 3924
rect 16347 3893 16359 3896
rect 16301 3887 16359 3893
rect 16390 3884 16396 3896
rect 16448 3924 16454 3936
rect 16592 3924 16620 3955
rect 17126 3952 17132 3964
rect 17184 3952 17190 4004
rect 18233 3995 18291 4001
rect 18233 3992 18245 3995
rect 17788 3964 18245 3992
rect 17788 3933 17816 3964
rect 18233 3961 18245 3964
rect 18279 3992 18291 3995
rect 18414 3992 18420 4004
rect 18279 3964 18420 3992
rect 18279 3961 18291 3964
rect 18233 3955 18291 3961
rect 18414 3952 18420 3964
rect 18472 3952 18478 4004
rect 21821 3995 21879 4001
rect 21821 3961 21833 3995
rect 21867 3961 21879 3995
rect 21821 3955 21879 3961
rect 17773 3927 17831 3933
rect 17773 3924 17785 3927
rect 16448 3896 17785 3924
rect 16448 3884 16454 3896
rect 17773 3893 17785 3896
rect 17819 3893 17831 3927
rect 17773 3887 17831 3893
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 20898 3924 20904 3936
rect 17920 3896 20904 3924
rect 17920 3884 17926 3896
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 21836 3924 21864 3955
rect 25148 3933 25176 4032
rect 21416 3896 21864 3924
rect 25133 3927 25191 3933
rect 21416 3884 21422 3896
rect 25133 3893 25145 3927
rect 25179 3924 25191 3927
rect 27614 3924 27620 3936
rect 25179 3896 27620 3924
rect 25179 3893 25191 3896
rect 25133 3887 25191 3893
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 5810 3680 5816 3732
rect 5868 3720 5874 3732
rect 8570 3720 8576 3732
rect 5868 3692 8576 3720
rect 5868 3680 5874 3692
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9582 3720 9588 3732
rect 9539 3692 9588 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 9582 3680 9588 3692
rect 9640 3720 9646 3732
rect 9950 3720 9956 3732
rect 9640 3692 9720 3720
rect 9911 3692 9956 3720
rect 9640 3680 9646 3692
rect 5261 3655 5319 3661
rect 5261 3621 5273 3655
rect 5307 3652 5319 3655
rect 7469 3655 7527 3661
rect 7469 3652 7481 3655
rect 5307 3624 7481 3652
rect 5307 3621 5319 3624
rect 5261 3615 5319 3621
rect 7469 3621 7481 3624
rect 7515 3652 7527 3655
rect 7742 3652 7748 3664
rect 7515 3624 7748 3652
rect 7515 3621 7527 3624
rect 7469 3615 7527 3621
rect 7742 3612 7748 3624
rect 7800 3612 7806 3664
rect 8389 3655 8447 3661
rect 8389 3621 8401 3655
rect 8435 3652 8447 3655
rect 8478 3652 8484 3664
rect 8435 3624 8484 3652
rect 8435 3621 8447 3624
rect 8389 3615 8447 3621
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 3694 3544 3700 3596
rect 3752 3584 3758 3596
rect 4513 3587 4571 3593
rect 4513 3584 4525 3587
rect 3752 3556 4525 3584
rect 3752 3544 3758 3556
rect 4513 3553 4525 3556
rect 4559 3553 4571 3587
rect 4513 3547 4571 3553
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3584 4859 3587
rect 5534 3584 5540 3596
rect 4847 3556 5540 3584
rect 4847 3553 4859 3556
rect 4801 3547 4859 3553
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 6178 3584 6184 3596
rect 6139 3556 6184 3584
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 6362 3544 6368 3596
rect 6420 3584 6426 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6420 3556 7113 3584
rect 6420 3544 6426 3556
rect 7101 3553 7113 3556
rect 7147 3584 7159 3587
rect 7190 3584 7196 3596
rect 7147 3556 7196 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 7653 3587 7711 3593
rect 7653 3553 7665 3587
rect 7699 3553 7711 3587
rect 7926 3584 7932 3596
rect 7887 3556 7932 3584
rect 7653 3547 7711 3553
rect 1578 3476 1584 3528
rect 1636 3516 1642 3528
rect 1636 3488 4154 3516
rect 1636 3476 1642 3488
rect 4126 3380 4154 3488
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 7668 3516 7696 3547
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 9692 3593 9720 3692
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 11330 3680 11336 3732
rect 11388 3720 11394 3732
rect 11425 3723 11483 3729
rect 11425 3720 11437 3723
rect 11388 3692 11437 3720
rect 11388 3680 11394 3692
rect 11425 3689 11437 3692
rect 11471 3689 11483 3723
rect 11425 3683 11483 3689
rect 11514 3680 11520 3732
rect 11572 3720 11578 3732
rect 12986 3720 12992 3732
rect 11572 3692 12664 3720
rect 12947 3692 12992 3720
rect 11572 3680 11578 3692
rect 10778 3652 10784 3664
rect 10428 3624 10784 3652
rect 10428 3593 10456 3624
rect 10778 3612 10784 3624
rect 10836 3612 10842 3664
rect 12084 3661 12112 3692
rect 12069 3655 12127 3661
rect 12069 3621 12081 3655
rect 12115 3621 12127 3655
rect 12069 3615 12127 3621
rect 12161 3655 12219 3661
rect 12161 3621 12173 3655
rect 12207 3652 12219 3655
rect 12342 3652 12348 3664
rect 12207 3624 12348 3652
rect 12207 3621 12219 3624
rect 12161 3615 12219 3621
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 12636 3652 12664 3692
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 14550 3720 14556 3732
rect 14511 3692 14556 3720
rect 14550 3680 14556 3692
rect 14608 3680 14614 3732
rect 18414 3720 18420 3732
rect 18375 3692 18420 3720
rect 18414 3680 18420 3692
rect 18472 3720 18478 3732
rect 20073 3723 20131 3729
rect 18472 3692 18736 3720
rect 18472 3680 18478 3692
rect 13262 3652 13268 3664
rect 12636 3624 13268 3652
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 13538 3652 13544 3664
rect 13499 3624 13544 3652
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 15651 3655 15709 3661
rect 15651 3621 15663 3655
rect 15697 3652 15709 3655
rect 15838 3652 15844 3664
rect 15697 3624 15844 3652
rect 15697 3621 15709 3624
rect 15651 3615 15709 3621
rect 15838 3612 15844 3624
rect 15896 3652 15902 3664
rect 16114 3652 16120 3664
rect 15896 3624 16120 3652
rect 15896 3612 15902 3624
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 16577 3655 16635 3661
rect 16577 3652 16589 3655
rect 16224 3624 16589 3652
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 10413 3587 10471 3593
rect 10413 3553 10425 3587
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3584 10563 3587
rect 10686 3584 10692 3596
rect 10551 3556 10692 3584
rect 10551 3553 10563 3556
rect 10505 3547 10563 3553
rect 8665 3519 8723 3525
rect 8665 3516 8677 3519
rect 7524 3488 8677 3516
rect 7524 3476 7530 3488
rect 8665 3485 8677 3488
rect 8711 3485 8723 3519
rect 8665 3479 8723 3485
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 10520 3516 10548 3547
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 11146 3584 11152 3596
rect 11103 3556 11152 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 9364 3488 10548 3516
rect 9364 3476 9370 3488
rect 4614 3448 4620 3460
rect 4575 3420 4620 3448
rect 4614 3408 4620 3420
rect 4672 3408 4678 3460
rect 6362 3448 6368 3460
rect 5368 3420 6368 3448
rect 5368 3380 5396 3420
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 7742 3448 7748 3460
rect 6564 3420 7748 3448
rect 6564 3392 6592 3420
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 8570 3408 8576 3460
rect 8628 3448 8634 3460
rect 10134 3448 10140 3460
rect 8628 3420 10140 3448
rect 8628 3408 8634 3420
rect 10134 3408 10140 3420
rect 10192 3448 10198 3460
rect 11072 3448 11100 3547
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 13630 3584 13636 3596
rect 13591 3556 13636 3584
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 16224 3593 16252 3624
rect 16577 3621 16589 3624
rect 16623 3652 16635 3655
rect 16758 3652 16764 3664
rect 16623 3624 16764 3652
rect 16623 3621 16635 3624
rect 16577 3615 16635 3621
rect 16758 3612 16764 3624
rect 16816 3652 16822 3664
rect 17218 3652 17224 3664
rect 16816 3624 17224 3652
rect 16816 3612 16822 3624
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 18708 3593 18736 3692
rect 20073 3689 20085 3723
rect 20119 3720 20131 3723
rect 20162 3720 20168 3732
rect 20119 3692 20168 3720
rect 20119 3689 20131 3692
rect 20073 3683 20131 3689
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20346 3680 20352 3732
rect 20404 3720 20410 3732
rect 21361 3723 21419 3729
rect 21361 3720 21373 3723
rect 20404 3692 21373 3720
rect 20404 3680 20410 3692
rect 21361 3689 21373 3692
rect 21407 3689 21419 3723
rect 21361 3683 21419 3689
rect 22646 3652 22652 3664
rect 21008 3624 22652 3652
rect 21008 3596 21036 3624
rect 22646 3612 22652 3624
rect 22704 3612 22710 3664
rect 16209 3587 16267 3593
rect 16209 3553 16221 3587
rect 16255 3553 16267 3587
rect 16209 3547 16267 3553
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3553 18751 3587
rect 20898 3584 20904 3596
rect 20859 3556 20904 3584
rect 18693 3547 18751 3553
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 20990 3544 20996 3596
rect 21048 3584 21054 3596
rect 21048 3556 21141 3584
rect 21048 3544 21054 3556
rect 21174 3544 21180 3596
rect 21232 3584 21238 3596
rect 22462 3584 22468 3596
rect 21232 3556 21277 3584
rect 22423 3556 22468 3584
rect 21232 3544 21238 3556
rect 22462 3544 22468 3556
rect 22520 3544 22526 3596
rect 23528 3587 23586 3593
rect 23528 3553 23540 3587
rect 23574 3584 23586 3587
rect 23842 3584 23848 3596
rect 23574 3556 23848 3584
rect 23574 3553 23586 3556
rect 23528 3547 23586 3553
rect 23842 3544 23848 3556
rect 23900 3544 23906 3596
rect 15289 3519 15347 3525
rect 15289 3485 15301 3519
rect 15335 3485 15347 3519
rect 17126 3516 17132 3528
rect 17087 3488 17132 3516
rect 15289 3479 15347 3485
rect 10192 3420 11100 3448
rect 10192 3408 10198 3420
rect 11698 3408 11704 3460
rect 11756 3448 11762 3460
rect 12621 3451 12679 3457
rect 12621 3448 12633 3451
rect 11756 3420 12633 3448
rect 11756 3408 11762 3420
rect 12621 3417 12633 3420
rect 12667 3448 12679 3451
rect 12802 3448 12808 3460
rect 12667 3420 12808 3448
rect 12667 3417 12679 3420
rect 12621 3411 12679 3417
rect 12802 3408 12808 3420
rect 12860 3408 12866 3460
rect 5534 3380 5540 3392
rect 4126 3352 5396 3380
rect 5495 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 6546 3380 6552 3392
rect 6507 3352 6552 3380
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 9122 3380 9128 3392
rect 9083 3352 9128 3380
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 11885 3383 11943 3389
rect 11885 3349 11897 3383
rect 11931 3380 11943 3383
rect 12158 3380 12164 3392
rect 11931 3352 12164 3380
rect 11931 3349 11943 3352
rect 11885 3343 11943 3349
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 13446 3380 13452 3392
rect 13407 3352 13452 3380
rect 13446 3340 13452 3352
rect 13504 3340 13510 3392
rect 15105 3383 15163 3389
rect 15105 3349 15117 3383
rect 15151 3380 15163 3383
rect 15304 3380 15332 3479
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 17402 3516 17408 3528
rect 17363 3488 17408 3516
rect 17402 3476 17408 3488
rect 17460 3516 17466 3528
rect 17770 3516 17776 3528
rect 17460 3488 17776 3516
rect 17460 3476 17466 3488
rect 17770 3476 17776 3488
rect 17828 3476 17834 3528
rect 18598 3516 18604 3528
rect 18559 3488 18604 3516
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 23615 3519 23673 3525
rect 23615 3516 23627 3519
rect 18892 3488 23627 3516
rect 16482 3408 16488 3460
rect 16540 3448 16546 3460
rect 16945 3451 17003 3457
rect 16945 3448 16957 3451
rect 16540 3420 16957 3448
rect 16540 3408 16546 3420
rect 16945 3417 16957 3420
rect 16991 3448 17003 3451
rect 18892 3448 18920 3488
rect 23615 3485 23627 3488
rect 23661 3485 23673 3519
rect 23615 3479 23673 3485
rect 16991 3420 18920 3448
rect 18984 3420 20944 3448
rect 16991 3417 17003 3420
rect 16945 3411 17003 3417
rect 15470 3380 15476 3392
rect 15151 3352 15476 3380
rect 15151 3349 15163 3352
rect 15105 3343 15163 3349
rect 15470 3340 15476 3352
rect 15528 3340 15534 3392
rect 18138 3380 18144 3392
rect 18099 3352 18144 3380
rect 18138 3340 18144 3352
rect 18196 3340 18202 3392
rect 18414 3340 18420 3392
rect 18472 3380 18478 3392
rect 18984 3380 19012 3420
rect 18472 3352 19012 3380
rect 19705 3383 19763 3389
rect 18472 3340 18478 3352
rect 19705 3349 19717 3383
rect 19751 3380 19763 3383
rect 20070 3380 20076 3392
rect 19751 3352 20076 3380
rect 19751 3349 19763 3352
rect 19705 3343 19763 3349
rect 20070 3340 20076 3352
rect 20128 3340 20134 3392
rect 20916 3380 20944 3420
rect 21266 3408 21272 3460
rect 21324 3448 21330 3460
rect 21913 3451 21971 3457
rect 21913 3448 21925 3451
rect 21324 3420 21925 3448
rect 21324 3408 21330 3420
rect 21913 3417 21925 3420
rect 21959 3417 21971 3451
rect 21913 3411 21971 3417
rect 22603 3383 22661 3389
rect 22603 3380 22615 3383
rect 20916 3352 22615 3380
rect 22603 3349 22615 3352
rect 22649 3349 22661 3383
rect 22603 3343 22661 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1535 3179 1593 3185
rect 1535 3145 1547 3179
rect 1581 3176 1593 3179
rect 1670 3176 1676 3188
rect 1581 3148 1676 3176
rect 1581 3145 1593 3148
rect 1535 3139 1593 3145
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 3694 3176 3700 3188
rect 3655 3148 3700 3176
rect 3694 3136 3700 3148
rect 3752 3176 3758 3188
rect 5258 3176 5264 3188
rect 3752 3148 5264 3176
rect 3752 3136 3758 3148
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 6546 3176 6552 3188
rect 6507 3148 6552 3176
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 12069 3179 12127 3185
rect 8536 3148 11002 3176
rect 8536 3136 8542 3148
rect 4295 3111 4353 3117
rect 4295 3077 4307 3111
rect 4341 3108 4353 3111
rect 9030 3108 9036 3120
rect 4341 3080 9036 3108
rect 4341 3077 4353 3080
rect 4295 3071 4353 3077
rect 9030 3068 9036 3080
rect 9088 3108 9094 3120
rect 10134 3108 10140 3120
rect 9088 3080 9168 3108
rect 10095 3080 10140 3108
rect 9088 3068 9094 3080
rect 106 3000 112 3052
rect 164 3040 170 3052
rect 5905 3043 5963 3049
rect 164 3012 1507 3040
rect 164 3000 170 3012
rect 1479 2981 1507 3012
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 7374 3040 7380 3052
rect 5951 3012 7380 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 7374 3000 7380 3012
rect 7432 3040 7438 3052
rect 7926 3040 7932 3052
rect 7432 3012 7932 3040
rect 7432 3000 7438 3012
rect 1464 2975 1522 2981
rect 1464 2941 1476 2975
rect 1510 2972 1522 2975
rect 1857 2975 1915 2981
rect 1857 2972 1869 2975
rect 1510 2944 1869 2972
rect 1510 2941 1522 2944
rect 1464 2935 1522 2941
rect 1857 2941 1869 2944
rect 1903 2941 1915 2975
rect 4062 2972 4068 2984
rect 3975 2944 4068 2972
rect 1857 2935 1915 2941
rect 4062 2932 4068 2944
rect 4120 2972 4126 2984
rect 4192 2975 4250 2981
rect 4192 2972 4204 2975
rect 4120 2944 4204 2972
rect 4120 2932 4126 2944
rect 4192 2941 4204 2944
rect 4238 2941 4250 2975
rect 4192 2935 4250 2941
rect 5077 2975 5135 2981
rect 5077 2941 5089 2975
rect 5123 2972 5135 2975
rect 5534 2972 5540 2984
rect 5123 2944 5540 2972
rect 5123 2941 5135 2944
rect 5077 2935 5135 2941
rect 5534 2932 5540 2944
rect 5592 2972 5598 2984
rect 5813 2975 5871 2981
rect 5813 2972 5825 2975
rect 5592 2944 5825 2972
rect 5592 2932 5598 2944
rect 5813 2941 5825 2944
rect 5859 2972 5871 2975
rect 5997 2975 6055 2981
rect 5997 2972 6009 2975
rect 5859 2944 6009 2972
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 5997 2941 6009 2944
rect 6043 2941 6055 2975
rect 7466 2972 7472 2984
rect 7427 2944 7472 2972
rect 5997 2935 6055 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 7760 2981 7788 3012
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 8202 3040 8208 3052
rect 8163 3012 8208 3040
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 9140 3049 9168 3080
rect 10134 3068 10140 3080
rect 10192 3068 10198 3120
rect 10505 3111 10563 3117
rect 10505 3077 10517 3111
rect 10551 3108 10563 3111
rect 10778 3108 10784 3120
rect 10551 3080 10784 3108
rect 10551 3077 10563 3080
rect 10505 3071 10563 3077
rect 10778 3068 10784 3080
rect 10836 3068 10842 3120
rect 10974 3108 11002 3148
rect 12069 3145 12081 3179
rect 12115 3176 12127 3179
rect 12342 3176 12348 3188
rect 12115 3148 12348 3176
rect 12115 3145 12127 3148
rect 12069 3139 12127 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 14274 3176 14280 3188
rect 12676 3148 14280 3176
rect 12676 3136 12682 3148
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 16298 3176 16304 3188
rect 16259 3148 16304 3176
rect 16298 3136 16304 3148
rect 16356 3176 16362 3188
rect 16574 3176 16580 3188
rect 16356 3148 16580 3176
rect 16356 3136 16362 3148
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17276 3148 17417 3176
rect 17276 3136 17282 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17405 3139 17463 3145
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 20898 3176 20904 3188
rect 17644 3148 19748 3176
rect 20859 3148 20904 3176
rect 17644 3136 17650 3148
rect 13541 3111 13599 3117
rect 13541 3108 13553 3111
rect 10974 3080 13553 3108
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3009 9183 3043
rect 9125 3003 9183 3009
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3040 10655 3043
rect 11330 3040 11336 3052
rect 10643 3012 11336 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 11330 3000 11336 3012
rect 11388 3000 11394 3052
rect 12526 3040 12532 3052
rect 12176 3012 12532 3040
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2972 7803 2975
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 7791 2944 8493 2972
rect 7791 2941 7803 2944
rect 7745 2935 7803 2941
rect 8481 2941 8493 2944
rect 8527 2941 8539 2975
rect 8481 2935 8539 2941
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2972 9827 2975
rect 12176 2972 12204 3012
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12802 3040 12808 3052
rect 12763 3012 12808 3040
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 9815 2944 12204 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 6178 2904 6184 2916
rect 4632 2876 6184 2904
rect 4632 2848 4660 2876
rect 6178 2864 6184 2876
rect 6236 2904 6242 2916
rect 7285 2907 7343 2913
rect 7285 2904 7297 2907
rect 6236 2876 7297 2904
rect 6236 2864 6242 2876
rect 7285 2873 7297 2876
rect 7331 2904 7343 2907
rect 7576 2904 7604 2935
rect 7331 2876 7604 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 9122 2864 9128 2916
rect 9180 2904 9186 2916
rect 9217 2907 9275 2913
rect 9217 2904 9229 2907
rect 9180 2876 9229 2904
rect 9180 2864 9186 2876
rect 9217 2873 9229 2876
rect 9263 2904 9275 2907
rect 10778 2904 10784 2916
rect 9263 2876 10784 2904
rect 9263 2873 9275 2876
rect 9217 2867 9275 2873
rect 10778 2864 10784 2876
rect 10836 2864 10842 2916
rect 12621 2907 12679 2913
rect 12621 2873 12633 2907
rect 12667 2904 12679 2907
rect 12986 2904 12992 2916
rect 12667 2876 12992 2904
rect 12667 2873 12679 2876
rect 12621 2867 12679 2873
rect 4614 2836 4620 2848
rect 4575 2808 4620 2836
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 5997 2839 6055 2845
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 7926 2836 7932 2848
rect 6043 2808 7932 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 8849 2839 8907 2845
rect 8849 2836 8861 2839
rect 8812 2808 8861 2836
rect 8812 2796 8818 2808
rect 8849 2805 8861 2808
rect 8895 2805 8907 2839
rect 10962 2836 10968 2848
rect 10923 2808 10968 2836
rect 8849 2799 8907 2805
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 12636 2836 12664 2867
rect 12986 2864 12992 2876
rect 13044 2864 13050 2916
rect 13372 2904 13400 3080
rect 13541 3077 13553 3080
rect 13587 3077 13599 3111
rect 15470 3108 15476 3120
rect 15431 3080 15476 3108
rect 13541 3071 13599 3077
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 18506 3108 18512 3120
rect 16500 3080 18512 3108
rect 13446 3000 13452 3052
rect 13504 3040 13510 3052
rect 16500 3049 16528 3080
rect 16485 3043 16543 3049
rect 16485 3040 16497 3043
rect 13504 3012 16497 3040
rect 13504 3000 13510 3012
rect 16485 3009 16497 3012
rect 16531 3009 16543 3043
rect 16485 3003 16543 3009
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3040 17187 3043
rect 17402 3040 17408 3052
rect 17175 3012 17408 3040
rect 17175 3009 17187 3012
rect 17129 3003 17187 3009
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 18138 3040 18144 3052
rect 18099 3012 18144 3040
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 18432 3049 18460 3080
rect 18506 3068 18512 3080
rect 18564 3068 18570 3120
rect 19720 3117 19748 3148
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 23750 3136 23756 3188
rect 23808 3176 23814 3188
rect 24719 3179 24777 3185
rect 24719 3176 24731 3179
rect 23808 3148 24731 3176
rect 23808 3136 23814 3148
rect 24719 3145 24731 3148
rect 24765 3145 24777 3179
rect 24719 3139 24777 3145
rect 19705 3111 19763 3117
rect 19705 3077 19717 3111
rect 19751 3108 19763 3111
rect 19978 3108 19984 3120
rect 19751 3080 19984 3108
rect 19751 3077 19763 3080
rect 19705 3071 19763 3077
rect 19978 3068 19984 3080
rect 20036 3108 20042 3120
rect 20990 3108 20996 3120
rect 20036 3080 20996 3108
rect 20036 3068 20042 3080
rect 20990 3068 20996 3080
rect 21048 3068 21054 3120
rect 21266 3108 21272 3120
rect 21227 3080 21272 3108
rect 21266 3068 21272 3080
rect 21324 3068 21330 3120
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 20070 3040 20076 3052
rect 19484 3012 19932 3040
rect 20031 3012 20076 3040
rect 19484 3000 19490 3012
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2972 14059 2975
rect 14090 2972 14096 2984
rect 14047 2944 14096 2972
rect 14047 2941 14059 2944
rect 14001 2935 14059 2941
rect 14090 2932 14096 2944
rect 14148 2932 14154 2984
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 14332 2944 14565 2972
rect 14332 2932 14338 2944
rect 14553 2941 14565 2944
rect 14599 2941 14611 2975
rect 14553 2935 14611 2941
rect 14921 2975 14979 2981
rect 14921 2941 14933 2975
rect 14967 2941 14979 2975
rect 14921 2935 14979 2941
rect 15473 2975 15531 2981
rect 15473 2941 15485 2975
rect 15519 2941 15531 2975
rect 15473 2935 15531 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2972 19211 2975
rect 19610 2972 19616 2984
rect 19199 2944 19616 2972
rect 19199 2941 19211 2944
rect 19153 2935 19211 2941
rect 14826 2904 14832 2916
rect 13372 2876 14832 2904
rect 14826 2864 14832 2876
rect 14884 2904 14890 2916
rect 14936 2904 14964 2935
rect 14884 2876 14964 2904
rect 14884 2864 14890 2876
rect 15010 2864 15016 2916
rect 15068 2904 15074 2916
rect 15488 2904 15516 2935
rect 16482 2904 16488 2916
rect 15068 2876 16488 2904
rect 15068 2864 15074 2876
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 17865 2907 17923 2913
rect 16632 2876 16677 2904
rect 16632 2864 16638 2876
rect 17865 2873 17877 2907
rect 17911 2904 17923 2907
rect 18233 2907 18291 2913
rect 18233 2904 18245 2907
rect 17911 2876 18245 2904
rect 17911 2873 17923 2876
rect 17865 2867 17923 2873
rect 18233 2873 18245 2876
rect 18279 2904 18291 2907
rect 18598 2904 18604 2916
rect 18279 2876 18604 2904
rect 18279 2873 18291 2876
rect 18233 2867 18291 2873
rect 18598 2864 18604 2876
rect 18656 2864 18662 2916
rect 11563 2808 12664 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 15028 2836 15056 2864
rect 15838 2836 15844 2848
rect 13964 2808 15056 2836
rect 15799 2808 15844 2836
rect 13964 2796 13970 2808
rect 15838 2796 15844 2808
rect 15896 2796 15902 2848
rect 16666 2796 16672 2848
rect 16724 2836 16730 2848
rect 19168 2836 19196 2935
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 19904 2981 19932 3012
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 21082 3000 21088 3052
rect 21140 3040 21146 3052
rect 21637 3043 21695 3049
rect 21637 3040 21649 3043
rect 21140 3012 21649 3040
rect 21140 3000 21146 3012
rect 21637 3009 21649 3012
rect 21683 3009 21695 3043
rect 21637 3003 21695 3009
rect 19889 2975 19947 2981
rect 19889 2941 19901 2975
rect 19935 2972 19947 2975
rect 20806 2972 20812 2984
rect 19935 2944 20812 2972
rect 19935 2941 19947 2944
rect 19889 2935 19947 2941
rect 20806 2932 20812 2944
rect 20864 2932 20870 2984
rect 20898 2932 20904 2984
rect 20956 2972 20962 2984
rect 21177 2975 21235 2981
rect 21177 2972 21189 2975
rect 20956 2944 21189 2972
rect 20956 2932 20962 2944
rect 21177 2941 21189 2944
rect 21223 2941 21235 2975
rect 21177 2935 21235 2941
rect 21266 2932 21272 2984
rect 21324 2972 21330 2984
rect 21453 2975 21511 2981
rect 21453 2972 21465 2975
rect 21324 2944 21465 2972
rect 21324 2932 21330 2944
rect 21453 2941 21465 2944
rect 21499 2972 21511 2975
rect 22189 2975 22247 2981
rect 22189 2972 22201 2975
rect 21499 2944 22201 2972
rect 21499 2941 21511 2944
rect 21453 2935 21511 2941
rect 22189 2941 22201 2944
rect 22235 2941 22247 2975
rect 22189 2935 22247 2941
rect 24648 2975 24706 2981
rect 24648 2941 24660 2975
rect 24694 2972 24706 2975
rect 24694 2944 25176 2972
rect 24694 2941 24706 2944
rect 24648 2935 24706 2941
rect 22462 2904 22468 2916
rect 20133 2876 22468 2904
rect 19426 2836 19432 2848
rect 16724 2808 19196 2836
rect 19387 2808 19432 2836
rect 16724 2796 16730 2808
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 19518 2796 19524 2848
rect 19576 2836 19582 2848
rect 20133 2836 20161 2876
rect 22462 2864 22468 2876
rect 22520 2904 22526 2916
rect 22925 2907 22983 2913
rect 22925 2904 22937 2907
rect 22520 2876 22937 2904
rect 22520 2864 22526 2876
rect 22925 2873 22937 2876
rect 22971 2873 22983 2907
rect 22925 2867 22983 2873
rect 22646 2836 22652 2848
rect 19576 2808 20161 2836
rect 22607 2808 22652 2836
rect 19576 2796 19582 2808
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 23842 2836 23848 2848
rect 23803 2808 23848 2836
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 25148 2845 25176 2944
rect 25133 2839 25191 2845
rect 25133 2805 25145 2839
rect 25179 2836 25191 2839
rect 26878 2836 26884 2848
rect 25179 2808 26884 2836
rect 25179 2805 25191 2808
rect 25133 2799 25191 2805
rect 26878 2796 26884 2808
rect 26936 2796 26942 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 3881 2635 3939 2641
rect 3881 2601 3893 2635
rect 3927 2632 3939 2635
rect 4338 2632 4344 2644
rect 3927 2604 4344 2632
rect 3927 2601 3939 2604
rect 3881 2595 3939 2601
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 4430 2592 4436 2644
rect 4488 2632 4494 2644
rect 4525 2635 4583 2641
rect 4525 2632 4537 2635
rect 4488 2604 4537 2632
rect 4488 2592 4494 2604
rect 4525 2601 4537 2604
rect 4571 2601 4583 2635
rect 5350 2632 5356 2644
rect 4525 2595 4583 2601
rect 4724 2604 5356 2632
rect 3513 2567 3571 2573
rect 3513 2564 3525 2567
rect 3043 2536 3525 2564
rect 3043 2505 3071 2536
rect 3513 2533 3525 2536
rect 3559 2564 3571 2567
rect 4724 2564 4752 2604
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 7101 2635 7159 2641
rect 7101 2601 7113 2635
rect 7147 2632 7159 2635
rect 13354 2632 13360 2644
rect 7147 2604 13360 2632
rect 7147 2601 7159 2604
rect 7101 2595 7159 2601
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 13630 2632 13636 2644
rect 13591 2604 13636 2632
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 14461 2635 14519 2641
rect 14461 2632 14473 2635
rect 13786 2604 14473 2632
rect 3559 2536 4752 2564
rect 4801 2567 4859 2573
rect 3559 2533 3571 2536
rect 3513 2527 3571 2533
rect 4801 2533 4813 2567
rect 4847 2564 4859 2567
rect 6638 2564 6644 2576
rect 4847 2536 6644 2564
rect 4847 2533 4859 2536
rect 4801 2527 4859 2533
rect 3028 2499 3086 2505
rect 3028 2465 3040 2499
rect 3074 2465 3086 2499
rect 3028 2459 3086 2465
rect 4316 2499 4374 2505
rect 4316 2465 4328 2499
rect 4362 2496 4374 2499
rect 4816 2496 4844 2527
rect 6638 2524 6644 2536
rect 6696 2524 6702 2576
rect 7374 2524 7380 2576
rect 7432 2564 7438 2576
rect 7469 2567 7527 2573
rect 7469 2564 7481 2567
rect 7432 2536 7481 2564
rect 7432 2524 7438 2536
rect 7469 2533 7481 2536
rect 7515 2533 7527 2567
rect 7926 2564 7932 2576
rect 7839 2536 7932 2564
rect 7469 2527 7527 2533
rect 7926 2524 7932 2536
rect 7984 2564 7990 2576
rect 8754 2564 8760 2576
rect 7984 2536 8340 2564
rect 8715 2536 8760 2564
rect 7984 2524 7990 2536
rect 8312 2508 8340 2536
rect 8754 2524 8760 2536
rect 8812 2524 8818 2576
rect 10182 2567 10240 2573
rect 10182 2564 10194 2567
rect 9508 2536 10194 2564
rect 4362 2468 4844 2496
rect 5169 2499 5227 2505
rect 4362 2465 4374 2468
rect 4316 2459 4374 2465
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5353 2499 5411 2505
rect 5353 2496 5365 2499
rect 5215 2468 5365 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5353 2465 5365 2468
rect 5399 2465 5411 2499
rect 6914 2496 6920 2508
rect 6875 2468 6920 2496
rect 5353 2459 5411 2465
rect 3099 2363 3157 2369
rect 3099 2329 3111 2363
rect 3145 2360 3157 2363
rect 3234 2360 3240 2372
rect 3145 2332 3240 2360
rect 3145 2329 3157 2332
rect 3099 2323 3157 2329
rect 3234 2320 3240 2332
rect 3292 2320 3298 2372
rect 5184 2360 5212 2459
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 7484 2468 8033 2496
rect 7484 2440 7512 2468
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 8294 2496 8300 2508
rect 8255 2468 8300 2496
rect 8021 2459 8079 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 6273 2431 6331 2437
rect 6273 2428 6285 2431
rect 5316 2400 6285 2428
rect 5316 2388 5322 2400
rect 6273 2397 6285 2400
rect 6319 2428 6331 2431
rect 6641 2431 6699 2437
rect 6641 2428 6653 2431
rect 6319 2400 6653 2428
rect 6319 2397 6331 2400
rect 6273 2391 6331 2397
rect 6641 2397 6653 2400
rect 6687 2428 6699 2431
rect 7466 2428 7472 2440
rect 6687 2400 7472 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7800 2400 8125 2428
rect 7800 2388 7806 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 4126 2332 5212 2360
rect 8128 2360 8156 2391
rect 9033 2363 9091 2369
rect 9033 2360 9045 2363
rect 8128 2332 9045 2360
rect 842 2252 848 2304
rect 900 2292 906 2304
rect 4126 2292 4154 2332
rect 9033 2329 9045 2332
rect 9079 2329 9091 2363
rect 9033 2323 9091 2329
rect 900 2264 4154 2292
rect 900 2252 906 2264
rect 7190 2252 7196 2304
rect 7248 2292 7254 2304
rect 9508 2301 9536 2536
rect 10182 2533 10194 2536
rect 10228 2564 10240 2567
rect 10962 2564 10968 2576
rect 10228 2536 10968 2564
rect 10228 2533 10240 2536
rect 10182 2527 10240 2533
rect 10962 2524 10968 2536
rect 11020 2564 11026 2576
rect 11057 2567 11115 2573
rect 11057 2564 11069 2567
rect 11020 2536 11069 2564
rect 11020 2524 11026 2536
rect 11057 2533 11069 2536
rect 11103 2533 11115 2567
rect 12713 2567 12771 2573
rect 12713 2564 12725 2567
rect 11057 2527 11115 2533
rect 11992 2536 12725 2564
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 9950 2496 9956 2508
rect 9907 2468 9956 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 9950 2456 9956 2468
rect 10008 2496 10014 2508
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 10008 2468 11437 2496
rect 10008 2456 10014 2468
rect 11425 2465 11437 2468
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 9766 2388 9772 2440
rect 9824 2428 9830 2440
rect 11992 2437 12020 2536
rect 12713 2533 12725 2536
rect 12759 2533 12771 2567
rect 12713 2527 12771 2533
rect 12802 2524 12808 2576
rect 12860 2564 12866 2576
rect 13786 2564 13814 2604
rect 14461 2601 14473 2604
rect 14507 2601 14519 2635
rect 14461 2595 14519 2601
rect 14921 2635 14979 2641
rect 14921 2601 14933 2635
rect 14967 2632 14979 2635
rect 15010 2632 15016 2644
rect 14967 2604 15016 2632
rect 14967 2601 14979 2604
rect 14921 2595 14979 2601
rect 15010 2592 15016 2604
rect 15068 2592 15074 2644
rect 16390 2632 16396 2644
rect 16351 2604 16396 2632
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 17221 2635 17279 2641
rect 17221 2601 17233 2635
rect 17267 2632 17279 2635
rect 18138 2632 18144 2644
rect 17267 2604 18144 2632
rect 17267 2601 17279 2604
rect 17221 2595 17279 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 19978 2632 19984 2644
rect 19751 2604 19984 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20530 2632 20536 2644
rect 20491 2604 20536 2632
rect 20530 2592 20536 2604
rect 20588 2592 20594 2644
rect 20898 2592 20904 2644
rect 20956 2632 20962 2644
rect 21361 2635 21419 2641
rect 21361 2632 21373 2635
rect 20956 2604 21373 2632
rect 20956 2592 20962 2604
rect 21361 2601 21373 2604
rect 21407 2601 21419 2635
rect 21361 2595 21419 2601
rect 14182 2564 14188 2576
rect 12860 2536 12905 2564
rect 13372 2536 13814 2564
rect 14143 2536 14188 2564
rect 12860 2524 12866 2536
rect 12434 2496 12440 2508
rect 12395 2468 12440 2496
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 9824 2400 11989 2428
rect 9824 2388 9830 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 12452 2428 12480 2456
rect 12802 2428 12808 2440
rect 12452 2400 12808 2428
rect 11977 2391 12035 2397
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 13372 2428 13400 2536
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 15838 2573 15844 2576
rect 15794 2567 15844 2573
rect 15794 2564 15806 2567
rect 15212 2536 15806 2564
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14277 2499 14335 2505
rect 14277 2496 14289 2499
rect 13872 2468 14289 2496
rect 13872 2456 13878 2468
rect 14277 2465 14289 2468
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 12912 2400 13400 2428
rect 10781 2363 10839 2369
rect 10781 2329 10793 2363
rect 10827 2360 10839 2363
rect 10870 2360 10876 2372
rect 10827 2332 10876 2360
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 10870 2320 10876 2332
rect 10928 2320 10934 2372
rect 10962 2320 10968 2372
rect 11020 2360 11026 2372
rect 12912 2360 12940 2400
rect 13262 2360 13268 2372
rect 11020 2332 12940 2360
rect 13223 2332 13268 2360
rect 11020 2320 11026 2332
rect 13262 2320 13268 2332
rect 13320 2320 13326 2372
rect 15212 2369 15240 2536
rect 15794 2533 15806 2536
rect 15840 2533 15844 2567
rect 15794 2527 15844 2533
rect 15838 2524 15844 2527
rect 15896 2524 15902 2576
rect 18049 2567 18107 2573
rect 18049 2533 18061 2567
rect 18095 2564 18107 2567
rect 18509 2567 18567 2573
rect 18509 2564 18521 2567
rect 18095 2536 18521 2564
rect 18095 2533 18107 2536
rect 18049 2527 18107 2533
rect 18509 2533 18521 2536
rect 18555 2564 18567 2567
rect 18598 2564 18604 2576
rect 18555 2536 18604 2564
rect 18555 2533 18567 2536
rect 18509 2527 18567 2533
rect 18598 2524 18604 2536
rect 18656 2524 18662 2576
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 15562 2496 15568 2508
rect 15519 2468 15568 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 15562 2456 15568 2468
rect 15620 2496 15626 2508
rect 16669 2499 16727 2505
rect 16669 2496 16681 2499
rect 15620 2468 16681 2496
rect 15620 2456 15626 2468
rect 16669 2465 16681 2468
rect 16715 2465 16727 2499
rect 16669 2459 16727 2465
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2496 17831 2499
rect 19889 2499 19947 2505
rect 17819 2468 18276 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 17126 2428 17132 2440
rect 17039 2400 17132 2428
rect 17126 2388 17132 2400
rect 17184 2428 17190 2440
rect 17865 2431 17923 2437
rect 17865 2428 17877 2431
rect 17184 2400 17877 2428
rect 17184 2388 17190 2400
rect 17865 2397 17877 2400
rect 17911 2397 17923 2431
rect 18248 2428 18276 2468
rect 19889 2465 19901 2499
rect 19935 2496 19947 2499
rect 20548 2496 20576 2592
rect 22554 2524 22560 2576
rect 22612 2564 22618 2576
rect 22612 2536 24624 2564
rect 22612 2524 22618 2536
rect 19935 2468 20576 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20806 2456 20812 2508
rect 20864 2496 20870 2508
rect 20901 2499 20959 2505
rect 20901 2496 20913 2499
rect 20864 2468 20913 2496
rect 20864 2456 20870 2468
rect 20901 2465 20913 2468
rect 20947 2496 20959 2499
rect 21174 2496 21180 2508
rect 20947 2468 21180 2496
rect 20947 2465 20959 2468
rect 20901 2459 20959 2465
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 21637 2499 21695 2505
rect 21637 2465 21649 2499
rect 21683 2496 21695 2499
rect 21726 2496 21732 2508
rect 21683 2468 21732 2496
rect 21683 2465 21695 2468
rect 21637 2459 21695 2465
rect 21726 2456 21732 2468
rect 21784 2496 21790 2508
rect 22189 2499 22247 2505
rect 22189 2496 22201 2499
rect 21784 2468 22201 2496
rect 21784 2456 21790 2468
rect 22189 2465 22201 2468
rect 22235 2465 22247 2499
rect 22189 2459 22247 2465
rect 22370 2456 22376 2508
rect 22428 2496 22434 2508
rect 24596 2505 24624 2536
rect 22776 2499 22834 2505
rect 22776 2496 22788 2499
rect 22428 2468 22788 2496
rect 22428 2456 22434 2468
rect 22776 2465 22788 2468
rect 22822 2496 22834 2499
rect 23201 2499 23259 2505
rect 23201 2496 23213 2499
rect 22822 2468 23213 2496
rect 22822 2465 22834 2468
rect 22776 2459 22834 2465
rect 23201 2465 23213 2468
rect 23247 2465 23259 2499
rect 23201 2459 23259 2465
rect 24581 2499 24639 2505
rect 24581 2465 24593 2499
rect 24627 2496 24639 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24627 2468 25145 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 18414 2428 18420 2440
rect 18248 2400 18420 2428
rect 17865 2391 17923 2397
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 18524 2400 19656 2428
rect 15197 2363 15255 2369
rect 15197 2329 15209 2363
rect 15243 2329 15255 2363
rect 15197 2323 15255 2329
rect 16022 2320 16028 2372
rect 16080 2360 16086 2372
rect 18524 2360 18552 2400
rect 18969 2363 19027 2369
rect 18969 2360 18981 2363
rect 16080 2332 18552 2360
rect 18708 2332 18981 2360
rect 16080 2320 16086 2332
rect 9493 2295 9551 2301
rect 9493 2292 9505 2295
rect 7248 2264 9505 2292
rect 7248 2252 7254 2264
rect 9493 2261 9505 2264
rect 9539 2261 9551 2295
rect 9493 2255 9551 2261
rect 17865 2295 17923 2301
rect 17865 2261 17877 2295
rect 17911 2292 17923 2295
rect 18708 2292 18736 2332
rect 18969 2329 18981 2332
rect 19015 2329 19027 2363
rect 19628 2360 19656 2400
rect 20073 2363 20131 2369
rect 20073 2360 20085 2363
rect 19628 2332 20085 2360
rect 18969 2323 19027 2329
rect 20073 2329 20085 2332
rect 20119 2329 20131 2363
rect 20073 2323 20131 2329
rect 21821 2363 21879 2369
rect 21821 2329 21833 2363
rect 21867 2360 21879 2363
rect 23014 2360 23020 2372
rect 21867 2332 23020 2360
rect 21867 2329 21879 2332
rect 21821 2323 21879 2329
rect 23014 2320 23020 2332
rect 23072 2320 23078 2372
rect 24765 2363 24823 2369
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 26050 2360 26056 2372
rect 24811 2332 26056 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 26050 2320 26056 2332
rect 26108 2320 26114 2372
rect 17911 2264 18736 2292
rect 17911 2261 17923 2264
rect 17865 2255 17923 2261
rect 21450 2252 21456 2304
rect 21508 2292 21514 2304
rect 22879 2295 22937 2301
rect 22879 2292 22891 2295
rect 21508 2264 22891 2292
rect 21508 2252 21514 2264
rect 22879 2261 22891 2264
rect 22925 2261 22937 2295
rect 22879 2255 22937 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 8300 27480 8352 27532
rect 9588 27480 9640 27532
rect 11060 27480 11112 27532
rect 11704 27480 11756 27532
rect 15752 27480 15804 27532
rect 18236 27480 18288 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 22836 24259 22888 24268
rect 22836 24225 22854 24259
rect 22854 24225 22888 24259
rect 22836 24216 22888 24225
rect 24676 24216 24728 24268
rect 21088 24012 21140 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 7472 23808 7524 23860
rect 22468 23808 22520 23860
rect 22836 23851 22888 23860
rect 22836 23817 22845 23851
rect 22845 23817 22879 23851
rect 22879 23817 22888 23851
rect 22836 23808 22888 23817
rect 24216 23851 24268 23860
rect 24216 23817 24225 23851
rect 24225 23817 24259 23851
rect 24259 23817 24268 23851
rect 24216 23808 24268 23817
rect 22744 23740 22796 23792
rect 6920 23604 6972 23656
rect 9588 23647 9640 23656
rect 9588 23613 9597 23647
rect 9597 23613 9631 23647
rect 9631 23613 9640 23647
rect 9588 23604 9640 23613
rect 10876 23647 10928 23656
rect 10876 23613 10885 23647
rect 10885 23613 10919 23647
rect 10919 23613 10928 23647
rect 10876 23604 10928 23613
rect 21548 23604 21600 23656
rect 24216 23604 24268 23656
rect 26792 23808 26844 23860
rect 22468 23536 22520 23588
rect 9404 23468 9456 23520
rect 10048 23468 10100 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5264 23264 5316 23316
rect 10048 23264 10100 23316
rect 10876 23264 10928 23316
rect 22836 23171 22888 23180
rect 22836 23137 22854 23171
rect 22854 23137 22888 23171
rect 22836 23128 22888 23137
rect 23204 23128 23256 23180
rect 10784 22967 10836 22976
rect 10784 22933 10793 22967
rect 10793 22933 10827 22967
rect 10827 22933 10836 22967
rect 10784 22924 10836 22933
rect 22100 22924 22152 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 22836 22763 22888 22772
rect 22836 22729 22845 22763
rect 22845 22729 22879 22763
rect 22879 22729 22888 22763
rect 22836 22720 22888 22729
rect 25136 22763 25188 22772
rect 25136 22729 25145 22763
rect 25145 22729 25179 22763
rect 25179 22729 25188 22763
rect 25136 22720 25188 22729
rect 1400 22559 1452 22568
rect 1400 22525 1409 22559
rect 1409 22525 1443 22559
rect 1443 22525 1452 22559
rect 1400 22516 1452 22525
rect 25136 22516 25188 22568
rect 18880 22448 18932 22500
rect 20 22380 72 22432
rect 10784 22380 10836 22432
rect 11612 22380 11664 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 2136 21292 2188 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 19984 21088 20036 21140
rect 19616 20995 19668 21004
rect 19616 20961 19625 20995
rect 19625 20961 19659 20995
rect 19659 20961 19668 20995
rect 19616 20952 19668 20961
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 19616 20519 19668 20528
rect 19616 20485 19625 20519
rect 19625 20485 19659 20519
rect 19659 20485 19668 20519
rect 19616 20476 19668 20485
rect 18420 20340 18472 20392
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 12256 19864 12308 19916
rect 13912 19864 13964 19916
rect 14556 19864 14608 19916
rect 13728 19796 13780 19848
rect 13636 19660 13688 19712
rect 15568 19660 15620 19712
rect 16488 19660 16540 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 12256 19499 12308 19508
rect 12256 19465 12265 19499
rect 12265 19465 12299 19499
rect 12299 19465 12308 19499
rect 12256 19456 12308 19465
rect 13636 19456 13688 19508
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 12900 19252 12952 19304
rect 16488 19295 16540 19304
rect 13452 19227 13504 19236
rect 13452 19193 13461 19227
rect 13461 19193 13495 19227
rect 13495 19193 13504 19227
rect 13452 19184 13504 19193
rect 15476 19184 15528 19236
rect 16488 19261 16497 19295
rect 16497 19261 16531 19295
rect 16531 19261 16540 19295
rect 16488 19252 16540 19261
rect 19064 19252 19116 19304
rect 16672 19227 16724 19236
rect 16672 19193 16681 19227
rect 16681 19193 16715 19227
rect 16715 19193 16724 19227
rect 16672 19184 16724 19193
rect 2412 19116 2464 19168
rect 14556 19116 14608 19168
rect 15660 19116 15712 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 9956 18955 10008 18964
rect 9956 18921 9965 18955
rect 9965 18921 9999 18955
rect 9999 18921 10008 18955
rect 9956 18912 10008 18921
rect 12808 18955 12860 18964
rect 12808 18921 12817 18955
rect 12817 18921 12851 18955
rect 12851 18921 12860 18955
rect 12808 18912 12860 18921
rect 10876 18844 10928 18896
rect 13636 18912 13688 18964
rect 13728 18912 13780 18964
rect 14280 18912 14332 18964
rect 13452 18844 13504 18896
rect 17224 18912 17276 18964
rect 21088 18912 21140 18964
rect 21548 18912 21600 18964
rect 24768 18955 24820 18964
rect 24768 18921 24777 18955
rect 24777 18921 24811 18955
rect 24811 18921 24820 18955
rect 24768 18912 24820 18921
rect 17132 18887 17184 18896
rect 17132 18853 17141 18887
rect 17141 18853 17175 18887
rect 17175 18853 17184 18887
rect 17132 18844 17184 18853
rect 1492 18776 1544 18828
rect 7932 18776 7984 18828
rect 8300 18776 8352 18828
rect 9864 18776 9916 18828
rect 15384 18819 15436 18828
rect 15384 18785 15393 18819
rect 15393 18785 15427 18819
rect 15427 18785 15436 18819
rect 15384 18776 15436 18785
rect 15844 18819 15896 18828
rect 15844 18785 15853 18819
rect 15853 18785 15887 18819
rect 15887 18785 15896 18819
rect 15844 18776 15896 18785
rect 21732 18776 21784 18828
rect 24676 18776 24728 18828
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 11980 18751 12032 18760
rect 11980 18717 11989 18751
rect 11989 18717 12023 18751
rect 12023 18717 12032 18751
rect 11980 18708 12032 18717
rect 13728 18751 13780 18760
rect 13728 18717 13737 18751
rect 13737 18717 13771 18751
rect 13771 18717 13780 18751
rect 13728 18708 13780 18717
rect 17408 18708 17460 18760
rect 17776 18708 17828 18760
rect 8024 18683 8076 18692
rect 8024 18649 8033 18683
rect 8033 18649 8067 18683
rect 8067 18649 8076 18683
rect 8024 18640 8076 18649
rect 16212 18640 16264 18692
rect 8300 18572 8352 18624
rect 16396 18615 16448 18624
rect 16396 18581 16405 18615
rect 16405 18581 16439 18615
rect 16439 18581 16448 18615
rect 16396 18572 16448 18581
rect 18052 18615 18104 18624
rect 18052 18581 18061 18615
rect 18061 18581 18095 18615
rect 18095 18581 18104 18615
rect 18052 18572 18104 18581
rect 21916 18615 21968 18624
rect 21916 18581 21925 18615
rect 21925 18581 21959 18615
rect 21959 18581 21968 18615
rect 21916 18572 21968 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1492 18368 1544 18420
rect 7932 18411 7984 18420
rect 7932 18377 7941 18411
rect 7941 18377 7975 18411
rect 7975 18377 7984 18411
rect 7932 18368 7984 18377
rect 1860 18232 1912 18284
rect 8944 18232 8996 18284
rect 12900 18368 12952 18420
rect 13452 18368 13504 18420
rect 14280 18275 14332 18284
rect 14280 18241 14289 18275
rect 14289 18241 14323 18275
rect 14323 18241 14332 18275
rect 14280 18232 14332 18241
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 16212 18275 16264 18284
rect 16212 18241 16221 18275
rect 16221 18241 16255 18275
rect 16255 18241 16264 18275
rect 16212 18232 16264 18241
rect 20812 18232 20864 18284
rect 24676 18232 24728 18284
rect 2412 18028 2464 18080
rect 9864 18028 9916 18080
rect 12716 18139 12768 18148
rect 12716 18105 12725 18139
rect 12725 18105 12759 18139
rect 12759 18105 12768 18139
rect 12716 18096 12768 18105
rect 12808 18139 12860 18148
rect 12808 18105 12817 18139
rect 12817 18105 12851 18139
rect 12851 18105 12860 18139
rect 12808 18096 12860 18105
rect 13728 18096 13780 18148
rect 14372 18139 14424 18148
rect 14372 18105 14381 18139
rect 14381 18105 14415 18139
rect 14415 18105 14424 18139
rect 14372 18096 14424 18105
rect 16396 18096 16448 18148
rect 16856 18139 16908 18148
rect 16856 18105 16865 18139
rect 16865 18105 16899 18139
rect 16899 18105 16908 18139
rect 16856 18096 16908 18105
rect 18144 18164 18196 18216
rect 18788 18096 18840 18148
rect 21732 18096 21784 18148
rect 21916 18139 21968 18148
rect 21916 18105 21925 18139
rect 21925 18105 21959 18139
rect 21959 18105 21968 18139
rect 21916 18096 21968 18105
rect 10784 18028 10836 18080
rect 10876 18028 10928 18080
rect 15384 18071 15436 18080
rect 15384 18037 15393 18071
rect 15393 18037 15427 18071
rect 15427 18037 15436 18071
rect 15384 18028 15436 18037
rect 15844 18071 15896 18080
rect 15844 18037 15853 18071
rect 15853 18037 15887 18071
rect 15887 18037 15896 18071
rect 15844 18028 15896 18037
rect 17040 18028 17092 18080
rect 17960 18028 18012 18080
rect 22192 18096 22244 18148
rect 24952 18096 25004 18148
rect 22928 18028 22980 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 12164 17867 12216 17876
rect 12164 17833 12173 17867
rect 12173 17833 12207 17867
rect 12207 17833 12216 17867
rect 12164 17824 12216 17833
rect 12808 17824 12860 17876
rect 15660 17824 15712 17876
rect 17224 17867 17276 17876
rect 17224 17833 17233 17867
rect 17233 17833 17267 17867
rect 17267 17833 17276 17867
rect 17224 17824 17276 17833
rect 22100 17867 22152 17876
rect 22100 17833 22109 17867
rect 22109 17833 22143 17867
rect 22143 17833 22152 17867
rect 22100 17824 22152 17833
rect 22468 17824 22520 17876
rect 24768 17867 24820 17876
rect 9404 17756 9456 17808
rect 10692 17756 10744 17808
rect 11980 17756 12032 17808
rect 13820 17799 13872 17808
rect 13820 17765 13829 17799
rect 13829 17765 13863 17799
rect 13863 17765 13872 17799
rect 13820 17756 13872 17765
rect 14556 17756 14608 17808
rect 16304 17799 16356 17808
rect 16304 17765 16313 17799
rect 16313 17765 16347 17799
rect 16347 17765 16356 17799
rect 16304 17756 16356 17765
rect 17868 17799 17920 17808
rect 17868 17765 17877 17799
rect 17877 17765 17911 17799
rect 17911 17765 17920 17799
rect 17868 17756 17920 17765
rect 18420 17799 18472 17808
rect 18420 17765 18429 17799
rect 18429 17765 18463 17799
rect 18463 17765 18472 17799
rect 18420 17756 18472 17765
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 23020 17756 23072 17808
rect 11704 17731 11756 17740
rect 11704 17697 11713 17731
rect 11713 17697 11747 17731
rect 11747 17697 11756 17731
rect 11704 17688 11756 17697
rect 11796 17663 11848 17672
rect 11796 17629 11805 17663
rect 11805 17629 11839 17663
rect 11839 17629 11848 17663
rect 11796 17620 11848 17629
rect 12716 17688 12768 17740
rect 25044 17688 25096 17740
rect 13544 17620 13596 17672
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 16856 17663 16908 17672
rect 16120 17552 16172 17604
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 17776 17663 17828 17672
rect 16856 17620 16908 17629
rect 17776 17629 17785 17663
rect 17785 17629 17819 17663
rect 17819 17629 17828 17663
rect 17776 17620 17828 17629
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 22836 17663 22888 17672
rect 22836 17629 22845 17663
rect 22845 17629 22879 17663
rect 22879 17629 22888 17663
rect 22836 17620 22888 17629
rect 11244 17527 11296 17536
rect 11244 17493 11253 17527
rect 11253 17493 11287 17527
rect 11287 17493 11296 17527
rect 11244 17484 11296 17493
rect 12808 17484 12860 17536
rect 20536 17484 20588 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 9404 17280 9456 17332
rect 17776 17280 17828 17332
rect 21456 17280 21508 17332
rect 22192 17280 22244 17332
rect 22284 17280 22336 17332
rect 23020 17323 23072 17332
rect 23020 17289 23029 17323
rect 23029 17289 23063 17323
rect 23063 17289 23072 17323
rect 23020 17280 23072 17289
rect 21180 17212 21232 17264
rect 11244 17144 11296 17196
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 15660 17144 15712 17196
rect 18236 17144 18288 17196
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 20996 17144 21048 17196
rect 21548 17144 21600 17196
rect 22100 17187 22152 17196
rect 22100 17153 22109 17187
rect 22109 17153 22143 17187
rect 22143 17153 22152 17187
rect 22100 17144 22152 17153
rect 22836 17212 22888 17264
rect 24216 17144 24268 17196
rect 12072 17076 12124 17128
rect 12808 17076 12860 17128
rect 13820 17076 13872 17128
rect 24860 17076 24912 17128
rect 11520 17051 11572 17060
rect 9864 16940 9916 16992
rect 10876 16940 10928 16992
rect 11520 17017 11529 17051
rect 11529 17017 11563 17051
rect 11563 17017 11572 17051
rect 11520 17008 11572 17017
rect 12164 17008 12216 17060
rect 13360 17008 13412 17060
rect 17040 17008 17092 17060
rect 16304 16940 16356 16992
rect 17316 16940 17368 16992
rect 17776 16983 17828 16992
rect 17776 16949 17785 16983
rect 17785 16949 17819 16983
rect 17819 16949 17828 16983
rect 18328 17008 18380 17060
rect 20996 17008 21048 17060
rect 22100 17008 22152 17060
rect 17776 16940 17828 16949
rect 22284 16940 22336 16992
rect 25044 16983 25096 16992
rect 25044 16949 25053 16983
rect 25053 16949 25087 16983
rect 25087 16949 25096 16983
rect 25044 16940 25096 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 13728 16779 13780 16788
rect 13728 16745 13737 16779
rect 13737 16745 13771 16779
rect 13771 16745 13780 16779
rect 13728 16736 13780 16745
rect 15660 16779 15712 16788
rect 15660 16745 15669 16779
rect 15669 16745 15703 16779
rect 15703 16745 15712 16779
rect 15660 16736 15712 16745
rect 16120 16779 16172 16788
rect 16120 16745 16129 16779
rect 16129 16745 16163 16779
rect 16163 16745 16172 16779
rect 16120 16736 16172 16745
rect 16948 16779 17000 16788
rect 16948 16745 16957 16779
rect 16957 16745 16991 16779
rect 16991 16745 17000 16779
rect 16948 16736 17000 16745
rect 17868 16736 17920 16788
rect 20536 16779 20588 16788
rect 20536 16745 20545 16779
rect 20545 16745 20579 16779
rect 20579 16745 20588 16779
rect 20536 16736 20588 16745
rect 22468 16779 22520 16788
rect 22468 16745 22477 16779
rect 22477 16745 22511 16779
rect 22511 16745 22520 16779
rect 22468 16736 22520 16745
rect 10232 16668 10284 16720
rect 10692 16668 10744 16720
rect 12900 16711 12952 16720
rect 12900 16677 12909 16711
rect 12909 16677 12943 16711
rect 12943 16677 12952 16711
rect 12900 16668 12952 16677
rect 17316 16668 17368 16720
rect 18328 16668 18380 16720
rect 21272 16711 21324 16720
rect 21272 16677 21281 16711
rect 21281 16677 21315 16711
rect 21315 16677 21324 16711
rect 21272 16668 21324 16677
rect 22744 16711 22796 16720
rect 22744 16677 22753 16711
rect 22753 16677 22787 16711
rect 22787 16677 22796 16711
rect 22744 16668 22796 16677
rect 22928 16668 22980 16720
rect 15568 16600 15620 16652
rect 16672 16600 16724 16652
rect 19064 16643 19116 16652
rect 19064 16609 19073 16643
rect 19073 16609 19107 16643
rect 19107 16609 19116 16643
rect 19064 16600 19116 16609
rect 19248 16643 19300 16652
rect 19248 16609 19257 16643
rect 19257 16609 19291 16643
rect 19291 16609 19300 16643
rect 19248 16600 19300 16609
rect 10140 16532 10192 16584
rect 11152 16575 11204 16584
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 11520 16532 11572 16584
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 19524 16575 19576 16584
rect 19524 16541 19533 16575
rect 19533 16541 19567 16575
rect 19567 16541 19576 16575
rect 19524 16532 19576 16541
rect 21180 16575 21232 16584
rect 21180 16541 21189 16575
rect 21189 16541 21223 16575
rect 21223 16541 21232 16575
rect 21180 16532 21232 16541
rect 21732 16507 21784 16516
rect 21732 16473 21741 16507
rect 21741 16473 21775 16507
rect 21775 16473 21784 16507
rect 21732 16464 21784 16473
rect 22284 16464 22336 16516
rect 24676 16668 24728 16720
rect 24952 16711 25004 16720
rect 24952 16677 24961 16711
rect 24961 16677 24995 16711
rect 24995 16677 25004 16711
rect 24952 16668 25004 16677
rect 24216 16464 24268 16516
rect 10232 16439 10284 16448
rect 10232 16405 10241 16439
rect 10241 16405 10275 16439
rect 10275 16405 10284 16439
rect 10232 16396 10284 16405
rect 11244 16396 11296 16448
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 11796 16396 11848 16405
rect 18144 16439 18196 16448
rect 18144 16405 18153 16439
rect 18153 16405 18187 16439
rect 18187 16405 18196 16439
rect 18144 16396 18196 16405
rect 22100 16439 22152 16448
rect 22100 16405 22109 16439
rect 22109 16405 22143 16439
rect 22143 16405 22152 16439
rect 22100 16396 22152 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 12808 16192 12860 16244
rect 15568 16235 15620 16244
rect 10232 16124 10284 16176
rect 13452 16124 13504 16176
rect 15568 16201 15577 16235
rect 15577 16201 15611 16235
rect 15611 16201 15620 16235
rect 15568 16192 15620 16201
rect 16672 16192 16724 16244
rect 21272 16192 21324 16244
rect 22744 16192 22796 16244
rect 24676 16235 24728 16244
rect 24676 16201 24685 16235
rect 24685 16201 24719 16235
rect 24719 16201 24728 16235
rect 24676 16192 24728 16201
rect 16212 16124 16264 16176
rect 22928 16124 22980 16176
rect 11152 16056 11204 16108
rect 12164 16056 12216 16108
rect 7656 15988 7708 16040
rect 13176 16031 13228 16040
rect 13176 15997 13185 16031
rect 13185 15997 13219 16031
rect 13219 15997 13228 16031
rect 13176 15988 13228 15997
rect 13544 16056 13596 16108
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 14924 16056 14976 16108
rect 19524 16056 19576 16108
rect 18052 16031 18104 16040
rect 10048 15920 10100 15972
rect 8208 15852 8260 15904
rect 13912 15920 13964 15972
rect 16120 15963 16172 15972
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 13176 15895 13228 15904
rect 13176 15861 13185 15895
rect 13185 15861 13219 15895
rect 13219 15861 13228 15895
rect 13176 15852 13228 15861
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 16120 15929 16129 15963
rect 16129 15929 16163 15963
rect 16163 15929 16172 15963
rect 16120 15920 16172 15929
rect 16212 15963 16264 15972
rect 16212 15929 16221 15963
rect 16221 15929 16255 15963
rect 16255 15929 16264 15963
rect 16212 15920 16264 15929
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 18144 15988 18196 16040
rect 18972 15988 19024 16040
rect 21088 15988 21140 16040
rect 22100 15988 22152 16040
rect 14280 15852 14332 15861
rect 16948 15852 17000 15904
rect 17868 15895 17920 15904
rect 17868 15861 17877 15895
rect 17877 15861 17911 15895
rect 17911 15861 17920 15895
rect 17868 15852 17920 15861
rect 18144 15895 18196 15904
rect 18144 15861 18153 15895
rect 18153 15861 18187 15895
rect 18187 15861 18196 15895
rect 18144 15852 18196 15861
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 20260 15852 20312 15904
rect 22468 15895 22520 15904
rect 22468 15861 22477 15895
rect 22477 15861 22511 15895
rect 22511 15861 22520 15895
rect 22468 15852 22520 15861
rect 24216 15895 24268 15904
rect 24216 15861 24225 15895
rect 24225 15861 24259 15895
rect 24259 15861 24268 15895
rect 24216 15852 24268 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 12900 15648 12952 15700
rect 14556 15691 14608 15700
rect 14556 15657 14565 15691
rect 14565 15657 14599 15691
rect 14599 15657 14608 15691
rect 14556 15648 14608 15657
rect 17776 15648 17828 15700
rect 19248 15691 19300 15700
rect 19248 15657 19257 15691
rect 19257 15657 19291 15691
rect 19291 15657 19300 15691
rect 19248 15648 19300 15657
rect 19524 15648 19576 15700
rect 21180 15691 21232 15700
rect 21180 15657 21189 15691
rect 21189 15657 21223 15691
rect 21223 15657 21232 15691
rect 21180 15648 21232 15657
rect 24216 15648 24268 15700
rect 8208 15623 8260 15632
rect 8208 15589 8217 15623
rect 8217 15589 8251 15623
rect 8251 15589 8260 15623
rect 8208 15580 8260 15589
rect 10416 15623 10468 15632
rect 10416 15589 10425 15623
rect 10425 15589 10459 15623
rect 10459 15589 10468 15623
rect 10416 15580 10468 15589
rect 13360 15580 13412 15632
rect 15936 15580 15988 15632
rect 16948 15580 17000 15632
rect 12256 15512 12308 15564
rect 17500 15580 17552 15632
rect 21640 15580 21692 15632
rect 22468 15580 22520 15632
rect 8208 15444 8260 15496
rect 8300 15444 8352 15496
rect 11060 15444 11112 15496
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 17224 15444 17276 15496
rect 17960 15444 18012 15496
rect 18236 15487 18288 15496
rect 18236 15453 18245 15487
rect 18245 15453 18279 15487
rect 18279 15453 18288 15487
rect 18236 15444 18288 15453
rect 18420 15444 18472 15496
rect 21456 15444 21508 15496
rect 21732 15444 21784 15496
rect 22836 15444 22888 15496
rect 10784 15376 10836 15428
rect 13452 15376 13504 15428
rect 16120 15376 16172 15428
rect 20076 15376 20128 15428
rect 12532 15308 12584 15360
rect 16212 15351 16264 15360
rect 16212 15317 16221 15351
rect 16221 15317 16255 15351
rect 16255 15317 16264 15351
rect 16212 15308 16264 15317
rect 20444 15351 20496 15360
rect 20444 15317 20453 15351
rect 20453 15317 20487 15351
rect 20487 15317 20496 15351
rect 20444 15308 20496 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 8116 15104 8168 15156
rect 10416 15104 10468 15156
rect 10692 15147 10744 15156
rect 10692 15113 10701 15147
rect 10701 15113 10735 15147
rect 10735 15113 10744 15147
rect 10692 15104 10744 15113
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 14280 15104 14332 15156
rect 15476 15147 15528 15156
rect 15476 15113 15485 15147
rect 15485 15113 15519 15147
rect 15519 15113 15528 15147
rect 15476 15104 15528 15113
rect 15752 15104 15804 15156
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 18236 15104 18288 15156
rect 21640 15147 21692 15156
rect 21640 15113 21649 15147
rect 21649 15113 21683 15147
rect 21683 15113 21692 15147
rect 21640 15104 21692 15113
rect 21916 15104 21968 15156
rect 22652 15147 22704 15156
rect 22652 15113 22661 15147
rect 22661 15113 22695 15147
rect 22695 15113 22704 15147
rect 22652 15104 22704 15113
rect 8300 15011 8352 15020
rect 8300 14977 8309 15011
rect 8309 14977 8343 15011
rect 8343 14977 8352 15011
rect 8300 14968 8352 14977
rect 8024 14875 8076 14884
rect 8024 14841 8033 14875
rect 8033 14841 8067 14875
rect 8067 14841 8076 14875
rect 8024 14832 8076 14841
rect 10140 14968 10192 15020
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 16212 14968 16264 15020
rect 17960 14968 18012 15020
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 21456 14968 21508 15020
rect 12256 14943 12308 14952
rect 12256 14909 12265 14943
rect 12265 14909 12299 14943
rect 12299 14909 12308 14943
rect 12256 14900 12308 14909
rect 14648 14900 14700 14952
rect 15752 14900 15804 14952
rect 19340 14900 19392 14952
rect 20444 14900 20496 14952
rect 22652 14900 22704 14952
rect 23296 14900 23348 14952
rect 8944 14807 8996 14816
rect 8944 14773 8953 14807
rect 8953 14773 8987 14807
rect 8987 14773 8996 14807
rect 8944 14764 8996 14773
rect 9680 14764 9732 14816
rect 10048 14764 10100 14816
rect 13360 14764 13412 14816
rect 16488 14832 16540 14884
rect 14004 14764 14056 14816
rect 15936 14764 15988 14816
rect 18328 14764 18380 14816
rect 20260 14807 20312 14816
rect 20260 14773 20269 14807
rect 20269 14773 20303 14807
rect 20303 14773 20312 14807
rect 20260 14764 20312 14773
rect 21824 14764 21876 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 10692 14560 10744 14612
rect 11520 14603 11572 14612
rect 11520 14569 11529 14603
rect 11529 14569 11563 14603
rect 11563 14569 11572 14603
rect 11520 14560 11572 14569
rect 12716 14560 12768 14612
rect 12900 14560 12952 14612
rect 13360 14603 13412 14612
rect 13360 14569 13369 14603
rect 13369 14569 13403 14603
rect 13403 14569 13412 14603
rect 13360 14560 13412 14569
rect 13912 14603 13964 14612
rect 13912 14569 13921 14603
rect 13921 14569 13955 14603
rect 13955 14569 13964 14603
rect 13912 14560 13964 14569
rect 15936 14560 15988 14612
rect 16488 14560 16540 14612
rect 16856 14603 16908 14612
rect 16856 14569 16865 14603
rect 16865 14569 16899 14603
rect 16899 14569 16908 14603
rect 16856 14560 16908 14569
rect 17224 14603 17276 14612
rect 17224 14569 17233 14603
rect 17233 14569 17267 14603
rect 17267 14569 17276 14603
rect 17224 14560 17276 14569
rect 17776 14603 17828 14612
rect 17776 14569 17785 14603
rect 17785 14569 17819 14603
rect 17819 14569 17828 14603
rect 17776 14560 17828 14569
rect 18328 14603 18380 14612
rect 18328 14569 18337 14603
rect 18337 14569 18371 14603
rect 18371 14569 18380 14603
rect 18328 14560 18380 14569
rect 21272 14603 21324 14612
rect 21272 14569 21281 14603
rect 21281 14569 21315 14603
rect 21315 14569 21324 14603
rect 21272 14560 21324 14569
rect 8944 14492 8996 14544
rect 9772 14492 9824 14544
rect 18236 14492 18288 14544
rect 21088 14492 21140 14544
rect 21824 14492 21876 14544
rect 23020 14492 23072 14544
rect 1676 14424 1728 14476
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 9128 14424 9180 14476
rect 11428 14467 11480 14476
rect 11428 14433 11437 14467
rect 11437 14433 11471 14467
rect 11471 14433 11480 14467
rect 11428 14424 11480 14433
rect 11796 14424 11848 14476
rect 12164 14424 12216 14476
rect 13268 14424 13320 14476
rect 18144 14424 18196 14476
rect 18788 14424 18840 14476
rect 19248 14424 19300 14476
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 12256 14356 12308 14408
rect 14464 14356 14516 14408
rect 17408 14399 17460 14408
rect 17408 14365 17417 14399
rect 17417 14365 17451 14399
rect 17451 14365 17460 14399
rect 17408 14356 17460 14365
rect 20628 14356 20680 14408
rect 22744 14399 22796 14408
rect 22744 14365 22753 14399
rect 22753 14365 22787 14399
rect 22787 14365 22796 14399
rect 22744 14356 22796 14365
rect 22836 14356 22888 14408
rect 7288 14220 7340 14272
rect 8208 14220 8260 14272
rect 9220 14220 9272 14272
rect 17224 14220 17276 14272
rect 20168 14263 20220 14272
rect 20168 14229 20177 14263
rect 20177 14229 20211 14263
rect 20211 14229 20220 14263
rect 20168 14220 20220 14229
rect 22284 14220 22336 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 7288 14016 7340 14068
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 9956 14016 10008 14068
rect 10416 14016 10468 14068
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 17408 14016 17460 14068
rect 20996 14016 21048 14068
rect 22192 14016 22244 14068
rect 23020 14059 23072 14068
rect 23020 14025 23029 14059
rect 23029 14025 23063 14059
rect 23063 14025 23072 14059
rect 23020 14016 23072 14025
rect 25412 14059 25464 14068
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 10140 13948 10192 14000
rect 11428 13991 11480 14000
rect 11428 13957 11437 13991
rect 11437 13957 11471 13991
rect 11471 13957 11480 13991
rect 11428 13948 11480 13957
rect 8300 13880 8352 13932
rect 8208 13812 8260 13864
rect 8852 13880 8904 13932
rect 9404 13923 9456 13932
rect 9404 13889 9413 13923
rect 9413 13889 9447 13923
rect 9447 13889 9456 13923
rect 9404 13880 9456 13889
rect 9680 13880 9732 13932
rect 10692 13880 10744 13932
rect 11520 13880 11572 13932
rect 9128 13855 9180 13864
rect 9128 13821 9137 13855
rect 9137 13821 9171 13855
rect 9171 13821 9180 13855
rect 9128 13812 9180 13821
rect 10876 13812 10928 13864
rect 13084 13855 13136 13864
rect 13084 13821 13093 13855
rect 13093 13821 13127 13855
rect 13127 13821 13136 13855
rect 13084 13812 13136 13821
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 13820 13812 13872 13864
rect 7196 13787 7248 13796
rect 7196 13753 7205 13787
rect 7205 13753 7239 13787
rect 7239 13753 7248 13787
rect 7196 13744 7248 13753
rect 7288 13787 7340 13796
rect 7288 13753 7297 13787
rect 7297 13753 7331 13787
rect 7331 13753 7340 13787
rect 7288 13744 7340 13753
rect 8024 13744 8076 13796
rect 10048 13744 10100 13796
rect 10416 13744 10468 13796
rect 14004 13880 14056 13932
rect 1676 13719 1728 13728
rect 1676 13685 1685 13719
rect 1685 13685 1719 13719
rect 1719 13685 1728 13719
rect 1676 13676 1728 13685
rect 8116 13719 8168 13728
rect 8116 13685 8125 13719
rect 8125 13685 8159 13719
rect 8159 13685 8168 13719
rect 8116 13676 8168 13685
rect 11796 13719 11848 13728
rect 11796 13685 11805 13719
rect 11805 13685 11839 13719
rect 11839 13685 11848 13719
rect 11796 13676 11848 13685
rect 12716 13676 12768 13728
rect 13360 13676 13412 13728
rect 20260 13948 20312 14000
rect 21272 13948 21324 14000
rect 22928 13948 22980 14000
rect 23848 13948 23900 14000
rect 19248 13880 19300 13932
rect 20168 13923 20220 13932
rect 20168 13889 20177 13923
rect 20177 13889 20211 13923
rect 20211 13889 20220 13923
rect 20168 13880 20220 13889
rect 22744 13923 22796 13932
rect 22744 13889 22753 13923
rect 22753 13889 22787 13923
rect 22787 13889 22796 13923
rect 22744 13880 22796 13889
rect 23388 13880 23440 13932
rect 14832 13855 14884 13864
rect 14832 13821 14841 13855
rect 14841 13821 14875 13855
rect 14875 13821 14884 13855
rect 14832 13812 14884 13821
rect 16764 13812 16816 13864
rect 16488 13744 16540 13796
rect 18328 13812 18380 13864
rect 18788 13812 18840 13864
rect 19156 13855 19208 13864
rect 19156 13821 19165 13855
rect 19165 13821 19199 13855
rect 19199 13821 19208 13855
rect 19156 13812 19208 13821
rect 19340 13855 19392 13864
rect 19340 13821 19349 13855
rect 19349 13821 19383 13855
rect 19383 13821 19392 13855
rect 19340 13812 19392 13821
rect 24952 13812 25004 13864
rect 20260 13744 20312 13796
rect 22100 13787 22152 13796
rect 14464 13719 14516 13728
rect 14464 13685 14473 13719
rect 14473 13685 14507 13719
rect 14507 13685 14516 13719
rect 14464 13676 14516 13685
rect 15844 13676 15896 13728
rect 17776 13676 17828 13728
rect 18696 13676 18748 13728
rect 22100 13753 22109 13787
rect 22109 13753 22143 13787
rect 22143 13753 22152 13787
rect 22100 13744 22152 13753
rect 22192 13787 22244 13796
rect 22192 13753 22201 13787
rect 22201 13753 22235 13787
rect 22235 13753 22244 13787
rect 22192 13744 22244 13753
rect 20720 13676 20772 13728
rect 21272 13676 21324 13728
rect 23664 13676 23716 13728
rect 23848 13787 23900 13796
rect 23848 13753 23857 13787
rect 23857 13753 23891 13787
rect 23891 13753 23900 13787
rect 23848 13744 23900 13753
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 1676 13472 1728 13524
rect 9404 13515 9456 13524
rect 9404 13481 9413 13515
rect 9413 13481 9447 13515
rect 9447 13481 9456 13515
rect 9404 13472 9456 13481
rect 10692 13472 10744 13524
rect 11428 13472 11480 13524
rect 2780 13404 2832 13456
rect 1676 13336 1728 13388
rect 5540 13336 5592 13388
rect 9220 13404 9272 13456
rect 7380 13336 7432 13388
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 8392 13336 8444 13388
rect 10508 13336 10560 13388
rect 9496 13268 9548 13320
rect 11888 13404 11940 13456
rect 13820 13472 13872 13524
rect 14832 13472 14884 13524
rect 19248 13472 19300 13524
rect 15568 13404 15620 13456
rect 17224 13447 17276 13456
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 13268 13336 13320 13388
rect 15384 13336 15436 13388
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 17224 13413 17233 13447
rect 17233 13413 17267 13447
rect 17267 13413 17276 13447
rect 17224 13404 17276 13413
rect 18788 13404 18840 13456
rect 18420 13336 18472 13388
rect 20720 13404 20772 13456
rect 22284 13404 22336 13456
rect 23204 13404 23256 13456
rect 23388 13447 23440 13456
rect 23388 13413 23397 13447
rect 23397 13413 23431 13447
rect 23431 13413 23440 13447
rect 23388 13404 23440 13413
rect 20260 13336 20312 13388
rect 21824 13336 21876 13388
rect 24768 13336 24820 13388
rect 7748 13132 7800 13184
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 9680 13132 9732 13184
rect 9772 13132 9824 13184
rect 10876 13268 10928 13320
rect 13452 13311 13504 13320
rect 13452 13277 13461 13311
rect 13461 13277 13495 13311
rect 13495 13277 13504 13311
rect 13452 13268 13504 13277
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 17960 13268 18012 13320
rect 18236 13268 18288 13320
rect 22744 13311 22796 13320
rect 22744 13277 22753 13311
rect 22753 13277 22787 13311
rect 22787 13277 22796 13311
rect 22744 13268 22796 13277
rect 11796 13243 11848 13252
rect 11796 13209 11805 13243
rect 11805 13209 11839 13243
rect 11839 13209 11848 13243
rect 11796 13200 11848 13209
rect 16672 13200 16724 13252
rect 17684 13200 17736 13252
rect 18696 13200 18748 13252
rect 22928 13200 22980 13252
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 16028 13132 16080 13184
rect 16488 13175 16540 13184
rect 16488 13141 16497 13175
rect 16497 13141 16531 13175
rect 16531 13141 16540 13175
rect 16488 13132 16540 13141
rect 18788 13132 18840 13184
rect 20628 13175 20680 13184
rect 20628 13141 20637 13175
rect 20637 13141 20671 13175
rect 20671 13141 20680 13175
rect 20628 13132 20680 13141
rect 22192 13175 22244 13184
rect 22192 13141 22201 13175
rect 22201 13141 22235 13175
rect 22235 13141 22244 13175
rect 22192 13132 22244 13141
rect 23664 13175 23716 13184
rect 23664 13141 23673 13175
rect 23673 13141 23707 13175
rect 23707 13141 23716 13175
rect 23664 13132 23716 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 6920 12928 6972 12980
rect 7380 12971 7432 12980
rect 7380 12937 7389 12971
rect 7389 12937 7423 12971
rect 7423 12937 7432 12971
rect 7380 12928 7432 12937
rect 8300 12928 8352 12980
rect 10140 12928 10192 12980
rect 10508 12971 10560 12980
rect 10508 12937 10517 12971
rect 10517 12937 10551 12971
rect 10551 12937 10560 12971
rect 10508 12928 10560 12937
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 13084 12928 13136 12980
rect 16672 12928 16724 12980
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 17224 12971 17276 12980
rect 17224 12937 17233 12971
rect 17233 12937 17267 12971
rect 17267 12937 17276 12971
rect 17224 12928 17276 12937
rect 18696 12928 18748 12980
rect 18972 12928 19024 12980
rect 21824 12971 21876 12980
rect 21824 12937 21833 12971
rect 21833 12937 21867 12971
rect 21867 12937 21876 12971
rect 21824 12928 21876 12937
rect 22192 12928 22244 12980
rect 23204 12971 23256 12980
rect 23204 12937 23213 12971
rect 23213 12937 23247 12971
rect 23247 12937 23256 12971
rect 23204 12928 23256 12937
rect 23664 12928 23716 12980
rect 7196 12860 7248 12912
rect 11520 12860 11572 12912
rect 15476 12903 15528 12912
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 7748 12792 7800 12844
rect 9404 12792 9456 12844
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 12532 12792 12584 12844
rect 15476 12869 15485 12903
rect 15485 12869 15519 12903
rect 15519 12869 15528 12903
rect 15476 12860 15528 12869
rect 15752 12860 15804 12912
rect 17868 12860 17920 12912
rect 22652 12860 22704 12912
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 15568 12792 15620 12844
rect 17500 12792 17552 12844
rect 18420 12835 18472 12844
rect 18420 12801 18429 12835
rect 18429 12801 18463 12835
rect 18463 12801 18472 12835
rect 18420 12792 18472 12801
rect 18604 12792 18656 12844
rect 7196 12724 7248 12776
rect 8208 12767 8260 12776
rect 8208 12733 8217 12767
rect 8217 12733 8251 12767
rect 8251 12733 8260 12767
rect 8208 12724 8260 12733
rect 8392 12767 8444 12776
rect 8392 12733 8401 12767
rect 8401 12733 8435 12767
rect 8435 12733 8444 12767
rect 8392 12724 8444 12733
rect 9220 12724 9272 12776
rect 15936 12767 15988 12776
rect 5540 12699 5592 12708
rect 5540 12665 5549 12699
rect 5549 12665 5583 12699
rect 5583 12665 5592 12699
rect 5540 12656 5592 12665
rect 8484 12656 8536 12708
rect 9588 12656 9640 12708
rect 9772 12656 9824 12708
rect 15936 12733 15945 12767
rect 15945 12733 15979 12767
rect 15979 12733 15988 12767
rect 15936 12724 15988 12733
rect 12716 12656 12768 12708
rect 14280 12699 14332 12708
rect 14280 12665 14289 12699
rect 14289 12665 14323 12699
rect 14323 12665 14332 12699
rect 14280 12656 14332 12665
rect 6276 12588 6328 12640
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 11612 12631 11664 12640
rect 11612 12597 11621 12631
rect 11621 12597 11655 12631
rect 11655 12597 11664 12631
rect 11612 12588 11664 12597
rect 14188 12588 14240 12640
rect 15844 12631 15896 12640
rect 15844 12597 15853 12631
rect 15853 12597 15887 12631
rect 15887 12597 15896 12631
rect 16304 12631 16356 12640
rect 15844 12588 15896 12597
rect 16304 12597 16313 12631
rect 16313 12597 16347 12631
rect 16347 12597 16356 12631
rect 16304 12588 16356 12597
rect 17132 12588 17184 12640
rect 18144 12588 18196 12640
rect 18696 12588 18748 12640
rect 19248 12724 19300 12776
rect 20628 12724 20680 12776
rect 20904 12699 20956 12708
rect 20904 12665 20913 12699
rect 20913 12665 20947 12699
rect 20947 12665 20956 12699
rect 20904 12656 20956 12665
rect 21180 12656 21232 12708
rect 21548 12699 21600 12708
rect 21548 12665 21557 12699
rect 21557 12665 21591 12699
rect 21591 12665 21600 12699
rect 21548 12656 21600 12665
rect 20352 12631 20404 12640
rect 20352 12597 20361 12631
rect 20361 12597 20395 12631
rect 20395 12597 20404 12631
rect 20352 12588 20404 12597
rect 20628 12631 20680 12640
rect 20628 12597 20637 12631
rect 20637 12597 20671 12631
rect 20671 12597 20680 12631
rect 20628 12588 20680 12597
rect 25136 12767 25188 12776
rect 25136 12733 25145 12767
rect 25145 12733 25179 12767
rect 25179 12733 25188 12767
rect 25136 12724 25188 12733
rect 25228 12656 25280 12708
rect 22928 12631 22980 12640
rect 22928 12597 22937 12631
rect 22937 12597 22971 12631
rect 22971 12597 22980 12631
rect 22928 12588 22980 12597
rect 24768 12588 24820 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 8392 12384 8444 12436
rect 9404 12427 9456 12436
rect 9404 12393 9413 12427
rect 9413 12393 9447 12427
rect 9447 12393 9456 12427
rect 9404 12384 9456 12393
rect 9956 12384 10008 12436
rect 11428 12384 11480 12436
rect 12532 12427 12584 12436
rect 6184 12316 6236 12368
rect 7840 12359 7892 12368
rect 7840 12325 7849 12359
rect 7849 12325 7883 12359
rect 7883 12325 7892 12359
rect 7840 12316 7892 12325
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 13636 12427 13688 12436
rect 13636 12393 13645 12427
rect 13645 12393 13679 12427
rect 13679 12393 13688 12427
rect 13636 12384 13688 12393
rect 15568 12427 15620 12436
rect 15568 12393 15577 12427
rect 15577 12393 15611 12427
rect 15611 12393 15620 12427
rect 15568 12384 15620 12393
rect 17040 12427 17092 12436
rect 17040 12393 17049 12427
rect 17049 12393 17083 12427
rect 17083 12393 17092 12427
rect 17040 12384 17092 12393
rect 17776 12384 17828 12436
rect 16304 12316 16356 12368
rect 18144 12384 18196 12436
rect 21548 12384 21600 12436
rect 21824 12384 21876 12436
rect 22744 12384 22796 12436
rect 18788 12316 18840 12368
rect 19248 12359 19300 12368
rect 19248 12325 19257 12359
rect 19257 12325 19291 12359
rect 19291 12325 19300 12359
rect 19248 12316 19300 12325
rect 21364 12359 21416 12368
rect 21364 12325 21373 12359
rect 21373 12325 21407 12359
rect 21407 12325 21416 12359
rect 21364 12316 21416 12325
rect 23112 12316 23164 12368
rect 1216 12248 1268 12300
rect 16120 12291 16172 12300
rect 16120 12257 16129 12291
rect 16129 12257 16163 12291
rect 16163 12257 16172 12291
rect 16120 12248 16172 12257
rect 19524 12248 19576 12300
rect 22744 12291 22796 12300
rect 22744 12257 22753 12291
rect 22753 12257 22787 12291
rect 22787 12257 22796 12291
rect 22744 12248 22796 12257
rect 24676 12248 24728 12300
rect 6276 12180 6328 12232
rect 6920 12180 6972 12232
rect 8208 12180 8260 12232
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 10048 12180 10100 12232
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 13728 12180 13780 12232
rect 17408 12180 17460 12232
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 21272 12223 21324 12232
rect 21272 12189 21281 12223
rect 21281 12189 21315 12223
rect 21315 12189 21324 12223
rect 21272 12180 21324 12189
rect 22192 12180 22244 12232
rect 7472 12112 7524 12164
rect 8484 12112 8536 12164
rect 14556 12112 14608 12164
rect 15936 12112 15988 12164
rect 25136 12180 25188 12232
rect 8576 12044 8628 12096
rect 9220 12044 9272 12096
rect 12440 12044 12492 12096
rect 13268 12044 13320 12096
rect 14004 12044 14056 12096
rect 14280 12044 14332 12096
rect 19984 12087 20036 12096
rect 19984 12053 19993 12087
rect 19993 12053 20027 12087
rect 20027 12053 20036 12087
rect 19984 12044 20036 12053
rect 22100 12044 22152 12096
rect 23756 12087 23808 12096
rect 23756 12053 23765 12087
rect 23765 12053 23799 12087
rect 23799 12053 23808 12087
rect 23756 12044 23808 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1216 11840 1268 11892
rect 7840 11883 7892 11892
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 7840 11840 7892 11849
rect 8208 11883 8260 11892
rect 8208 11849 8217 11883
rect 8217 11849 8251 11883
rect 8251 11849 8260 11883
rect 8208 11840 8260 11849
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 7196 11747 7248 11756
rect 7196 11713 7205 11747
rect 7205 11713 7239 11747
rect 7239 11713 7248 11747
rect 7196 11704 7248 11713
rect 9312 11840 9364 11892
rect 9680 11840 9732 11892
rect 11428 11883 11480 11892
rect 11428 11849 11437 11883
rect 11437 11849 11471 11883
rect 11471 11849 11480 11883
rect 11428 11840 11480 11849
rect 11520 11840 11572 11892
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 14188 11840 14240 11849
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 20076 11840 20128 11892
rect 23204 11840 23256 11892
rect 24952 11840 25004 11892
rect 9036 11772 9088 11824
rect 19524 11815 19576 11824
rect 19524 11781 19533 11815
rect 19533 11781 19567 11815
rect 19567 11781 19576 11815
rect 19524 11772 19576 11781
rect 24676 11772 24728 11824
rect 25228 11815 25280 11824
rect 25228 11781 25237 11815
rect 25237 11781 25271 11815
rect 25271 11781 25280 11815
rect 25228 11772 25280 11781
rect 9496 11704 9548 11756
rect 13452 11704 13504 11756
rect 18236 11704 18288 11756
rect 13728 11636 13780 11688
rect 15752 11636 15804 11688
rect 18328 11679 18380 11688
rect 18328 11645 18337 11679
rect 18337 11645 18371 11679
rect 18371 11645 18380 11679
rect 19892 11704 19944 11756
rect 21824 11747 21876 11756
rect 21824 11713 21833 11747
rect 21833 11713 21867 11747
rect 21867 11713 21876 11747
rect 21824 11704 21876 11713
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 22744 11747 22796 11756
rect 22744 11713 22753 11747
rect 22753 11713 22787 11747
rect 22787 11713 22796 11747
rect 22744 11704 22796 11713
rect 23112 11747 23164 11756
rect 23112 11713 23121 11747
rect 23121 11713 23155 11747
rect 23155 11713 23164 11747
rect 23112 11704 23164 11713
rect 18328 11636 18380 11645
rect 18512 11636 18564 11688
rect 19524 11636 19576 11688
rect 19984 11679 20036 11688
rect 19984 11645 19993 11679
rect 19993 11645 20027 11679
rect 20027 11645 20036 11679
rect 19984 11636 20036 11645
rect 6184 11611 6236 11620
rect 6184 11577 6193 11611
rect 6193 11577 6227 11611
rect 6227 11577 6236 11611
rect 6184 11568 6236 11577
rect 6920 11611 6972 11620
rect 6920 11577 6929 11611
rect 6929 11577 6963 11611
rect 6963 11577 6972 11611
rect 6920 11568 6972 11577
rect 6552 11543 6604 11552
rect 6552 11509 6561 11543
rect 6561 11509 6595 11543
rect 6595 11509 6604 11543
rect 6552 11500 6604 11509
rect 7932 11500 7984 11552
rect 9312 11543 9364 11552
rect 9312 11509 9321 11543
rect 9321 11509 9355 11543
rect 9355 11509 9364 11543
rect 9956 11568 10008 11620
rect 13268 11568 13320 11620
rect 13636 11611 13688 11620
rect 13636 11577 13639 11611
rect 13639 11577 13673 11611
rect 13673 11577 13688 11611
rect 16488 11611 16540 11620
rect 13636 11568 13688 11577
rect 16488 11577 16497 11611
rect 16497 11577 16531 11611
rect 16531 11577 16540 11611
rect 16488 11568 16540 11577
rect 16856 11568 16908 11620
rect 19156 11611 19208 11620
rect 19156 11577 19165 11611
rect 19165 11577 19199 11611
rect 19199 11577 19208 11611
rect 19156 11568 19208 11577
rect 9312 11500 9364 11509
rect 9772 11500 9824 11552
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 19248 11500 19300 11552
rect 20628 11568 20680 11620
rect 20812 11500 20864 11552
rect 21364 11500 21416 11552
rect 23756 11636 23808 11688
rect 24676 11500 24728 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6276 11296 6328 11305
rect 8208 11296 8260 11348
rect 10876 11296 10928 11348
rect 5080 11228 5132 11280
rect 6920 11228 6972 11280
rect 7012 11271 7064 11280
rect 7012 11237 7021 11271
rect 7021 11237 7055 11271
rect 7055 11237 7064 11271
rect 7012 11228 7064 11237
rect 9496 11228 9548 11280
rect 11336 11296 11388 11348
rect 13268 11339 13320 11348
rect 13268 11305 13277 11339
rect 13277 11305 13311 11339
rect 13311 11305 13320 11339
rect 13268 11296 13320 11305
rect 16120 11296 16172 11348
rect 16856 11296 16908 11348
rect 20352 11296 20404 11348
rect 11428 11228 11480 11280
rect 11796 11228 11848 11280
rect 4252 11160 4304 11212
rect 8484 11160 8536 11212
rect 10692 11160 10744 11212
rect 4712 11092 4764 11144
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 7472 11024 7524 11076
rect 14004 11228 14056 11280
rect 14556 11228 14608 11280
rect 15476 11271 15528 11280
rect 15476 11237 15485 11271
rect 15485 11237 15519 11271
rect 15519 11237 15528 11271
rect 15476 11228 15528 11237
rect 16488 11228 16540 11280
rect 19248 11228 19300 11280
rect 21180 11228 21232 11280
rect 23572 11271 23624 11280
rect 23572 11237 23581 11271
rect 23581 11237 23615 11271
rect 23615 11237 23624 11271
rect 23572 11228 23624 11237
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 18512 11160 18564 11212
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 19064 11135 19116 11144
rect 12992 10999 13044 11008
rect 12992 10965 13001 10999
rect 13001 10965 13035 10999
rect 13035 10965 13044 10999
rect 12992 10956 13044 10965
rect 19064 11101 19073 11135
rect 19073 11101 19107 11135
rect 19107 11101 19116 11135
rect 19064 11092 19116 11101
rect 21916 11135 21968 11144
rect 21916 11101 21925 11135
rect 21925 11101 21959 11135
rect 21959 11101 21968 11135
rect 21916 11092 21968 11101
rect 23756 11135 23808 11144
rect 21548 11024 21600 11076
rect 18512 10999 18564 11008
rect 18512 10965 18521 10999
rect 18521 10965 18555 10999
rect 18555 10965 18564 10999
rect 18512 10956 18564 10965
rect 21272 10999 21324 11008
rect 21272 10965 21281 10999
rect 21281 10965 21315 10999
rect 21315 10965 21324 10999
rect 21272 10956 21324 10965
rect 21364 10956 21416 11008
rect 23756 11101 23765 11135
rect 23765 11101 23799 11135
rect 23799 11101 23808 11135
rect 23756 11092 23808 11101
rect 24676 10956 24728 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 4252 10795 4304 10804
rect 4252 10761 4261 10795
rect 4261 10761 4295 10795
rect 4295 10761 4304 10795
rect 4252 10752 4304 10761
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 5080 10795 5132 10804
rect 5080 10761 5089 10795
rect 5089 10761 5123 10795
rect 5123 10761 5132 10795
rect 5080 10752 5132 10761
rect 6184 10752 6236 10804
rect 7932 10795 7984 10804
rect 7932 10761 7941 10795
rect 7941 10761 7975 10795
rect 7975 10761 7984 10795
rect 7932 10752 7984 10761
rect 11060 10752 11112 10804
rect 11796 10752 11848 10804
rect 15384 10752 15436 10804
rect 16488 10752 16540 10804
rect 17224 10752 17276 10804
rect 17500 10795 17552 10804
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 20812 10795 20864 10804
rect 20812 10761 20821 10795
rect 20821 10761 20855 10795
rect 20855 10761 20864 10795
rect 20812 10752 20864 10761
rect 21180 10795 21232 10804
rect 21180 10761 21189 10795
rect 21189 10761 21223 10795
rect 21223 10761 21232 10795
rect 21180 10752 21232 10761
rect 21916 10752 21968 10804
rect 23572 10752 23624 10804
rect 24676 10752 24728 10804
rect 7472 10727 7524 10736
rect 6552 10616 6604 10668
rect 7472 10693 7481 10727
rect 7481 10693 7515 10727
rect 7515 10693 7524 10727
rect 7472 10684 7524 10693
rect 12716 10684 12768 10736
rect 13636 10684 13688 10736
rect 15476 10684 15528 10736
rect 8484 10659 8536 10668
rect 8484 10625 8493 10659
rect 8493 10625 8527 10659
rect 8527 10625 8536 10659
rect 8484 10616 8536 10625
rect 12992 10616 13044 10668
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 13544 10616 13596 10625
rect 13728 10616 13780 10668
rect 18788 10659 18840 10668
rect 18788 10625 18797 10659
rect 18797 10625 18831 10659
rect 18831 10625 18840 10659
rect 18788 10616 18840 10625
rect 19156 10616 19208 10668
rect 20168 10616 20220 10668
rect 11612 10548 11664 10600
rect 11796 10548 11848 10600
rect 9772 10523 9824 10532
rect 9772 10489 9781 10523
rect 9781 10489 9815 10523
rect 9815 10489 9824 10523
rect 9772 10480 9824 10489
rect 11520 10480 11572 10532
rect 6276 10455 6328 10464
rect 6276 10421 6285 10455
rect 6285 10421 6319 10455
rect 6319 10421 6328 10455
rect 6276 10412 6328 10421
rect 9036 10455 9088 10464
rect 9036 10421 9045 10455
rect 9045 10421 9079 10455
rect 9079 10421 9088 10455
rect 9036 10412 9088 10421
rect 10692 10455 10744 10464
rect 10692 10421 10701 10455
rect 10701 10421 10735 10455
rect 10735 10421 10744 10455
rect 10692 10412 10744 10421
rect 11428 10412 11480 10464
rect 13636 10523 13688 10532
rect 13636 10489 13645 10523
rect 13645 10489 13679 10523
rect 13679 10489 13688 10523
rect 13636 10480 13688 10489
rect 14188 10523 14240 10532
rect 14188 10489 14197 10523
rect 14197 10489 14231 10523
rect 14231 10489 14240 10523
rect 14188 10480 14240 10489
rect 15108 10548 15160 10600
rect 15568 10480 15620 10532
rect 21364 10548 21416 10600
rect 22928 10548 22980 10600
rect 18144 10523 18196 10532
rect 18144 10489 18153 10523
rect 18153 10489 18187 10523
rect 18187 10489 18196 10523
rect 18144 10480 18196 10489
rect 13084 10412 13136 10464
rect 14004 10412 14056 10464
rect 17132 10455 17184 10464
rect 17132 10421 17141 10455
rect 17141 10421 17175 10455
rect 17175 10421 17184 10455
rect 17132 10412 17184 10421
rect 18328 10480 18380 10532
rect 19248 10412 19300 10464
rect 23388 10480 23440 10532
rect 24216 10523 24268 10532
rect 24216 10489 24225 10523
rect 24225 10489 24259 10523
rect 24259 10489 24268 10523
rect 24216 10480 24268 10489
rect 22560 10455 22612 10464
rect 22560 10421 22569 10455
rect 22569 10421 22603 10455
rect 22603 10421 22612 10455
rect 22560 10412 22612 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 6276 10208 6328 10260
rect 7288 10208 7340 10260
rect 7472 10208 7524 10260
rect 11060 10251 11112 10260
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 12440 10251 12492 10260
rect 12440 10217 12449 10251
rect 12449 10217 12483 10251
rect 12483 10217 12492 10251
rect 12440 10208 12492 10217
rect 12992 10208 13044 10260
rect 11336 10183 11388 10192
rect 11336 10149 11345 10183
rect 11345 10149 11379 10183
rect 11379 10149 11388 10183
rect 11336 10140 11388 10149
rect 11428 10183 11480 10192
rect 11428 10149 11437 10183
rect 11437 10149 11471 10183
rect 11471 10149 11480 10183
rect 13268 10183 13320 10192
rect 11428 10140 11480 10149
rect 13268 10149 13271 10183
rect 13271 10149 13305 10183
rect 13305 10149 13320 10183
rect 13268 10140 13320 10149
rect 13636 10208 13688 10260
rect 15108 10251 15160 10260
rect 15108 10217 15117 10251
rect 15117 10217 15151 10251
rect 15151 10217 15160 10251
rect 15108 10208 15160 10217
rect 15568 10208 15620 10260
rect 16120 10208 16172 10260
rect 16028 10183 16080 10192
rect 16028 10149 16037 10183
rect 16037 10149 16071 10183
rect 16071 10149 16080 10183
rect 16028 10140 16080 10149
rect 17316 10140 17368 10192
rect 19064 10208 19116 10260
rect 20168 10251 20220 10260
rect 20168 10217 20177 10251
rect 20177 10217 20211 10251
rect 20211 10217 20220 10251
rect 20168 10208 20220 10217
rect 23020 10208 23072 10260
rect 23756 10208 23808 10260
rect 19340 10140 19392 10192
rect 21364 10140 21416 10192
rect 21640 10183 21692 10192
rect 21640 10149 21649 10183
rect 21649 10149 21683 10183
rect 21683 10149 21692 10183
rect 21640 10140 21692 10149
rect 22560 10140 22612 10192
rect 7840 10072 7892 10124
rect 6460 10047 6512 10056
rect 6460 10013 6469 10047
rect 6469 10013 6503 10047
rect 6503 10013 6512 10047
rect 6460 10004 6512 10013
rect 10048 10047 10100 10056
rect 4436 9936 4488 9988
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 11520 10004 11572 10056
rect 14188 10072 14240 10124
rect 15292 10115 15344 10124
rect 15292 10081 15301 10115
rect 15301 10081 15335 10115
rect 15335 10081 15344 10115
rect 15292 10072 15344 10081
rect 15568 10115 15620 10124
rect 15568 10081 15577 10115
rect 15577 10081 15611 10115
rect 15611 10081 15620 10115
rect 15568 10072 15620 10081
rect 19064 10115 19116 10124
rect 19064 10081 19073 10115
rect 19073 10081 19107 10115
rect 19107 10081 19116 10115
rect 19064 10072 19116 10081
rect 19156 10072 19208 10124
rect 22192 10115 22244 10124
rect 22192 10081 22201 10115
rect 22201 10081 22235 10115
rect 22235 10081 22244 10115
rect 23112 10115 23164 10124
rect 22192 10072 22244 10081
rect 23112 10081 23121 10115
rect 23121 10081 23155 10115
rect 23155 10081 23164 10115
rect 23112 10072 23164 10081
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 16948 10047 17000 10056
rect 10692 9936 10744 9988
rect 11980 9936 12032 9988
rect 15384 9979 15436 9988
rect 15384 9945 15393 9979
rect 15393 9945 15427 9979
rect 15427 9945 15436 9979
rect 15384 9936 15436 9945
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 17592 10047 17644 10056
rect 17592 10013 17601 10047
rect 17601 10013 17635 10047
rect 17635 10013 17644 10047
rect 17592 10004 17644 10013
rect 21548 10047 21600 10056
rect 21548 10013 21557 10047
rect 21557 10013 21591 10047
rect 21591 10013 21600 10047
rect 21548 10004 21600 10013
rect 18144 9936 18196 9988
rect 18328 9936 18380 9988
rect 8116 9868 8168 9920
rect 12164 9868 12216 9920
rect 14556 9911 14608 9920
rect 14556 9877 14565 9911
rect 14565 9877 14599 9911
rect 14599 9877 14608 9911
rect 14556 9868 14608 9877
rect 18512 9868 18564 9920
rect 19156 9868 19208 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 6276 9664 6328 9716
rect 7012 9664 7064 9716
rect 9864 9664 9916 9716
rect 7288 9596 7340 9648
rect 9312 9639 9364 9648
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 10692 9639 10744 9648
rect 10692 9605 10701 9639
rect 10701 9605 10735 9639
rect 10735 9605 10744 9639
rect 10692 9596 10744 9605
rect 11336 9664 11388 9716
rect 12164 9707 12216 9716
rect 12164 9673 12173 9707
rect 12173 9673 12207 9707
rect 12207 9673 12216 9707
rect 12164 9664 12216 9673
rect 13268 9664 13320 9716
rect 15292 9664 15344 9716
rect 17408 9664 17460 9716
rect 11428 9596 11480 9648
rect 1676 9528 1728 9580
rect 9036 9528 9088 9580
rect 11980 9528 12032 9580
rect 18696 9664 18748 9716
rect 21640 9707 21692 9716
rect 21640 9673 21649 9707
rect 21649 9673 21683 9707
rect 21683 9673 21692 9707
rect 21640 9664 21692 9673
rect 21916 9664 21968 9716
rect 22652 9707 22704 9716
rect 22652 9673 22661 9707
rect 22661 9673 22695 9707
rect 22695 9673 22704 9707
rect 22652 9664 22704 9673
rect 23112 9707 23164 9716
rect 23112 9673 23121 9707
rect 23121 9673 23155 9707
rect 23155 9673 23164 9707
rect 23112 9664 23164 9673
rect 7288 9392 7340 9444
rect 5908 9367 5960 9376
rect 5908 9333 5917 9367
rect 5917 9333 5951 9367
rect 5951 9333 5960 9367
rect 5908 9324 5960 9333
rect 8116 9367 8168 9376
rect 8116 9333 8125 9367
rect 8125 9333 8159 9367
rect 8159 9333 8168 9367
rect 8116 9324 8168 9333
rect 12992 9503 13044 9512
rect 12992 9469 13001 9503
rect 13001 9469 13035 9503
rect 13035 9469 13044 9503
rect 12992 9460 13044 9469
rect 18604 9596 18656 9648
rect 17592 9528 17644 9580
rect 18788 9571 18840 9580
rect 18788 9537 18797 9571
rect 18797 9537 18831 9571
rect 18831 9537 18840 9571
rect 18788 9528 18840 9537
rect 14556 9460 14608 9512
rect 15200 9503 15252 9512
rect 15200 9469 15209 9503
rect 15209 9469 15243 9503
rect 15243 9469 15252 9503
rect 15200 9460 15252 9469
rect 15292 9392 15344 9444
rect 13544 9324 13596 9376
rect 14648 9324 14700 9376
rect 15660 9435 15712 9444
rect 15660 9401 15669 9435
rect 15669 9401 15703 9435
rect 15703 9401 15712 9435
rect 15660 9392 15712 9401
rect 15568 9324 15620 9376
rect 16672 9392 16724 9444
rect 23112 9528 23164 9580
rect 23204 9528 23256 9580
rect 23940 9528 23992 9580
rect 22008 9460 22060 9512
rect 22652 9460 22704 9512
rect 20628 9435 20680 9444
rect 20628 9401 20637 9435
rect 20637 9401 20671 9435
rect 20671 9401 20680 9435
rect 20628 9392 20680 9401
rect 20720 9435 20772 9444
rect 20720 9401 20729 9435
rect 20729 9401 20763 9435
rect 20763 9401 20772 9435
rect 21272 9435 21324 9444
rect 20720 9392 20772 9401
rect 21272 9401 21281 9435
rect 21281 9401 21315 9435
rect 21315 9401 21324 9435
rect 21272 9392 21324 9401
rect 23020 9392 23072 9444
rect 17040 9367 17092 9376
rect 17040 9333 17049 9367
rect 17049 9333 17083 9367
rect 17083 9333 17092 9367
rect 17040 9324 17092 9333
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 19064 9367 19116 9376
rect 19064 9333 19073 9367
rect 19073 9333 19107 9367
rect 19107 9333 19116 9367
rect 19064 9324 19116 9333
rect 19156 9324 19208 9376
rect 21548 9324 21600 9376
rect 22192 9324 22244 9376
rect 25136 9367 25188 9376
rect 25136 9333 25145 9367
rect 25145 9333 25179 9367
rect 25179 9333 25188 9367
rect 25136 9324 25188 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 5908 9120 5960 9172
rect 6460 9120 6512 9172
rect 11244 9120 11296 9172
rect 12900 9163 12952 9172
rect 12900 9129 12909 9163
rect 12909 9129 12943 9163
rect 12943 9129 12952 9163
rect 12900 9120 12952 9129
rect 14648 9120 14700 9172
rect 15384 9120 15436 9172
rect 16672 9120 16724 9172
rect 21180 9120 21232 9172
rect 6092 9052 6144 9104
rect 12992 9052 13044 9104
rect 5080 9027 5132 9036
rect 5080 8993 5089 9027
rect 5089 8993 5123 9027
rect 5123 8993 5132 9027
rect 5080 8984 5132 8993
rect 5172 8984 5224 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 7380 9027 7432 9036
rect 7380 8993 7389 9027
rect 7389 8993 7423 9027
rect 7423 8993 7432 9027
rect 7380 8984 7432 8993
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 11152 9027 11204 9036
rect 5540 8848 5592 8900
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 11796 8984 11848 9036
rect 11980 8984 12032 9036
rect 12256 9027 12308 9036
rect 12256 8993 12265 9027
rect 12265 8993 12299 9027
rect 12299 8993 12308 9027
rect 12256 8984 12308 8993
rect 13360 9027 13412 9036
rect 13360 8993 13369 9027
rect 13369 8993 13403 9027
rect 13403 8993 13412 9027
rect 13360 8984 13412 8993
rect 14372 9052 14424 9104
rect 14556 9052 14608 9104
rect 16304 9052 16356 9104
rect 17500 9052 17552 9104
rect 22836 9095 22888 9104
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 18696 8984 18748 9036
rect 16948 8916 17000 8968
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9404 8780 9456 8789
rect 9864 8780 9916 8832
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 17592 8916 17644 8968
rect 19156 8984 19208 9036
rect 22836 9061 22845 9095
rect 22845 9061 22879 9095
rect 22879 9061 22888 9095
rect 22836 9052 22888 9061
rect 24124 9052 24176 9104
rect 19340 8916 19392 8968
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 19708 8916 19760 8925
rect 20904 8959 20956 8968
rect 20904 8925 20913 8959
rect 20913 8925 20947 8959
rect 20947 8925 20956 8959
rect 20904 8916 20956 8925
rect 22744 8959 22796 8968
rect 22744 8925 22753 8959
rect 22753 8925 22787 8959
rect 22787 8925 22796 8959
rect 22744 8916 22796 8925
rect 23020 8959 23072 8968
rect 23020 8925 23029 8959
rect 23029 8925 23063 8959
rect 23063 8925 23072 8959
rect 23020 8916 23072 8925
rect 23388 8916 23440 8968
rect 18236 8848 18288 8900
rect 14464 8780 14516 8832
rect 15292 8780 15344 8832
rect 15844 8780 15896 8832
rect 20628 8780 20680 8832
rect 22192 8780 22244 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 5080 8576 5132 8628
rect 7564 8576 7616 8628
rect 5172 8551 5224 8560
rect 5172 8517 5181 8551
rect 5181 8517 5215 8551
rect 5215 8517 5224 8551
rect 9680 8576 9732 8628
rect 9956 8576 10008 8628
rect 11612 8576 11664 8628
rect 13360 8576 13412 8628
rect 15660 8576 15712 8628
rect 16488 8576 16540 8628
rect 5172 8508 5224 8517
rect 8116 8508 8168 8560
rect 8668 8508 8720 8560
rect 10968 8551 11020 8560
rect 9128 8440 9180 8492
rect 10968 8517 10977 8551
rect 10977 8517 11011 8551
rect 11011 8517 11020 8551
rect 10968 8508 11020 8517
rect 12256 8508 12308 8560
rect 16212 8508 16264 8560
rect 6828 8372 6880 8424
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 7656 8372 7708 8424
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 8116 8372 8168 8381
rect 9404 8415 9456 8424
rect 9404 8381 9413 8415
rect 9413 8381 9447 8415
rect 9447 8381 9456 8415
rect 9404 8372 9456 8381
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 10048 8372 10100 8424
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 14372 8415 14424 8424
rect 12624 8372 12676 8381
rect 8484 8304 8536 8356
rect 10784 8304 10836 8356
rect 12532 8304 12584 8356
rect 13268 8347 13320 8356
rect 13268 8313 13277 8347
rect 13277 8313 13311 8347
rect 13311 8313 13320 8347
rect 13268 8304 13320 8313
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 14648 8415 14700 8424
rect 14648 8381 14657 8415
rect 14657 8381 14691 8415
rect 14691 8381 14700 8415
rect 14648 8372 14700 8381
rect 17684 8508 17736 8560
rect 20720 8508 20772 8560
rect 21640 8508 21692 8560
rect 22744 8576 22796 8628
rect 23388 8619 23440 8628
rect 23388 8585 23397 8619
rect 23397 8585 23431 8619
rect 23431 8585 23440 8619
rect 23388 8576 23440 8585
rect 19524 8440 19576 8492
rect 19708 8483 19760 8492
rect 19708 8449 19717 8483
rect 19717 8449 19751 8483
rect 19751 8449 19760 8483
rect 19708 8440 19760 8449
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 22836 8440 22888 8492
rect 18604 8372 18656 8424
rect 19156 8372 19208 8424
rect 19248 8372 19300 8424
rect 15292 8304 15344 8356
rect 15476 8304 15528 8356
rect 17500 8304 17552 8356
rect 5540 8279 5592 8288
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 5540 8236 5592 8245
rect 6460 8236 6512 8288
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 6644 8236 6696 8245
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 10048 8236 10100 8288
rect 11152 8236 11204 8288
rect 11520 8236 11572 8288
rect 11888 8279 11940 8288
rect 11888 8245 11897 8279
rect 11897 8245 11931 8279
rect 11931 8245 11940 8279
rect 11888 8236 11940 8245
rect 15108 8236 15160 8288
rect 16304 8236 16356 8288
rect 18144 8236 18196 8288
rect 21180 8304 21232 8356
rect 19340 8236 19392 8288
rect 20996 8236 21048 8288
rect 21640 8347 21692 8356
rect 21640 8313 21649 8347
rect 21649 8313 21683 8347
rect 21683 8313 21692 8347
rect 21640 8304 21692 8313
rect 24124 8304 24176 8356
rect 24216 8236 24268 8288
rect 24676 8236 24728 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 6920 8075 6972 8084
rect 6920 8041 6929 8075
rect 6929 8041 6963 8075
rect 6963 8041 6972 8075
rect 6920 8032 6972 8041
rect 7656 8032 7708 8084
rect 8024 7964 8076 8016
rect 10968 8032 11020 8084
rect 12072 8032 12124 8084
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 6000 7896 6052 7948
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 7380 7939 7432 7948
rect 7380 7905 7389 7939
rect 7389 7905 7423 7939
rect 7423 7905 7432 7939
rect 7380 7896 7432 7905
rect 7564 7896 7616 7948
rect 12992 7964 13044 8016
rect 15476 7964 15528 8016
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 11520 7939 11572 7948
rect 8116 7828 8168 7880
rect 11520 7905 11529 7939
rect 11529 7905 11563 7939
rect 11563 7905 11572 7939
rect 11520 7896 11572 7905
rect 11888 7939 11940 7948
rect 11888 7905 11897 7939
rect 11897 7905 11931 7939
rect 11931 7905 11940 7939
rect 11888 7896 11940 7905
rect 12072 7939 12124 7948
rect 12072 7905 12081 7939
rect 12081 7905 12115 7939
rect 12115 7905 12124 7939
rect 12072 7896 12124 7905
rect 13544 7896 13596 7948
rect 13912 7939 13964 7948
rect 13912 7905 13921 7939
rect 13921 7905 13955 7939
rect 13955 7905 13964 7939
rect 13912 7896 13964 7905
rect 21640 8032 21692 8084
rect 22744 8032 22796 8084
rect 16304 7964 16356 8016
rect 17500 7964 17552 8016
rect 20904 7964 20956 8016
rect 22560 7964 22612 8016
rect 22836 7964 22888 8016
rect 17408 7896 17460 7948
rect 14556 7828 14608 7880
rect 17684 7828 17736 7880
rect 17868 7871 17920 7880
rect 17868 7837 17877 7871
rect 17877 7837 17911 7871
rect 17911 7837 17920 7871
rect 17868 7828 17920 7837
rect 18972 7896 19024 7948
rect 19248 7896 19300 7948
rect 22468 7896 22520 7948
rect 23020 7896 23072 7948
rect 9772 7803 9824 7812
rect 9772 7769 9781 7803
rect 9781 7769 9815 7803
rect 9815 7769 9824 7803
rect 9772 7760 9824 7769
rect 9864 7760 9916 7812
rect 14372 7760 14424 7812
rect 15936 7760 15988 7812
rect 19156 7760 19208 7812
rect 6184 7692 6236 7744
rect 6460 7692 6512 7744
rect 7380 7692 7432 7744
rect 8668 7692 8720 7744
rect 10784 7692 10836 7744
rect 13912 7692 13964 7744
rect 17316 7692 17368 7744
rect 20260 7735 20312 7744
rect 20260 7701 20269 7735
rect 20269 7701 20303 7735
rect 20303 7701 20312 7735
rect 20260 7692 20312 7701
rect 21916 7828 21968 7880
rect 24676 7828 24728 7880
rect 23664 7760 23716 7812
rect 22836 7735 22888 7744
rect 22836 7701 22845 7735
rect 22845 7701 22879 7735
rect 22879 7701 22888 7735
rect 22836 7692 22888 7701
rect 22928 7692 22980 7744
rect 23848 7735 23900 7744
rect 23848 7701 23857 7735
rect 23857 7701 23891 7735
rect 23891 7701 23900 7735
rect 23848 7692 23900 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 6000 7488 6052 7540
rect 7564 7488 7616 7540
rect 7748 7488 7800 7540
rect 9680 7488 9732 7540
rect 9864 7488 9916 7540
rect 11520 7488 11572 7540
rect 13912 7531 13964 7540
rect 13912 7497 13921 7531
rect 13921 7497 13955 7531
rect 13955 7497 13964 7531
rect 13912 7488 13964 7497
rect 14464 7488 14516 7540
rect 16304 7531 16356 7540
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 18144 7488 18196 7540
rect 18972 7488 19024 7540
rect 20076 7488 20128 7540
rect 21824 7488 21876 7540
rect 22560 7531 22612 7540
rect 22560 7497 22569 7531
rect 22569 7497 22603 7531
rect 22603 7497 22612 7531
rect 22560 7488 22612 7497
rect 23020 7531 23072 7540
rect 23020 7497 23029 7531
rect 23029 7497 23063 7531
rect 23063 7497 23072 7531
rect 23020 7488 23072 7497
rect 25780 7531 25832 7540
rect 25780 7497 25789 7531
rect 25789 7497 25823 7531
rect 25823 7497 25832 7531
rect 25780 7488 25832 7497
rect 6184 7420 6236 7472
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 10692 7352 10744 7404
rect 10784 7352 10836 7404
rect 12072 7352 12124 7404
rect 12992 7420 13044 7472
rect 13268 7420 13320 7472
rect 15476 7420 15528 7472
rect 17500 7420 17552 7472
rect 19248 7420 19300 7472
rect 22192 7463 22244 7472
rect 22192 7429 22201 7463
rect 22201 7429 22235 7463
rect 22235 7429 22244 7463
rect 22192 7420 22244 7429
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 3424 7284 3476 7336
rect 6644 7327 6696 7336
rect 6644 7293 6653 7327
rect 6653 7293 6687 7327
rect 6687 7293 6696 7327
rect 6644 7284 6696 7293
rect 8024 7284 8076 7336
rect 9404 7327 9456 7336
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 9404 7284 9456 7293
rect 12348 7284 12400 7336
rect 14464 7284 14516 7336
rect 14832 7284 14884 7336
rect 18236 7352 18288 7404
rect 20720 7352 20772 7404
rect 22928 7352 22980 7404
rect 23756 7395 23808 7404
rect 23756 7361 23765 7395
rect 23765 7361 23799 7395
rect 23799 7361 23808 7395
rect 23756 7352 23808 7361
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 15660 7284 15712 7336
rect 15936 7327 15988 7336
rect 15936 7293 15945 7327
rect 15945 7293 15979 7327
rect 15979 7293 15988 7327
rect 15936 7284 15988 7293
rect 16672 7284 16724 7336
rect 17040 7284 17092 7336
rect 19984 7327 20036 7336
rect 19984 7293 19993 7327
rect 19993 7293 20027 7327
rect 20027 7293 20036 7327
rect 19984 7284 20036 7293
rect 20260 7284 20312 7336
rect 20628 7327 20680 7336
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 20628 7284 20680 7293
rect 22560 7284 22612 7336
rect 23296 7284 23348 7336
rect 23664 7327 23716 7336
rect 23664 7293 23673 7327
rect 23673 7293 23707 7327
rect 23707 7293 23716 7327
rect 23664 7284 23716 7293
rect 23848 7284 23900 7336
rect 25780 7284 25832 7336
rect 4896 7148 4948 7200
rect 6460 7148 6512 7200
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 7840 7191 7892 7200
rect 7840 7157 7849 7191
rect 7849 7157 7883 7191
rect 7883 7157 7892 7191
rect 7840 7148 7892 7157
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 12440 7148 12492 7200
rect 15660 7148 15712 7200
rect 16856 7148 16908 7200
rect 18512 7259 18564 7268
rect 18512 7225 18521 7259
rect 18521 7225 18555 7259
rect 18555 7225 18564 7259
rect 18512 7216 18564 7225
rect 21824 7216 21876 7268
rect 19984 7148 20036 7200
rect 21088 7148 21140 7200
rect 24676 7191 24728 7200
rect 24676 7157 24685 7191
rect 24685 7157 24719 7191
rect 24719 7157 24728 7191
rect 24676 7148 24728 7157
rect 24768 7148 24820 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 6920 6944 6972 6996
rect 8116 6944 8168 6996
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 4896 6876 4948 6928
rect 5172 6919 5224 6928
rect 5172 6885 5181 6919
rect 5181 6885 5215 6919
rect 5215 6885 5224 6919
rect 6736 6919 6788 6928
rect 5172 6876 5224 6885
rect 6736 6885 6745 6919
rect 6745 6885 6779 6919
rect 6779 6885 6788 6919
rect 6736 6876 6788 6885
rect 9680 6944 9732 6996
rect 9956 6944 10008 6996
rect 10692 6944 10744 6996
rect 11888 6987 11940 6996
rect 11888 6953 11897 6987
rect 11897 6953 11931 6987
rect 11931 6953 11940 6987
rect 11888 6944 11940 6953
rect 12348 6944 12400 6996
rect 16856 6987 16908 6996
rect 8208 6808 8260 6860
rect 4068 6740 4120 6792
rect 6000 6740 6052 6792
rect 6644 6783 6696 6792
rect 6644 6749 6653 6783
rect 6653 6749 6687 6783
rect 6687 6749 6696 6783
rect 6644 6740 6696 6749
rect 7196 6715 7248 6724
rect 7196 6681 7205 6715
rect 7205 6681 7239 6715
rect 7239 6681 7248 6715
rect 7196 6672 7248 6681
rect 9864 6876 9916 6928
rect 12256 6876 12308 6928
rect 12992 6919 13044 6928
rect 12992 6885 13001 6919
rect 13001 6885 13035 6919
rect 13035 6885 13044 6919
rect 12992 6876 13044 6885
rect 9772 6808 9824 6860
rect 10416 6851 10468 6860
rect 10416 6817 10425 6851
rect 10425 6817 10459 6851
rect 10459 6817 10468 6851
rect 10416 6808 10468 6817
rect 10692 6851 10744 6860
rect 10692 6817 10701 6851
rect 10701 6817 10735 6851
rect 10735 6817 10744 6851
rect 10692 6808 10744 6817
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 10048 6740 10100 6792
rect 11520 6740 11572 6792
rect 12716 6783 12768 6792
rect 12716 6749 12725 6783
rect 12725 6749 12759 6783
rect 12759 6749 12768 6783
rect 12716 6740 12768 6749
rect 16856 6953 16865 6987
rect 16865 6953 16899 6987
rect 16899 6953 16908 6987
rect 16856 6944 16908 6953
rect 17408 6987 17460 6996
rect 17408 6953 17417 6987
rect 17417 6953 17451 6987
rect 17451 6953 17460 6987
rect 17408 6944 17460 6953
rect 18144 6987 18196 6996
rect 18144 6953 18153 6987
rect 18153 6953 18187 6987
rect 18187 6953 18196 6987
rect 18144 6944 18196 6953
rect 18512 6944 18564 6996
rect 19524 6987 19576 6996
rect 19524 6953 19533 6987
rect 19533 6953 19567 6987
rect 19567 6953 19576 6987
rect 19524 6944 19576 6953
rect 20720 6987 20772 6996
rect 20720 6953 20729 6987
rect 20729 6953 20763 6987
rect 20763 6953 20772 6987
rect 20720 6944 20772 6953
rect 20996 6987 21048 6996
rect 20996 6953 21005 6987
rect 21005 6953 21039 6987
rect 21039 6953 21048 6987
rect 20996 6944 21048 6953
rect 22836 6944 22888 6996
rect 14556 6876 14608 6928
rect 17040 6876 17092 6928
rect 19156 6919 19208 6928
rect 19156 6885 19165 6919
rect 19165 6885 19199 6919
rect 19199 6885 19208 6919
rect 19156 6876 19208 6885
rect 22192 6919 22244 6928
rect 22192 6885 22201 6919
rect 22201 6885 22235 6919
rect 22235 6885 22244 6919
rect 22192 6876 22244 6885
rect 24032 6876 24084 6928
rect 13544 6808 13596 6860
rect 13728 6808 13780 6860
rect 15384 6851 15436 6860
rect 15384 6817 15393 6851
rect 15393 6817 15427 6851
rect 15427 6817 15436 6851
rect 15384 6808 15436 6817
rect 15660 6851 15712 6860
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 17868 6808 17920 6860
rect 19616 6808 19668 6860
rect 25228 6808 25280 6860
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 21272 6740 21324 6792
rect 22100 6783 22152 6792
rect 22100 6749 22109 6783
rect 22109 6749 22143 6783
rect 22143 6749 22152 6783
rect 22100 6740 22152 6749
rect 23664 6783 23716 6792
rect 16580 6672 16632 6724
rect 23664 6749 23673 6783
rect 23673 6749 23707 6783
rect 23707 6749 23716 6783
rect 23664 6740 23716 6749
rect 23020 6672 23072 6724
rect 4896 6647 4948 6656
rect 4896 6613 4905 6647
rect 4905 6613 4939 6647
rect 4939 6613 4948 6647
rect 4896 6604 4948 6613
rect 6828 6604 6880 6656
rect 7288 6604 7340 6656
rect 8116 6604 8168 6656
rect 11244 6604 11296 6656
rect 13544 6604 13596 6656
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 21456 6604 21508 6656
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1400 6400 1452 6452
rect 1952 6400 2004 6452
rect 4068 6443 4120 6452
rect 4068 6409 4077 6443
rect 4077 6409 4111 6443
rect 4111 6409 4120 6443
rect 4068 6400 4120 6409
rect 5172 6400 5224 6452
rect 6736 6400 6788 6452
rect 8300 6400 8352 6452
rect 9128 6332 9180 6384
rect 9220 6375 9272 6384
rect 9220 6341 9229 6375
rect 9229 6341 9263 6375
rect 9263 6341 9272 6375
rect 9220 6332 9272 6341
rect 4896 6264 4948 6316
rect 7380 6264 7432 6316
rect 10048 6196 10100 6248
rect 10416 6332 10468 6384
rect 11888 6332 11940 6384
rect 15476 6400 15528 6452
rect 18696 6400 18748 6452
rect 23112 6400 23164 6452
rect 23664 6400 23716 6452
rect 24768 6443 24820 6452
rect 24768 6409 24777 6443
rect 24777 6409 24811 6443
rect 24811 6409 24820 6443
rect 24768 6400 24820 6409
rect 25228 6443 25280 6452
rect 25228 6409 25237 6443
rect 25237 6409 25271 6443
rect 25271 6409 25280 6443
rect 25228 6400 25280 6409
rect 27620 6400 27672 6452
rect 15384 6332 15436 6384
rect 19524 6332 19576 6384
rect 22192 6332 22244 6384
rect 24400 6332 24452 6384
rect 11520 6264 11572 6316
rect 12808 6307 12860 6316
rect 12808 6273 12817 6307
rect 12817 6273 12851 6307
rect 12851 6273 12860 6307
rect 12808 6264 12860 6273
rect 13176 6264 13228 6316
rect 16856 6264 16908 6316
rect 21640 6307 21692 6316
rect 21640 6273 21649 6307
rect 21649 6273 21683 6307
rect 21683 6273 21692 6307
rect 21640 6264 21692 6273
rect 10692 6196 10744 6248
rect 11244 6196 11296 6248
rect 17684 6196 17736 6248
rect 20260 6196 20312 6248
rect 5356 6171 5408 6180
rect 5356 6137 5365 6171
rect 5365 6137 5399 6171
rect 5399 6137 5408 6171
rect 5356 6128 5408 6137
rect 5908 6171 5960 6180
rect 5908 6137 5917 6171
rect 5917 6137 5951 6171
rect 5951 6137 5960 6171
rect 5908 6128 5960 6137
rect 7196 6171 7248 6180
rect 2228 6103 2280 6112
rect 2228 6069 2237 6103
rect 2237 6069 2271 6103
rect 2271 6069 2280 6103
rect 2228 6060 2280 6069
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 7196 6137 7205 6171
rect 7205 6137 7239 6171
rect 7239 6137 7248 6171
rect 7196 6128 7248 6137
rect 7932 6128 7984 6180
rect 8760 6128 8812 6180
rect 10876 6128 10928 6180
rect 12256 6128 12308 6180
rect 12532 6171 12584 6180
rect 12532 6137 12541 6171
rect 12541 6137 12575 6171
rect 12575 6137 12584 6171
rect 12532 6128 12584 6137
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 8576 6103 8628 6112
rect 8576 6069 8585 6103
rect 8585 6069 8619 6103
rect 8619 6069 8628 6103
rect 8576 6060 8628 6069
rect 9956 6103 10008 6112
rect 9956 6069 9965 6103
rect 9965 6069 9999 6103
rect 9999 6069 10008 6103
rect 9956 6060 10008 6069
rect 10692 6060 10744 6112
rect 12072 6060 12124 6112
rect 13912 6128 13964 6180
rect 13728 6103 13780 6112
rect 13728 6069 13737 6103
rect 13737 6069 13771 6103
rect 13771 6069 13780 6103
rect 13728 6060 13780 6069
rect 14188 6171 14240 6180
rect 14188 6137 14197 6171
rect 14197 6137 14231 6171
rect 14231 6137 14240 6171
rect 14188 6128 14240 6137
rect 16580 6171 16632 6180
rect 16580 6137 16589 6171
rect 16589 6137 16623 6171
rect 16623 6137 16632 6171
rect 16580 6128 16632 6137
rect 18236 6128 18288 6180
rect 14556 6060 14608 6112
rect 15384 6103 15436 6112
rect 15384 6069 15393 6103
rect 15393 6069 15427 6103
rect 15427 6069 15436 6103
rect 15384 6060 15436 6069
rect 15660 6060 15712 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 18144 6060 18196 6112
rect 19984 6128 20036 6180
rect 22284 6171 22336 6180
rect 18972 6103 19024 6112
rect 18972 6069 18981 6103
rect 18981 6069 19015 6103
rect 19015 6069 19024 6103
rect 18972 6060 19024 6069
rect 19524 6060 19576 6112
rect 22284 6137 22293 6171
rect 22293 6137 22327 6171
rect 22327 6137 22336 6171
rect 22284 6128 22336 6137
rect 24032 6128 24084 6180
rect 24860 6128 24912 6180
rect 21824 6060 21876 6112
rect 23112 6103 23164 6112
rect 23112 6069 23121 6103
rect 23121 6069 23155 6103
rect 23155 6069 23164 6103
rect 23112 6060 23164 6069
rect 23388 6103 23440 6112
rect 23388 6069 23397 6103
rect 23397 6069 23431 6103
rect 23431 6069 23440 6103
rect 23388 6060 23440 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 6644 5899 6696 5908
rect 6644 5865 6653 5899
rect 6653 5865 6687 5899
rect 6687 5865 6696 5899
rect 6644 5856 6696 5865
rect 7932 5856 7984 5908
rect 8116 5899 8168 5908
rect 8116 5865 8125 5899
rect 8125 5865 8159 5899
rect 8159 5865 8168 5899
rect 8116 5856 8168 5865
rect 8576 5856 8628 5908
rect 9772 5856 9824 5908
rect 10048 5856 10100 5908
rect 11520 5899 11572 5908
rect 11520 5865 11529 5899
rect 11529 5865 11563 5899
rect 11563 5865 11572 5899
rect 11520 5856 11572 5865
rect 12532 5856 12584 5908
rect 17040 5899 17092 5908
rect 6736 5788 6788 5840
rect 7104 5788 7156 5840
rect 9864 5788 9916 5840
rect 11060 5788 11112 5840
rect 12164 5831 12216 5840
rect 12164 5797 12173 5831
rect 12173 5797 12207 5831
rect 12207 5797 12216 5831
rect 12164 5788 12216 5797
rect 12256 5788 12308 5840
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 4528 5720 4580 5772
rect 5356 5720 5408 5772
rect 6276 5720 6328 5772
rect 8392 5720 8444 5772
rect 9956 5720 10008 5772
rect 13636 5763 13688 5772
rect 13636 5729 13645 5763
rect 13645 5729 13679 5763
rect 13679 5729 13688 5763
rect 13636 5720 13688 5729
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 17040 5865 17049 5899
rect 17049 5865 17083 5899
rect 17083 5865 17092 5899
rect 17040 5856 17092 5865
rect 17408 5856 17460 5908
rect 21824 5899 21876 5908
rect 17684 5788 17736 5840
rect 21824 5865 21833 5899
rect 21833 5865 21867 5899
rect 21867 5865 21876 5899
rect 21824 5856 21876 5865
rect 22100 5899 22152 5908
rect 22100 5865 22109 5899
rect 22109 5865 22143 5899
rect 22143 5865 22152 5899
rect 22100 5856 22152 5865
rect 23112 5856 23164 5908
rect 24032 5899 24084 5908
rect 24032 5865 24041 5899
rect 24041 5865 24075 5899
rect 24075 5865 24084 5899
rect 24032 5856 24084 5865
rect 18972 5788 19024 5840
rect 19432 5831 19484 5840
rect 19432 5797 19441 5831
rect 19441 5797 19475 5831
rect 19475 5797 19484 5831
rect 19432 5788 19484 5797
rect 19984 5788 20036 5840
rect 21456 5788 21508 5840
rect 22744 5831 22796 5840
rect 22744 5797 22753 5831
rect 22753 5797 22787 5831
rect 22787 5797 22796 5831
rect 22744 5788 22796 5797
rect 22836 5831 22888 5840
rect 22836 5797 22845 5831
rect 22845 5797 22879 5831
rect 22879 5797 22888 5831
rect 24400 5831 24452 5840
rect 22836 5788 22888 5797
rect 24400 5797 24409 5831
rect 24409 5797 24443 5831
rect 24443 5797 24452 5831
rect 24400 5788 24452 5797
rect 24676 5788 24728 5840
rect 20628 5720 20680 5772
rect 5908 5652 5960 5704
rect 7380 5695 7432 5704
rect 1584 5627 1636 5636
rect 1584 5593 1593 5627
rect 1593 5593 1627 5627
rect 1627 5593 1636 5627
rect 1584 5584 1636 5593
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 13176 5652 13228 5704
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 18236 5652 18288 5704
rect 7932 5584 7984 5636
rect 11336 5584 11388 5636
rect 5080 5516 5132 5568
rect 11152 5559 11204 5568
rect 11152 5525 11161 5559
rect 11161 5525 11195 5559
rect 11195 5525 11204 5559
rect 11152 5516 11204 5525
rect 12532 5516 12584 5568
rect 12716 5584 12768 5636
rect 17868 5584 17920 5636
rect 18328 5584 18380 5636
rect 22284 5652 22336 5704
rect 23020 5695 23072 5704
rect 23020 5661 23029 5695
rect 23029 5661 23063 5695
rect 23063 5661 23072 5695
rect 23020 5652 23072 5661
rect 25044 5652 25096 5704
rect 20720 5584 20772 5636
rect 22468 5584 22520 5636
rect 24860 5627 24912 5636
rect 24860 5593 24869 5627
rect 24869 5593 24903 5627
rect 24903 5593 24912 5627
rect 24860 5584 24912 5593
rect 13544 5516 13596 5568
rect 13912 5516 13964 5568
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 14740 5516 14792 5568
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 23848 5516 23900 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1400 5312 1452 5364
rect 7380 5312 7432 5364
rect 8392 5312 8444 5364
rect 9220 5312 9272 5364
rect 9680 5355 9732 5364
rect 9680 5321 9689 5355
rect 9689 5321 9723 5355
rect 9723 5321 9732 5355
rect 9680 5312 9732 5321
rect 11152 5312 11204 5364
rect 12164 5312 12216 5364
rect 13636 5312 13688 5364
rect 16120 5312 16172 5364
rect 19432 5355 19484 5364
rect 19432 5321 19441 5355
rect 19441 5321 19475 5355
rect 19475 5321 19484 5355
rect 19432 5312 19484 5321
rect 19984 5312 20036 5364
rect 22744 5312 22796 5364
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 25044 5355 25096 5364
rect 25044 5321 25053 5355
rect 25053 5321 25087 5355
rect 25087 5321 25096 5355
rect 25044 5312 25096 5321
rect 7196 5244 7248 5296
rect 6184 5176 6236 5228
rect 6276 5219 6328 5228
rect 6276 5185 6285 5219
rect 6285 5185 6319 5219
rect 6319 5185 6328 5219
rect 6276 5176 6328 5185
rect 4528 5151 4580 5160
rect 4528 5117 4537 5151
rect 4537 5117 4571 5151
rect 4571 5117 4580 5151
rect 4528 5108 4580 5117
rect 8116 5176 8168 5228
rect 9220 5108 9272 5160
rect 12440 5244 12492 5296
rect 12072 5176 12124 5228
rect 13176 5219 13228 5228
rect 13176 5185 13185 5219
rect 13185 5185 13219 5219
rect 13219 5185 13228 5219
rect 13176 5176 13228 5185
rect 17224 5244 17276 5296
rect 20352 5244 20404 5296
rect 23756 5287 23808 5296
rect 23756 5253 23765 5287
rect 23765 5253 23799 5287
rect 23799 5253 23808 5287
rect 23756 5244 23808 5253
rect 7840 5040 7892 5092
rect 9404 5040 9456 5092
rect 10968 5040 11020 5092
rect 12532 5083 12584 5092
rect 12532 5049 12541 5083
rect 12541 5049 12575 5083
rect 12575 5049 12584 5083
rect 12532 5040 12584 5049
rect 6644 5015 6696 5024
rect 6644 4981 6653 5015
rect 6653 4981 6687 5015
rect 6687 4981 6696 5015
rect 6644 4972 6696 4981
rect 7288 4972 7340 5024
rect 12440 4972 12492 5024
rect 14004 5108 14056 5160
rect 17500 5176 17552 5228
rect 18236 5176 18288 5228
rect 23388 5176 23440 5228
rect 23848 5176 23900 5228
rect 24124 5219 24176 5228
rect 17040 5108 17092 5160
rect 20444 5151 20496 5160
rect 20444 5117 20453 5151
rect 20453 5117 20487 5151
rect 20487 5117 20496 5151
rect 20444 5108 20496 5117
rect 16764 5040 16816 5092
rect 17316 5040 17368 5092
rect 18144 5083 18196 5092
rect 18144 5049 18153 5083
rect 18153 5049 18187 5083
rect 18187 5049 18196 5083
rect 18144 5040 18196 5049
rect 18420 5040 18472 5092
rect 22376 5108 22428 5160
rect 22836 5108 22888 5160
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 20904 5040 20956 5092
rect 27620 5108 27672 5160
rect 13728 4972 13780 5024
rect 16120 4972 16172 5024
rect 17408 4972 17460 5024
rect 19984 4972 20036 5024
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 21364 4972 21416 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1400 4768 1452 4820
rect 6644 4768 6696 4820
rect 7104 4768 7156 4820
rect 7932 4768 7984 4820
rect 9956 4768 10008 4820
rect 14832 4811 14884 4820
rect 7196 4743 7248 4752
rect 7196 4709 7205 4743
rect 7205 4709 7239 4743
rect 7239 4709 7248 4743
rect 7196 4700 7248 4709
rect 14832 4777 14841 4811
rect 14841 4777 14875 4811
rect 14875 4777 14884 4811
rect 14832 4768 14884 4777
rect 17316 4768 17368 4820
rect 17500 4811 17552 4820
rect 17500 4777 17509 4811
rect 17509 4777 17543 4811
rect 17543 4777 17552 4811
rect 17500 4768 17552 4777
rect 18144 4768 18196 4820
rect 20628 4768 20680 4820
rect 23756 4811 23808 4820
rect 23756 4777 23765 4811
rect 23765 4777 23799 4811
rect 23799 4777 23808 4811
rect 23756 4768 23808 4777
rect 10968 4743 11020 4752
rect 10968 4709 10977 4743
rect 10977 4709 11011 4743
rect 11011 4709 11020 4743
rect 10968 4700 11020 4709
rect 11520 4743 11572 4752
rect 11520 4709 11529 4743
rect 11529 4709 11563 4743
rect 11563 4709 11572 4743
rect 11520 4700 11572 4709
rect 13820 4743 13872 4752
rect 13820 4709 13829 4743
rect 13829 4709 13863 4743
rect 13863 4709 13872 4743
rect 13820 4700 13872 4709
rect 20444 4743 20496 4752
rect 20444 4709 20453 4743
rect 20453 4709 20487 4743
rect 20487 4709 20496 4743
rect 20444 4700 20496 4709
rect 22376 4743 22428 4752
rect 22376 4709 22385 4743
rect 22385 4709 22419 4743
rect 22419 4709 22428 4743
rect 22376 4700 22428 4709
rect 6184 4632 6236 4684
rect 9404 4632 9456 4684
rect 9588 4632 9640 4684
rect 9680 4632 9732 4684
rect 12992 4675 13044 4684
rect 12992 4641 13001 4675
rect 13001 4641 13035 4675
rect 13035 4641 13044 4675
rect 12992 4632 13044 4641
rect 14556 4632 14608 4684
rect 15752 4632 15804 4684
rect 16764 4675 16816 4684
rect 16764 4641 16773 4675
rect 16773 4641 16807 4675
rect 16807 4641 16816 4675
rect 16764 4632 16816 4641
rect 18328 4632 18380 4684
rect 18604 4632 18656 4684
rect 19248 4675 19300 4684
rect 19248 4641 19257 4675
rect 19257 4641 19291 4675
rect 19291 4641 19300 4675
rect 19248 4632 19300 4641
rect 20168 4632 20220 4684
rect 7012 4564 7064 4616
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 12348 4607 12400 4616
rect 12348 4573 12357 4607
rect 12357 4573 12391 4607
rect 12391 4573 12400 4607
rect 12348 4564 12400 4573
rect 16304 4607 16356 4616
rect 16304 4573 16313 4607
rect 16313 4573 16347 4607
rect 16347 4573 16356 4607
rect 16304 4564 16356 4573
rect 17776 4564 17828 4616
rect 23020 4564 23072 4616
rect 6828 4471 6880 4480
rect 6828 4437 6837 4471
rect 6837 4437 6871 4471
rect 6871 4437 6880 4471
rect 6828 4428 6880 4437
rect 9036 4471 9088 4480
rect 9036 4437 9045 4471
rect 9045 4437 9079 4471
rect 9079 4437 9088 4471
rect 9036 4428 9088 4437
rect 10324 4471 10376 4480
rect 10324 4437 10333 4471
rect 10333 4437 10367 4471
rect 10367 4437 10376 4471
rect 10324 4428 10376 4437
rect 11336 4496 11388 4548
rect 14648 4496 14700 4548
rect 15292 4496 15344 4548
rect 22468 4496 22520 4548
rect 24860 4496 24912 4548
rect 12532 4428 12584 4480
rect 14280 4428 14332 4480
rect 17040 4428 17092 4480
rect 18144 4428 18196 4480
rect 18880 4428 18932 4480
rect 22652 4428 22704 4480
rect 23756 4428 23808 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 6184 4267 6236 4276
rect 6184 4233 6193 4267
rect 6193 4233 6227 4267
rect 6227 4233 6236 4267
rect 6184 4224 6236 4233
rect 11152 4224 11204 4276
rect 15752 4224 15804 4276
rect 16948 4224 17000 4276
rect 18328 4224 18380 4276
rect 19248 4267 19300 4276
rect 19248 4233 19257 4267
rect 19257 4233 19291 4267
rect 19291 4233 19300 4267
rect 19248 4224 19300 4233
rect 21364 4224 21416 4276
rect 22376 4224 22428 4276
rect 23020 4267 23072 4276
rect 23020 4233 23029 4267
rect 23029 4233 23063 4267
rect 23063 4233 23072 4267
rect 23020 4224 23072 4233
rect 12532 4156 12584 4208
rect 14740 4156 14792 4208
rect 6460 4088 6512 4140
rect 5816 4063 5868 4072
rect 3332 3884 3384 3936
rect 5816 4029 5825 4063
rect 5825 4029 5859 4063
rect 5859 4029 5868 4063
rect 5816 4020 5868 4029
rect 6828 4020 6880 4072
rect 7748 4063 7800 4072
rect 7748 4029 7757 4063
rect 7757 4029 7791 4063
rect 7791 4029 7800 4063
rect 7748 4020 7800 4029
rect 10324 4088 10376 4140
rect 9588 4020 9640 4072
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 10968 4088 11020 4140
rect 13636 4088 13688 4140
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 11244 4020 11296 4029
rect 14096 4063 14148 4072
rect 14096 4029 14105 4063
rect 14105 4029 14139 4063
rect 14139 4029 14148 4063
rect 14096 4020 14148 4029
rect 14280 4020 14332 4072
rect 14832 4020 14884 4072
rect 17868 4088 17920 4140
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 18512 4131 18564 4140
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 19984 4020 20036 4072
rect 20168 4156 20220 4208
rect 22284 4199 22336 4208
rect 22284 4165 22293 4199
rect 22293 4165 22327 4199
rect 22327 4165 22336 4199
rect 22284 4156 22336 4165
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 22468 4088 22520 4140
rect 10784 3952 10836 4004
rect 11336 3995 11388 4004
rect 11336 3961 11345 3995
rect 11345 3961 11379 3995
rect 11379 3961 11388 3995
rect 11336 3952 11388 3961
rect 12164 3952 12216 4004
rect 15568 3995 15620 4004
rect 6460 3884 6512 3936
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 8760 3884 8812 3936
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 12440 3884 12492 3936
rect 15568 3961 15577 3995
rect 15577 3961 15611 3995
rect 15611 3961 15620 3995
rect 15568 3952 15620 3961
rect 16488 3995 16540 4004
rect 16488 3961 16497 3995
rect 16497 3961 16531 3995
rect 16531 3961 16540 3995
rect 16488 3952 16540 3961
rect 17132 3995 17184 4004
rect 13544 3884 13596 3936
rect 16396 3884 16448 3936
rect 17132 3961 17141 3995
rect 17141 3961 17175 3995
rect 17175 3961 17184 3995
rect 17132 3952 17184 3961
rect 18420 3952 18472 4004
rect 17868 3884 17920 3936
rect 20904 3884 20956 3936
rect 21364 3884 21416 3936
rect 27620 3884 27672 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5816 3680 5868 3732
rect 8576 3680 8628 3732
rect 9588 3680 9640 3732
rect 9956 3723 10008 3732
rect 7748 3612 7800 3664
rect 8484 3612 8536 3664
rect 3700 3544 3752 3596
rect 5540 3544 5592 3596
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 6368 3544 6420 3596
rect 7196 3544 7248 3596
rect 7932 3587 7984 3596
rect 1584 3476 1636 3528
rect 7472 3476 7524 3528
rect 7932 3553 7941 3587
rect 7941 3553 7975 3587
rect 7975 3553 7984 3587
rect 7932 3544 7984 3553
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 11336 3680 11388 3732
rect 11520 3680 11572 3732
rect 12992 3723 13044 3732
rect 10784 3612 10836 3664
rect 12348 3612 12400 3664
rect 12992 3689 13001 3723
rect 13001 3689 13035 3723
rect 13035 3689 13044 3723
rect 12992 3680 13044 3689
rect 14556 3723 14608 3732
rect 14556 3689 14565 3723
rect 14565 3689 14599 3723
rect 14599 3689 14608 3723
rect 14556 3680 14608 3689
rect 18420 3723 18472 3732
rect 18420 3689 18429 3723
rect 18429 3689 18463 3723
rect 18463 3689 18472 3723
rect 18420 3680 18472 3689
rect 13268 3612 13320 3664
rect 13544 3655 13596 3664
rect 13544 3621 13553 3655
rect 13553 3621 13587 3655
rect 13587 3621 13596 3655
rect 13544 3612 13596 3621
rect 15844 3612 15896 3664
rect 16120 3612 16172 3664
rect 9312 3476 9364 3528
rect 10692 3544 10744 3596
rect 4620 3451 4672 3460
rect 4620 3417 4629 3451
rect 4629 3417 4663 3451
rect 4663 3417 4672 3451
rect 4620 3408 4672 3417
rect 6368 3408 6420 3460
rect 7748 3451 7800 3460
rect 7748 3417 7757 3451
rect 7757 3417 7791 3451
rect 7791 3417 7800 3451
rect 7748 3408 7800 3417
rect 8576 3408 8628 3460
rect 10140 3408 10192 3460
rect 11152 3544 11204 3596
rect 13636 3587 13688 3596
rect 13636 3553 13645 3587
rect 13645 3553 13679 3587
rect 13679 3553 13688 3587
rect 13636 3544 13688 3553
rect 16764 3612 16816 3664
rect 17224 3655 17276 3664
rect 17224 3621 17233 3655
rect 17233 3621 17267 3655
rect 17267 3621 17276 3655
rect 17224 3612 17276 3621
rect 20168 3680 20220 3732
rect 20352 3680 20404 3732
rect 22652 3612 22704 3664
rect 20904 3587 20956 3596
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 20996 3587 21048 3596
rect 20996 3553 21005 3587
rect 21005 3553 21039 3587
rect 21039 3553 21048 3587
rect 20996 3544 21048 3553
rect 21180 3587 21232 3596
rect 21180 3553 21189 3587
rect 21189 3553 21223 3587
rect 21223 3553 21232 3587
rect 22468 3587 22520 3596
rect 21180 3544 21232 3553
rect 22468 3553 22477 3587
rect 22477 3553 22511 3587
rect 22511 3553 22520 3587
rect 22468 3544 22520 3553
rect 23848 3544 23900 3596
rect 17132 3519 17184 3528
rect 11704 3408 11756 3460
rect 12808 3408 12860 3460
rect 5540 3383 5592 3392
rect 5540 3349 5549 3383
rect 5549 3349 5583 3383
rect 5583 3349 5592 3383
rect 5540 3340 5592 3349
rect 6552 3383 6604 3392
rect 6552 3349 6561 3383
rect 6561 3349 6595 3383
rect 6595 3349 6604 3383
rect 6552 3340 6604 3349
rect 9128 3383 9180 3392
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 12164 3340 12216 3392
rect 13452 3383 13504 3392
rect 13452 3349 13461 3383
rect 13461 3349 13495 3383
rect 13495 3349 13504 3383
rect 13452 3340 13504 3349
rect 17132 3485 17141 3519
rect 17141 3485 17175 3519
rect 17175 3485 17184 3519
rect 17132 3476 17184 3485
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 17776 3476 17828 3528
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 16488 3408 16540 3460
rect 15476 3340 15528 3392
rect 18144 3383 18196 3392
rect 18144 3349 18153 3383
rect 18153 3349 18187 3383
rect 18187 3349 18196 3383
rect 18144 3340 18196 3349
rect 18420 3340 18472 3392
rect 20076 3340 20128 3392
rect 21272 3408 21324 3460
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1676 3136 1728 3188
rect 3700 3179 3752 3188
rect 3700 3145 3709 3179
rect 3709 3145 3743 3179
rect 3743 3145 3752 3179
rect 3700 3136 3752 3145
rect 5264 3136 5316 3188
rect 6552 3179 6604 3188
rect 6552 3145 6561 3179
rect 6561 3145 6595 3179
rect 6595 3145 6604 3179
rect 6552 3136 6604 3145
rect 8484 3136 8536 3188
rect 9036 3068 9088 3120
rect 10140 3111 10192 3120
rect 112 3000 164 3052
rect 7380 3000 7432 3052
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 5540 2932 5592 2984
rect 7472 2975 7524 2984
rect 7472 2941 7481 2975
rect 7481 2941 7515 2975
rect 7515 2941 7524 2975
rect 7472 2932 7524 2941
rect 7932 3000 7984 3052
rect 8208 3043 8260 3052
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 10140 3077 10149 3111
rect 10149 3077 10183 3111
rect 10183 3077 10192 3111
rect 10140 3068 10192 3077
rect 10784 3068 10836 3120
rect 12348 3136 12400 3188
rect 12624 3136 12676 3188
rect 14280 3136 14332 3188
rect 16304 3179 16356 3188
rect 16304 3145 16313 3179
rect 16313 3145 16347 3179
rect 16347 3145 16356 3179
rect 16304 3136 16356 3145
rect 16580 3136 16632 3188
rect 17224 3136 17276 3188
rect 17592 3136 17644 3188
rect 20904 3179 20956 3188
rect 11336 3000 11388 3052
rect 12532 3043 12584 3052
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 12808 3043 12860 3052
rect 12808 3009 12817 3043
rect 12817 3009 12851 3043
rect 12851 3009 12860 3043
rect 12808 3000 12860 3009
rect 6184 2907 6236 2916
rect 6184 2873 6193 2907
rect 6193 2873 6227 2907
rect 6227 2873 6236 2907
rect 6184 2864 6236 2873
rect 9128 2864 9180 2916
rect 10784 2864 10836 2916
rect 4620 2839 4672 2848
rect 4620 2805 4629 2839
rect 4629 2805 4663 2839
rect 4663 2805 4672 2839
rect 4620 2796 4672 2805
rect 7932 2796 7984 2848
rect 8760 2796 8812 2848
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 12992 2864 13044 2916
rect 15476 3111 15528 3120
rect 15476 3077 15485 3111
rect 15485 3077 15519 3111
rect 15519 3077 15528 3111
rect 15476 3068 15528 3077
rect 13452 3000 13504 3052
rect 17408 3000 17460 3052
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 18512 3068 18564 3120
rect 20904 3145 20913 3179
rect 20913 3145 20947 3179
rect 20947 3145 20956 3179
rect 20904 3136 20956 3145
rect 23756 3136 23808 3188
rect 19984 3068 20036 3120
rect 20996 3068 21048 3120
rect 21272 3111 21324 3120
rect 21272 3077 21281 3111
rect 21281 3077 21315 3111
rect 21315 3077 21324 3111
rect 21272 3068 21324 3077
rect 19432 3000 19484 3052
rect 20076 3043 20128 3052
rect 14096 2975 14148 2984
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 14280 2932 14332 2984
rect 19616 2975 19668 2984
rect 14832 2864 14884 2916
rect 15016 2864 15068 2916
rect 16488 2864 16540 2916
rect 16580 2907 16632 2916
rect 16580 2873 16589 2907
rect 16589 2873 16623 2907
rect 16623 2873 16632 2907
rect 16580 2864 16632 2873
rect 18604 2864 18656 2916
rect 13912 2796 13964 2848
rect 15844 2839 15896 2848
rect 15844 2805 15853 2839
rect 15853 2805 15887 2839
rect 15887 2805 15896 2839
rect 15844 2796 15896 2805
rect 16672 2796 16724 2848
rect 19616 2941 19625 2975
rect 19625 2941 19659 2975
rect 19659 2941 19668 2975
rect 19616 2932 19668 2941
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 21088 3000 21140 3052
rect 20812 2932 20864 2984
rect 20904 2932 20956 2984
rect 21272 2932 21324 2984
rect 19432 2839 19484 2848
rect 19432 2805 19441 2839
rect 19441 2805 19475 2839
rect 19475 2805 19484 2839
rect 19432 2796 19484 2805
rect 19524 2796 19576 2848
rect 22468 2864 22520 2916
rect 22652 2839 22704 2848
rect 22652 2805 22661 2839
rect 22661 2805 22695 2839
rect 22695 2805 22704 2839
rect 22652 2796 22704 2805
rect 23848 2839 23900 2848
rect 23848 2805 23857 2839
rect 23857 2805 23891 2839
rect 23891 2805 23900 2839
rect 23848 2796 23900 2805
rect 26884 2796 26936 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 4344 2592 4396 2644
rect 4436 2592 4488 2644
rect 5356 2592 5408 2644
rect 13360 2592 13412 2644
rect 13636 2635 13688 2644
rect 13636 2601 13645 2635
rect 13645 2601 13679 2635
rect 13679 2601 13688 2635
rect 13636 2592 13688 2601
rect 6644 2524 6696 2576
rect 7380 2524 7432 2576
rect 7932 2567 7984 2576
rect 7932 2533 7941 2567
rect 7941 2533 7975 2567
rect 7975 2533 7984 2567
rect 8760 2567 8812 2576
rect 7932 2524 7984 2533
rect 8760 2533 8769 2567
rect 8769 2533 8803 2567
rect 8803 2533 8812 2567
rect 8760 2524 8812 2533
rect 6920 2499 6972 2508
rect 3240 2320 3292 2372
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 8300 2499 8352 2508
rect 8300 2465 8309 2499
rect 8309 2465 8343 2499
rect 8343 2465 8352 2499
rect 8300 2456 8352 2465
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 7472 2388 7524 2440
rect 7748 2388 7800 2440
rect 848 2252 900 2304
rect 7196 2252 7248 2304
rect 10968 2524 11020 2576
rect 9956 2456 10008 2508
rect 9772 2388 9824 2440
rect 12808 2567 12860 2576
rect 12808 2533 12817 2567
rect 12817 2533 12851 2567
rect 12851 2533 12860 2567
rect 15016 2592 15068 2644
rect 16396 2635 16448 2644
rect 16396 2601 16405 2635
rect 16405 2601 16439 2635
rect 16439 2601 16448 2635
rect 16396 2592 16448 2601
rect 18144 2592 18196 2644
rect 19984 2592 20036 2644
rect 20536 2635 20588 2644
rect 20536 2601 20545 2635
rect 20545 2601 20579 2635
rect 20579 2601 20588 2635
rect 20536 2592 20588 2601
rect 20904 2592 20956 2644
rect 14188 2567 14240 2576
rect 12808 2524 12860 2533
rect 12440 2499 12492 2508
rect 12440 2465 12449 2499
rect 12449 2465 12483 2499
rect 12483 2465 12492 2499
rect 12440 2456 12492 2465
rect 12808 2388 12860 2440
rect 14188 2533 14197 2567
rect 14197 2533 14231 2567
rect 14231 2533 14240 2567
rect 14188 2524 14240 2533
rect 13820 2456 13872 2508
rect 10876 2320 10928 2372
rect 10968 2320 11020 2372
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 15844 2524 15896 2576
rect 18604 2524 18656 2576
rect 15568 2456 15620 2508
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 22560 2524 22612 2576
rect 20812 2456 20864 2508
rect 21180 2456 21232 2508
rect 21732 2456 21784 2508
rect 22376 2456 22428 2508
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 16028 2320 16080 2372
rect 23020 2320 23072 2372
rect 26056 2320 26108 2372
rect 21456 2252 21508 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 1030 27520 1086 28000
rect 2792 27526 3096 27554
rect 1044 23474 1072 27520
rect 1490 25936 1546 25945
rect 1490 25871 1546 25880
rect 1398 23488 1454 23497
rect 1044 23446 1256 23474
rect 20 22432 72 22438
rect 20 22374 72 22380
rect 32 5273 60 22374
rect 110 13424 166 13433
rect 110 13359 166 13368
rect 124 12481 152 13359
rect 110 12472 166 12481
rect 110 12407 166 12416
rect 1228 12306 1256 23446
rect 1398 23423 1454 23432
rect 1412 22574 1440 23423
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 1504 18834 1532 25871
rect 1858 24712 1914 24721
rect 1858 24647 1914 24656
rect 1582 22264 1638 22273
rect 1582 22199 1638 22208
rect 1596 21690 1624 22199
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1582 21040 1638 21049
rect 1582 20975 1638 20984
rect 1596 19514 1624 20975
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1492 18828 1544 18834
rect 1492 18770 1544 18776
rect 1504 18426 1532 18770
rect 1492 18420 1544 18426
rect 1492 18362 1544 18368
rect 1872 18290 1900 24647
rect 2136 21344 2188 21350
rect 2136 21286 2188 21292
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1582 16416 1638 16425
rect 1582 16351 1638 16360
rect 1596 14618 1624 16351
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1582 14240 1638 14249
rect 1582 14175 1638 14184
rect 1596 13530 1624 14175
rect 1688 13734 1716 14418
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1688 13530 1716 13670
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1688 12850 1716 13330
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1688 12753 1716 12786
rect 1674 12744 1730 12753
rect 1674 12679 1730 12688
rect 1216 12300 1268 12306
rect 1216 12242 1268 12248
rect 1228 11898 1256 12242
rect 1216 11892 1268 11898
rect 1216 11834 1268 11840
rect 2148 10713 2176 21286
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2424 18086 2452 19110
rect 2412 18080 2464 18086
rect 2412 18022 2464 18028
rect 2792 13462 2820 27526
rect 3068 27418 3096 27526
rect 3146 27520 3202 28000
rect 5262 27520 5318 28000
rect 7470 27520 7526 28000
rect 8300 27532 8352 27538
rect 3160 27418 3188 27520
rect 3068 27390 3188 27418
rect 5276 23322 5304 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 7484 23866 7512 27520
rect 9586 27532 9642 28000
rect 9586 27520 9588 27532
rect 8300 27474 8352 27480
rect 9640 27520 9642 27532
rect 11060 27532 11112 27538
rect 9588 27474 9640 27480
rect 11702 27532 11758 28000
rect 11702 27520 11704 27532
rect 11060 27474 11112 27480
rect 11756 27520 11758 27532
rect 13910 27520 13966 28000
rect 15752 27532 15804 27538
rect 11704 27474 11756 27480
rect 7472 23860 7524 23866
rect 7472 23802 7524 23808
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 5264 23316 5316 23322
rect 5264 23258 5316 23264
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5998 19408 6054 19417
rect 5998 19343 6054 19352
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 3422 17504 3478 17513
rect 3422 17439 3478 17448
rect 2780 13456 2832 13462
rect 2780 13398 2832 13404
rect 2134 10704 2190 10713
rect 2134 10639 2190 10648
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1596 8090 1624 8191
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1582 7168 1638 7177
rect 1582 7103 1638 7112
rect 1596 7002 1624 7103
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 6458 1440 6802
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1582 5944 1638 5953
rect 1582 5879 1638 5888
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5370 1440 5714
rect 1596 5642 1624 5879
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 18 5264 74 5273
rect 18 5199 74 5208
rect 1412 4826 1440 5306
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 112 3052 164 3058
rect 112 2994 164 3000
rect 124 2961 152 2994
rect 110 2952 166 2961
rect 110 2887 166 2896
rect 848 2304 900 2310
rect 848 2246 900 2252
rect 570 82 626 480
rect 860 82 888 2246
rect 570 54 888 82
rect 1596 82 1624 3470
rect 1688 3194 1716 9522
rect 3436 7342 3464 17439
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5552 12714 5580 13330
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5080 11688 5132 11694
rect 4250 11656 4306 11665
rect 5080 11630 5132 11636
rect 4250 11591 4306 11600
rect 4264 11218 4292 11591
rect 5092 11286 5120 11630
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4264 10810 4292 11154
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4724 10810 4752 11086
rect 5092 10810 5120 11222
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4080 6458 4108 6734
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 1964 5914 1992 6394
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2240 5681 2268 6054
rect 2226 5672 2282 5681
rect 2226 5607 2282 5616
rect 4066 4040 4122 4049
rect 4066 3975 4122 3984
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 3146 2408 3202 2417
rect 3240 2372 3292 2378
rect 3202 2352 3240 2360
rect 3146 2343 3240 2352
rect 3160 2332 3240 2343
rect 3240 2314 3292 2320
rect 1766 82 1822 480
rect 1596 54 1822 82
rect 570 0 626 54
rect 1766 0 1822 54
rect 3054 82 3110 480
rect 3344 82 3372 3878
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3712 3194 3740 3538
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 4080 2990 4108 3975
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4448 2650 4476 9930
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 9178 5948 9318
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5092 8634 5120 8978
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5184 8566 5212 8978
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5552 8294 5580 8842
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 6012 7954 6040 19343
rect 6932 12986 6960 23598
rect 8022 19000 8078 19009
rect 8022 18935 8078 18944
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7944 18426 7972 18770
rect 8036 18698 8064 18935
rect 8312 18834 8340 27474
rect 9600 27443 9628 27474
rect 9586 26888 9642 26897
rect 9586 26823 9642 26832
rect 9600 23662 9628 26823
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 9588 23656 9640 23662
rect 9588 23598 9640 23604
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 9404 23520 9456 23526
rect 9404 23462 9456 23468
rect 10048 23520 10100 23526
rect 10048 23462 10100 23468
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8024 18692 8076 18698
rect 8024 18634 8076 18640
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 8312 17105 8340 18566
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8956 18193 8984 18226
rect 8942 18184 8998 18193
rect 8942 18119 8998 18128
rect 9416 17814 9444 23462
rect 10060 23322 10088 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10888 23322 10916 23598
rect 10048 23316 10100 23322
rect 10048 23258 10100 23264
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10796 22438 10824 22918
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 9954 19816 10010 19825
rect 9954 19751 10010 19760
rect 9968 18970 9996 19751
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9876 18086 9904 18770
rect 10888 18086 10916 18838
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 9404 17808 9456 17814
rect 9310 17776 9366 17785
rect 9404 17750 9456 17756
rect 9310 17711 9366 17720
rect 8298 17096 8354 17105
rect 8298 17031 8354 17040
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 14074 7328 14214
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7300 13802 7328 14010
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 7208 12918 7236 13738
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7392 12986 7420 13330
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6090 11656 6146 11665
rect 6196 11626 6224 12310
rect 6288 12238 6316 12582
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6090 11591 6146 11600
rect 6184 11620 6236 11626
rect 6104 9110 6132 11591
rect 6184 11562 6236 11568
rect 6196 10810 6224 11562
rect 6288 11354 6316 12174
rect 6932 11626 6960 12174
rect 7208 11762 7236 12718
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6564 10674 6592 11494
rect 6932 11286 6960 11562
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6288 10266 6316 10406
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6288 9722 6316 10202
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6472 9178 6500 9998
rect 7024 9722 7052 11222
rect 7208 11150 7236 11698
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7484 11082 7512 12106
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7484 10742 7512 11018
rect 7472 10736 7524 10742
rect 7668 10713 7696 15982
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8220 15638 8248 15846
rect 8208 15632 8260 15638
rect 8128 15592 8208 15620
rect 8128 15162 8156 15592
rect 8208 15574 8260 15580
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 8036 13802 8064 14826
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 8128 13734 8156 14418
rect 8220 14278 8248 15438
rect 8312 15026 8340 15438
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8312 13938 8340 14962
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8956 14550 8984 14758
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8208 13864 8260 13870
rect 8864 13841 8892 13874
rect 9140 13870 9168 14418
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9128 13864 9180 13870
rect 8208 13806 8260 13812
rect 8850 13832 8906 13841
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12850 7788 13126
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 7852 11898 7880 12310
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7472 10678 7524 10684
rect 7654 10704 7710 10713
rect 7484 10266 7512 10678
rect 7654 10639 7710 10648
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7300 9654 7328 10202
rect 7852 10130 7880 11834
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7944 10810 7972 11494
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 8128 9926 8156 13670
rect 8220 12782 8248 13806
rect 9128 13806 9180 13812
rect 8850 13767 8906 13776
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8312 12986 8340 13330
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8404 12782 8432 13330
rect 9140 13190 9168 13806
rect 9232 13462 9260 14214
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8404 12442 8432 12718
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11898 8248 12174
rect 8496 12170 8524 12650
rect 9034 12472 9090 12481
rect 9034 12407 9090 12416
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8220 11354 8248 11834
rect 8588 11801 8616 12038
rect 9048 11830 9076 12407
rect 9036 11824 9088 11830
rect 8574 11792 8630 11801
rect 9036 11766 9088 11772
rect 8574 11727 8630 11736
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8390 10704 8446 10713
rect 8496 10674 8524 11154
rect 8390 10639 8446 10648
rect 8484 10668 8536 10674
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7300 9450 7328 9590
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8430 6868 8978
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6012 7546 6040 7890
rect 6472 7750 6500 8230
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6196 7478 6224 7686
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6472 7206 6500 7686
rect 6656 7342 6684 8230
rect 6840 7954 6868 8366
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 4908 6934 4936 7142
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 6322 4936 6598
rect 5184 6458 5212 6870
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5908 6180 5960 6186
rect 6012 6168 6040 6734
rect 5960 6140 6040 6168
rect 5908 6122 5960 6128
rect 5368 5778 5396 6122
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 4540 5273 4568 5714
rect 5920 5710 5948 6122
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4526 5264 4582 5273
rect 4526 5199 4582 5208
rect 4540 5166 4568 5199
rect 4528 5160 4580 5166
rect 5092 5137 5120 5510
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6196 5234 6224 6054
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6288 5234 6316 5714
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 4528 5102 4580 5108
rect 5078 5128 5134 5137
rect 5078 5063 5134 5072
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6196 4282 6224 4626
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6472 4146 6500 7142
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6656 5914 6684 6734
rect 6748 6458 6776 6870
rect 6840 6662 6868 7890
rect 6932 7410 6960 8026
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6932 7002 6960 7346
rect 7300 7206 7328 9386
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7392 8430 7420 8978
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 7954 7420 8366
rect 7576 7954 7604 8570
rect 7668 8430 7696 8978
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7668 8090 7696 8366
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 8036 8022 8064 8978
rect 8128 8566 8156 9318
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7392 7750 7420 7890
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7576 7546 7604 7890
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6748 5846 6776 6394
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4826 6684 4966
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6840 4486 6868 6598
rect 7208 6186 7236 6666
rect 7300 6662 7328 7142
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 7116 4826 7144 5782
rect 7208 5302 7236 6122
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7300 5030 7328 6598
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7392 5710 7420 6258
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7392 5370 7420 5646
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7196 4752 7248 4758
rect 7300 4740 7328 4966
rect 7248 4712 7328 4740
rect 7196 4694 7248 4700
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5828 3738 5856 4014
rect 6472 3942 6500 4082
rect 6840 4078 6868 4422
rect 6828 4072 6880 4078
rect 6826 4040 6828 4049
rect 6880 4040 6882 4049
rect 6826 3975 6882 3984
rect 7024 3942 7052 4558
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4632 2854 4660 3402
rect 5552 3398 5580 3538
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4356 2553 4384 2586
rect 4342 2544 4398 2553
rect 4342 2479 4398 2488
rect 3054 54 3372 82
rect 4342 82 4398 480
rect 4632 82 4660 2790
rect 5276 2446 5304 3130
rect 5552 2990 5580 3334
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 6196 2922 6224 3538
rect 6380 3466 6408 3538
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6184 2916 6236 2922
rect 6184 2858 6236 2864
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 4342 54 4660 82
rect 5368 82 5396 2586
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6472 2009 6500 3878
rect 7208 3602 7236 4694
rect 7760 4078 7788 7482
rect 8036 7342 8064 7958
rect 8128 7886 8156 8366
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7852 5098 7880 7142
rect 8128 7002 8156 7822
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7944 5914 7972 6122
rect 8128 5914 8156 6598
rect 8220 6118 8248 6802
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7944 4826 7972 5578
rect 8128 5234 8156 5850
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8220 4457 8248 6054
rect 8206 4448 8262 4457
rect 8206 4383 8262 4392
rect 8312 4154 8340 6394
rect 8404 5778 8432 10639
rect 8484 10610 8536 10616
rect 8496 10577 8524 10610
rect 8482 10568 8538 10577
rect 8482 10503 8538 10512
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9048 9586 9076 10406
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8404 5370 8432 5714
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8390 4312 8446 4321
rect 8390 4247 8446 4256
rect 8220 4126 8340 4154
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7760 3670 7788 4014
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6564 3194 6592 3334
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6918 2544 6974 2553
rect 6458 2000 6514 2009
rect 6458 1935 6514 1944
rect 5630 82 5686 480
rect 5368 54 5686 82
rect 6656 82 6684 2518
rect 6918 2479 6920 2488
rect 6972 2479 6974 2488
rect 6920 2450 6972 2456
rect 6932 2009 6960 2450
rect 7208 2310 7236 3538
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7392 2582 7420 2994
rect 7484 2990 7512 3470
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 7484 2446 7512 2926
rect 7760 2446 7788 3402
rect 7944 3058 7972 3538
rect 8220 3058 8248 4126
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7944 2582 7972 2790
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 6918 2000 6974 2009
rect 6918 1935 6974 1944
rect 8312 1465 8340 2450
rect 8298 1456 8354 1465
rect 8298 1391 8354 1400
rect 6918 82 6974 480
rect 6656 54 6974 82
rect 3054 0 3110 54
rect 4342 0 4398 54
rect 5630 0 5686 54
rect 6918 0 6974 54
rect 8114 82 8170 480
rect 8404 82 8432 4247
rect 8496 3670 8524 8298
rect 8680 8294 8708 8502
rect 9140 8498 9168 13126
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9232 12102 9260 12718
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9324 11898 9352 17711
rect 9416 17338 9444 17750
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9876 16998 9904 18022
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10692 17808 10744 17814
rect 10692 17750 10744 17756
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9680 14816 9732 14822
rect 9732 14776 9812 14804
rect 9680 14758 9732 14764
rect 9784 14550 9812 14776
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 13938 9720 14350
rect 9784 14074 9812 14486
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9416 13530 9444 13874
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9678 13424 9734 13433
rect 9678 13359 9734 13368
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9416 12442 9444 12786
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9508 11762 9536 13262
rect 9692 13190 9720 13359
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9784 12714 9812 13126
rect 9588 12708 9640 12714
rect 9772 12708 9824 12714
rect 9640 12668 9720 12696
rect 9588 12650 9640 12656
rect 9692 12238 9720 12668
rect 9772 12650 9824 12656
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9692 11898 9720 12174
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9324 9654 9352 11494
rect 9508 11286 9536 11698
rect 9784 11558 9812 12650
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9784 10538 9812 11494
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9876 10282 9904 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16726 10732 17750
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 16250 10180 16526
rect 10244 16454 10272 16662
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10244 16182 10272 16390
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10244 16028 10272 16118
rect 10152 16000 10272 16028
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10060 15706 10088 15914
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10152 15026 10180 16000
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10428 15162 10456 15574
rect 10796 15434 10824 18022
rect 10888 16998 10916 18022
rect 11072 17785 11100 27474
rect 11716 27443 11744 27474
rect 11612 22432 11664 22438
rect 11612 22374 11664 22380
rect 11058 17776 11114 17785
rect 11058 17711 11114 17720
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 11256 17202 11284 17478
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9968 12442 9996 14010
rect 10060 13802 10088 14758
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14618 10732 15098
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10152 12986 10180 13942
rect 10428 13802 10456 14010
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13530 10732 13874
rect 10888 13870 10916 16934
rect 11532 16590 11560 17002
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11164 16114 11192 16526
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11072 15162 11100 15438
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10520 12986 10548 13330
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9968 11626 9996 12378
rect 10060 12238 10088 12786
rect 10888 12646 10916 13262
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9876 10254 9996 10282
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9876 9722 9904 10134
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9416 8430 9444 8774
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9692 8430 9720 8570
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8680 7750 8708 8230
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 9692 7546 9720 7890
rect 9876 7818 9904 8774
rect 9968 8634 9996 10254
rect 10060 10062 10088 12174
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10888 11354 10916 12582
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10704 10470 10732 11154
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10810 11100 11086
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10169 10732 10406
rect 11072 10266 11100 10746
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10690 10160 10746 10169
rect 10690 10095 10746 10104
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10704 9654 10732 9930
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 11256 9178 11284 16390
rect 11334 15600 11390 15609
rect 11334 15535 11390 15544
rect 11348 11354 11376 15535
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11440 14006 11468 14418
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 11440 13530 11468 13942
rect 11532 13938 11560 14554
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11624 13814 11652 22374
rect 13924 19922 13952 27520
rect 16026 27520 16082 28000
rect 18234 27532 18290 28000
rect 18234 27520 18236 27532
rect 15752 27474 15804 27480
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 12268 19514 12296 19858
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13648 19514 13676 19654
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12820 18970 12848 19246
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11716 17746 11744 18702
rect 11992 17814 12020 18702
rect 12820 18154 12848 18906
rect 12912 18426 12940 19246
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13464 18902 13492 19178
rect 13648 18970 13676 19450
rect 13740 18970 13768 19790
rect 14568 19174 14596 19858
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15476 19236 15528 19242
rect 15396 19196 15476 19224
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13464 18426 13492 18838
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13740 18154 13768 18702
rect 14292 18290 14320 18906
rect 14568 18290 14596 19110
rect 15396 18834 15424 19196
rect 15476 19178 15528 19184
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 14372 18148 14424 18154
rect 14372 18090 14424 18096
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 11980 17808 12032 17814
rect 11980 17750 12032 17756
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17649 11744 17682
rect 11796 17672 11848 17678
rect 11702 17640 11758 17649
rect 11796 17614 11848 17620
rect 11702 17575 11758 17584
rect 11808 16454 11836 17614
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11624 13786 11744 13814
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11440 11898 11468 12378
rect 11532 12238 11560 12854
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11532 11898 11560 12174
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11440 10470 11468 11222
rect 11624 10606 11652 12582
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11440 10198 11468 10406
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11348 9722 11376 10134
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11440 9654 11468 10134
rect 11532 10062 11560 10474
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11428 9648 11480 9654
rect 11428 9590 11480 9596
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 10060 8294 10088 8366
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9864 7812 9916 7818
rect 9916 7772 9996 7800
rect 9864 7754 9916 7760
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9220 6384 9272 6390
rect 9416 6361 9444 7278
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9220 6326 9272 6332
rect 9402 6352 9458 6361
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 5914 8616 6054
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8772 4154 8800 6122
rect 8942 5808 8998 5817
rect 8942 5743 8998 5752
rect 8956 4729 8984 5743
rect 9140 4729 9168 6326
rect 9232 5370 9260 6326
rect 9402 6287 9458 6296
rect 9494 6216 9550 6225
rect 9494 6151 9550 6160
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9232 5166 9260 5306
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 8942 4720 8998 4729
rect 8942 4655 8998 4664
rect 9126 4720 9182 4729
rect 9416 4690 9444 5034
rect 9126 4655 9182 4664
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 8588 4126 8800 4154
rect 8588 3738 8616 4126
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8496 3194 8524 3606
rect 8588 3466 8616 3674
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8772 2854 8800 3878
rect 9048 3126 9076 4422
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3534 9352 3878
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 9140 2922 9168 3334
rect 9128 2916 9180 2922
rect 9128 2858 9180 2864
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8772 2582 8800 2790
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 8114 54 8432 82
rect 9402 82 9458 480
rect 9508 82 9536 6151
rect 9692 5370 9720 6938
rect 9784 6866 9812 7754
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9876 7206 9904 7482
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6934 9904 7142
rect 9968 7002 9996 7772
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9784 5914 9812 6802
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9876 5846 9904 6870
rect 10060 6798 10088 8230
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 7410 10732 8774
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10796 7750 10824 8298
rect 10980 8090 11008 8502
rect 11164 8294 11192 8978
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 7410 10824 7686
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10704 7002 10732 7346
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6254 10088 6734
rect 10428 6390 10456 6802
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10704 6254 10732 6802
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9968 5778 9996 6054
rect 10060 5914 10088 6190
rect 10704 6118 10732 6190
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9692 4690 9720 5306
rect 9968 4826 9996 5714
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9600 4078 9628 4626
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9588 4072 9640 4078
rect 9586 4040 9588 4049
rect 9640 4040 9642 4049
rect 9586 3975 9642 3984
rect 9600 3738 9628 3975
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9784 2446 9812 4558
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10336 4146 10364 4422
rect 10796 4196 10824 7346
rect 10980 6866 11008 8026
rect 11532 7954 11560 8230
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11532 7546 11560 7890
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 10968 6860 11020 6866
rect 10888 6820 10968 6848
rect 10888 6186 10916 6820
rect 10968 6802 11020 6808
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11256 6254 11284 6598
rect 11532 6322 11560 6734
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10980 4865 11008 5034
rect 10966 4856 11022 4865
rect 10966 4791 11022 4800
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10704 4168 10824 4196
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10704 4078 10732 4168
rect 10980 4146 11008 4694
rect 10968 4140 11020 4146
rect 10888 4100 10968 4128
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9968 2514 9996 3674
rect 10704 3602 10732 4014
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10796 3670 10824 3946
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 10152 3126 10180 3402
rect 10796 3126 10824 3606
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 10784 2916 10836 2922
rect 10888 2904 10916 4100
rect 10968 4082 11020 4088
rect 10836 2876 10916 2904
rect 10784 2858 10836 2864
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 10888 2378 10916 2876
rect 10968 2848 11020 2854
rect 11072 2836 11100 5782
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11164 5370 11192 5510
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11164 3602 11192 4218
rect 11256 4078 11284 6190
rect 11532 5914 11560 6258
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11348 4554 11376 5578
rect 11624 5273 11652 8570
rect 11610 5264 11666 5273
rect 11610 5199 11666 5208
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11348 3738 11376 3946
rect 11532 3738 11560 4694
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11348 3058 11376 3674
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11020 2808 11100 2836
rect 10968 2790 11020 2796
rect 10980 2582 11008 2790
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 9402 54 9536 82
rect 10690 82 10746 480
rect 10980 82 11008 2314
rect 10690 54 11008 82
rect 11624 82 11652 5199
rect 11716 3466 11744 13786
rect 11808 13734 11836 14418
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13433 11836 13670
rect 11888 13456 11940 13462
rect 11794 13424 11850 13433
rect 11888 13398 11940 13404
rect 11794 13359 11850 13368
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11808 11286 11836 13194
rect 11900 12986 11928 13398
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11808 10810 11836 11222
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11794 10704 11850 10713
rect 11794 10639 11850 10648
rect 11808 10606 11836 10639
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11992 9586 12020 9930
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11796 9036 11848 9042
rect 11980 9036 12032 9042
rect 11848 8996 11928 9024
rect 11796 8978 11848 8984
rect 11900 8294 11928 8996
rect 11980 8978 12032 8984
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11900 7954 11928 8230
rect 11888 7948 11940 7954
rect 11992 7936 12020 8978
rect 12084 8090 12112 17070
rect 12176 17066 12204 17818
rect 12728 17746 12756 18090
rect 12820 17882 12848 18090
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 13740 17678 13768 18090
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12820 17134 12848 17478
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 13360 17060 13412 17066
rect 13360 17002 13412 17008
rect 12900 16720 12952 16726
rect 12900 16662 12952 16668
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12820 16250 12848 16526
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12176 15910 12204 16050
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 14482 12204 15846
rect 12912 15706 12940 16662
rect 13174 16144 13230 16153
rect 13174 16079 13230 16088
rect 13188 16046 13216 16079
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12268 15065 12296 15506
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12254 15056 12310 15065
rect 12254 14991 12310 15000
rect 12268 14958 12296 14991
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12268 14074 12296 14350
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12544 12850 12572 15302
rect 12912 14618 12940 15438
rect 13188 15026 13216 15846
rect 13372 15638 13400 17002
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13464 16182 13492 16526
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13372 14822 13400 15574
rect 13464 15434 13492 16118
rect 13556 16114 13584 17614
rect 13740 16794 13768 17614
rect 13832 17134 13860 17750
rect 14384 17202 14412 18090
rect 14568 17814 14596 18226
rect 15396 18086 15424 18770
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 14556 16108 14608 16114
rect 14924 16108 14976 16114
rect 14608 16068 14924 16096
rect 14556 16050 14608 16056
rect 14924 16050 14976 16056
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13372 14618 13400 14758
rect 13924 14618 13952 15914
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14292 15162 14320 15846
rect 14568 15706 14596 16050
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 12728 13734 12756 14554
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13280 13870 13308 14418
rect 14016 13938 14044 14758
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 13096 13394 13124 13806
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12544 12442 12572 12786
rect 12728 12714 12756 13126
rect 13096 12986 13124 13330
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 10266 12480 12038
rect 12728 10742 12756 12650
rect 13280 12102 13308 13330
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13280 11354 13308 11562
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 13004 10674 13032 10950
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 9722 12204 9862
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12912 9178 12940 9998
rect 13004 9518 13032 10202
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13004 9110 13032 9454
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12268 8566 12296 8978
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12072 7948 12124 7954
rect 11992 7908 12072 7936
rect 11888 7890 11940 7896
rect 12072 7890 12124 7896
rect 11900 7002 11928 7890
rect 12084 7410 12112 7890
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12360 7002 12388 7278
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 11900 6390 11928 6938
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 12268 6186 12296 6870
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12084 5234 12112 6054
rect 12268 5846 12296 6122
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 12176 5370 12204 5782
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12452 5302 12480 7142
rect 12544 6186 12572 8298
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12544 5914 12572 6122
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12530 5672 12586 5681
rect 12530 5607 12586 5616
rect 12544 5574 12572 5607
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12452 5030 12480 5238
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 12176 3398 12204 3946
rect 12360 3670 12388 4558
rect 12544 4486 12572 5034
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12176 1737 12204 3334
rect 12360 3194 12388 3606
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12452 2514 12480 3878
rect 12544 3058 12572 4150
rect 12636 3194 12664 8366
rect 13004 8022 13032 9046
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12728 5642 12756 6734
rect 12820 6322 12848 7346
rect 13004 6934 13032 7414
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 13096 4865 13124 10406
rect 13280 10198 13308 11290
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13280 9722 13308 10134
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13372 9042 13400 13670
rect 13832 13530 13860 13806
rect 14476 13734 14504 14350
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13464 11762 13492 13262
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13648 11626 13676 12378
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11694 13768 12174
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13556 10169 13584 10610
rect 13648 10538 13676 10678
rect 13740 10674 13768 11630
rect 14016 11286 14044 12038
rect 14200 11898 14228 12582
rect 14292 12102 14320 12650
rect 14568 12170 14596 12786
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13648 10266 13676 10474
rect 14016 10470 14044 11222
rect 14188 10532 14240 10538
rect 14292 10520 14320 12038
rect 14568 11286 14596 12106
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14240 10492 14320 10520
rect 14188 10474 14240 10480
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13542 10160 13598 10169
rect 14200 10130 14228 10474
rect 13542 10095 13598 10104
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14660 10010 14688 14894
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14844 13530 14872 13806
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 15396 13394 15424 18022
rect 15580 16658 15608 19654
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15672 17882 15700 19110
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15672 17202 15700 17818
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15672 16697 15700 16730
rect 15658 16688 15714 16697
rect 15568 16652 15620 16658
rect 15658 16623 15714 16632
rect 15568 16594 15620 16600
rect 15580 16250 15608 16594
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15474 15464 15530 15473
rect 15474 15399 15530 15408
rect 15488 15162 15516 15399
rect 15764 15162 15792 27474
rect 16040 19417 16068 27520
rect 18288 27520 18290 27532
rect 20350 27520 20406 28000
rect 22466 27520 22522 28000
rect 24674 27520 24730 28000
rect 26790 27520 26846 28000
rect 18236 27474 18288 27480
rect 18248 27443 18276 27474
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19982 22536 20038 22545
rect 18880 22500 18932 22506
rect 19982 22471 20038 22480
rect 18880 22442 18932 22448
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16026 19408 16082 19417
rect 16026 19343 16082 19352
rect 16500 19310 16528 19654
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15856 18086 15884 18770
rect 16212 18692 16264 18698
rect 16212 18634 16264 18640
rect 16224 18290 16252 18634
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16224 18193 16252 18226
rect 16210 18184 16266 18193
rect 16408 18154 16436 18566
rect 16210 18119 16266 18128
rect 16396 18148 16448 18154
rect 16396 18090 16448 18096
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15764 14958 15792 15098
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15856 13841 15884 18022
rect 16304 17808 16356 17814
rect 16304 17750 16356 17756
rect 16120 17604 16172 17610
rect 16120 17546 16172 17552
rect 16132 17105 16160 17546
rect 16118 17096 16174 17105
rect 16118 17031 16174 17040
rect 16132 16794 16160 17031
rect 16316 16998 16344 17750
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16212 16176 16264 16182
rect 16212 16118 16264 16124
rect 16224 15978 16252 16118
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 15948 14822 15976 15574
rect 16132 15434 16160 15914
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 16224 15026 16252 15302
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15948 14618 15976 14758
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15842 13832 15898 13841
rect 15842 13767 15898 13776
rect 15844 13728 15896 13734
rect 15948 13716 15976 14554
rect 15896 13688 15976 13716
rect 15844 13670 15896 13676
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15488 11665 15516 12854
rect 15580 12850 15608 13398
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15764 12918 15792 13330
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 12442 15608 12786
rect 15856 12646 15884 13670
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15948 12170 15976 12718
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15752 11688 15804 11694
rect 15474 11656 15530 11665
rect 15752 11630 15804 11636
rect 15474 11591 15530 11600
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15396 10810 15424 11086
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15488 10742 15516 11222
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15120 10266 15148 10542
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 10266 15608 10474
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 14476 9982 14688 10010
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13372 8634 13400 8978
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13280 7478 13308 8298
rect 13556 7954 13584 9318
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14384 8430 14412 9046
rect 14476 8838 14504 9982
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14568 9674 14596 9862
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 10066
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15292 9716 15344 9722
rect 15212 9676 15292 9704
rect 14568 9646 14688 9674
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14568 9110 14596 9454
rect 14660 9382 14688 9646
rect 15212 9518 15240 9676
rect 15292 9658 15344 9664
rect 15304 9593 15332 9658
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 13556 6866 13584 7890
rect 13924 7750 13952 7890
rect 14384 7818 14412 8366
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13924 7546 13952 7686
rect 14476 7546 14504 8774
rect 14660 8430 14688 9114
rect 15212 8820 15240 9454
rect 15292 9444 15344 9450
rect 15396 9432 15424 9930
rect 15344 9404 15424 9432
rect 15292 9386 15344 9392
rect 15396 9178 15424 9404
rect 15580 9382 15608 10066
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15292 8832 15344 8838
rect 15212 8792 15292 8820
rect 15292 8774 15344 8780
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 15304 8362 15332 8774
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15120 8090 15148 8230
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14476 7342 14504 7482
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14568 6934 14596 7822
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14556 6928 14608 6934
rect 14556 6870 14608 6876
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13556 6662 13584 6802
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13188 5710 13216 6258
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13188 5234 13216 5646
rect 13556 5574 13584 6598
rect 13740 6118 13768 6802
rect 13924 6186 14228 6202
rect 13912 6180 14240 6186
rect 13964 6174 14188 6180
rect 13912 6122 13964 6128
rect 14188 6122 14240 6128
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13648 5370 13676 5714
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13740 5030 13768 6054
rect 14568 5574 14596 6054
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13082 4856 13138 4865
rect 13082 4791 13138 4800
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 13004 3738 13032 4626
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12820 3058 12848 3402
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 13004 2922 13032 3674
rect 13556 3670 13584 3878
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 12992 2916 13044 2922
rect 12992 2858 13044 2864
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12820 2446 12848 2518
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 13280 2378 13308 3606
rect 13648 3602 13676 4082
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13464 3058 13492 3334
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13648 2650 13676 3538
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12162 1728 12218 1737
rect 12162 1663 12218 1672
rect 11978 82 12034 480
rect 11624 54 12034 82
rect 8114 0 8170 54
rect 9402 0 9458 54
rect 10690 0 10746 54
rect 11978 0 12034 54
rect 13266 82 13322 480
rect 13372 82 13400 2586
rect 13832 2514 13860 4694
rect 13924 2854 13952 5510
rect 14462 5264 14518 5273
rect 14462 5199 14518 5208
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 14016 2961 14044 5102
rect 14280 4480 14332 4486
rect 14476 4457 14504 5199
rect 14568 5137 14596 5510
rect 14554 5128 14610 5137
rect 14554 5063 14610 5072
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14568 4593 14596 4626
rect 14554 4584 14610 4593
rect 14554 4519 14610 4528
rect 14648 4548 14700 4554
rect 14280 4422 14332 4428
rect 14462 4448 14518 4457
rect 14292 4078 14320 4422
rect 14462 4383 14518 4392
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14108 3097 14136 4014
rect 14292 3194 14320 4014
rect 14568 3738 14596 4519
rect 14648 4490 14700 4496
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14094 3088 14150 3097
rect 14094 3023 14150 3032
rect 14108 2990 14136 3023
rect 14292 2990 14320 3130
rect 14096 2984 14148 2990
rect 14002 2952 14058 2961
rect 14280 2984 14332 2990
rect 14096 2926 14148 2932
rect 14200 2944 14280 2972
rect 14002 2887 14058 2896
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 14016 649 14044 2887
rect 14200 2582 14228 2944
rect 14280 2926 14332 2932
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 14002 640 14058 649
rect 14002 575 14058 584
rect 13266 54 13400 82
rect 14554 82 14610 480
rect 14660 82 14688 4490
rect 14752 4214 14780 5510
rect 14844 4826 14872 7278
rect 15304 6848 15332 8298
rect 15488 8022 15516 8298
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15384 6860 15436 6866
rect 15304 6820 15384 6848
rect 15384 6802 15436 6808
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15396 6390 15424 6802
rect 15488 6798 15516 7414
rect 15580 7324 15608 9318
rect 15672 9042 15700 9386
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8634 15700 8978
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15660 7336 15712 7342
rect 15580 7296 15660 7324
rect 15660 7278 15712 7284
rect 15672 7206 15700 7278
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15672 6866 15700 7142
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15488 6458 15516 6734
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 15672 6118 15700 6802
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14844 4078 14872 4762
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14844 2922 14872 4014
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 15028 2650 15056 2858
rect 15016 2644 15068 2650
rect 15016 2586 15068 2592
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15304 2009 15332 4490
rect 15396 3097 15424 6054
rect 15764 4690 15792 11630
rect 16040 10198 16068 13126
rect 16132 12306 16160 13262
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16132 11354 16160 12242
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15764 4282 15792 4626
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15856 4154 15884 8774
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15948 7342 15976 7754
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 16132 5778 16160 10202
rect 16224 8566 16252 14962
rect 16408 14872 16436 18090
rect 16684 16658 16712 19178
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17132 18896 17184 18902
rect 17052 18856 17132 18884
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 16868 17678 16896 18090
rect 17052 18086 17080 18856
rect 17132 18838 17184 18844
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 17052 17066 17080 18022
rect 17236 17882 17264 18906
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16684 16250 16712 16594
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16960 15910 16988 16730
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16960 15638 16988 15846
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 16488 14884 16540 14890
rect 16408 14844 16488 14872
rect 16488 14826 16540 14832
rect 16500 14618 16528 14826
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16500 13190 16528 13738
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16684 12986 16712 13194
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16776 12889 16804 13806
rect 16868 12986 16896 14554
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16762 12880 16818 12889
rect 16762 12815 16818 12824
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16316 12374 16344 12582
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16316 11558 16344 12310
rect 16868 11626 16896 12922
rect 17052 12442 17080 17002
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17328 16726 17356 16934
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17236 14618 17264 15438
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17224 14272 17276 14278
rect 17328 14260 17356 16662
rect 17420 14414 17448 18702
rect 17788 17678 17816 18702
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 18064 18204 18092 18566
rect 18144 18216 18196 18222
rect 18064 18176 18144 18204
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17788 17338 17816 17614
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17788 15706 17816 16934
rect 17880 16794 17908 17750
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17512 15162 17540 15574
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17276 14232 17356 14260
rect 17224 14214 17276 14220
rect 17236 13462 17264 14214
rect 17420 14074 17448 14350
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17788 13734 17816 14554
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17144 12646 17172 13262
rect 17236 12986 17264 13398
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16316 9110 16344 11494
rect 16500 11286 16528 11562
rect 16868 11354 16896 11562
rect 17420 11558 17448 12174
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16500 10810 16528 11222
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 16948 10056 17000 10062
rect 16486 10024 16542 10033
rect 16948 9998 17000 10004
rect 16486 9959 16542 9968
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16316 8294 16344 9046
rect 16500 8634 16528 9959
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16684 9178 16712 9386
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16960 8974 16988 9998
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 8022 16344 8230
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 16316 7546 16344 7958
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 17052 7342 17080 9318
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16592 6186 16620 6666
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 16132 5370 16160 5714
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 15764 4126 15884 4154
rect 15568 4004 15620 4010
rect 15568 3946 15620 3952
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15488 3126 15516 3334
rect 15476 3120 15528 3126
rect 15382 3088 15438 3097
rect 15476 3062 15528 3068
rect 15382 3023 15438 3032
rect 15580 2514 15608 3946
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15764 2417 15792 4126
rect 16132 3670 16160 4966
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 15856 2854 15884 3606
rect 16316 3194 16344 4558
rect 16684 4185 16712 7278
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16868 7002 16896 7142
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16868 6322 16896 6938
rect 17040 6928 17092 6934
rect 17040 6870 17092 6876
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 17052 5914 17080 6870
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17052 5166 17080 5850
rect 17144 5817 17172 10406
rect 17130 5808 17186 5817
rect 17130 5743 17186 5752
rect 17236 5302 17264 10746
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17328 9382 17356 10134
rect 17420 9722 17448 11494
rect 17512 11218 17540 12786
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17512 10810 17540 11154
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17604 9586 17632 9998
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 7750 17356 9318
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17512 8362 17540 9046
rect 17604 8974 17632 9522
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17696 8566 17724 13194
rect 17880 12918 17908 15846
rect 17972 15502 18000 18022
rect 18064 16046 18092 18176
rect 18144 18158 18196 18164
rect 18432 17814 18460 20334
rect 18788 18148 18840 18154
rect 18788 18090 18840 18096
rect 18420 17808 18472 17814
rect 18420 17750 18472 17756
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18156 16046 18184 16390
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17972 13326 18000 14962
rect 18156 14482 18184 15846
rect 18248 15502 18276 17138
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 18340 16726 18368 17002
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18432 15502 18460 17750
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18248 15162 18276 15438
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 18248 14550 18276 15098
rect 18432 15026 18460 15438
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18340 14618 18368 14758
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18236 14544 18288 14550
rect 18236 14486 18288 14492
rect 18800 14482 18828 18090
rect 18144 14476 18196 14482
rect 18788 14476 18840 14482
rect 18144 14418 18196 14424
rect 18708 14436 18788 14464
rect 18340 13870 18368 13901
rect 18328 13864 18380 13870
rect 18326 13832 18328 13841
rect 18380 13832 18382 13841
rect 18326 13767 18382 13776
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18156 12442 18184 12582
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 17788 11898 17816 12378
rect 18248 12238 18276 13262
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 18248 11762 18276 12174
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18340 11694 18368 13767
rect 18708 13734 18736 14436
rect 18788 14418 18840 14424
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18432 12850 18460 13330
rect 18708 13258 18736 13670
rect 18800 13462 18828 13806
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18800 13190 18828 13398
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18616 12753 18644 12786
rect 18602 12744 18658 12753
rect 18602 12679 18658 12688
rect 18708 12646 18736 12922
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18524 11218 18552 11630
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18524 11014 18552 11154
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 18156 9994 18184 10474
rect 18340 9994 18368 10474
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18524 9926 18552 10950
rect 18602 10160 18658 10169
rect 18602 10095 18658 10104
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18616 9654 18644 10095
rect 18708 9722 18736 12582
rect 18800 12374 18828 13126
rect 18788 12368 18840 12374
rect 18788 12310 18840 12316
rect 18786 11248 18842 11257
rect 18786 11183 18842 11192
rect 18800 10674 18828 11183
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18708 9042 18736 9658
rect 18800 9586 18828 10610
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18236 8900 18288 8906
rect 18236 8842 18288 8848
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17420 7002 17448 7890
rect 17512 7478 17540 7958
rect 17696 7886 17724 8502
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17500 7472 17552 7478
rect 17500 7414 17552 7420
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17880 6866 17908 7822
rect 18156 7546 18184 8230
rect 18248 7993 18276 8842
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18234 7984 18290 7993
rect 18234 7919 18290 7928
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18156 7002 18184 7482
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17590 6352 17646 6361
rect 17590 6287 17646 6296
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17420 5914 17448 6054
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 17040 5160 17092 5166
rect 16854 5128 16910 5137
rect 16764 5092 16816 5098
rect 16816 5072 16854 5080
rect 17040 5102 17092 5108
rect 16816 5063 16910 5072
rect 16816 5052 16896 5063
rect 16764 5034 16816 5040
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16670 4176 16726 4185
rect 16670 4111 16726 4120
rect 16488 4004 16540 4010
rect 16488 3946 16540 3952
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 15856 2582 15884 2790
rect 16408 2650 16436 3878
rect 16500 3466 16528 3946
rect 16776 3670 16804 4626
rect 17052 4486 17080 5102
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 17328 4826 17356 5034
rect 17420 5030 17448 5850
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17512 5234 17540 5646
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17512 4826 17540 5170
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16592 2922 16620 3130
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16500 2666 16528 2858
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16684 2666 16712 2790
rect 16396 2644 16448 2650
rect 16500 2638 16712 2666
rect 16396 2586 16448 2592
rect 15844 2576 15896 2582
rect 15844 2518 15896 2524
rect 15750 2408 15806 2417
rect 15750 2343 15806 2352
rect 16028 2372 16080 2378
rect 16028 2314 16080 2320
rect 15290 2000 15346 2009
rect 15290 1935 15346 1944
rect 14554 54 14688 82
rect 15750 82 15806 480
rect 16040 82 16068 2314
rect 16960 2009 16988 4218
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 17144 3534 17172 3946
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17144 2446 17172 3470
rect 17236 3194 17264 3606
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17420 3058 17448 3470
rect 17604 3194 17632 6287
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17696 5846 17724 6190
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17880 5642 17908 6802
rect 18156 6118 18184 6938
rect 18248 6186 18276 7346
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 18524 7002 18552 7210
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18248 5710 18276 6122
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 18248 5234 18276 5646
rect 18328 5636 18380 5642
rect 18328 5578 18380 5584
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18156 4826 18184 5034
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18340 4690 18368 5578
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18432 5098 18460 5510
rect 18420 5092 18472 5098
rect 18420 5034 18472 5040
rect 18616 4690 18644 8366
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18708 6458 18736 6598
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 17788 3534 17816 4558
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18156 4146 18184 4422
rect 18340 4282 18368 4626
rect 18892 4486 18920 22442
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19996 21146 20024 22471
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 19628 20534 19656 20946
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19076 16658 19104 19246
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19076 16153 19104 16594
rect 19062 16144 19118 16153
rect 19062 16079 19118 16088
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18984 12986 19012 15982
rect 19076 15910 19104 16079
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18970 12880 19026 12889
rect 18970 12815 19026 12824
rect 18984 7954 19012 12815
rect 19076 12220 19104 15846
rect 19260 15706 19288 16594
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19536 16114 19564 16526
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19536 15706 19564 16050
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19260 14482 19288 15642
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19248 14476 19300 14482
rect 19168 14436 19248 14464
rect 19168 13870 19196 14436
rect 19248 14418 19300 14424
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19260 13530 19288 13874
rect 19352 13870 19380 14894
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 19260 12374 19288 12718
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19076 12192 19380 12220
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 19076 10266 19104 11086
rect 19168 10674 19196 11562
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19260 11286 19288 11494
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19260 10470 19288 11222
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19076 9382 19104 10066
rect 19168 9926 19196 10066
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19168 9382 19196 9862
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18984 7546 19012 7890
rect 19076 7857 19104 9318
rect 19168 9042 19196 9318
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19168 8430 19196 8978
rect 19260 8430 19288 10406
rect 19352 10198 19380 12192
rect 19536 11830 19564 12242
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19168 7936 19196 8366
rect 19352 8294 19380 8910
rect 19536 8498 19564 11630
rect 19904 11540 19932 11698
rect 19996 11694 20024 12038
rect 20088 11898 20116 15370
rect 20272 14822 20300 15846
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20180 13938 20208 14214
rect 20272 14006 20300 14758
rect 20260 14000 20312 14006
rect 20260 13942 20312 13948
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20364 13814 20392 27520
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 21100 18970 21128 24006
rect 22480 23866 22508 27520
rect 23202 26888 23258 26897
rect 23202 26823 23258 26832
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22848 23866 22876 24210
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 22744 23792 22796 23798
rect 22744 23734 22796 23740
rect 21548 23656 21600 23662
rect 21548 23598 21600 23604
rect 21560 18970 21588 23598
rect 22468 23588 22520 23594
rect 22468 23530 22520 23536
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 21732 18828 21784 18834
rect 21732 18770 21784 18776
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20548 17202 20576 17478
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20548 16794 20576 17138
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20456 14958 20484 15302
rect 20444 14952 20496 14958
rect 20444 14894 20496 14900
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20260 13796 20312 13802
rect 20364 13786 20576 13814
rect 20260 13738 20312 13744
rect 20272 13394 20300 13738
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19904 11512 20024 11540
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19720 8498 19748 8910
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19248 7948 19300 7954
rect 19168 7908 19248 7936
rect 19062 7848 19118 7857
rect 19168 7818 19196 7908
rect 19248 7890 19300 7896
rect 19062 7783 19118 7792
rect 19156 7812 19208 7818
rect 19156 7754 19208 7760
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 19168 6934 19196 7754
rect 19248 7472 19300 7478
rect 19352 7460 19380 8230
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19300 7432 19380 7460
rect 19248 7414 19300 7420
rect 19156 6928 19208 6934
rect 19156 6870 19208 6876
rect 19352 6361 19380 7432
rect 19996 7342 20024 11512
rect 20364 11354 20392 12582
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 20180 10266 20208 10610
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19996 7206 20024 7278
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19536 6390 19564 6938
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19524 6384 19576 6390
rect 19338 6352 19394 6361
rect 19524 6326 19576 6332
rect 19338 6287 19394 6296
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 19524 6112 19576 6118
rect 19628 6100 19656 6802
rect 19984 6180 20036 6186
rect 19984 6122 20036 6128
rect 19576 6072 19656 6100
rect 19524 6054 19576 6060
rect 18984 5846 19012 6054
rect 18972 5840 19024 5846
rect 18972 5782 19024 5788
rect 19432 5840 19484 5846
rect 19536 5817 19564 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19996 5846 20024 6122
rect 19984 5840 20036 5846
rect 19432 5782 19484 5788
rect 19522 5808 19578 5817
rect 19444 5370 19472 5782
rect 19984 5782 20036 5788
rect 19522 5743 19578 5752
rect 19996 5370 20024 5782
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19996 5030 20024 5306
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 19260 4282 19288 4626
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 20088 4154 20116 7482
rect 20272 7342 20300 7686
rect 20260 7336 20312 7342
rect 20180 7296 20260 7324
rect 20180 4690 20208 7296
rect 20260 7278 20312 7284
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20272 5574 20300 6190
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20168 4684 20220 4690
rect 20168 4626 20220 4632
rect 20180 4214 20208 4626
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 19904 4126 20116 4154
rect 20168 4208 20220 4214
rect 20168 4150 20220 4156
rect 17880 3942 17908 4082
rect 18050 4040 18106 4049
rect 18050 3975 18106 3984
rect 18420 4004 18472 4010
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 16946 2000 17002 2009
rect 16946 1935 17002 1944
rect 15750 54 16068 82
rect 16960 82 16988 1935
rect 17038 82 17094 480
rect 16960 54 17094 82
rect 18064 82 18092 3975
rect 18420 3946 18472 3952
rect 18432 3738 18460 3946
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18156 3058 18184 3334
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18156 2650 18184 2994
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18432 2446 18460 3334
rect 18524 3126 18552 4082
rect 19904 4060 19932 4126
rect 19984 4072 20036 4078
rect 19904 4032 19984 4060
rect 20036 4032 20116 4060
rect 19984 4014 20036 4020
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18512 3120 18564 3126
rect 18512 3062 18564 3068
rect 18616 2922 18644 3470
rect 20088 3398 20116 4032
rect 20180 3738 20208 4150
rect 20272 4146 20300 5510
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20364 3738 20392 5238
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20456 4758 20484 5102
rect 20444 4752 20496 4758
rect 20548 4729 20576 13786
rect 20640 13190 20668 14350
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20732 13462 20760 13670
rect 20720 13456 20772 13462
rect 20720 13398 20772 13404
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20640 12782 20668 13126
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20628 12640 20680 12646
rect 20732 12628 20760 13398
rect 20680 12600 20760 12628
rect 20628 12582 20680 12588
rect 20640 11626 20668 12582
rect 20824 11642 20852 18226
rect 21744 18154 21772 18770
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21928 18154 21956 18566
rect 21732 18148 21784 18154
rect 21732 18090 21784 18096
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 20994 17776 21050 17785
rect 20994 17711 21050 17720
rect 21008 17678 21036 17711
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17202 21036 17614
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 21008 14074 21036 17002
rect 21192 16590 21220 17206
rect 21272 16720 21324 16726
rect 21272 16662 21324 16668
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21100 14550 21128 15982
rect 21192 15706 21220 16526
rect 21284 16250 21312 16662
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21468 15502 21496 17274
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21468 15026 21496 15438
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21284 14006 21312 14554
rect 21272 14000 21324 14006
rect 21272 13942 21324 13948
rect 21284 13734 21312 13942
rect 21560 13814 21588 17138
rect 21744 16522 21772 18090
rect 21732 16516 21784 16522
rect 21732 16458 21784 16464
rect 21640 15632 21692 15638
rect 21640 15574 21692 15580
rect 21652 15162 21680 15574
rect 21744 15502 21772 16458
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 21928 15162 21956 18090
rect 22112 17882 22140 22918
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22112 17202 22140 17818
rect 22204 17338 22232 18090
rect 22480 17882 22508 23530
rect 22558 21040 22614 21049
rect 22558 20975 22614 20984
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22296 17082 22324 17274
rect 22112 17066 22324 17082
rect 22100 17060 22324 17066
rect 22152 17054 22324 17060
rect 22100 17002 22152 17008
rect 22284 16992 22336 16998
rect 22284 16934 22336 16940
rect 22296 16522 22324 16934
rect 22480 16794 22508 17818
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 22112 16046 22140 16390
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 21640 15156 21692 15162
rect 21640 15098 21692 15104
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21836 14550 21864 14758
rect 21824 14544 21876 14550
rect 21824 14486 21876 14492
rect 22296 14278 22324 16458
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22480 15638 22508 15846
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 21560 13786 21772 13814
rect 22204 13802 22232 14010
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 20916 11801 20944 12650
rect 20902 11792 20958 11801
rect 20902 11727 20958 11736
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20732 11614 20852 11642
rect 20732 10577 20760 11614
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20824 10810 20852 11494
rect 21192 11286 21220 12650
rect 21560 12442 21588 12650
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 21192 10810 21220 11222
rect 21284 11014 21312 12174
rect 21376 11558 21404 12310
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 20718 10568 20774 10577
rect 20718 10503 20774 10512
rect 21284 9450 21312 10950
rect 21376 10606 21404 10950
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21376 10198 21404 10542
rect 21364 10192 21416 10198
rect 21364 10134 21416 10140
rect 21560 10062 21588 11018
rect 21640 10192 21692 10198
rect 21640 10134 21692 10140
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 21272 9444 21324 9450
rect 21272 9386 21324 9392
rect 20640 8838 20668 9386
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20732 8566 20760 9386
rect 21560 9382 21588 9998
rect 21652 9722 21680 10134
rect 21640 9716 21692 9722
rect 21640 9658 21692 9664
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20916 8022 20944 8910
rect 21192 8362 21220 9114
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21652 8362 21680 8502
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 21640 8356 21692 8362
rect 21640 8298 21692 8304
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 20904 8016 20956 8022
rect 20904 7958 20956 7964
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20640 5778 20668 7278
rect 20732 7002 20760 7346
rect 21008 7002 21036 8230
rect 21652 8090 21680 8298
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20640 4826 20668 5714
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20444 4694 20496 4700
rect 20534 4720 20590 4729
rect 20534 4655 20590 4664
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 19614 3224 19670 3233
rect 19614 3159 19670 3168
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 2961 19472 2994
rect 19628 2990 19656 3159
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 19616 2984 19668 2990
rect 19430 2952 19486 2961
rect 18604 2916 18656 2922
rect 19616 2926 19668 2932
rect 19430 2887 19486 2896
rect 18604 2858 18656 2864
rect 18616 2582 18644 2858
rect 19444 2854 19472 2887
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18326 82 18382 480
rect 18064 54 18382 82
rect 19536 82 19564 2790
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19996 2650 20024 3062
rect 20088 3058 20116 3334
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20548 2650 20576 4655
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 19614 82 19670 480
rect 19536 54 19670 82
rect 20732 82 20760 5578
rect 20904 5092 20956 5098
rect 20904 5034 20956 5040
rect 20916 3942 20944 5034
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20916 3602 20944 3878
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 20916 3194 20944 3538
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20916 2990 20944 3130
rect 21008 3126 21036 3538
rect 20996 3120 21048 3126
rect 20996 3062 21048 3068
rect 21100 3058 21128 7142
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 21192 2972 21220 3538
rect 21284 3466 21312 6734
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21468 5846 21496 6598
rect 21652 6322 21680 6598
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 21456 5840 21508 5846
rect 21456 5782 21508 5788
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21376 4282 21404 4966
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21376 3942 21404 4218
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21272 3460 21324 3466
rect 21272 3402 21324 3408
rect 21284 3126 21312 3402
rect 21272 3120 21324 3126
rect 21272 3062 21324 3068
rect 21272 2984 21324 2990
rect 21192 2944 21272 2972
rect 20824 2514 20852 2926
rect 20916 2650 20944 2926
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 21192 2514 21220 2944
rect 21272 2926 21324 2932
rect 21744 2514 21772 13786
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21836 12986 21864 13330
rect 22112 13172 22140 13738
rect 22296 13462 22324 14214
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22192 13184 22244 13190
rect 22112 13144 22192 13172
rect 22192 13126 22244 13132
rect 22204 12986 22232 13126
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 21824 12436 21876 12442
rect 21824 12378 21876 12384
rect 21836 11762 21864 12378
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 21836 8498 21864 11698
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21928 10810 21956 11086
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 21928 9722 21956 10746
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21836 7868 21864 8434
rect 21916 7880 21968 7886
rect 21836 7840 21916 7868
rect 21916 7822 21968 7828
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21836 7274 21864 7482
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21836 5914 21864 6054
rect 21824 5908 21876 5914
rect 21824 5850 21876 5856
rect 22020 4593 22048 9454
rect 22112 6798 22140 12038
rect 22204 11762 22232 12174
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22204 10130 22232 11698
rect 22466 10568 22522 10577
rect 22572 10554 22600 20975
rect 22650 17776 22706 17785
rect 22650 17711 22706 17720
rect 22664 15162 22692 17711
rect 22756 16726 22784 23734
rect 23216 23186 23244 26823
rect 24214 25664 24270 25673
rect 24214 25599 24270 25608
rect 24228 23866 24256 25599
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24688 24274 24716 27520
rect 24858 24576 24914 24585
rect 24858 24511 24914 24520
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24216 23860 24268 23866
rect 24216 23802 24268 23808
rect 24228 23662 24256 23802
rect 24216 23656 24268 23662
rect 24216 23598 24268 23604
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 23204 23180 23256 23186
rect 23204 23122 23256 23128
rect 22848 22778 22876 23122
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24766 19816 24822 19825
rect 24766 19751 24822 19760
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24780 18970 24808 19751
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18290 24716 18770
rect 24766 18728 24822 18737
rect 24766 18663 24822 18672
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 22928 18080 22980 18086
rect 22928 18022 22980 18028
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 22848 17270 22876 17614
rect 22836 17264 22888 17270
rect 22836 17206 22888 17212
rect 22940 16726 22968 18022
rect 24780 17882 24808 18663
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 23032 17338 23060 17750
rect 24214 17640 24270 17649
rect 24214 17575 24270 17584
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 24228 17202 24256 17575
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24872 17134 24900 24511
rect 26804 23866 26832 27520
rect 26792 23860 26844 23866
rect 26792 23802 26844 23808
rect 25134 23488 25190 23497
rect 25134 23423 25190 23432
rect 25148 22778 25176 23423
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25148 22574 25176 22714
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 24952 18148 25004 18154
rect 24952 18090 25004 18096
rect 24860 17128 24912 17134
rect 24860 17070 24912 17076
rect 24964 16726 24992 18090
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25056 16998 25084 17682
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 22744 16720 22796 16726
rect 22744 16662 22796 16668
rect 22928 16720 22980 16726
rect 22928 16662 22980 16668
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24952 16720 25004 16726
rect 24952 16662 25004 16668
rect 22756 16250 22784 16662
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22940 16182 22968 16662
rect 24216 16516 24268 16522
rect 24216 16458 24268 16464
rect 22928 16176 22980 16182
rect 22928 16118 22980 16124
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22664 14958 22692 15098
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22848 14414 22876 15438
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22756 13938 22784 14350
rect 22940 14006 22968 16118
rect 24228 15910 24256 16458
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16250 24716 16662
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24216 15904 24268 15910
rect 24216 15846 24268 15852
rect 24228 15706 24256 15846
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 25056 15609 25084 16934
rect 25042 15600 25098 15609
rect 25042 15535 25098 15544
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 25410 15192 25466 15201
rect 25410 15127 25466 15136
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23020 14544 23072 14550
rect 23020 14486 23072 14492
rect 23032 14074 23060 14486
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22652 12912 22704 12918
rect 22652 12854 22704 12860
rect 22664 12288 22692 12854
rect 22756 12442 22784 13262
rect 22940 13258 22968 13942
rect 23204 13456 23256 13462
rect 23204 13398 23256 13404
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 23216 12986 23244 13398
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23110 12880 23166 12889
rect 23110 12815 23166 12824
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22744 12300 22796 12306
rect 22664 12260 22744 12288
rect 22744 12242 22796 12248
rect 22756 11762 22784 12242
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22940 10606 22968 12582
rect 23124 12374 23152 12815
rect 23112 12368 23164 12374
rect 23112 12310 23164 12316
rect 23124 11762 23152 12310
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 23112 11756 23164 11762
rect 23112 11698 23164 11704
rect 22928 10600 22980 10606
rect 22572 10526 22692 10554
rect 22928 10542 22980 10548
rect 22466 10503 22522 10512
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 22204 8838 22232 9318
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22204 7478 22232 8774
rect 22480 7954 22508 10503
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22572 10198 22600 10406
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 22664 9722 22692 10526
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22664 9518 22692 9658
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 23032 9450 23060 10202
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23124 9722 23152 10066
rect 23112 9716 23164 9722
rect 23112 9658 23164 9664
rect 23124 9586 23152 9658
rect 23216 9586 23244 11834
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23020 9444 23072 9450
rect 23020 9386 23072 9392
rect 22836 9104 22888 9110
rect 22836 9046 22888 9052
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22756 8634 22784 8910
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22756 8090 22784 8570
rect 22848 8498 22876 9046
rect 23032 8974 23060 9386
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 22744 8084 22796 8090
rect 22744 8026 22796 8032
rect 22848 8022 22876 8434
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22836 8016 22888 8022
rect 22836 7958 22888 7964
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 22192 6928 22244 6934
rect 22192 6870 22244 6876
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22112 5914 22140 6734
rect 22204 6390 22232 6870
rect 22192 6384 22244 6390
rect 22192 6326 22244 6332
rect 22284 6180 22336 6186
rect 22284 6122 22336 6128
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22296 5710 22324 6122
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22006 4584 22062 4593
rect 22006 4519 22062 4528
rect 22296 4214 22324 5646
rect 22480 5642 22508 7890
rect 22572 7546 22600 7958
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22468 5636 22520 5642
rect 22468 5578 22520 5584
rect 22572 5273 22600 7278
rect 22848 7002 22876 7686
rect 22940 7410 22968 7686
rect 23032 7546 23060 7890
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 23308 7342 23336 14894
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 25424 14074 25452 15127
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 23848 14000 23900 14006
rect 23848 13942 23900 13948
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23400 13462 23428 13874
rect 23860 13802 23888 13942
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23388 13456 23440 13462
rect 23388 13398 23440 13404
rect 23676 13190 23704 13670
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23676 12986 23704 13126
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 24674 12880 24730 12889
rect 24674 12815 24730 12824
rect 24688 12306 24716 12815
rect 24780 12646 24808 13330
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24676 12300 24728 12306
rect 24676 12242 24728 12248
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23768 11694 23796 12038
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11830 24716 12242
rect 24676 11824 24728 11830
rect 24676 11766 24728 11772
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 23572 11280 23624 11286
rect 23768 11257 23796 11630
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 23572 11222 23624 11228
rect 23754 11248 23810 11257
rect 23584 10810 23612 11222
rect 23754 11183 23810 11192
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23388 10532 23440 10538
rect 23388 10474 23440 10480
rect 23400 8974 23428 10474
rect 23768 10266 23796 11086
rect 24688 11014 24716 11494
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10810 24716 10950
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24216 10532 24268 10538
rect 24216 10474 24268 10480
rect 24228 10441 24256 10474
rect 24214 10432 24270 10441
rect 24214 10367 24270 10376
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23400 8634 23428 8910
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23664 7812 23716 7818
rect 23664 7754 23716 7760
rect 23676 7342 23704 7754
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23296 7336 23348 7342
rect 23664 7336 23716 7342
rect 23296 7278 23348 7284
rect 23584 7296 23664 7324
rect 22836 6996 22888 7002
rect 22836 6938 22888 6944
rect 23020 6724 23072 6730
rect 23020 6666 23072 6672
rect 22744 5840 22796 5846
rect 22744 5782 22796 5788
rect 22836 5840 22888 5846
rect 22836 5782 22888 5788
rect 22756 5370 22784 5782
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22558 5264 22614 5273
rect 22558 5199 22614 5208
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 22388 4758 22416 5102
rect 22376 4752 22428 4758
rect 22376 4694 22428 4700
rect 22388 4282 22416 4694
rect 22468 4548 22520 4554
rect 22468 4490 22520 4496
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22480 4146 22508 4490
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22480 2922 22508 3538
rect 22468 2916 22520 2922
rect 22468 2858 22520 2864
rect 22572 2582 22600 5199
rect 22848 5166 22876 5782
rect 23032 5710 23060 6666
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23124 6118 23152 6394
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23124 5914 23152 6054
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 23400 5234 23428 6054
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 22836 5160 22888 5166
rect 22836 5102 22888 5108
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22664 3670 22692 4422
rect 23032 4282 23060 4558
rect 23020 4276 23072 4282
rect 23020 4218 23072 4224
rect 22652 3664 22704 3670
rect 22652 3606 22704 3612
rect 22664 2854 22692 3606
rect 23584 3233 23612 7296
rect 23664 7278 23716 7284
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23676 6458 23704 6734
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23768 5302 23796 7346
rect 23860 7342 23888 7686
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23860 5574 23888 7278
rect 23848 5568 23900 5574
rect 23848 5510 23900 5516
rect 23756 5296 23808 5302
rect 23756 5238 23808 5244
rect 23768 4826 23796 5238
rect 23860 5234 23888 5510
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23860 5137 23888 5170
rect 23846 5128 23902 5137
rect 23846 5063 23902 5072
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23768 4486 23796 4762
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23952 4154 23980 9522
rect 24124 9104 24176 9110
rect 24124 9046 24176 9052
rect 24136 8362 24164 9046
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24124 8356 24176 8362
rect 24124 8298 24176 8304
rect 24216 8288 24268 8294
rect 24216 8230 24268 8236
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24122 7848 24178 7857
rect 24122 7783 24178 7792
rect 24136 7410 24164 7783
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24032 6928 24084 6934
rect 24032 6870 24084 6876
rect 24044 6186 24072 6870
rect 24122 6352 24178 6361
rect 24122 6287 24178 6296
rect 24032 6180 24084 6186
rect 24032 6122 24084 6128
rect 24044 5914 24072 6122
rect 24032 5908 24084 5914
rect 24032 5850 24084 5856
rect 24136 5234 24164 6287
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 23768 4126 23980 4154
rect 23570 3224 23626 3233
rect 23768 3194 23796 4126
rect 23848 3596 23900 3602
rect 23848 3538 23900 3544
rect 23570 3159 23626 3168
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23860 2854 23888 3538
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 22560 2576 22612 2582
rect 22560 2518 22612 2524
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21732 2508 21784 2514
rect 21732 2450 21784 2456
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 21456 2304 21508 2310
rect 21456 2246 21508 2252
rect 21468 1737 21496 2246
rect 21454 1728 21510 1737
rect 21454 1663 21510 1672
rect 20902 82 20958 480
rect 20732 54 20958 82
rect 13266 0 13322 54
rect 14554 0 14610 54
rect 15750 0 15806 54
rect 17038 0 17094 54
rect 18326 0 18382 54
rect 19614 0 19670 54
rect 20902 0 20958 54
rect 22098 82 22154 480
rect 22388 82 22416 2450
rect 22664 1193 22692 2790
rect 23020 2372 23072 2378
rect 23020 2314 23072 2320
rect 22650 1184 22706 1193
rect 22650 1119 22706 1128
rect 22098 54 22416 82
rect 23032 82 23060 2314
rect 23860 2009 23888 2790
rect 23846 2000 23902 2009
rect 23846 1935 23902 1944
rect 23386 82 23442 480
rect 23032 54 23442 82
rect 24228 82 24256 8230
rect 24688 7993 24716 8230
rect 24674 7984 24730 7993
rect 24674 7919 24730 7928
rect 24676 7880 24728 7886
rect 24780 7834 24808 12582
rect 24964 11898 24992 13806
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 25148 12238 25176 12718
rect 25228 12708 25280 12714
rect 25228 12650 25280 12656
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 25240 11937 25268 12650
rect 25226 11928 25282 11937
rect 24952 11892 25004 11898
rect 25226 11863 25282 11872
rect 24952 11834 25004 11840
rect 25240 11830 25268 11863
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 25148 8129 25176 9318
rect 25778 8256 25834 8265
rect 25778 8191 25834 8200
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 24728 7828 24808 7834
rect 24676 7822 24808 7828
rect 24688 7806 24808 7822
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7206 24716 7806
rect 25792 7546 25820 8191
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 25792 7342 25820 7482
rect 25780 7336 25832 7342
rect 25780 7278 25832 7284
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24400 6384 24452 6390
rect 24400 6326 24452 6332
rect 24412 5846 24440 6326
rect 24688 6225 24716 7142
rect 24780 6458 24808 7142
rect 25228 6860 25280 6866
rect 25228 6802 25280 6808
rect 25240 6458 25268 6802
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 27620 6452 27672 6458
rect 27620 6394 27672 6400
rect 27632 6361 27660 6394
rect 27618 6352 27674 6361
rect 27618 6287 27674 6296
rect 24674 6216 24730 6225
rect 24674 6151 24730 6160
rect 24860 6180 24912 6186
rect 24860 6122 24912 6128
rect 24400 5840 24452 5846
rect 24400 5782 24452 5788
rect 24676 5840 24728 5846
rect 24676 5782 24728 5788
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5370 24716 5782
rect 24872 5642 24900 6122
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24872 4554 24900 5578
rect 25056 5370 25084 5646
rect 25044 5364 25096 5370
rect 25044 5306 25096 5312
rect 27618 5264 27674 5273
rect 27618 5199 27674 5208
rect 27632 5166 27660 5199
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 24860 4548 24912 4554
rect 24860 4490 24912 4496
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 27618 4040 27674 4049
rect 27618 3975 27674 3984
rect 27632 3942 27660 3975
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 26884 2848 26936 2854
rect 26884 2790 26936 2796
rect 26056 2372 26108 2378
rect 26056 2314 26108 2320
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24674 82 24730 480
rect 24228 54 24730 82
rect 22098 0 22154 54
rect 23386 0 23442 54
rect 24674 0 24730 54
rect 25962 82 26018 480
rect 26068 82 26096 2314
rect 25962 54 26096 82
rect 26896 82 26924 2790
rect 27250 82 27306 480
rect 26896 54 27306 82
rect 25962 0 26018 54
rect 27250 0 27306 54
<< via2 >>
rect 1490 25880 1546 25936
rect 110 13368 166 13424
rect 110 12416 166 12472
rect 1398 23432 1454 23488
rect 1858 24656 1914 24712
rect 1582 22208 1638 22264
rect 1582 20984 1638 21040
rect 1582 16360 1638 16416
rect 1582 14184 1638 14240
rect 1674 12688 1730 12744
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5998 19352 6054 19408
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 3422 17448 3478 17504
rect 2134 10648 2190 10704
rect 1582 8200 1638 8256
rect 1582 7112 1638 7168
rect 1582 5888 1638 5944
rect 18 5208 74 5264
rect 110 2896 166 2952
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 4250 11600 4306 11656
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 2226 5616 2282 5672
rect 4066 3984 4122 4040
rect 3146 2352 3202 2408
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 8022 18944 8078 19000
rect 9586 26832 9642 26888
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 8942 18128 8998 18184
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9954 19760 10010 19816
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 9310 17720 9366 17776
rect 8298 17040 8354 17096
rect 6090 11600 6146 11656
rect 7654 10648 7710 10704
rect 8850 13776 8906 13832
rect 9034 12416 9090 12472
rect 8574 11736 8630 11792
rect 8390 10648 8446 10704
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 4526 5208 4582 5264
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5078 5072 5134 5128
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6826 4020 6828 4040
rect 6828 4020 6880 4040
rect 6880 4020 6882 4040
rect 6826 3984 6882 4020
rect 4342 2488 4398 2544
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 8206 4392 8262 4448
rect 8482 10512 8538 10568
rect 8390 4256 8446 4312
rect 6458 1944 6514 2000
rect 6918 2508 6974 2544
rect 6918 2488 6920 2508
rect 6920 2488 6972 2508
rect 6972 2488 6974 2508
rect 6918 1944 6974 2000
rect 8298 1400 8354 1456
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 9678 13368 9734 13424
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 11058 17720 11114 17776
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10690 10104 10746 10160
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 11334 15544 11390 15600
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 11702 17584 11758 17640
rect 8942 5752 8998 5808
rect 9402 6296 9458 6352
rect 9494 6160 9550 6216
rect 8942 4664 8998 4720
rect 9126 4664 9182 4720
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 9586 4020 9588 4040
rect 9588 4020 9640 4040
rect 9640 4020 9642 4040
rect 9586 3984 9642 4020
rect 10966 4800 11022 4856
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11610 5208 11666 5264
rect 11794 13368 11850 13424
rect 11794 10648 11850 10704
rect 13174 16088 13230 16144
rect 12254 15000 12310 15056
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 12530 5616 12586 5672
rect 13542 10104 13598 10160
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15658 16632 15714 16688
rect 15474 15408 15530 15464
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19982 22480 20038 22536
rect 16026 19352 16082 19408
rect 16210 18128 16266 18184
rect 16118 17040 16174 17096
rect 15842 13776 15898 13832
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15474 11600 15530 11656
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 13082 4800 13138 4856
rect 12162 1672 12218 1728
rect 14462 5208 14518 5264
rect 14554 5072 14610 5128
rect 14554 4528 14610 4584
rect 14462 4392 14518 4448
rect 14094 3032 14150 3088
rect 14002 2896 14058 2952
rect 14002 584 14058 640
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16762 12824 16818 12880
rect 16486 9968 16542 10024
rect 15382 3032 15438 3088
rect 17130 5752 17186 5808
rect 18326 13812 18328 13832
rect 18328 13812 18380 13832
rect 18380 13812 18382 13832
rect 18326 13776 18382 13812
rect 18602 12688 18658 12744
rect 18602 10104 18658 10160
rect 18786 11192 18842 11248
rect 18234 7928 18290 7984
rect 17590 6296 17646 6352
rect 16854 5072 16910 5128
rect 16670 4120 16726 4176
rect 15750 2352 15806 2408
rect 15290 1944 15346 2000
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19062 16088 19118 16144
rect 18970 12824 19026 12880
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 23202 26832 23258 26888
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19062 7792 19118 7848
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19338 6296 19394 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19522 5752 19578 5808
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 18050 3984 18106 4040
rect 16946 1944 17002 2000
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20994 17720 21050 17776
rect 22558 20984 22614 21040
rect 20902 11736 20958 11792
rect 20718 10512 20774 10568
rect 20534 4664 20590 4720
rect 19614 3168 19670 3224
rect 19430 2896 19486 2952
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 22466 10512 22522 10568
rect 22650 17720 22706 17776
rect 24214 25608 24270 25664
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24858 24520 24914 24576
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24766 19760 24822 19816
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24766 18672 24822 18728
rect 24214 17584 24270 17640
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 25134 23432 25190 23488
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 25042 15544 25098 15600
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 25410 15136 25466 15192
rect 23110 12824 23166 12880
rect 22006 4528 22062 4584
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24674 12824 24730 12880
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 23754 11192 23810 11248
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24214 10376 24270 10432
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 22558 5208 22614 5264
rect 23846 5072 23902 5128
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24122 7792 24178 7848
rect 24122 6296 24178 6352
rect 23570 3168 23626 3224
rect 21454 1672 21510 1728
rect 22650 1128 22706 1184
rect 23846 1944 23902 2000
rect 24674 7928 24730 7984
rect 25226 11872 25282 11928
rect 25778 8200 25834 8256
rect 25134 8064 25190 8120
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 27618 6296 27674 6352
rect 24674 6160 24730 6216
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 27618 5208 27674 5264
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 27618 3984 27674 4040
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
<< metal3 >>
rect 0 27344 480 27464
rect 27520 27344 28000 27464
rect 62 26890 122 27344
rect 9581 26890 9647 26893
rect 62 26888 9647 26890
rect 62 26832 9586 26888
rect 9642 26832 9647 26888
rect 62 26830 9647 26832
rect 9581 26827 9647 26830
rect 23197 26890 23263 26893
rect 27662 26890 27722 27344
rect 23197 26888 27722 26890
rect 23197 26832 23202 26888
rect 23258 26832 27722 26888
rect 23197 26830 27722 26832
rect 23197 26827 23263 26830
rect 0 26120 480 26240
rect 27520 26120 28000 26240
rect 62 25938 122 26120
rect 1485 25938 1551 25941
rect 62 25936 1551 25938
rect 62 25880 1490 25936
rect 1546 25880 1551 25936
rect 62 25878 1551 25880
rect 1485 25875 1551 25878
rect 24209 25666 24275 25669
rect 27662 25666 27722 26120
rect 24209 25664 27722 25666
rect 24209 25608 24214 25664
rect 24270 25608 27722 25664
rect 24209 25606 27722 25608
rect 24209 25603 24275 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25032 480 25152
rect 27520 25124 28000 25152
rect 27520 25060 27660 25124
rect 27724 25060 28000 25124
rect 5610 25056 5930 25057
rect 62 24714 122 25032
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 27520 25032 28000 25060
rect 24277 24991 24597 24992
rect 1853 24714 1919 24717
rect 62 24712 1919 24714
rect 62 24656 1858 24712
rect 1914 24656 1919 24712
rect 62 24654 1919 24656
rect 1853 24651 1919 24654
rect 24853 24578 24919 24581
rect 27654 24578 27660 24580
rect 24853 24576 27660 24578
rect 24853 24520 24858 24576
rect 24914 24520 27660 24576
rect 24853 24518 27660 24520
rect 24853 24515 24919 24518
rect 27654 24516 27660 24518
rect 27724 24516 27730 24580
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 5610 23968 5930 23969
rect 0 23808 480 23928
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 27520 23808 28000 23928
rect 62 23490 122 23808
rect 1393 23490 1459 23493
rect 62 23488 1459 23490
rect 62 23432 1398 23488
rect 1454 23432 1459 23488
rect 62 23430 1459 23432
rect 1393 23427 1459 23430
rect 25129 23490 25195 23493
rect 27662 23490 27722 23808
rect 25129 23488 27722 23490
rect 25129 23432 25134 23488
rect 25190 23432 27722 23488
rect 25129 23430 27722 23432
rect 25129 23427 25195 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 5610 22880 5930 22881
rect 0 22720 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 27520 22720 28000 22840
rect 62 22266 122 22720
rect 19977 22538 20043 22541
rect 27662 22538 27722 22720
rect 19977 22536 27722 22538
rect 19977 22480 19982 22536
rect 20038 22480 27722 22536
rect 19977 22478 27722 22480
rect 19977 22475 20043 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 1577 22266 1643 22269
rect 62 22264 1643 22266
rect 62 22208 1582 22264
rect 1638 22208 1643 22264
rect 62 22206 1643 22208
rect 1577 22203 1643 22206
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21496 480 21616
rect 27520 21496 28000 21616
rect 62 21042 122 21496
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1577 21042 1643 21045
rect 62 21040 1643 21042
rect 62 20984 1582 21040
rect 1638 20984 1643 21040
rect 62 20982 1643 20984
rect 1577 20979 1643 20982
rect 22553 21042 22619 21045
rect 27662 21042 27722 21496
rect 22553 21040 27722 21042
rect 22553 20984 22558 21040
rect 22614 20984 27722 21040
rect 22553 20982 27722 20984
rect 22553 20979 22619 20982
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 0 20272 480 20392
rect 27520 20272 28000 20392
rect 62 19818 122 20272
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 9949 19818 10015 19821
rect 62 19816 10015 19818
rect 62 19760 9954 19816
rect 10010 19760 10015 19816
rect 62 19758 10015 19760
rect 9949 19755 10015 19758
rect 24761 19818 24827 19821
rect 27662 19818 27722 20272
rect 24761 19816 27722 19818
rect 24761 19760 24766 19816
rect 24822 19760 27722 19816
rect 24761 19758 27722 19760
rect 24761 19755 24827 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 5993 19410 6059 19413
rect 16021 19410 16087 19413
rect 5993 19408 16087 19410
rect 5993 19352 5998 19408
rect 6054 19352 16026 19408
rect 16082 19352 16087 19408
rect 5993 19350 16087 19352
rect 5993 19347 6059 19350
rect 16021 19347 16087 19350
rect 0 19184 480 19304
rect 27520 19184 28000 19304
rect 62 19002 122 19184
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 8017 19002 8083 19005
rect 62 19000 8083 19002
rect 62 18944 8022 19000
rect 8078 18944 8083 19000
rect 62 18942 8083 18944
rect 8017 18939 8083 18942
rect 24761 18730 24827 18733
rect 27662 18730 27722 19184
rect 24761 18728 27722 18730
rect 24761 18672 24766 18728
rect 24822 18672 27722 18728
rect 24761 18670 27722 18672
rect 24761 18667 24827 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 8937 18186 9003 18189
rect 16205 18186 16271 18189
rect 8937 18184 16271 18186
rect 8937 18128 8942 18184
rect 8998 18128 16210 18184
rect 16266 18128 16271 18184
rect 8937 18126 16271 18128
rect 8937 18123 9003 18126
rect 16205 18123 16271 18126
rect 0 17960 480 18080
rect 10277 17984 10597 17985
rect 62 17506 122 17960
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 18080
rect 19610 17919 19930 17920
rect 9305 17778 9371 17781
rect 11053 17778 11119 17781
rect 20989 17778 21055 17781
rect 9305 17776 21055 17778
rect 9305 17720 9310 17776
rect 9366 17720 11058 17776
rect 11114 17720 20994 17776
rect 21050 17720 21055 17776
rect 9305 17718 21055 17720
rect 9305 17715 9371 17718
rect 11053 17715 11119 17718
rect 20989 17715 21055 17718
rect 22645 17778 22711 17781
rect 27662 17778 27722 17960
rect 22645 17776 27722 17778
rect 22645 17720 22650 17776
rect 22706 17720 27722 17776
rect 22645 17718 27722 17720
rect 22645 17715 22711 17718
rect 11697 17642 11763 17645
rect 24209 17642 24275 17645
rect 11697 17640 24275 17642
rect 11697 17584 11702 17640
rect 11758 17584 24214 17640
rect 24270 17584 24275 17640
rect 11697 17582 24275 17584
rect 11697 17579 11763 17582
rect 24209 17579 24275 17582
rect 3417 17506 3483 17509
rect 62 17504 3483 17506
rect 62 17448 3422 17504
rect 3478 17448 3483 17504
rect 62 17446 3483 17448
rect 3417 17443 3483 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 8293 17098 8359 17101
rect 16113 17098 16179 17101
rect 8293 17096 16179 17098
rect 8293 17040 8298 17096
rect 8354 17040 16118 17096
rect 16174 17040 16179 17096
rect 8293 17038 16179 17040
rect 8293 17035 8359 17038
rect 16113 17035 16179 17038
rect 0 16872 480 16992
rect 10277 16896 10597 16897
rect 62 16418 122 16872
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 27520 16872 28000 16992
rect 19610 16831 19930 16832
rect 15653 16690 15719 16693
rect 27662 16690 27722 16872
rect 15653 16688 27722 16690
rect 15653 16632 15658 16688
rect 15714 16632 27722 16688
rect 15653 16630 27722 16632
rect 15653 16627 15719 16630
rect 1577 16418 1643 16421
rect 62 16416 1643 16418
rect 62 16360 1582 16416
rect 1638 16360 1643 16416
rect 62 16358 1643 16360
rect 1577 16355 1643 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 13169 16146 13235 16149
rect 19057 16146 19123 16149
rect 13169 16144 19123 16146
rect 13169 16088 13174 16144
rect 13230 16088 19062 16144
rect 19118 16088 19123 16144
rect 13169 16086 19123 16088
rect 13169 16083 13235 16086
rect 19057 16083 19123 16086
rect 10277 15808 10597 15809
rect 0 15648 480 15768
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 27520 15648 28000 15768
rect 62 15466 122 15648
rect 11329 15602 11395 15605
rect 25037 15602 25103 15605
rect 11329 15600 25103 15602
rect 11329 15544 11334 15600
rect 11390 15544 25042 15600
rect 25098 15544 25103 15600
rect 11329 15542 25103 15544
rect 11329 15539 11395 15542
rect 25037 15539 25103 15542
rect 15469 15466 15535 15469
rect 62 15464 15535 15466
rect 62 15408 15474 15464
rect 15530 15408 15535 15464
rect 62 15406 15535 15408
rect 15469 15403 15535 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 25405 15194 25471 15197
rect 27662 15194 27722 15648
rect 25405 15192 27722 15194
rect 25405 15136 25410 15192
rect 25466 15136 27722 15192
rect 25405 15134 27722 15136
rect 25405 15131 25471 15134
rect 12249 15058 12315 15061
rect 12249 15056 27722 15058
rect 12249 15000 12254 15056
rect 12310 15000 27722 15056
rect 12249 14998 27722 15000
rect 12249 14995 12315 14998
rect 10277 14720 10597 14721
rect 0 14560 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 27662 14680 27722 14998
rect 19610 14655 19930 14656
rect 27520 14560 28000 14680
rect 62 14242 122 14560
rect 1577 14242 1643 14245
rect 62 14240 1643 14242
rect 62 14184 1582 14240
rect 1638 14184 1643 14240
rect 62 14182 1643 14184
rect 1577 14179 1643 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 8845 13834 8911 13837
rect 15837 13834 15903 13837
rect 18321 13834 18387 13837
rect 8845 13832 18387 13834
rect 8845 13776 8850 13832
rect 8906 13776 15842 13832
rect 15898 13776 18326 13832
rect 18382 13776 18387 13832
rect 8845 13774 18387 13776
rect 8845 13771 8911 13774
rect 15837 13771 15903 13774
rect 18321 13771 18387 13774
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 0 13424 480 13456
rect 0 13368 110 13424
rect 166 13368 480 13424
rect 0 13336 480 13368
rect 9673 13426 9739 13429
rect 11789 13426 11855 13429
rect 9673 13424 11855 13426
rect 9673 13368 9678 13424
rect 9734 13368 11794 13424
rect 11850 13368 11855 13424
rect 9673 13366 11855 13368
rect 9673 13363 9739 13366
rect 11789 13363 11855 13366
rect 27520 13336 28000 13456
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 16757 12882 16823 12885
rect 18965 12882 19031 12885
rect 23105 12882 23171 12885
rect 16757 12880 23171 12882
rect 16757 12824 16762 12880
rect 16818 12824 18970 12880
rect 19026 12824 23110 12880
rect 23166 12824 23171 12880
rect 16757 12822 23171 12824
rect 16757 12819 16823 12822
rect 18965 12819 19031 12822
rect 23105 12819 23171 12822
rect 24669 12882 24735 12885
rect 27662 12882 27722 13336
rect 24669 12880 27722 12882
rect 24669 12824 24674 12880
rect 24730 12824 27722 12880
rect 24669 12822 27722 12824
rect 24669 12819 24735 12822
rect 1669 12746 1735 12749
rect 18597 12746 18663 12749
rect 1669 12744 18663 12746
rect 1669 12688 1674 12744
rect 1730 12688 18602 12744
rect 18658 12688 18663 12744
rect 1669 12686 18663 12688
rect 1669 12683 1735 12686
rect 18597 12683 18663 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 105 12474 171 12477
rect 9029 12474 9095 12477
rect 105 12472 9095 12474
rect 105 12416 110 12472
rect 166 12416 9034 12472
rect 9090 12416 9095 12472
rect 105 12414 9095 12416
rect 105 12411 171 12414
rect 9029 12411 9095 12414
rect 0 12112 480 12232
rect 27520 12112 28000 12232
rect 62 11658 122 12112
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 25221 11930 25287 11933
rect 27662 11930 27722 12112
rect 25221 11928 27722 11930
rect 25221 11872 25226 11928
rect 25282 11872 27722 11928
rect 25221 11870 27722 11872
rect 25221 11867 25287 11870
rect 8569 11794 8635 11797
rect 20897 11794 20963 11797
rect 8569 11792 20963 11794
rect 8569 11736 8574 11792
rect 8630 11736 20902 11792
rect 20958 11736 20963 11792
rect 8569 11734 20963 11736
rect 8569 11731 8635 11734
rect 20897 11731 20963 11734
rect 4245 11658 4311 11661
rect 62 11656 4311 11658
rect 62 11600 4250 11656
rect 4306 11600 4311 11656
rect 62 11598 4311 11600
rect 4245 11595 4311 11598
rect 6085 11658 6151 11661
rect 15469 11658 15535 11661
rect 6085 11656 15535 11658
rect 6085 11600 6090 11656
rect 6146 11600 15474 11656
rect 15530 11600 15535 11656
rect 6085 11598 15535 11600
rect 6085 11595 6151 11598
rect 15469 11595 15535 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 18781 11250 18847 11253
rect 23749 11250 23815 11253
rect 18781 11248 23815 11250
rect 18781 11192 18786 11248
rect 18842 11192 23754 11248
rect 23810 11192 23815 11248
rect 18781 11190 23815 11192
rect 18781 11187 18847 11190
rect 23749 11187 23815 11190
rect 0 11024 480 11144
rect 27520 11024 28000 11144
rect 62 10706 122 11024
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 2129 10706 2195 10709
rect 7649 10706 7715 10709
rect 8385 10706 8451 10709
rect 62 10704 8451 10706
rect 62 10648 2134 10704
rect 2190 10648 7654 10704
rect 7710 10648 8390 10704
rect 8446 10648 8451 10704
rect 62 10646 8451 10648
rect 2129 10643 2195 10646
rect 7649 10643 7715 10646
rect 8385 10643 8451 10646
rect 11789 10706 11855 10709
rect 27662 10706 27722 11024
rect 11789 10704 27722 10706
rect 11789 10648 11794 10704
rect 11850 10648 27722 10704
rect 11789 10646 27722 10648
rect 11789 10643 11855 10646
rect 8477 10570 8543 10573
rect 20713 10570 20779 10573
rect 22461 10570 22527 10573
rect 8477 10568 22527 10570
rect 8477 10512 8482 10568
rect 8538 10512 20718 10568
rect 20774 10512 22466 10568
rect 22522 10512 22527 10568
rect 8477 10510 22527 10512
rect 8477 10507 8543 10510
rect 20713 10507 20779 10510
rect 22461 10507 22527 10510
rect 24209 10434 24275 10437
rect 24209 10432 27722 10434
rect 24209 10376 24214 10432
rect 24270 10376 27722 10432
rect 24209 10374 27722 10376
rect 24209 10371 24275 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 54 10100 60 10164
rect 124 10162 130 10164
rect 124 10102 674 10162
rect 124 10100 130 10102
rect 614 10026 674 10102
rect 9254 10100 9260 10164
rect 9324 10162 9330 10164
rect 10685 10162 10751 10165
rect 9324 10160 10751 10162
rect 9324 10104 10690 10160
rect 10746 10104 10751 10160
rect 9324 10102 10751 10104
rect 9324 10100 9330 10102
rect 10685 10099 10751 10102
rect 13537 10162 13603 10165
rect 18597 10162 18663 10165
rect 13537 10160 18663 10162
rect 13537 10104 13542 10160
rect 13598 10104 18602 10160
rect 18658 10104 18663 10160
rect 13537 10102 18663 10104
rect 13537 10099 13603 10102
rect 18597 10099 18663 10102
rect 16481 10026 16547 10029
rect 614 10024 16547 10026
rect 614 9968 16486 10024
rect 16542 9968 16547 10024
rect 614 9966 16547 9968
rect 16481 9963 16547 9966
rect 27662 9920 27722 10374
rect 0 9892 480 9920
rect 0 9828 60 9892
rect 124 9828 480 9892
rect 0 9800 480 9828
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9920
rect 24277 9759 24597 9760
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 0 8712 480 8832
rect 5610 8736 5930 8737
rect 62 8258 122 8712
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8832
rect 24277 8671 24597 8672
rect 1577 8258 1643 8261
rect 62 8256 1643 8258
rect 62 8200 1582 8256
rect 1638 8200 1643 8256
rect 62 8198 1643 8200
rect 1577 8195 1643 8198
rect 25773 8258 25839 8261
rect 27662 8258 27722 8712
rect 25773 8256 27722 8258
rect 25773 8200 25778 8256
rect 25834 8200 27722 8256
rect 25773 8198 27722 8200
rect 25773 8195 25839 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 25129 8122 25195 8125
rect 25129 8120 27722 8122
rect 25129 8064 25134 8120
rect 25190 8064 27722 8120
rect 25129 8062 27722 8064
rect 25129 8059 25195 8062
rect 18229 7986 18295 7989
rect 24669 7986 24735 7989
rect 18229 7984 24735 7986
rect 18229 7928 18234 7984
rect 18290 7928 24674 7984
rect 24730 7928 24735 7984
rect 18229 7926 24735 7928
rect 18229 7923 18295 7926
rect 24669 7923 24735 7926
rect 19057 7850 19123 7853
rect 24117 7850 24183 7853
rect 19057 7848 24183 7850
rect 19057 7792 19062 7848
rect 19118 7792 24122 7848
rect 24178 7792 24183 7848
rect 19057 7790 24183 7792
rect 19057 7787 19123 7790
rect 24117 7787 24183 7790
rect 5610 7648 5930 7649
rect 0 7488 480 7608
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27662 7608 27722 8062
rect 24277 7583 24597 7584
rect 27520 7488 28000 7608
rect 62 7170 122 7488
rect 1577 7170 1643 7173
rect 62 7168 1643 7170
rect 62 7112 1582 7168
rect 1638 7112 1643 7168
rect 62 7110 1643 7112
rect 1577 7107 1643 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6264 480 6384
rect 9397 6354 9463 6357
rect 17585 6354 17651 6357
rect 9397 6352 17651 6354
rect 9397 6296 9402 6352
rect 9458 6296 17590 6352
rect 17646 6296 17651 6352
rect 9397 6294 17651 6296
rect 9397 6291 9463 6294
rect 17585 6291 17651 6294
rect 19333 6354 19399 6357
rect 24117 6354 24183 6357
rect 19333 6352 24183 6354
rect 19333 6296 19338 6352
rect 19394 6296 24122 6352
rect 24178 6296 24183 6352
rect 19333 6294 24183 6296
rect 19333 6291 19399 6294
rect 24117 6291 24183 6294
rect 27520 6352 28000 6384
rect 27520 6296 27618 6352
rect 27674 6296 28000 6352
rect 27520 6264 28000 6296
rect 62 5946 122 6264
rect 9489 6218 9555 6221
rect 24669 6218 24735 6221
rect 9489 6216 24735 6218
rect 9489 6160 9494 6216
rect 9550 6160 24674 6216
rect 24730 6160 24735 6216
rect 9489 6158 24735 6160
rect 9489 6155 9555 6158
rect 24669 6155 24735 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 1577 5946 1643 5949
rect 62 5944 1643 5946
rect 62 5888 1582 5944
rect 1638 5888 1643 5944
rect 62 5886 1643 5888
rect 1577 5883 1643 5886
rect 8937 5810 9003 5813
rect 17125 5810 17191 5813
rect 19517 5810 19583 5813
rect 8937 5808 19583 5810
rect 8937 5752 8942 5808
rect 8998 5752 17130 5808
rect 17186 5752 19522 5808
rect 19578 5752 19583 5808
rect 8937 5750 19583 5752
rect 8937 5747 9003 5750
rect 17125 5747 17191 5750
rect 19517 5747 19583 5750
rect 2221 5674 2287 5677
rect 12525 5674 12591 5677
rect 2221 5672 12591 5674
rect 2221 5616 2226 5672
rect 2282 5616 12530 5672
rect 12586 5616 12591 5672
rect 2221 5614 12591 5616
rect 2221 5611 2287 5614
rect 12525 5611 12591 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 0 5264 480 5296
rect 0 5208 18 5264
rect 74 5208 480 5264
rect 0 5176 480 5208
rect 4521 5266 4587 5269
rect 11605 5266 11671 5269
rect 4521 5264 11671 5266
rect 4521 5208 4526 5264
rect 4582 5208 11610 5264
rect 11666 5208 11671 5264
rect 4521 5206 11671 5208
rect 4521 5203 4587 5206
rect 11605 5203 11671 5206
rect 14457 5266 14523 5269
rect 22553 5266 22619 5269
rect 14457 5264 22619 5266
rect 14457 5208 14462 5264
rect 14518 5208 22558 5264
rect 22614 5208 22619 5264
rect 14457 5206 22619 5208
rect 14457 5203 14523 5206
rect 22553 5203 22619 5206
rect 27520 5264 28000 5296
rect 27520 5208 27618 5264
rect 27674 5208 28000 5264
rect 27520 5176 28000 5208
rect 5073 5130 5139 5133
rect 14549 5130 14615 5133
rect 5073 5128 14615 5130
rect 5073 5072 5078 5128
rect 5134 5072 14554 5128
rect 14610 5072 14615 5128
rect 5073 5070 14615 5072
rect 5073 5067 5139 5070
rect 14549 5067 14615 5070
rect 16849 5130 16915 5133
rect 23841 5130 23907 5133
rect 16849 5128 23907 5130
rect 16849 5072 16854 5128
rect 16910 5072 23846 5128
rect 23902 5072 23907 5128
rect 16849 5070 23907 5072
rect 16849 5067 16915 5070
rect 23841 5067 23907 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 10961 4858 11027 4861
rect 13077 4858 13143 4861
rect 10961 4856 15946 4858
rect 10961 4800 10966 4856
rect 11022 4800 13082 4856
rect 13138 4800 15946 4856
rect 10961 4798 15946 4800
rect 10961 4795 11027 4798
rect 13077 4795 13143 4798
rect 8937 4722 9003 4725
rect 62 4720 9003 4722
rect 62 4664 8942 4720
rect 8998 4664 9003 4720
rect 62 4662 9003 4664
rect 62 4072 122 4662
rect 8937 4659 9003 4662
rect 9121 4722 9187 4725
rect 15886 4722 15946 4798
rect 20529 4722 20595 4725
rect 9121 4720 13830 4722
rect 9121 4664 9126 4720
rect 9182 4664 13830 4720
rect 9121 4662 13830 4664
rect 15886 4720 20595 4722
rect 15886 4664 20534 4720
rect 20590 4664 20595 4720
rect 15886 4662 20595 4664
rect 9121 4659 9187 4662
rect 13770 4586 13830 4662
rect 20529 4659 20595 4662
rect 14549 4586 14615 4589
rect 22001 4586 22067 4589
rect 13770 4584 22067 4586
rect 13770 4528 14554 4584
rect 14610 4528 22006 4584
rect 22062 4528 22067 4584
rect 13770 4526 22067 4528
rect 14549 4523 14615 4526
rect 22001 4523 22067 4526
rect 8201 4450 8267 4453
rect 14457 4450 14523 4453
rect 8201 4448 14523 4450
rect 8201 4392 8206 4448
rect 8262 4392 14462 4448
rect 14518 4392 14523 4448
rect 8201 4390 14523 4392
rect 8201 4387 8267 4390
rect 14457 4387 14523 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 8385 4314 8451 4317
rect 8385 4312 13830 4314
rect 8385 4256 8390 4312
rect 8446 4256 13830 4312
rect 8385 4254 13830 4256
rect 8385 4251 8451 4254
rect 13770 4178 13830 4254
rect 16665 4178 16731 4181
rect 13770 4176 16731 4178
rect 13770 4120 16670 4176
rect 16726 4120 16731 4176
rect 13770 4118 16731 4120
rect 16665 4115 16731 4118
rect 0 3952 480 4072
rect 4061 4042 4127 4045
rect 6821 4042 6887 4045
rect 9581 4042 9647 4045
rect 18045 4042 18111 4045
rect 4061 4040 6746 4042
rect 4061 3984 4066 4040
rect 4122 3984 6746 4040
rect 4061 3982 6746 3984
rect 4061 3979 4127 3982
rect 6686 3906 6746 3982
rect 6821 4040 9647 4042
rect 6821 3984 6826 4040
rect 6882 3984 9586 4040
rect 9642 3984 9647 4040
rect 6821 3982 9647 3984
rect 6821 3979 6887 3982
rect 9581 3979 9647 3982
rect 9814 4040 18111 4042
rect 9814 3984 18050 4040
rect 18106 3984 18111 4040
rect 9814 3982 18111 3984
rect 9254 3906 9260 3908
rect 6686 3846 9260 3906
rect 9254 3844 9260 3846
rect 9324 3906 9330 3908
rect 9814 3906 9874 3982
rect 18045 3979 18111 3982
rect 27520 4040 28000 4072
rect 27520 3984 27618 4040
rect 27674 3984 28000 4040
rect 27520 3952 28000 3984
rect 9324 3846 9874 3906
rect 9324 3844 9330 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 19609 3226 19675 3229
rect 23565 3226 23631 3229
rect 27654 3226 27660 3228
rect 19609 3224 23631 3226
rect 19609 3168 19614 3224
rect 19670 3168 23570 3224
rect 23626 3168 23631 3224
rect 19609 3166 23631 3168
rect 19609 3163 19675 3166
rect 23565 3163 23631 3166
rect 27294 3166 27660 3226
rect 14089 3090 14155 3093
rect 15377 3090 15443 3093
rect 27294 3090 27354 3166
rect 27654 3164 27660 3166
rect 27724 3164 27730 3228
rect 14089 3088 27354 3090
rect 14089 3032 14094 3088
rect 14150 3032 15382 3088
rect 15438 3032 27354 3088
rect 14089 3030 27354 3032
rect 14089 3027 14155 3030
rect 15377 3027 15443 3030
rect 0 2952 480 2984
rect 0 2896 110 2952
rect 166 2896 480 2952
rect 0 2864 480 2896
rect 13997 2954 14063 2957
rect 19425 2954 19491 2957
rect 13997 2952 19491 2954
rect 13997 2896 14002 2952
rect 14058 2896 19430 2952
rect 19486 2896 19491 2952
rect 13997 2894 19491 2896
rect 13997 2891 14063 2894
rect 19425 2891 19491 2894
rect 27520 2956 28000 2984
rect 27520 2892 27660 2956
rect 27724 2892 28000 2956
rect 27520 2864 28000 2892
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 4337 2546 4403 2549
rect 6913 2546 6979 2549
rect 4337 2544 6979 2546
rect 4337 2488 4342 2544
rect 4398 2488 6918 2544
rect 6974 2488 6979 2544
rect 4337 2486 6979 2488
rect 4337 2483 4403 2486
rect 6913 2483 6979 2486
rect 3141 2410 3207 2413
rect 15745 2410 15811 2413
rect 3141 2408 15811 2410
rect 3141 2352 3146 2408
rect 3202 2352 15750 2408
rect 15806 2352 15811 2408
rect 3141 2350 15811 2352
rect 3141 2347 3207 2350
rect 15745 2347 15811 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6453 2002 6519 2005
rect 62 2000 6519 2002
rect 62 1944 6458 2000
rect 6514 1944 6519 2000
rect 62 1942 6519 1944
rect 62 1760 122 1942
rect 6453 1939 6519 1942
rect 6913 2002 6979 2005
rect 15285 2002 15351 2005
rect 6913 2000 15351 2002
rect 6913 1944 6918 2000
rect 6974 1944 15290 2000
rect 15346 1944 15351 2000
rect 6913 1942 15351 1944
rect 6913 1939 6979 1942
rect 15285 1939 15351 1942
rect 16941 2002 17007 2005
rect 23841 2002 23907 2005
rect 16941 2000 23907 2002
rect 16941 1944 16946 2000
rect 17002 1944 23846 2000
rect 23902 1944 23907 2000
rect 16941 1942 23907 1944
rect 16941 1939 17007 1942
rect 23841 1939 23907 1942
rect 0 1640 480 1760
rect 12157 1730 12223 1733
rect 21449 1730 21515 1733
rect 12157 1728 21515 1730
rect 12157 1672 12162 1728
rect 12218 1672 21454 1728
rect 21510 1672 21515 1728
rect 12157 1670 21515 1672
rect 12157 1667 12223 1670
rect 21449 1667 21515 1670
rect 27520 1640 28000 1760
rect 8293 1458 8359 1461
rect 27662 1458 27722 1640
rect 8293 1456 27722 1458
rect 8293 1400 8298 1456
rect 8354 1400 27722 1456
rect 8293 1398 27722 1400
rect 8293 1395 8359 1398
rect 22645 1186 22711 1189
rect 22645 1184 27722 1186
rect 22645 1128 22650 1184
rect 22706 1128 27722 1184
rect 22645 1126 27722 1128
rect 22645 1123 22711 1126
rect 54 852 60 916
rect 124 914 130 916
rect 124 854 9690 914
rect 124 852 130 854
rect 0 644 480 672
rect 0 580 60 644
rect 124 580 480 644
rect 9630 642 9690 854
rect 27662 672 27722 1126
rect 13997 642 14063 645
rect 9630 640 14063 642
rect 9630 584 14002 640
rect 14058 584 14063 640
rect 9630 582 14063 584
rect 0 552 480 580
rect 13997 579 14063 582
rect 27520 552 28000 672
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 27660 25060 27724 25124
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 27660 24516 27724 24580
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 60 10100 124 10164
rect 9260 10100 9324 10164
rect 60 9828 124 9892
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 9260 3844 9324 3908
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 27660 3164 27724 3228
rect 27660 2892 27724 2956
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 60 852 124 916
rect 60 580 124 644
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 59 10164 125 10165
rect 59 10100 60 10164
rect 124 10100 125 10164
rect 59 10099 125 10100
rect 62 9893 122 10099
rect 59 9892 125 9893
rect 59 9828 60 9892
rect 124 9828 125 9892
rect 59 9827 125 9828
rect 5610 9824 5931 10848
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9259 10164 9325 10165
rect 9259 10100 9260 10164
rect 9324 10100 9325 10164
rect 9259 10099 9325 10100
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 9262 3909 9322 10099
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 9259 3908 9325 3909
rect 9259 3844 9260 3908
rect 9324 3844 9325 3908
rect 9259 3843 9325 3844
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 27659 25124 27725 25125
rect 27659 25060 27660 25124
rect 27724 25060 27725 25124
rect 27659 25059 27725 25060
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 27662 24581 27722 25059
rect 27659 24580 27725 24581
rect 27659 24516 27660 24580
rect 27724 24516 27725 24580
rect 27659 24515 27725 24516
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 27659 3228 27725 3229
rect 27659 3164 27660 3228
rect 27724 3164 27725 3228
rect 27659 3163 27725 3164
rect 27662 2957 27722 3163
rect 27659 2956 27725 2957
rect 27659 2892 27660 2956
rect 27724 2892 27725 2956
rect 27659 2891 27725 2892
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 59 916 125 917
rect 59 852 60 916
rect 124 852 125 916
rect 59 851 125 852
rect 62 645 122 851
rect 59 644 125 645
rect 59 580 60 644
rect 124 580 125 644
rect 59 579 125 580
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_10
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_22
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_19 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__C
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _058_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _056_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__C
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _169_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_or3_4  _095_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_78
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_82
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 866 592
use scs8hd_or3_4  _087_
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9844 0 -1 2720
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_110
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_120
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_137
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__C
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_nor4_4  _125_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 1602 592
use scs8hd_buf_2  _159_
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__D
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_158
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_162
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_167
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_171
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _145_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _162_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_222
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__C
timestamp 1586364061
transform 1 0 21344 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_231
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_227
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _175_
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 406 592
use scs8hd_or3_4  _077_
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_235
timestamp 1586364061
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_238
timestamp 1586364061
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_243
timestamp 1586364061
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_239
timestamp 1586364061
transform 1 0 23092 0 1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_0_242 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_1_249
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _171_
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_262
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_274
timestamp 1586364061
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_or3_4  _074_
timestamp 1586364061
transform 1 0 4508 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_50
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_8  _057_
timestamp 1586364061
transform 1 0 6072 0 -1 3808
box -38 -48 866 592
use scs8hd_or3_4  _110_
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_63
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _130_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_110
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_114
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _064_
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_165
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _060_
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_203
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_207
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_or3_4  _085_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_235 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22724 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_246
timestamp 1586364061
transform 1 0 23736 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_270
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_8  _053_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _127_
timestamp 1586364061
transform 1 0 6900 0 1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__C
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__D
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_84
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 130 592
use scs8hd_nor4_4  _129_
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_91
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _126_
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_137
timestamp 1586364061
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_158
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_210
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_253
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_262
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_274
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_55
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_74
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_conb_1  _147_
timestamp 1586364061
transform 1 0 9752 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__D
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_101
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _063_
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_118
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _167_
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_135
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_151
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_157
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_8  _059_
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 15916 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_174
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_188
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_192
timestamp 1586364061
transform 1 0 18768 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_196
timestamp 1586364061
transform 1 0 19136 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_212
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21344 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_218
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_222
timestamp 1586364061
transform 1 0 21528 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_226
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_238
timestamp 1586364061
transform 1 0 23000 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_244
timestamp 1586364061
transform 1 0 23552 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_259
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_271
timestamp 1586364061
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_9
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_13
timestamp 1586364061
transform 1 0 2300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_25
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_33
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 314 592
use scs8hd_inv_8  _061_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_inv_8  _054_
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_76
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_80
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 314 592
use scs8hd_inv_8  _068_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_97
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_137
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_141
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 130 592
use scs8hd_inv_8  _051_
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_163
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_180
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_201
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_205
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 314 592
use scs8hd_conb_1  _139_
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 406 592
use scs8hd_or3_4  _081_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__081__C
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_265
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 314 592
use scs8hd_buf_2  _158_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_9
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_13
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_11
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_7_25
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_43
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_39
timestamp 1586364061
transform 1 0 4692 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _062_
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_73
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_78
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_77
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_85
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_conb_1  _146_
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_89
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _133_
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__C
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_114
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _067_
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__C
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_131
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_148
timestamp 1586364061
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_157
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_160
timestamp 1586364061
transform 1 0 15824 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__C
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_165
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_161
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_174
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_170
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_189
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_193
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_199
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_214
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_226
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_230
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_231
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_235
timestamp 1586364061
transform 1 0 22724 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_243
timestamp 1586364061
transform 1 0 23460 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_260
timestamp 1586364061
transform 1 0 25024 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _154_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _134_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__D
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__D
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_114
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use scs8hd_or3_4  _073_
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_131
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 314 592
use scs8hd_or3_4  _103_
timestamp 1586364061
transform 1 0 15364 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_164
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_168
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_172
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_192
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 590 592
use scs8hd_conb_1  _141_
timestamp 1586364061
transform 1 0 20976 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_219
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23552 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_236
timestamp 1586364061
transform 1 0 22816 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25116 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_253
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_8  FILLER_8_264
timestamp 1586364061
transform 1 0 25392 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_272
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_44
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6900 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use scs8hd_inv_8  _052_
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__C
timestamp 1586364061
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_78
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_96
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_or3_4  _111_
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_145
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__C
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_166
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_200
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_213
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_or3_4  _079_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_265
timestamp 1586364061
transform 1 0 25484 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_buf_2  _152_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use scs8hd_nor4_4  _128_
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__132__C
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__D
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_58
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_79
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_85
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_or3_4  _118_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__C
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use scs8hd_nor4_4  _137_
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_10_108
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _070_
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_168
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_185
timestamp 1586364061
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_209
timestamp 1586364061
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_219
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_223
timestamp 1586364061
transform 1 0 21620 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23276 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 23736 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_233
timestamp 1586364061
transform 1 0 22540 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_237
timestamp 1586364061
transform 1 0 22908 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_244
timestamp 1586364061
transform 1 0 23552 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_248
timestamp 1586364061
transform 1 0 23920 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24288 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__C
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_255
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_45
timestamp 1586364061
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_49
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _131_
timestamp 1586364061
transform 1 0 6900 0 1 8160
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_84
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 406 592
use scs8hd_or3_4  _088_
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__D
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _055_
timestamp 1586364061
transform 1 0 12512 0 1 8160
box -38 -48 866 592
use scs8hd_conb_1  _143_
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 130 592
use scs8hd_nor4_4  _136_
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__136__D
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_133
timestamp 1586364061
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_137
timestamp 1586364061
transform 1 0 13708 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_163
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_170
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_194
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_198
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_230
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _173_
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_249
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 24196 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_253
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_260
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_264
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_52
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _132_
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__131__C
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 6072 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_77
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 130 592
use scs8hd_nor4_4  _138_
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 1602 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__C
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_98
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_123
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_130
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__C
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17388 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_173
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_207
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_12_226
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_243
timestamp 1586364061
transform 1 0 23460 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_12_260
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_272
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_73
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_87
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _140_
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_109
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _148_
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_nor4_4  _135_
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_139
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 314 592
use scs8hd_or3_4  _096_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__D
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_148
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_163
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__C
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_184
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_180
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_188
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_201
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22080 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_224
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_230
timestamp 1586364061
transform 1 0 22264 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_8  _069_
timestamp 1586364061
transform 1 0 23000 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_235
timestamp 1586364061
transform 1 0 22724 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_253
timestamp 1586364061
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_262
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_274
timestamp 1586364061
transform 1 0 26312 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 130 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_15_81
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_85
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_126
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_130
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_201
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_215
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_219
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_234
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_238
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_248
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_252
timestamp 1586364061
transform 1 0 24288 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_256
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_268
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_37
timestamp 1586364061
transform 1 0 4508 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_54
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_58
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_99
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_103
timestamp 1586364061
transform 1 0 10580 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_116
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_175
timestamp 1586364061
transform 1 0 17204 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21804 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21620 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_220
timestamp 1586364061
transform 1 0 21344 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_234
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 774 592
use scs8hd_inv_8  _066_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_90
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_109
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_128
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _168_
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_216
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 23092 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_233
timestamp 1586364061
transform 1 0 22540 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_237
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_241
timestamp 1586364061
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_248
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24288 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_263
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_18
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_52
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_63
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_104
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_143
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_147
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_158
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_174
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_191
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_195
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_18_207
timestamp 1586364061
transform 1 0 20148 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_231
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22540 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_244
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_248
timestamp 1586364061
transform 1 0 23920 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_255
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_267
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_2  _165_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_31
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_conb_1  _142_
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_43
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_49
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_50
timestamp 1586364061
transform 1 0 5704 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_70
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_87
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_96
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_100
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_104
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_100
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_108
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_124
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_127
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_6  FILLER_20_146
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_143
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_157
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_176
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_169
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_192
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_190
timestamp 1586364061
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 18952 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_210
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_223
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_227
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_226
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_238
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_243
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_248
timestamp 1586364061
transform 1 0 23920 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_242
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_252
timestamp 1586364061
transform 1 0 24288 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_266
timestamp 1586364061
transform 1 0 25576 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_254
timestamp 1586364061
transform 1 0 24472 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_19
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_43
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_78
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_140
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20148 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_199
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_203
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_218
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_222
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _156_
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 406 592
use scs8hd_decap_8  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_266
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_270
timestamp 1586364061
transform 1 0 25944 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use scs8hd_buf_2  _161_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 590 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 17388 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17204 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_169
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_173
timestamp 1586364061
transform 1 0 17020 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 19136 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_188
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_192
timestamp 1586364061
transform 1 0 18768 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_205
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_209
timestamp 1586364061
transform 1 0 20332 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_22_226
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_243
timestamp 1586364061
transform 1 0 23460 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_255
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_267
timestamp 1586364061
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_70
timestamp 1586364061
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_83
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_102
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_106
timestamp 1586364061
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_127
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_142
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _164_
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_146
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20332 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_205
timestamp 1586364061
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_224
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_235
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_243
timestamp 1586364061
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_116
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_120
timestamp 1586364061
transform 1 0 12144 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_139
timestamp 1586364061
transform 1 0 13892 0 -1 15776
box -38 -48 590 592
use scs8hd_conb_1  _149_
timestamp 1586364061
transform 1 0 15364 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_147
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_158
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_162
timestamp 1586364061
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_177
timestamp 1586364061
transform 1 0 17388 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 19136 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_194
timestamp 1586364061
transform 1 0 18952 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19780 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20332 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_198
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_205
timestamp 1586364061
transform 1 0 19964 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_24_211
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_219
timestamp 1586364061
transform 1 0 21252 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_231
timestamp 1586364061
transform 1 0 22356 0 -1 15776
box -38 -48 774 592
use scs8hd_conb_1  _150_
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_242
timestamp 1586364061
transform 1 0 23368 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_254
timestamp 1586364061
transform 1 0 24472 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_266
timestamp 1586364061
transform 1 0 25576 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_137
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_141
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_154
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21528 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_218
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22724 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23092 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_233
timestamp 1586364061
transform 1 0 22540 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_237
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_241
timestamp 1586364061
transform 1 0 23276 0 1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_conb_1  _151_
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_110
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_8  FILLER_26_118
timestamp 1586364061
transform 1 0 11960 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12604 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_135
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_139
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_151
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_160
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_157
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_160
timestamp 1586364061
transform 1 0 15824 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_2  _153_
timestamp 1586364061
transform 1 0 15456 0 -1 16864
box -38 -48 406 592
use scs8hd_inv_8  _071_
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_165
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_173
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_183
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_179
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_201
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_209
timestamp 1586364061
transform 1 0 20332 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_205
timestamp 1586364061
transform 1 0 19964 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_230
timestamp 1586364061
transform 1 0 22264 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_226
timestamp 1586364061
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_243
timestamp 1586364061
transform 1 0 23460 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_260
timestamp 1586364061
transform 1 0 25024 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_262
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_266
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_272
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_274
timestamp 1586364061
transform 1 0 26312 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_127
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_6  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_160
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_172
timestamp 1586364061
transform 1 0 16928 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_176
timestamp 1586364061
transform 1 0 17296 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_189
timestamp 1586364061
transform 1 0 18492 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_201
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21068 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_220
timestamp 1586364061
transform 1 0 21344 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_226
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_229
timestamp 1586364061
transform 1 0 22172 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_241
timestamp 1586364061
transform 1 0 23276 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _166_
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_253
timestamp 1586364061
transform 1 0 24380 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_259
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_14
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_26
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_58
timestamp 1586364061
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_75
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_91
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_103
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 17952
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_134
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_138
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_151
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_157
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_161
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_176
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_205
timestamp 1586364061
transform 1 0 19964 0 1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_221
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_29_234
timestamp 1586364061
transform 1 0 22632 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_242
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_253
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 406 592
use scs8hd_buf_2  _177_
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_72
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_77
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_30_89
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_2  _176_
timestamp 1586364061
transform 1 0 9752 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_98
timestamp 1586364061
transform 1 0 10120 0 -1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_4  FILLER_30_110
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  FILLER_30_123
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_140
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 15364 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_144
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16928 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_164
timestamp 1586364061
transform 1 0 16192 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_168
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_181
timestamp 1586364061
transform 1 0 17756 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_198
timestamp 1586364061
transform 1 0 19320 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_210
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_219
timestamp 1586364061
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_223
timestamp 1586364061
transform 1 0 21620 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_buf_2  _163_
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_259
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_271
timestamp 1586364061
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _174_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_35
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_47
timestamp 1586364061
transform 1 0 5428 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_inv_8  _072_
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_139
timestamp 1586364061
transform 1 0 13892 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_153
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_157
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 866 592
use scs8hd_decap_12  FILLER_31_170
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_123
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 130 592
use scs8hd_conb_1  _144_
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_127
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_151
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_157
timestamp 1586364061
transform 1 0 15548 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 15916 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_175
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_187
timestamp 1586364061
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_199
timestamp 1586364061
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_32_211
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_193
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 774 592
use scs8hd_buf_2  _178_
timestamp 1586364061
transform 1 0 19596 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_197
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_33_203
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_34_198
timestamp 1586364061
transform 1 0 19320 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_205
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_215
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_227
timestamp 1586364061
transform 1 0 21988 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_239
timestamp 1586364061
transform 1 0 23092 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_243
timestamp 1586364061
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _172_
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_11
timestamp 1586364061
transform 1 0 2116 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_23
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_47
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _160_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_23
timestamp 1586364061
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_35
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_47
timestamp 1586364061
transform 1 0 5428 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_108
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_37_120
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_37_237
timestamp 1586364061
transform 1 0 22908 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_243
timestamp 1586364061
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_262
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_274
timestamp 1586364061
transform 1 0 26312 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_109
timestamp 1586364061
transform 1 0 11132 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_121
timestamp 1586364061
transform 1 0 12236 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_133
timestamp 1586364061
transform 1 0 13340 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22724 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_238
timestamp 1586364061
transform 1 0 23000 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_250
timestamp 1586364061
transform 1 0 24104 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_262
timestamp 1586364061
transform 1 0 25208 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_274
timestamp 1586364061
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _155_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_70
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _157_
timestamp 1586364061
transform 1 0 10304 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 10856 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_90
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_94
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_104
timestamp 1586364061
transform 1 0 10672 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_108
timestamp 1586364061
transform 1 0 11040 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_120
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _170_
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_228
timestamp 1586364061
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_39_237
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_248
timestamp 1586364061
transform 1 0 23920 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_238
timestamp 1586364061
transform 1 0 23000 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_252
timestamp 1586364061
transform 1 0 24288 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_250
timestamp 1586364061
transform 1 0 24104 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_262
timestamp 1586364061
transform 1 0 25208 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 3054 0 3110 480 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 552 480 672 6 address[1]
port 1 nsew default input
rlabel metal3 s 27520 552 28000 672 6 address[2]
port 2 nsew default input
rlabel metal2 s 4342 0 4398 480 6 address[3]
port 3 nsew default input
rlabel metal3 s 27520 1640 28000 1760 6 address[4]
port 4 nsew default input
rlabel metal3 s 27520 2864 28000 2984 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 1640 480 1760 6 address[6]
port 6 nsew default input
rlabel metal3 s 27520 5176 28000 5296 6 bottom_left_grid_pin_11_
port 7 nsew default input
rlabel metal3 s 27520 6264 28000 6384 6 bottom_left_grid_pin_13_
port 8 nsew default input
rlabel metal3 s 27520 7488 28000 7608 6 bottom_left_grid_pin_15_
port 9 nsew default input
rlabel metal2 s 5630 0 5686 480 6 bottom_left_grid_pin_1_
port 10 nsew default input
rlabel metal2 s 6918 0 6974 480 6 bottom_left_grid_pin_3_
port 11 nsew default input
rlabel metal3 s 27520 3952 28000 4072 6 bottom_left_grid_pin_5_
port 12 nsew default input
rlabel metal2 s 1030 27520 1086 28000 6 bottom_left_grid_pin_7_
port 13 nsew default input
rlabel metal3 s 0 2864 480 2984 6 bottom_left_grid_pin_9_
port 14 nsew default input
rlabel metal3 s 27520 8712 28000 8832 6 bottom_right_grid_pin_11_
port 15 nsew default input
rlabel metal3 s 27520 9800 28000 9920 6 chanx_right_in[0]
port 16 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chanx_right_in[1]
port 17 nsew default input
rlabel metal3 s 27520 11024 28000 11144 6 chanx_right_in[2]
port 18 nsew default input
rlabel metal3 s 27520 12112 28000 12232 6 chanx_right_in[3]
port 19 nsew default input
rlabel metal3 s 0 3952 480 4072 6 chanx_right_in[4]
port 20 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 chanx_right_in[5]
port 21 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chanx_right_in[6]
port 22 nsew default input
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_in[7]
port 23 nsew default input
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_in[8]
port 24 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_right_out[0]
port 25 nsew default tristate
rlabel metal2 s 10690 0 10746 480 6 chanx_right_out[1]
port 26 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_right_out[2]
port 27 nsew default tristate
rlabel metal2 s 5262 27520 5318 28000 6 chanx_right_out[3]
port 28 nsew default tristate
rlabel metal3 s 27520 15648 28000 15768 6 chanx_right_out[4]
port 29 nsew default tristate
rlabel metal2 s 7470 27520 7526 28000 6 chanx_right_out[5]
port 30 nsew default tristate
rlabel metal3 s 0 7488 480 7608 6 chanx_right_out[6]
port 31 nsew default tristate
rlabel metal3 s 27520 16872 28000 16992 6 chanx_right_out[7]
port 32 nsew default tristate
rlabel metal3 s 0 8712 480 8832 6 chanx_right_out[8]
port 33 nsew default tristate
rlabel metal2 s 9586 27520 9642 28000 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal3 s 27520 17960 28000 18080 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal2 s 13266 0 13322 480 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal3 s 27520 19184 28000 19304 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal3 s 0 15648 480 15768 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_top_in[0]
port 52 nsew default input
rlabel metal3 s 27520 21496 28000 21616 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 18326 0 18382 480 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 19614 0 19670 480 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 18234 27520 18290 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 20902 0 20958 480 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 20350 27520 20406 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal3 s 0 17960 480 18080 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 22098 0 22154 480 6 chany_top_in[8]
port 60 nsew default input
rlabel metal3 s 27520 22720 28000 22840 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal2 s 23386 0 23442 480 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal2 s 24674 0 24730 480 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 data_in
port 70 nsew default input
rlabel metal2 s 570 0 626 480 6 enable
port 71 nsew default input
rlabel metal3 s 27520 23808 28000 23928 6 right_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal3 s 0 23808 480 23928 6 right_top_grid_pin_10_
port 73 nsew default input
rlabel metal2 s 26790 27520 26846 28000 6 top_left_grid_pin_11_
port 74 nsew default input
rlabel metal3 s 0 26120 480 26240 6 top_left_grid_pin_13_
port 75 nsew default input
rlabel metal3 s 0 27344 480 27464 6 top_left_grid_pin_15_
port 76 nsew default input
rlabel metal2 s 24674 27520 24730 28000 6 top_left_grid_pin_1_
port 77 nsew default input
rlabel metal3 s 27520 25032 28000 25152 6 top_left_grid_pin_3_
port 78 nsew default input
rlabel metal3 s 27520 26120 28000 26240 6 top_left_grid_pin_5_
port 79 nsew default input
rlabel metal3 s 0 25032 480 25152 6 top_left_grid_pin_7_
port 80 nsew default input
rlabel metal2 s 27250 0 27306 480 6 top_left_grid_pin_9_
port 81 nsew default input
rlabel metal3 s 27520 27344 28000 27464 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
